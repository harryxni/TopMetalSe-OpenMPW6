magic
tech sky130A
magscale 1 2
timestamp 1608072956
<< nwell >>
rect -1947 -819 1947 819
<< pmos >>
rect -1751 -600 -1631 600
rect -1573 -600 -1453 600
rect -1395 -600 -1275 600
rect -1217 -600 -1097 600
rect -1039 -600 -919 600
rect -861 -600 -741 600
rect -683 -600 -563 600
rect -505 -600 -385 600
rect -327 -600 -207 600
rect -149 -600 -29 600
rect 29 -600 149 600
rect 207 -600 327 600
rect 385 -600 505 600
rect 563 -600 683 600
rect 741 -600 861 600
rect 919 -600 1039 600
rect 1097 -600 1217 600
rect 1275 -600 1395 600
rect 1453 -600 1573 600
rect 1631 -600 1751 600
<< pdiff >>
rect -1809 588 -1751 600
rect -1809 -588 -1797 588
rect -1763 -588 -1751 588
rect -1809 -600 -1751 -588
rect -1631 588 -1573 600
rect -1631 -588 -1619 588
rect -1585 -588 -1573 588
rect -1631 -600 -1573 -588
rect -1453 588 -1395 600
rect -1453 -588 -1441 588
rect -1407 -588 -1395 588
rect -1453 -600 -1395 -588
rect -1275 588 -1217 600
rect -1275 -588 -1263 588
rect -1229 -588 -1217 588
rect -1275 -600 -1217 -588
rect -1097 588 -1039 600
rect -1097 -588 -1085 588
rect -1051 -588 -1039 588
rect -1097 -600 -1039 -588
rect -919 588 -861 600
rect -919 -588 -907 588
rect -873 -588 -861 588
rect -919 -600 -861 -588
rect -741 588 -683 600
rect -741 -588 -729 588
rect -695 -588 -683 588
rect -741 -600 -683 -588
rect -563 588 -505 600
rect -563 -588 -551 588
rect -517 -588 -505 588
rect -563 -600 -505 -588
rect -385 588 -327 600
rect -385 -588 -373 588
rect -339 -588 -327 588
rect -385 -600 -327 -588
rect -207 588 -149 600
rect -207 -588 -195 588
rect -161 -588 -149 588
rect -207 -600 -149 -588
rect -29 588 29 600
rect -29 -588 -17 588
rect 17 -588 29 588
rect -29 -600 29 -588
rect 149 588 207 600
rect 149 -588 161 588
rect 195 -588 207 588
rect 149 -600 207 -588
rect 327 588 385 600
rect 327 -588 339 588
rect 373 -588 385 588
rect 327 -600 385 -588
rect 505 588 563 600
rect 505 -588 517 588
rect 551 -588 563 588
rect 505 -600 563 -588
rect 683 588 741 600
rect 683 -588 695 588
rect 729 -588 741 588
rect 683 -600 741 -588
rect 861 588 919 600
rect 861 -588 873 588
rect 907 -588 919 588
rect 861 -600 919 -588
rect 1039 588 1097 600
rect 1039 -588 1051 588
rect 1085 -588 1097 588
rect 1039 -600 1097 -588
rect 1217 588 1275 600
rect 1217 -588 1229 588
rect 1263 -588 1275 588
rect 1217 -600 1275 -588
rect 1395 588 1453 600
rect 1395 -588 1407 588
rect 1441 -588 1453 588
rect 1395 -600 1453 -588
rect 1573 588 1631 600
rect 1573 -588 1585 588
rect 1619 -588 1631 588
rect 1573 -600 1631 -588
rect 1751 588 1809 600
rect 1751 -588 1763 588
rect 1797 -588 1809 588
rect 1751 -600 1809 -588
<< pdiffc >>
rect -1797 -588 -1763 588
rect -1619 -588 -1585 588
rect -1441 -588 -1407 588
rect -1263 -588 -1229 588
rect -1085 -588 -1051 588
rect -907 -588 -873 588
rect -729 -588 -695 588
rect -551 -588 -517 588
rect -373 -588 -339 588
rect -195 -588 -161 588
rect -17 -588 17 588
rect 161 -588 195 588
rect 339 -588 373 588
rect 517 -588 551 588
rect 695 -588 729 588
rect 873 -588 907 588
rect 1051 -588 1085 588
rect 1229 -588 1263 588
rect 1407 -588 1441 588
rect 1585 -588 1619 588
rect 1763 -588 1797 588
<< nsubdiff >>
rect -1911 749 -1815 783
rect 1815 749 1911 783
rect -1911 687 -1877 749
rect 1877 687 1911 749
rect -1911 -749 -1877 -687
rect 1877 -749 1911 -687
rect -1911 -783 -1815 -749
rect 1815 -783 1911 -749
<< nsubdiffcont >>
rect -1815 749 1815 783
rect -1911 -687 -1877 687
rect 1877 -687 1911 687
rect -1815 -783 1815 -749
<< poly >>
rect -1751 600 -1631 688
rect -1573 600 -1453 688
rect -1395 600 -1275 688
rect -1217 600 -1097 688
rect -1039 600 -919 688
rect -861 600 -741 688
rect -683 600 -563 688
rect -505 600 -385 688
rect -327 600 -207 688
rect -149 600 -29 688
rect 29 600 149 688
rect 207 600 327 688
rect 385 600 505 688
rect 563 600 683 688
rect 741 600 861 688
rect 919 600 1039 688
rect 1097 600 1217 688
rect 1275 600 1395 688
rect 1453 600 1573 688
rect 1631 600 1751 688
rect -1751 -647 -1631 -600
rect -1751 -681 -1735 -647
rect -1647 -681 -1631 -647
rect -1751 -697 -1631 -681
rect -1573 -647 -1453 -600
rect -1573 -681 -1557 -647
rect -1469 -681 -1453 -647
rect -1573 -697 -1453 -681
rect -1395 -647 -1275 -600
rect -1395 -681 -1379 -647
rect -1291 -681 -1275 -647
rect -1395 -697 -1275 -681
rect -1217 -647 -1097 -600
rect -1217 -681 -1201 -647
rect -1113 -681 -1097 -647
rect -1217 -697 -1097 -681
rect -1039 -647 -919 -600
rect -1039 -681 -1023 -647
rect -935 -681 -919 -647
rect -1039 -697 -919 -681
rect -861 -647 -741 -600
rect -861 -681 -845 -647
rect -757 -681 -741 -647
rect -861 -697 -741 -681
rect -683 -647 -563 -600
rect -683 -681 -667 -647
rect -579 -681 -563 -647
rect -683 -697 -563 -681
rect -505 -647 -385 -600
rect -505 -681 -489 -647
rect -401 -681 -385 -647
rect -505 -697 -385 -681
rect -327 -647 -207 -600
rect -327 -681 -311 -647
rect -223 -681 -207 -647
rect -327 -697 -207 -681
rect -149 -647 -29 -600
rect -149 -681 -133 -647
rect -45 -681 -29 -647
rect -149 -697 -29 -681
rect 29 -647 149 -600
rect 29 -681 45 -647
rect 133 -681 149 -647
rect 29 -697 149 -681
rect 207 -647 327 -600
rect 207 -681 223 -647
rect 311 -681 327 -647
rect 207 -697 327 -681
rect 385 -647 505 -600
rect 385 -681 401 -647
rect 489 -681 505 -647
rect 385 -697 505 -681
rect 563 -647 683 -600
rect 563 -681 579 -647
rect 667 -681 683 -647
rect 563 -697 683 -681
rect 741 -647 861 -600
rect 741 -681 757 -647
rect 845 -681 861 -647
rect 741 -697 861 -681
rect 919 -647 1039 -600
rect 919 -681 935 -647
rect 1023 -681 1039 -647
rect 919 -697 1039 -681
rect 1097 -647 1217 -600
rect 1097 -681 1113 -647
rect 1201 -681 1217 -647
rect 1097 -697 1217 -681
rect 1275 -647 1395 -600
rect 1275 -681 1291 -647
rect 1379 -681 1395 -647
rect 1275 -697 1395 -681
rect 1453 -647 1573 -600
rect 1453 -681 1469 -647
rect 1557 -681 1573 -647
rect 1453 -697 1573 -681
rect 1631 -647 1751 -600
rect 1631 -681 1647 -647
rect 1735 -681 1751 -647
rect 1631 -697 1751 -681
<< polycont >>
rect -1735 -681 -1647 -647
rect -1557 -681 -1469 -647
rect -1379 -681 -1291 -647
rect -1201 -681 -1113 -647
rect -1023 -681 -935 -647
rect -845 -681 -757 -647
rect -667 -681 -579 -647
rect -489 -681 -401 -647
rect -311 -681 -223 -647
rect -133 -681 -45 -647
rect 45 -681 133 -647
rect 223 -681 311 -647
rect 401 -681 489 -647
rect 579 -681 667 -647
rect 757 -681 845 -647
rect 935 -681 1023 -647
rect 1113 -681 1201 -647
rect 1291 -681 1379 -647
rect 1469 -681 1557 -647
rect 1647 -681 1735 -647
<< locali >>
rect -1911 749 -1815 783
rect 1815 749 1911 783
rect -1911 687 -1877 749
rect 1877 687 1911 749
rect -1797 588 -1763 604
rect -1797 -604 -1763 -588
rect -1619 588 -1585 604
rect -1619 -604 -1585 -588
rect -1441 588 -1407 604
rect -1441 -604 -1407 -588
rect -1263 588 -1229 604
rect -1263 -604 -1229 -588
rect -1085 588 -1051 604
rect -1085 -604 -1051 -588
rect -907 588 -873 604
rect -907 -604 -873 -588
rect -729 588 -695 604
rect -729 -604 -695 -588
rect -551 588 -517 604
rect -551 -604 -517 -588
rect -373 588 -339 604
rect -373 -604 -339 -588
rect -195 588 -161 604
rect -195 -604 -161 -588
rect -17 588 17 604
rect -17 -604 17 -588
rect 161 588 195 604
rect 161 -604 195 -588
rect 339 588 373 604
rect 339 -604 373 -588
rect 517 588 551 604
rect 517 -604 551 -588
rect 695 588 729 604
rect 695 -604 729 -588
rect 873 588 907 604
rect 873 -604 907 -588
rect 1051 588 1085 604
rect 1051 -604 1085 -588
rect 1229 588 1263 604
rect 1229 -604 1263 -588
rect 1407 588 1441 604
rect 1407 -604 1441 -588
rect 1585 588 1619 604
rect 1585 -604 1619 -588
rect 1763 588 1797 604
rect 1763 -604 1797 -588
rect -1751 -681 -1735 -647
rect -1647 -681 -1631 -647
rect -1573 -681 -1557 -647
rect -1469 -681 -1453 -647
rect -1395 -681 -1379 -647
rect -1291 -681 -1275 -647
rect -1217 -681 -1201 -647
rect -1113 -681 -1097 -647
rect -1039 -681 -1023 -647
rect -935 -681 -919 -647
rect -861 -681 -845 -647
rect -757 -681 -741 -647
rect -683 -681 -667 -647
rect -579 -681 -563 -647
rect -505 -681 -489 -647
rect -401 -681 -385 -647
rect -327 -681 -311 -647
rect -223 -681 -207 -647
rect -149 -681 -133 -647
rect -45 -681 -29 -647
rect 29 -681 45 -647
rect 133 -681 149 -647
rect 207 -681 223 -647
rect 311 -681 327 -647
rect 385 -681 401 -647
rect 489 -681 505 -647
rect 563 -681 579 -647
rect 667 -681 683 -647
rect 741 -681 757 -647
rect 845 -681 861 -647
rect 919 -681 935 -647
rect 1023 -681 1039 -647
rect 1097 -681 1113 -647
rect 1201 -681 1217 -647
rect 1275 -681 1291 -647
rect 1379 -681 1395 -647
rect 1453 -681 1469 -647
rect 1557 -681 1573 -647
rect 1631 -681 1647 -647
rect 1735 -681 1751 -647
rect -1911 -749 -1877 -687
rect 1877 -749 1911 -687
rect -1911 -783 -1815 -749
rect 1815 -783 1911 -749
<< viali >>
rect -1797 -588 -1763 588
rect -1619 -588 -1585 588
rect -1441 -588 -1407 588
rect -1263 -588 -1229 588
rect -1085 -588 -1051 588
rect -907 -588 -873 588
rect -729 -588 -695 588
rect -551 -588 -517 588
rect -373 -588 -339 588
rect -195 -588 -161 588
rect -17 -588 17 588
rect 161 -588 195 588
rect 339 -588 373 588
rect 517 -588 551 588
rect 695 -588 729 588
rect 873 -588 907 588
rect 1051 -588 1085 588
rect 1229 -588 1263 588
rect 1407 -588 1441 588
rect 1585 -588 1619 588
rect 1763 -588 1797 588
rect -1735 -681 -1647 -647
rect -1557 -681 -1469 -647
rect -1379 -681 -1291 -647
rect -1201 -681 -1113 -647
rect -1023 -681 -935 -647
rect -845 -681 -757 -647
rect -667 -681 -579 -647
rect -489 -681 -401 -647
rect -311 -681 -223 -647
rect -133 -681 -45 -647
rect 45 -681 133 -647
rect 223 -681 311 -647
rect 401 -681 489 -647
rect 579 -681 667 -647
rect 757 -681 845 -647
rect 935 -681 1023 -647
rect 1113 -681 1201 -647
rect 1291 -681 1379 -647
rect 1469 -681 1557 -647
rect 1647 -681 1735 -647
<< metal1 >>
rect -1803 588 -1757 600
rect -1803 -588 -1797 588
rect -1763 -588 -1757 588
rect -1803 -600 -1757 -588
rect -1625 588 -1579 600
rect -1625 -588 -1619 588
rect -1585 -588 -1579 588
rect -1625 -600 -1579 -588
rect -1447 588 -1401 600
rect -1447 -588 -1441 588
rect -1407 -588 -1401 588
rect -1447 -600 -1401 -588
rect -1269 588 -1223 600
rect -1269 -588 -1263 588
rect -1229 -588 -1223 588
rect -1269 -600 -1223 -588
rect -1091 588 -1045 600
rect -1091 -588 -1085 588
rect -1051 -588 -1045 588
rect -1091 -600 -1045 -588
rect -913 588 -867 600
rect -913 -588 -907 588
rect -873 -588 -867 588
rect -913 -600 -867 -588
rect -735 588 -689 600
rect -735 -588 -729 588
rect -695 -588 -689 588
rect -735 -600 -689 -588
rect -557 588 -511 600
rect -557 -588 -551 588
rect -517 -588 -511 588
rect -557 -600 -511 -588
rect -379 588 -333 600
rect -379 -588 -373 588
rect -339 -588 -333 588
rect -379 -600 -333 -588
rect -201 588 -155 600
rect -201 -588 -195 588
rect -161 -588 -155 588
rect -201 -600 -155 -588
rect -23 588 23 600
rect -23 -588 -17 588
rect 17 -588 23 588
rect -23 -600 23 -588
rect 155 588 201 600
rect 155 -588 161 588
rect 195 -588 201 588
rect 155 -600 201 -588
rect 333 588 379 600
rect 333 -588 339 588
rect 373 -588 379 588
rect 333 -600 379 -588
rect 511 588 557 600
rect 511 -588 517 588
rect 551 -588 557 588
rect 511 -600 557 -588
rect 689 588 735 600
rect 689 -588 695 588
rect 729 -588 735 588
rect 689 -600 735 -588
rect 867 588 913 600
rect 867 -588 873 588
rect 907 -588 913 588
rect 867 -600 913 -588
rect 1045 588 1091 600
rect 1045 -588 1051 588
rect 1085 -588 1091 588
rect 1045 -600 1091 -588
rect 1223 588 1269 600
rect 1223 -588 1229 588
rect 1263 -588 1269 588
rect 1223 -600 1269 -588
rect 1401 588 1447 600
rect 1401 -588 1407 588
rect 1441 -588 1447 588
rect 1401 -600 1447 -588
rect 1579 588 1625 600
rect 1579 -588 1585 588
rect 1619 -588 1625 588
rect 1579 -600 1625 -588
rect 1757 588 1803 600
rect 1757 -588 1763 588
rect 1797 -588 1803 588
rect 1757 -600 1803 -588
rect -1747 -647 -1635 -641
rect -1747 -681 -1735 -647
rect -1647 -681 -1635 -647
rect -1747 -687 -1635 -681
rect -1569 -647 -1457 -641
rect -1569 -681 -1557 -647
rect -1469 -681 -1457 -647
rect -1569 -687 -1457 -681
rect -1391 -647 -1279 -641
rect -1391 -681 -1379 -647
rect -1291 -681 -1279 -647
rect -1391 -687 -1279 -681
rect -1213 -647 -1101 -641
rect -1213 -681 -1201 -647
rect -1113 -681 -1101 -647
rect -1213 -687 -1101 -681
rect -1035 -647 -923 -641
rect -1035 -681 -1023 -647
rect -935 -681 -923 -647
rect -1035 -687 -923 -681
rect -857 -647 -745 -641
rect -857 -681 -845 -647
rect -757 -681 -745 -647
rect -857 -687 -745 -681
rect -679 -647 -567 -641
rect -679 -681 -667 -647
rect -579 -681 -567 -647
rect -679 -687 -567 -681
rect -501 -647 -389 -641
rect -501 -681 -489 -647
rect -401 -681 -389 -647
rect -501 -687 -389 -681
rect -323 -647 -211 -641
rect -323 -681 -311 -647
rect -223 -681 -211 -647
rect -323 -687 -211 -681
rect -145 -647 -33 -641
rect -145 -681 -133 -647
rect -45 -681 -33 -647
rect -145 -687 -33 -681
rect 33 -647 145 -641
rect 33 -681 45 -647
rect 133 -681 145 -647
rect 33 -687 145 -681
rect 211 -647 323 -641
rect 211 -681 223 -647
rect 311 -681 323 -647
rect 211 -687 323 -681
rect 389 -647 501 -641
rect 389 -681 401 -647
rect 489 -681 501 -647
rect 389 -687 501 -681
rect 567 -647 679 -641
rect 567 -681 579 -647
rect 667 -681 679 -647
rect 567 -687 679 -681
rect 745 -647 857 -641
rect 745 -681 757 -647
rect 845 -681 857 -647
rect 745 -687 857 -681
rect 923 -647 1035 -641
rect 923 -681 935 -647
rect 1023 -681 1035 -647
rect 923 -687 1035 -681
rect 1101 -647 1213 -641
rect 1101 -681 1113 -647
rect 1201 -681 1213 -647
rect 1101 -687 1213 -681
rect 1279 -647 1391 -641
rect 1279 -681 1291 -647
rect 1379 -681 1391 -647
rect 1279 -687 1391 -681
rect 1457 -647 1569 -641
rect 1457 -681 1469 -647
rect 1557 -681 1569 -647
rect 1457 -687 1569 -681
rect 1635 -647 1747 -641
rect 1635 -681 1647 -647
rect 1735 -681 1747 -647
rect 1635 -687 1747 -681
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -1894 -766 1894 766
string parameters w 6 l 0.6 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
