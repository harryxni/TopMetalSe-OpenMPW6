magic
tech sky130A
magscale 1 2
timestamp 1608356159
<< nwell >>
rect -5124 5197 6792 5532
rect -5124 5195 5831 5197
rect -5124 5190 5094 5195
rect 3800 4122 5514 4893
rect 6289 4441 6792 5197
rect 4280 4023 4727 4122
rect 4280 3871 4475 4023
rect 6289 3947 6785 4441
<< pwell >>
rect 5563 3908 5957 3913
rect 5556 3689 5957 3908
rect 5761 3427 5957 3689
rect 5553 3253 5957 3427
rect 5563 3251 5957 3253
rect 5582 3225 5957 3251
rect 6159 3225 6802 3911
rect 5689 2805 6802 3225
rect 5650 2804 6802 2805
rect 4729 2800 6802 2804
rect -5124 2469 6802 2800
rect -5124 2464 6798 2469
<< psubdiff >>
rect 5707 3159 5767 3195
rect 6631 3159 6717 3195
rect 5711 3057 5771 3093
rect 6635 3057 6721 3093
rect 5713 2963 5773 2999
rect 6637 2963 6723 2999
rect 5713 2851 5773 2887
rect 6637 2851 6723 2887
rect -4962 2652 -4902 2692
rect -3534 2652 -3488 2692
rect -3072 2666 -3012 2706
rect -1644 2666 -1598 2706
rect -440 2676 -380 2716
rect 988 2676 1034 2716
rect 2298 2666 2358 2706
rect 3726 2666 3772 2706
rect 5265 2699 5325 2739
rect 6693 2699 6739 2739
rect -4964 2556 -4904 2596
rect -3536 2556 -3490 2596
rect -3074 2570 -3014 2610
rect -1646 2570 -1600 2610
rect -442 2580 -382 2620
rect 986 2580 1032 2620
rect 2296 2570 2356 2610
rect 3724 2570 3770 2610
rect 5263 2603 5323 2643
rect 6691 2603 6737 2643
<< nsubdiff >>
rect -4908 5400 -4866 5440
rect -3574 5400 -3540 5440
rect -2724 5404 -2682 5444
rect -1390 5404 -1356 5444
rect -92 5394 -50 5434
rect 1242 5394 1276 5434
rect 2266 5422 2308 5462
rect 3600 5422 3634 5462
rect 4795 5427 4837 5467
rect 6129 5427 6163 5467
rect -4912 5304 -4870 5344
rect -3578 5304 -3544 5344
rect -2728 5308 -2686 5348
rect -1394 5308 -1360 5348
rect -96 5298 -54 5338
rect 1238 5298 1272 5338
rect 2262 5326 2304 5366
rect 3596 5326 3630 5366
rect 4791 5331 4833 5371
rect 6125 5331 6159 5371
rect 6345 5296 6369 5375
rect 6721 5296 6745 5375
rect 6342 5142 6366 5221
rect 6718 5142 6742 5221
rect 6336 5001 6360 5080
rect 6712 5001 6736 5080
rect 6334 4845 6358 4924
rect 6710 4845 6734 4924
rect 6326 4697 6350 4776
rect 6702 4697 6726 4776
<< psubdiffcont >>
rect 5767 3159 6631 3195
rect 5771 3057 6635 3093
rect 5773 2963 6637 2999
rect 5773 2851 6637 2887
rect -4902 2652 -3534 2692
rect -3012 2666 -1644 2706
rect -380 2676 988 2716
rect 2358 2666 3726 2706
rect 5325 2699 6693 2739
rect -4904 2556 -3536 2596
rect -3014 2570 -1646 2610
rect -382 2580 986 2620
rect 2356 2570 3724 2610
rect 5323 2603 6691 2643
<< nsubdiffcont >>
rect -4866 5400 -3574 5440
rect -2682 5404 -1390 5444
rect -50 5394 1242 5434
rect 2308 5422 3600 5462
rect 4837 5427 6129 5467
rect -4870 5304 -3578 5344
rect -2686 5308 -1394 5348
rect -54 5298 1238 5338
rect 2304 5326 3596 5366
rect 4833 5331 6125 5371
rect 6369 5296 6721 5375
rect 6366 5142 6718 5221
rect 6360 5001 6712 5080
rect 6358 4845 6710 4924
rect 6350 4697 6702 4776
<< poly >>
rect 5698 4268 5728 4325
rect 5794 4268 5824 4326
rect 5698 4234 5824 4268
rect 5496 3942 5610 3958
rect 5496 3902 5512 3942
rect 5592 3925 5610 3942
rect 5773 3925 5803 4234
rect 6216 3943 6246 3958
rect 5592 3902 5803 3925
rect 5496 3891 5803 3902
rect 5496 3884 5610 3891
rect 5773 3376 5803 3891
rect 6167 3927 6246 3943
rect 6167 3893 6183 3927
rect 6217 3925 6246 3927
rect 6565 3925 6595 4408
rect 6217 3893 6595 3925
rect 6167 3891 6595 3893
rect 6167 3877 6246 3891
rect 6181 3875 6246 3877
rect 6216 3862 6246 3875
rect 6565 3490 6595 3891
<< polycont >>
rect 5512 3902 5592 3942
rect 6183 3893 6217 3927
<< locali >>
rect -4908 5400 -4866 5440
rect -3574 5400 -3540 5440
rect -2724 5410 -2710 5444
rect -1380 5410 -1342 5444
rect -1308 5410 -1278 5444
rect -2724 5404 -2682 5410
rect -1390 5404 -1356 5410
rect -92 5400 -78 5434
rect 1252 5400 1290 5434
rect 1324 5400 1354 5434
rect 2266 5428 2280 5462
rect 3610 5428 3648 5462
rect 3682 5428 3712 5462
rect 4795 5433 4809 5467
rect 6139 5433 6177 5467
rect 6211 5433 6241 5467
rect 2266 5422 2308 5428
rect 3600 5422 3634 5428
rect 4795 5427 4837 5433
rect 6129 5427 6163 5433
rect -92 5394 -50 5400
rect 1242 5394 1276 5400
rect 4791 5367 4833 5371
rect 6125 5367 6159 5371
rect 2262 5362 2304 5366
rect 3596 5362 3630 5366
rect -2728 5344 -2686 5348
rect -1394 5344 -1360 5348
rect -4912 5304 -4870 5344
rect -3578 5304 -3544 5344
rect -2728 5310 -2718 5344
rect -1388 5310 -1350 5344
rect -1316 5310 -1286 5344
rect -96 5334 -54 5338
rect 1238 5334 1272 5338
rect -2728 5308 -2686 5310
rect -1394 5308 -1360 5310
rect -96 5300 -86 5334
rect 1244 5300 1282 5334
rect 1316 5300 1346 5334
rect 2262 5328 2272 5362
rect 3602 5328 3640 5362
rect 3674 5328 3704 5362
rect 4791 5333 4801 5367
rect 6131 5333 6169 5367
rect 6203 5333 6233 5367
rect 4791 5331 4833 5333
rect 6125 5331 6159 5333
rect 2262 5326 2304 5328
rect 3596 5326 3630 5328
rect -96 5298 -54 5300
rect 1238 5298 1272 5300
rect 6353 5296 6369 5375
rect 6721 5296 6737 5375
rect 6350 5142 6366 5221
rect 6718 5142 6734 5221
rect 6344 5001 6360 5080
rect 6712 5001 6728 5080
rect 6342 4845 6358 4924
rect 6710 4845 6726 4924
rect 6334 4697 6350 4776
rect 6702 4697 6718 4776
rect 5496 3942 5610 3958
rect 5496 3902 5512 3942
rect 5592 3902 5610 3942
rect 5496 3884 5610 3902
rect 6167 3893 6183 3927
rect 6217 3893 6233 3927
rect 5707 3159 5767 3195
rect 6631 3159 6717 3195
rect 5711 3059 5721 3093
rect 5755 3059 5771 3093
rect 6635 3059 6657 3093
rect 6691 3059 6721 3093
rect 5711 3057 5771 3059
rect 6635 3057 6721 3059
rect 5713 2965 5723 2999
rect 5757 2965 5773 2999
rect 6637 2965 6659 2999
rect 6693 2965 6723 2999
rect 5713 2963 5773 2965
rect 6637 2963 6723 2965
rect 5713 2853 5723 2887
rect 5757 2853 5773 2887
rect 6637 2853 6659 2887
rect 6693 2853 6723 2887
rect 5713 2851 5773 2853
rect 6637 2851 6723 2853
rect 5265 2737 5325 2739
rect 6693 2737 6739 2739
rect -440 2714 -380 2716
rect 988 2714 1034 2716
rect -3072 2704 -3012 2706
rect -1644 2704 -1598 2706
rect -4962 2652 -4902 2692
rect -3534 2652 -3488 2692
rect -3072 2670 -3040 2704
rect -1638 2670 -1598 2704
rect -440 2680 -408 2714
rect 994 2680 1034 2714
rect -440 2676 -380 2680
rect 988 2676 1034 2680
rect 2298 2704 2358 2706
rect 3726 2704 3772 2706
rect -3072 2666 -3012 2670
rect -1644 2666 -1598 2670
rect 2298 2670 2330 2704
rect 3732 2670 3772 2704
rect 5265 2703 5297 2737
rect 6699 2703 6739 2737
rect 5265 2699 5325 2703
rect 6693 2699 6739 2703
rect 2298 2666 2358 2670
rect 3726 2666 3772 2670
rect 5263 2637 5323 2643
rect 6691 2637 6737 2643
rect -442 2614 -382 2620
rect 986 2614 1032 2620
rect -3074 2604 -3014 2610
rect -1646 2604 -1600 2610
rect -4964 2556 -4904 2596
rect -3536 2556 -3490 2596
rect -3074 2570 -3040 2604
rect -1638 2570 -1600 2604
rect -442 2580 -408 2614
rect 994 2580 1032 2614
rect 2296 2604 2356 2610
rect 3724 2604 3770 2610
rect 2296 2570 2330 2604
rect 3732 2570 3770 2604
rect 5263 2603 5297 2637
rect 6699 2603 6737 2637
<< viali >>
rect -2710 5410 -2682 5444
rect -2682 5410 -2676 5444
rect -2638 5410 -2604 5444
rect -2566 5410 -2532 5444
rect -2494 5410 -2460 5444
rect -2422 5410 -2388 5444
rect -2350 5410 -2316 5444
rect -2278 5410 -2244 5444
rect -2206 5410 -2172 5444
rect -2134 5410 -2100 5444
rect -2062 5410 -2028 5444
rect -1990 5410 -1956 5444
rect -1918 5410 -1884 5444
rect -1846 5410 -1812 5444
rect -1774 5410 -1740 5444
rect -1702 5410 -1668 5444
rect -1630 5410 -1596 5444
rect -1558 5410 -1524 5444
rect -1486 5410 -1452 5444
rect -1414 5410 -1390 5444
rect -1390 5410 -1380 5444
rect -1342 5410 -1308 5444
rect -78 5400 -50 5434
rect -50 5400 -44 5434
rect -6 5400 28 5434
rect 66 5400 100 5434
rect 138 5400 172 5434
rect 210 5400 244 5434
rect 282 5400 316 5434
rect 354 5400 388 5434
rect 426 5400 460 5434
rect 498 5400 532 5434
rect 570 5400 604 5434
rect 642 5400 676 5434
rect 714 5400 748 5434
rect 786 5400 820 5434
rect 858 5400 892 5434
rect 930 5400 964 5434
rect 1002 5400 1036 5434
rect 1074 5400 1108 5434
rect 1146 5400 1180 5434
rect 1218 5400 1242 5434
rect 1242 5400 1252 5434
rect 1290 5400 1324 5434
rect 2280 5428 2308 5462
rect 2308 5428 2314 5462
rect 2352 5428 2386 5462
rect 2424 5428 2458 5462
rect 2496 5428 2530 5462
rect 2568 5428 2602 5462
rect 2640 5428 2674 5462
rect 2712 5428 2746 5462
rect 2784 5428 2818 5462
rect 2856 5428 2890 5462
rect 2928 5428 2962 5462
rect 3000 5428 3034 5462
rect 3072 5428 3106 5462
rect 3144 5428 3178 5462
rect 3216 5428 3250 5462
rect 3288 5428 3322 5462
rect 3360 5428 3394 5462
rect 3432 5428 3466 5462
rect 3504 5428 3538 5462
rect 3576 5428 3600 5462
rect 3600 5428 3610 5462
rect 3648 5428 3682 5462
rect 4809 5433 4837 5467
rect 4837 5433 4843 5467
rect 4881 5433 4915 5467
rect 4953 5433 4987 5467
rect 5025 5433 5059 5467
rect 5097 5433 5131 5467
rect 5169 5433 5203 5467
rect 5241 5433 5275 5467
rect 5313 5433 5347 5467
rect 5385 5433 5419 5467
rect 5457 5433 5491 5467
rect 5529 5433 5563 5467
rect 5601 5433 5635 5467
rect 5673 5433 5707 5467
rect 5745 5433 5779 5467
rect 5817 5433 5851 5467
rect 5889 5433 5923 5467
rect 5961 5433 5995 5467
rect 6033 5433 6067 5467
rect 6105 5433 6129 5467
rect 6129 5433 6139 5467
rect 6177 5433 6211 5467
rect -2718 5310 -2686 5344
rect -2686 5310 -2684 5344
rect -2646 5310 -2612 5344
rect -2574 5310 -2540 5344
rect -2502 5310 -2468 5344
rect -2430 5310 -2396 5344
rect -2358 5310 -2324 5344
rect -2286 5310 -2252 5344
rect -2214 5310 -2180 5344
rect -2142 5310 -2108 5344
rect -2070 5310 -2036 5344
rect -1998 5310 -1964 5344
rect -1926 5310 -1892 5344
rect -1854 5310 -1820 5344
rect -1782 5310 -1748 5344
rect -1710 5310 -1676 5344
rect -1638 5310 -1604 5344
rect -1566 5310 -1532 5344
rect -1494 5310 -1460 5344
rect -1422 5310 -1394 5344
rect -1394 5310 -1388 5344
rect -1350 5310 -1316 5344
rect -86 5300 -54 5334
rect -54 5300 -52 5334
rect -14 5300 20 5334
rect 58 5300 92 5334
rect 130 5300 164 5334
rect 202 5300 236 5334
rect 274 5300 308 5334
rect 346 5300 380 5334
rect 418 5300 452 5334
rect 490 5300 524 5334
rect 562 5300 596 5334
rect 634 5300 668 5334
rect 706 5300 740 5334
rect 778 5300 812 5334
rect 850 5300 884 5334
rect 922 5300 956 5334
rect 994 5300 1028 5334
rect 1066 5300 1100 5334
rect 1138 5300 1172 5334
rect 1210 5300 1238 5334
rect 1238 5300 1244 5334
rect 1282 5300 1316 5334
rect 2272 5328 2304 5362
rect 2304 5328 2306 5362
rect 2344 5328 2378 5362
rect 2416 5328 2450 5362
rect 2488 5328 2522 5362
rect 2560 5328 2594 5362
rect 2632 5328 2666 5362
rect 2704 5328 2738 5362
rect 2776 5328 2810 5362
rect 2848 5328 2882 5362
rect 2920 5328 2954 5362
rect 2992 5328 3026 5362
rect 3064 5328 3098 5362
rect 3136 5328 3170 5362
rect 3208 5328 3242 5362
rect 3280 5328 3314 5362
rect 3352 5328 3386 5362
rect 3424 5328 3458 5362
rect 3496 5328 3530 5362
rect 3568 5328 3596 5362
rect 3596 5328 3602 5362
rect 3640 5328 3674 5362
rect 4801 5333 4833 5367
rect 4833 5333 4835 5367
rect 4873 5333 4907 5367
rect 4945 5333 4979 5367
rect 5017 5333 5051 5367
rect 5089 5333 5123 5367
rect 5161 5333 5195 5367
rect 5233 5333 5267 5367
rect 5305 5333 5339 5367
rect 5377 5333 5411 5367
rect 5449 5333 5483 5367
rect 5521 5333 5555 5367
rect 5593 5333 5627 5367
rect 5665 5333 5699 5367
rect 5737 5333 5771 5367
rect 5809 5333 5843 5367
rect 5881 5333 5915 5367
rect 5953 5333 5987 5367
rect 6025 5333 6059 5367
rect 6097 5333 6125 5367
rect 6125 5333 6131 5367
rect 6169 5333 6203 5367
rect 5534 4714 5984 4811
rect 5512 3902 5592 3942
rect 6183 3893 6217 3927
rect 5721 3059 5755 3093
rect 5793 3059 5827 3093
rect 5865 3059 5899 3093
rect 5937 3059 5971 3093
rect 6009 3059 6043 3093
rect 6081 3059 6115 3093
rect 6153 3059 6187 3093
rect 6225 3059 6259 3093
rect 6297 3059 6331 3093
rect 6369 3059 6403 3093
rect 6441 3059 6475 3093
rect 6513 3059 6547 3093
rect 6585 3059 6619 3093
rect 6657 3059 6691 3093
rect 5723 2965 5757 2999
rect 5795 2965 5829 2999
rect 5867 2965 5901 2999
rect 5939 2965 5973 2999
rect 6011 2965 6045 2999
rect 6083 2965 6117 2999
rect 6155 2965 6189 2999
rect 6227 2965 6261 2999
rect 6299 2965 6333 2999
rect 6371 2965 6405 2999
rect 6443 2965 6477 2999
rect 6515 2965 6549 2999
rect 6587 2965 6621 2999
rect 6659 2965 6693 2999
rect 5723 2853 5757 2887
rect 5795 2853 5829 2887
rect 5867 2853 5901 2887
rect 5939 2853 5973 2887
rect 6011 2853 6045 2887
rect 6083 2853 6117 2887
rect 6155 2853 6189 2887
rect 6227 2853 6261 2887
rect 6299 2853 6333 2887
rect 6371 2853 6405 2887
rect 6443 2853 6477 2887
rect 6515 2853 6549 2887
rect 6587 2853 6621 2887
rect 6659 2853 6693 2887
rect -3040 2670 -3012 2704
rect -3012 2670 -3006 2704
rect -2968 2670 -2934 2704
rect -2896 2670 -2862 2704
rect -2824 2670 -2790 2704
rect -2752 2670 -2718 2704
rect -2680 2670 -2646 2704
rect -2608 2670 -2574 2704
rect -2536 2670 -2502 2704
rect -2464 2670 -2430 2704
rect -2392 2670 -2358 2704
rect -2320 2670 -2286 2704
rect -2248 2670 -2214 2704
rect -2176 2670 -2142 2704
rect -2104 2670 -2070 2704
rect -2032 2670 -1998 2704
rect -1960 2670 -1926 2704
rect -1888 2670 -1854 2704
rect -1816 2670 -1782 2704
rect -1744 2670 -1710 2704
rect -1672 2670 -1644 2704
rect -1644 2670 -1638 2704
rect -408 2680 -380 2714
rect -380 2680 -374 2714
rect -336 2680 -302 2714
rect -264 2680 -230 2714
rect -192 2680 -158 2714
rect -120 2680 -86 2714
rect -48 2680 -14 2714
rect 24 2680 58 2714
rect 96 2680 130 2714
rect 168 2680 202 2714
rect 240 2680 274 2714
rect 312 2680 346 2714
rect 384 2680 418 2714
rect 456 2680 490 2714
rect 528 2680 562 2714
rect 600 2680 634 2714
rect 672 2680 706 2714
rect 744 2680 778 2714
rect 816 2680 850 2714
rect 888 2680 922 2714
rect 960 2680 988 2714
rect 988 2680 994 2714
rect 2330 2670 2358 2704
rect 2358 2670 2364 2704
rect 2402 2670 2436 2704
rect 2474 2670 2508 2704
rect 2546 2670 2580 2704
rect 2618 2670 2652 2704
rect 2690 2670 2724 2704
rect 2762 2670 2796 2704
rect 2834 2670 2868 2704
rect 2906 2670 2940 2704
rect 2978 2670 3012 2704
rect 3050 2670 3084 2704
rect 3122 2670 3156 2704
rect 3194 2670 3228 2704
rect 3266 2670 3300 2704
rect 3338 2670 3372 2704
rect 3410 2670 3444 2704
rect 3482 2670 3516 2704
rect 3554 2670 3588 2704
rect 3626 2670 3660 2704
rect 3698 2670 3726 2704
rect 3726 2670 3732 2704
rect 5297 2703 5325 2737
rect 5325 2703 5331 2737
rect 5369 2703 5403 2737
rect 5441 2703 5475 2737
rect 5513 2703 5547 2737
rect 5585 2703 5619 2737
rect 5657 2703 5691 2737
rect 5729 2703 5763 2737
rect 5801 2703 5835 2737
rect 5873 2703 5907 2737
rect 5945 2703 5979 2737
rect 6017 2703 6051 2737
rect 6089 2703 6123 2737
rect 6161 2703 6195 2737
rect 6233 2703 6267 2737
rect 6305 2703 6339 2737
rect 6377 2703 6411 2737
rect 6449 2703 6483 2737
rect 6521 2703 6555 2737
rect 6593 2703 6627 2737
rect 6665 2703 6693 2737
rect 6693 2703 6699 2737
rect -3040 2570 -3014 2604
rect -3014 2570 -3006 2604
rect -2968 2570 -2934 2604
rect -2896 2570 -2862 2604
rect -2824 2570 -2790 2604
rect -2752 2570 -2718 2604
rect -2680 2570 -2646 2604
rect -2608 2570 -2574 2604
rect -2536 2570 -2502 2604
rect -2464 2570 -2430 2604
rect -2392 2570 -2358 2604
rect -2320 2570 -2286 2604
rect -2248 2570 -2214 2604
rect -2176 2570 -2142 2604
rect -2104 2570 -2070 2604
rect -2032 2570 -1998 2604
rect -1960 2570 -1926 2604
rect -1888 2570 -1854 2604
rect -1816 2570 -1782 2604
rect -1744 2570 -1710 2604
rect -1672 2570 -1646 2604
rect -1646 2570 -1638 2604
rect -408 2580 -382 2614
rect -382 2580 -374 2614
rect -336 2580 -302 2614
rect -264 2580 -230 2614
rect -192 2580 -158 2614
rect -120 2580 -86 2614
rect -48 2580 -14 2614
rect 24 2580 58 2614
rect 96 2580 130 2614
rect 168 2580 202 2614
rect 240 2580 274 2614
rect 312 2580 346 2614
rect 384 2580 418 2614
rect 456 2580 490 2614
rect 528 2580 562 2614
rect 600 2580 634 2614
rect 672 2580 706 2614
rect 744 2580 778 2614
rect 816 2580 850 2614
rect 888 2580 922 2614
rect 960 2580 986 2614
rect 986 2580 994 2614
rect 2330 2570 2356 2604
rect 2356 2570 2364 2604
rect 2402 2570 2436 2604
rect 2474 2570 2508 2604
rect 2546 2570 2580 2604
rect 2618 2570 2652 2604
rect 2690 2570 2724 2604
rect 2762 2570 2796 2604
rect 2834 2570 2868 2604
rect 2906 2570 2940 2604
rect 2978 2570 3012 2604
rect 3050 2570 3084 2604
rect 3122 2570 3156 2604
rect 3194 2570 3228 2604
rect 3266 2570 3300 2604
rect 3338 2570 3372 2604
rect 3410 2570 3444 2604
rect 3482 2570 3516 2604
rect 3554 2570 3588 2604
rect 3626 2570 3660 2604
rect 3698 2570 3724 2604
rect 3724 2570 3732 2604
rect 5297 2603 5323 2637
rect 5323 2603 5331 2637
rect 5369 2603 5403 2637
rect 5441 2603 5475 2637
rect 5513 2603 5547 2637
rect 5585 2603 5619 2637
rect 5657 2603 5691 2637
rect 5729 2603 5763 2637
rect 5801 2603 5835 2637
rect 5873 2603 5907 2637
rect 5945 2603 5979 2637
rect 6017 2603 6051 2637
rect 6089 2603 6123 2637
rect 6161 2603 6195 2637
rect 6233 2603 6267 2637
rect 6305 2603 6339 2637
rect 6377 2603 6411 2637
rect 6449 2603 6483 2637
rect 6521 2603 6555 2637
rect 6593 2603 6627 2637
rect 6665 2603 6691 2637
rect 6691 2603 6699 2637
<< metal1 >>
rect -5122 5467 6790 5516
rect -5122 5462 4809 5467
rect -5122 5444 2280 5462
rect -5122 5410 -2710 5444
rect -2676 5410 -2638 5444
rect -2604 5410 -2566 5444
rect -2532 5410 -2494 5444
rect -2460 5410 -2422 5444
rect -2388 5410 -2350 5444
rect -2316 5410 -2278 5444
rect -2244 5410 -2206 5444
rect -2172 5410 -2134 5444
rect -2100 5410 -2062 5444
rect -2028 5410 -1990 5444
rect -1956 5410 -1918 5444
rect -1884 5410 -1846 5444
rect -1812 5410 -1774 5444
rect -1740 5410 -1702 5444
rect -1668 5410 -1630 5444
rect -1596 5410 -1558 5444
rect -1524 5410 -1486 5444
rect -1452 5410 -1414 5444
rect -1380 5410 -1342 5444
rect -1308 5434 2280 5444
rect -1308 5410 -78 5434
rect -5122 5400 -78 5410
rect -44 5400 -6 5434
rect 28 5400 66 5434
rect 100 5400 138 5434
rect 172 5400 210 5434
rect 244 5400 282 5434
rect 316 5400 354 5434
rect 388 5400 426 5434
rect 460 5400 498 5434
rect 532 5400 570 5434
rect 604 5400 642 5434
rect 676 5400 714 5434
rect 748 5400 786 5434
rect 820 5400 858 5434
rect 892 5400 930 5434
rect 964 5400 1002 5434
rect 1036 5400 1074 5434
rect 1108 5400 1146 5434
rect 1180 5400 1218 5434
rect 1252 5400 1290 5434
rect 1324 5428 2280 5434
rect 2314 5428 2352 5462
rect 2386 5428 2424 5462
rect 2458 5428 2496 5462
rect 2530 5428 2568 5462
rect 2602 5428 2640 5462
rect 2674 5428 2712 5462
rect 2746 5428 2784 5462
rect 2818 5428 2856 5462
rect 2890 5428 2928 5462
rect 2962 5428 3000 5462
rect 3034 5428 3072 5462
rect 3106 5428 3144 5462
rect 3178 5428 3216 5462
rect 3250 5428 3288 5462
rect 3322 5428 3360 5462
rect 3394 5428 3432 5462
rect 3466 5428 3504 5462
rect 3538 5428 3576 5462
rect 3610 5428 3648 5462
rect 3682 5433 4809 5462
rect 4843 5433 4881 5467
rect 4915 5433 4953 5467
rect 4987 5433 5025 5467
rect 5059 5433 5097 5467
rect 5131 5433 5169 5467
rect 5203 5433 5241 5467
rect 5275 5433 5313 5467
rect 5347 5433 5385 5467
rect 5419 5433 5457 5467
rect 5491 5433 5529 5467
rect 5563 5433 5601 5467
rect 5635 5433 5673 5467
rect 5707 5433 5745 5467
rect 5779 5433 5817 5467
rect 5851 5433 5889 5467
rect 5923 5433 5961 5467
rect 5995 5433 6033 5467
rect 6067 5433 6105 5467
rect 6139 5433 6177 5467
rect 6211 5433 6790 5467
rect 3682 5428 6790 5433
rect 1324 5400 6790 5428
rect -5122 5367 6790 5400
rect -5122 5362 4801 5367
rect -5122 5344 2272 5362
rect -5122 5310 -2718 5344
rect -2684 5310 -2646 5344
rect -2612 5310 -2574 5344
rect -2540 5310 -2502 5344
rect -2468 5310 -2430 5344
rect -2396 5310 -2358 5344
rect -2324 5310 -2286 5344
rect -2252 5310 -2214 5344
rect -2180 5310 -2142 5344
rect -2108 5310 -2070 5344
rect -2036 5310 -1998 5344
rect -1964 5310 -1926 5344
rect -1892 5310 -1854 5344
rect -1820 5310 -1782 5344
rect -1748 5310 -1710 5344
rect -1676 5310 -1638 5344
rect -1604 5310 -1566 5344
rect -1532 5310 -1494 5344
rect -1460 5310 -1422 5344
rect -1388 5310 -1350 5344
rect -1316 5334 2272 5344
rect -1316 5310 -86 5334
rect -5122 5300 -86 5310
rect -52 5300 -14 5334
rect 20 5300 58 5334
rect 92 5300 130 5334
rect 164 5300 202 5334
rect 236 5300 274 5334
rect 308 5300 346 5334
rect 380 5300 418 5334
rect 452 5300 490 5334
rect 524 5300 562 5334
rect 596 5300 634 5334
rect 668 5300 706 5334
rect 740 5300 778 5334
rect 812 5300 850 5334
rect 884 5300 922 5334
rect 956 5300 994 5334
rect 1028 5300 1066 5334
rect 1100 5300 1138 5334
rect 1172 5300 1210 5334
rect 1244 5300 1282 5334
rect 1316 5328 2272 5334
rect 2306 5328 2344 5362
rect 2378 5328 2416 5362
rect 2450 5328 2488 5362
rect 2522 5328 2560 5362
rect 2594 5328 2632 5362
rect 2666 5328 2704 5362
rect 2738 5328 2776 5362
rect 2810 5328 2848 5362
rect 2882 5328 2920 5362
rect 2954 5328 2992 5362
rect 3026 5328 3064 5362
rect 3098 5328 3136 5362
rect 3170 5328 3208 5362
rect 3242 5328 3280 5362
rect 3314 5328 3352 5362
rect 3386 5328 3424 5362
rect 3458 5328 3496 5362
rect 3530 5328 3568 5362
rect 3602 5328 3640 5362
rect 3674 5333 4801 5362
rect 4835 5333 4873 5367
rect 4907 5333 4945 5367
rect 4979 5333 5017 5367
rect 5051 5333 5089 5367
rect 5123 5333 5161 5367
rect 5195 5333 5233 5367
rect 5267 5333 5305 5367
rect 5339 5333 5377 5367
rect 5411 5333 5449 5367
rect 5483 5333 5521 5367
rect 5555 5333 5593 5367
rect 5627 5333 5665 5367
rect 5699 5333 5737 5367
rect 5771 5333 5809 5367
rect 5843 5333 5881 5367
rect 5915 5333 5953 5367
rect 5987 5333 6025 5367
rect 6059 5333 6097 5367
rect 6131 5333 6169 5367
rect 6203 5333 6790 5367
rect 3674 5328 6790 5333
rect 1316 5300 6790 5328
rect -5122 5199 6790 5300
rect -5122 5198 -3779 5199
rect -3442 5198 6790 5199
rect -4874 5053 -4832 5198
rect -4804 5082 -4794 5142
rect -4734 5082 -4724 5142
rect -4874 5051 -4804 5053
rect -4874 4888 -4790 5051
rect -210 5049 -134 5198
rect -103 5077 -93 5137
rect -33 5077 -23 5137
rect -4726 5040 -4470 5046
rect -4736 5032 -4470 5040
rect -4740 4882 -4730 5032
rect -4674 4882 -4470 5032
rect -4896 3112 -4822 3114
rect -4898 2932 -4822 3112
rect -4736 3109 -4470 4882
rect -210 5036 -106 5049
rect -210 4761 -87 5036
rect -32 5035 -1 5039
rect -32 4220 135 5035
rect -29 4207 135 4220
rect 3939 4817 5989 4818
rect 3939 4811 5996 4817
rect 3939 4714 5534 4811
rect 5984 4714 5996 4811
rect 3939 4708 5996 4714
rect 6298 4711 6790 5198
rect 3939 4680 5989 4708
rect 3939 4570 5422 4680
rect 5738 4597 5784 4680
rect 3939 4121 4311 4570
rect 6298 4456 6788 4711
rect 5642 4229 5688 4355
rect 5836 4347 5875 4352
rect 5833 4229 5878 4347
rect 5642 4183 5878 4229
rect 5833 4065 5878 4183
rect 6517 4165 6551 4456
rect 4936 3930 4946 4016
rect 5118 4002 5128 4016
rect 5118 3958 5605 4002
rect 5118 3944 5610 3958
rect 5118 3930 5128 3944
rect 5494 3942 5610 3944
rect 5494 3902 5512 3942
rect 5592 3902 5610 3942
rect 5494 3884 5610 3902
rect 5815 3927 5878 4065
rect 6089 3927 6099 3944
rect 6220 3943 6230 3944
rect 6221 3927 6231 3943
rect 5815 3891 6099 3927
rect 6221 3925 6246 3927
rect 6607 3925 6639 4355
rect 5504 3881 5562 3884
rect -4077 3714 -4067 3864
rect -3917 3828 -3907 3864
rect -3917 3754 -3803 3828
rect 4209 3754 4628 3828
rect -3917 3714 -3907 3754
rect 4231 3660 4498 3691
rect 4231 3645 4254 3660
rect 4227 3590 4254 3645
rect 4244 3574 4254 3590
rect 4340 3636 4498 3660
rect 4340 3590 4351 3636
rect 4340 3574 4350 3590
rect 5352 3519 5756 3583
rect -4767 2937 -4470 3109
rect -4736 2935 -4470 2937
rect -179 2943 -89 3157
rect -47 2959 -37 3157
rect 76 2959 86 3157
rect -4898 2804 -4862 2932
rect -4834 2848 -4824 2902
rect -4764 2848 -4754 2902
rect -3768 2804 -3732 2805
rect -179 2804 -137 2943
rect -94 2906 -20 2912
rect -94 2854 -84 2906
rect -32 2866 -20 2906
rect -32 2854 -22 2866
rect 204 2804 379 3501
rect 4650 2804 5165 3414
rect 5352 3155 5416 3519
rect 5815 3479 5849 3891
rect 6089 3874 6099 3891
rect 6221 3891 6250 3925
rect 6607 3891 6897 3925
rect 6221 3875 6231 3891
rect 6220 3874 6230 3875
rect 6607 3531 6639 3891
rect 5900 3356 5957 3424
rect 6513 3422 6559 3531
rect 5649 3225 5957 3356
rect 6159 3225 6800 3422
rect 5342 2979 5352 3155
rect 5416 2979 5426 3155
rect 5650 3093 6802 3225
rect 5650 3059 5721 3093
rect 5755 3059 5793 3093
rect 5827 3059 5865 3093
rect 5899 3059 5937 3093
rect 5971 3059 6009 3093
rect 6043 3059 6081 3093
rect 6115 3059 6153 3093
rect 6187 3059 6225 3093
rect 6259 3059 6297 3093
rect 6331 3059 6369 3093
rect 6403 3059 6441 3093
rect 6475 3059 6513 3093
rect 6547 3059 6585 3093
rect 6619 3059 6657 3093
rect 6691 3059 6802 3093
rect 5650 2999 6802 3059
rect 5650 2965 5723 2999
rect 5757 2965 5795 2999
rect 5829 2965 5867 2999
rect 5901 2965 5939 2999
rect 5973 2965 6011 2999
rect 6045 2965 6083 2999
rect 6117 2965 6155 2999
rect 6189 2965 6227 2999
rect 6261 2965 6299 2999
rect 6333 2965 6371 2999
rect 6405 2965 6443 2999
rect 6477 2965 6515 2999
rect 6549 2965 6587 2999
rect 6621 2965 6659 2999
rect 6693 2965 6802 2999
rect 5650 2887 6802 2965
rect 5650 2853 5723 2887
rect 5757 2853 5795 2887
rect 5829 2853 5867 2887
rect 5901 2853 5939 2887
rect 5973 2853 6011 2887
rect 6045 2853 6083 2887
rect 6117 2853 6155 2887
rect 6189 2853 6227 2887
rect 6261 2853 6299 2887
rect 6333 2853 6371 2887
rect 6405 2853 6443 2887
rect 6477 2853 6515 2887
rect 6549 2853 6587 2887
rect 6621 2853 6659 2887
rect 6693 2853 6802 2887
rect 5650 2804 6802 2853
rect -5118 2737 6804 2804
rect -5118 2714 5297 2737
rect -5118 2704 -408 2714
rect -5118 2670 -3040 2704
rect -3006 2670 -2968 2704
rect -2934 2670 -2896 2704
rect -2862 2670 -2824 2704
rect -2790 2670 -2752 2704
rect -2718 2670 -2680 2704
rect -2646 2670 -2608 2704
rect -2574 2670 -2536 2704
rect -2502 2670 -2464 2704
rect -2430 2670 -2392 2704
rect -2358 2670 -2320 2704
rect -2286 2670 -2248 2704
rect -2214 2670 -2176 2704
rect -2142 2670 -2104 2704
rect -2070 2670 -2032 2704
rect -1998 2670 -1960 2704
rect -1926 2670 -1888 2704
rect -1854 2670 -1816 2704
rect -1782 2670 -1744 2704
rect -1710 2670 -1672 2704
rect -1638 2680 -408 2704
rect -374 2680 -336 2714
rect -302 2680 -264 2714
rect -230 2680 -192 2714
rect -158 2680 -120 2714
rect -86 2680 -48 2714
rect -14 2680 24 2714
rect 58 2680 96 2714
rect 130 2680 168 2714
rect 202 2680 240 2714
rect 274 2680 312 2714
rect 346 2680 384 2714
rect 418 2680 456 2714
rect 490 2680 528 2714
rect 562 2680 600 2714
rect 634 2680 672 2714
rect 706 2680 744 2714
rect 778 2680 816 2714
rect 850 2680 888 2714
rect 922 2680 960 2714
rect 994 2704 5297 2714
rect 994 2680 2330 2704
rect -1638 2670 2330 2680
rect 2364 2670 2402 2704
rect 2436 2670 2474 2704
rect 2508 2670 2546 2704
rect 2580 2670 2618 2704
rect 2652 2670 2690 2704
rect 2724 2670 2762 2704
rect 2796 2670 2834 2704
rect 2868 2670 2906 2704
rect 2940 2670 2978 2704
rect 3012 2670 3050 2704
rect 3084 2670 3122 2704
rect 3156 2670 3194 2704
rect 3228 2670 3266 2704
rect 3300 2670 3338 2704
rect 3372 2670 3410 2704
rect 3444 2670 3482 2704
rect 3516 2670 3554 2704
rect 3588 2670 3626 2704
rect 3660 2670 3698 2704
rect 3732 2703 5297 2704
rect 5331 2703 5369 2737
rect 5403 2703 5441 2737
rect 5475 2703 5513 2737
rect 5547 2703 5585 2737
rect 5619 2703 5657 2737
rect 5691 2703 5729 2737
rect 5763 2703 5801 2737
rect 5835 2703 5873 2737
rect 5907 2703 5945 2737
rect 5979 2703 6017 2737
rect 6051 2703 6089 2737
rect 6123 2703 6161 2737
rect 6195 2703 6233 2737
rect 6267 2703 6305 2737
rect 6339 2703 6377 2737
rect 6411 2703 6449 2737
rect 6483 2703 6521 2737
rect 6555 2703 6593 2737
rect 6627 2703 6665 2737
rect 6699 2703 6804 2737
rect 3732 2670 6804 2703
rect -5118 2637 6804 2670
rect -5118 2624 5297 2637
rect -5114 2614 5297 2624
rect -5114 2604 -408 2614
rect -5114 2570 -3040 2604
rect -3006 2570 -2968 2604
rect -2934 2570 -2896 2604
rect -2862 2570 -2824 2604
rect -2790 2570 -2752 2604
rect -2718 2570 -2680 2604
rect -2646 2570 -2608 2604
rect -2574 2570 -2536 2604
rect -2502 2570 -2464 2604
rect -2430 2570 -2392 2604
rect -2358 2570 -2320 2604
rect -2286 2570 -2248 2604
rect -2214 2570 -2176 2604
rect -2142 2570 -2104 2604
rect -2070 2570 -2032 2604
rect -1998 2570 -1960 2604
rect -1926 2570 -1888 2604
rect -1854 2570 -1816 2604
rect -1782 2570 -1744 2604
rect -1710 2570 -1672 2604
rect -1638 2580 -408 2604
rect -374 2580 -336 2614
rect -302 2580 -264 2614
rect -230 2580 -192 2614
rect -158 2580 -120 2614
rect -86 2580 -48 2614
rect -14 2580 24 2614
rect 58 2580 96 2614
rect 130 2580 168 2614
rect 202 2580 240 2614
rect 274 2580 312 2614
rect 346 2580 384 2614
rect 418 2580 456 2614
rect 490 2580 528 2614
rect 562 2580 600 2614
rect 634 2580 672 2614
rect 706 2580 744 2614
rect 778 2580 816 2614
rect 850 2580 888 2614
rect 922 2580 960 2614
rect 994 2604 5297 2614
rect 994 2580 2330 2604
rect -1638 2570 2330 2580
rect 2364 2570 2402 2604
rect 2436 2570 2474 2604
rect 2508 2570 2546 2604
rect 2580 2570 2618 2604
rect 2652 2570 2690 2604
rect 2724 2570 2762 2604
rect 2796 2570 2834 2604
rect 2868 2570 2906 2604
rect 2940 2570 2978 2604
rect 3012 2570 3050 2604
rect 3084 2570 3122 2604
rect 3156 2570 3194 2604
rect 3228 2570 3266 2604
rect 3300 2570 3338 2604
rect 3372 2570 3410 2604
rect 3444 2570 3482 2604
rect 3516 2570 3554 2604
rect 3588 2570 3626 2604
rect 3660 2570 3698 2604
rect 3732 2603 5297 2604
rect 5331 2603 5369 2637
rect 5403 2603 5441 2637
rect 5475 2603 5513 2637
rect 5547 2603 5585 2637
rect 5619 2603 5657 2637
rect 5691 2603 5729 2637
rect 5763 2603 5801 2637
rect 5835 2603 5873 2637
rect 5907 2603 5945 2637
rect 5979 2603 6017 2637
rect 6051 2603 6089 2637
rect 6123 2603 6161 2637
rect 6195 2603 6233 2637
rect 6267 2603 6305 2637
rect 6339 2603 6377 2637
rect 6411 2603 6449 2637
rect 6483 2603 6521 2637
rect 6555 2603 6593 2637
rect 6627 2603 6665 2637
rect 6699 2603 6804 2637
rect 3732 2570 6804 2603
rect -5114 2462 6804 2570
<< via1 >>
rect -4794 5082 -4734 5142
rect -93 5077 -33 5137
rect -4730 4882 -4674 5032
rect 4946 3930 5118 4016
rect 6099 3943 6220 3944
rect 6099 3927 6221 3943
rect 6099 3893 6183 3927
rect 6183 3893 6217 3927
rect 6217 3893 6221 3927
rect -4067 3714 -3917 3864
rect 4254 3574 4340 3660
rect -37 2959 76 3157
rect -4824 2848 -4764 2902
rect -84 2854 -32 2906
rect 6099 3875 6221 3893
rect 6099 3874 6220 3875
rect 5352 2979 5416 3155
<< metal2 >>
rect -4794 5148 -4734 5152
rect -4802 5144 -4734 5148
rect -93 5144 -33 5147
rect -4802 5142 -31 5144
rect -4802 5090 -4794 5142
rect -4796 5086 -4794 5090
rect -4734 5137 -31 5142
rect -4734 5086 -93 5137
rect -4794 5072 -4734 5082
rect -4696 5042 -4658 5086
rect -33 5086 -31 5137
rect -93 5067 -33 5077
rect -4730 5032 -4658 5042
rect -4674 4884 -4658 5032
rect -4730 4872 -4674 4882
rect 979 4879 6229 5029
rect 979 4558 1148 4879
rect -4067 4408 1148 4558
rect -4067 3864 -3917 4408
rect 4946 4016 5118 4026
rect 4946 3920 5118 3930
rect 6079 3959 6229 4879
rect 6079 3944 6233 3959
rect 6079 3874 6099 3944
rect 6220 3943 6233 3944
rect 6221 3875 6233 3943
rect 6220 3874 6233 3875
rect 6079 3850 6233 3874
rect 6151 3847 6233 3850
rect -4067 3704 -3917 3714
rect 4254 3660 4340 3670
rect 3 3624 105 3660
rect -39 3157 105 3624
rect 4163 3574 4254 3660
rect 4197 3564 4340 3574
rect -39 2959 -37 3157
rect 76 2959 104 3157
rect 4197 3112 4283 3564
rect 4499 3314 4555 3753
rect 4499 3258 6895 3314
rect 5352 3155 5416 3165
rect 4197 3026 5352 3112
rect 5352 2969 5416 2979
rect -39 2952 104 2959
rect -37 2949 76 2952
rect -4824 2910 -4764 2912
rect -4836 2909 -4764 2910
rect -84 2909 -32 2916
rect -4836 2906 -22 2909
rect -4836 2902 -84 2906
rect -4836 2848 -4824 2902
rect -4764 2854 -84 2902
rect -32 2854 -22 2906
rect -4764 2853 -22 2854
rect -4824 2838 -4764 2848
rect -84 2844 -32 2853
use sky130_fd_pr__nfet_01v8_X8MMG7  sky130_fd_pr__nfet_01v8_X8MMG7_0
timestamp 1608352057
transform -1 0 -64 0 -1 3066
box -211 -329 211 329
use via_li_m1  via_li_m1_1
array 0 19 72 0 0 74
timestamp 1606675505
transform 1 0 -4942 0 1 2536
box 4 0 76 74
use via_li_m1  via_li_m1_0
array 0 19 72 0 0 74
timestamp 1606675505
transform 1 0 -4942 0 1 2636
box 4 0 76 74
use sky130_fd_pr__nfet_01v8_YK3456  sky130_fd_pr__nfet_01v8_YK3456_0
timestamp 1608249442
transform -1 0 -4795 0 -1 3024
box -211 -300 211 300
use sky130_fd_pr__nfet_01v8_8GKXY7  sky130_fd_pr__nfet_01v8_8GKXY7_0
timestamp 1608351071
transform 1 0 6580 0 1 3561
box -211 -208 211 208
use sky130_fd_pr__pfet_01v8_5UMBUD  sky130_fd_pr__pfet_01v8_5UMBUD_0
timestamp 1608350919
transform 1 0 6580 0 1 4245
box -211 -298 211 298
use via_li_m1  via_li_m1_4
array 0 13 72 0 0 74
timestamp 1606675505
transform 1 0 5705 0 1 3141
box 4 0 76 74
use sky130_fd_pr__nfet_01v8_R7545W  sky130_fd_pr__nfet_01v8_R7545W_0
timestamp 1608229183
transform 1 0 5788 0 1 3563
box -211 -330 211 330
use inverter  inverter_1
array 0 18 430 0 0 936
timestamp 1608352248
transform 1 0 1365 0 1 3178
box -5252 188 -4822 1124
use sky130_fd_pr__pfet_01v8_5U9U2E  sky130_fd_pr__pfet_01v8_5U9U2E_0
timestamp 1608350448
transform 1 0 5761 0 1 4476
box -263 -369 263 369
use via_li_m1  via_li_m1_3
array 0 19 72 0 0 74
timestamp 1606675505
transform 1 0 -4914 0 1 5286
box 4 0 76 74
use via_li_m1  via_li_m1_2
array 0 19 72 0 0 74
timestamp 1606675505
transform 1 0 -4906 0 1 5386
box 4 0 76 74
use sky130_fd_pr__pfet_01v8_JRPBUD  sky130_fd_pr__pfet_01v8_JRPBUD_0
timestamp 1608343268
transform 1 0 -57 0 1 4935
box -211 -334 211 334
use sky130_fd_pr__pfet_01v8_35M7SP  sky130_fd_pr__pfet_01v8_35M7SP_0
timestamp 1608253040
transform 1 0 -4755 0 1 4963
box -211 -309 211 309
use nand  nand_0
timestamp 1608325973
transform 1 0 4710 0 1 4083
box -267 -910 511 767
<< labels >>
rlabel metal1 -5114 2462 -3040 2804 1 vss
rlabel metal1 -5122 5198 -2718 5516 1 vdd
rlabel metal2 -4734 5086 -93 5144 1 5
rlabel space -32 4122 135 5035 1 10
rlabel space 5815 3891 6246 3927 1 out_ring
rlabel metal1 6607 3891 6897 3925 1 out_vco
rlabel metal2 4499 3258 6895 3314 1 en
rlabel space 204 2714 379 3510 1 9
rlabel metal2 -4764 2853 -99 2909 1 in
<< end >>
