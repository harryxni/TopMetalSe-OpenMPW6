magic
tech sky130A
magscale 1 2
timestamp 1654643737
<< error_p >>
rect -1445 71 -1387 77
rect -1327 71 -1269 77
rect -1209 71 -1151 77
rect -1091 71 -1033 77
rect -973 71 -915 77
rect -855 71 -797 77
rect -737 71 -679 77
rect -619 71 -561 77
rect -501 71 -443 77
rect -383 71 -325 77
rect -265 71 -207 77
rect -147 71 -89 77
rect -29 71 29 77
rect 89 71 147 77
rect 207 71 265 77
rect 325 71 383 77
rect 443 71 501 77
rect 561 71 619 77
rect 679 71 737 77
rect 797 71 855 77
rect 915 71 973 77
rect 1033 71 1091 77
rect 1151 71 1209 77
rect 1269 71 1327 77
rect 1387 71 1445 77
rect -1445 37 -1433 71
rect -1327 37 -1315 71
rect -1209 37 -1197 71
rect -1091 37 -1079 71
rect -973 37 -961 71
rect -855 37 -843 71
rect -737 37 -725 71
rect -619 37 -607 71
rect -501 37 -489 71
rect -383 37 -371 71
rect -265 37 -253 71
rect -147 37 -135 71
rect -29 37 -17 71
rect 89 37 101 71
rect 207 37 219 71
rect 325 37 337 71
rect 443 37 455 71
rect 561 37 573 71
rect 679 37 691 71
rect 797 37 809 71
rect 915 37 927 71
rect 1033 37 1045 71
rect 1151 37 1163 71
rect 1269 37 1281 71
rect 1387 37 1399 71
rect -1445 31 -1387 37
rect -1327 31 -1269 37
rect -1209 31 -1151 37
rect -1091 31 -1033 37
rect -973 31 -915 37
rect -855 31 -797 37
rect -737 31 -679 37
rect -619 31 -561 37
rect -501 31 -443 37
rect -383 31 -325 37
rect -265 31 -207 37
rect -147 31 -89 37
rect -29 31 29 37
rect 89 31 147 37
rect 207 31 265 37
rect 325 31 383 37
rect 443 31 501 37
rect 561 31 619 37
rect 679 31 737 37
rect 797 31 855 37
rect 915 31 973 37
rect 1033 31 1091 37
rect 1151 31 1209 37
rect 1269 31 1327 37
rect 1387 31 1445 37
rect -1445 -37 -1387 -31
rect -1327 -37 -1269 -31
rect -1209 -37 -1151 -31
rect -1091 -37 -1033 -31
rect -973 -37 -915 -31
rect -855 -37 -797 -31
rect -737 -37 -679 -31
rect -619 -37 -561 -31
rect -501 -37 -443 -31
rect -383 -37 -325 -31
rect -265 -37 -207 -31
rect -147 -37 -89 -31
rect -29 -37 29 -31
rect 89 -37 147 -31
rect 207 -37 265 -31
rect 325 -37 383 -31
rect 443 -37 501 -31
rect 561 -37 619 -31
rect 679 -37 737 -31
rect 797 -37 855 -31
rect 915 -37 973 -31
rect 1033 -37 1091 -31
rect 1151 -37 1209 -31
rect 1269 -37 1327 -31
rect 1387 -37 1445 -31
rect -1445 -71 -1433 -37
rect -1327 -71 -1315 -37
rect -1209 -71 -1197 -37
rect -1091 -71 -1079 -37
rect -973 -71 -961 -37
rect -855 -71 -843 -37
rect -737 -71 -725 -37
rect -619 -71 -607 -37
rect -501 -71 -489 -37
rect -383 -71 -371 -37
rect -265 -71 -253 -37
rect -147 -71 -135 -37
rect -29 -71 -17 -37
rect 89 -71 101 -37
rect 207 -71 219 -37
rect 325 -71 337 -37
rect 443 -71 455 -37
rect 561 -71 573 -37
rect 679 -71 691 -37
rect 797 -71 809 -37
rect 915 -71 927 -37
rect 1033 -71 1045 -37
rect 1151 -71 1163 -37
rect 1269 -71 1281 -37
rect 1387 -71 1399 -37
rect -1445 -77 -1387 -71
rect -1327 -77 -1269 -71
rect -1209 -77 -1151 -71
rect -1091 -77 -1033 -71
rect -973 -77 -915 -71
rect -855 -77 -797 -71
rect -737 -77 -679 -71
rect -619 -77 -561 -71
rect -501 -77 -443 -71
rect -383 -77 -325 -71
rect -265 -77 -207 -71
rect -147 -77 -89 -71
rect -29 -77 29 -71
rect 89 -77 147 -71
rect 207 -77 265 -71
rect 325 -77 383 -71
rect 443 -77 501 -71
rect 561 -77 619 -71
rect 679 -77 737 -71
rect 797 -77 855 -71
rect 915 -77 973 -71
rect 1033 -77 1091 -71
rect 1151 -77 1209 -71
rect 1269 -77 1327 -71
rect 1387 -77 1445 -71
<< nwell >>
rect -1642 -937 1642 937
<< pmos >>
rect -1446 118 -1386 718
rect -1328 118 -1268 718
rect -1210 118 -1150 718
rect -1092 118 -1032 718
rect -974 118 -914 718
rect -856 118 -796 718
rect -738 118 -678 718
rect -620 118 -560 718
rect -502 118 -442 718
rect -384 118 -324 718
rect -266 118 -206 718
rect -148 118 -88 718
rect -30 118 30 718
rect 88 118 148 718
rect 206 118 266 718
rect 324 118 384 718
rect 442 118 502 718
rect 560 118 620 718
rect 678 118 738 718
rect 796 118 856 718
rect 914 118 974 718
rect 1032 118 1092 718
rect 1150 118 1210 718
rect 1268 118 1328 718
rect 1386 118 1446 718
rect -1446 -718 -1386 -118
rect -1328 -718 -1268 -118
rect -1210 -718 -1150 -118
rect -1092 -718 -1032 -118
rect -974 -718 -914 -118
rect -856 -718 -796 -118
rect -738 -718 -678 -118
rect -620 -718 -560 -118
rect -502 -718 -442 -118
rect -384 -718 -324 -118
rect -266 -718 -206 -118
rect -148 -718 -88 -118
rect -30 -718 30 -118
rect 88 -718 148 -118
rect 206 -718 266 -118
rect 324 -718 384 -118
rect 442 -718 502 -118
rect 560 -718 620 -118
rect 678 -718 738 -118
rect 796 -718 856 -118
rect 914 -718 974 -118
rect 1032 -718 1092 -118
rect 1150 -718 1210 -118
rect 1268 -718 1328 -118
rect 1386 -718 1446 -118
<< pdiff >>
rect -1504 673 -1446 718
rect -1504 639 -1492 673
rect -1458 639 -1446 673
rect -1504 605 -1446 639
rect -1504 571 -1492 605
rect -1458 571 -1446 605
rect -1504 537 -1446 571
rect -1504 503 -1492 537
rect -1458 503 -1446 537
rect -1504 469 -1446 503
rect -1504 435 -1492 469
rect -1458 435 -1446 469
rect -1504 401 -1446 435
rect -1504 367 -1492 401
rect -1458 367 -1446 401
rect -1504 333 -1446 367
rect -1504 299 -1492 333
rect -1458 299 -1446 333
rect -1504 265 -1446 299
rect -1504 231 -1492 265
rect -1458 231 -1446 265
rect -1504 197 -1446 231
rect -1504 163 -1492 197
rect -1458 163 -1446 197
rect -1504 118 -1446 163
rect -1386 673 -1328 718
rect -1386 639 -1374 673
rect -1340 639 -1328 673
rect -1386 605 -1328 639
rect -1386 571 -1374 605
rect -1340 571 -1328 605
rect -1386 537 -1328 571
rect -1386 503 -1374 537
rect -1340 503 -1328 537
rect -1386 469 -1328 503
rect -1386 435 -1374 469
rect -1340 435 -1328 469
rect -1386 401 -1328 435
rect -1386 367 -1374 401
rect -1340 367 -1328 401
rect -1386 333 -1328 367
rect -1386 299 -1374 333
rect -1340 299 -1328 333
rect -1386 265 -1328 299
rect -1386 231 -1374 265
rect -1340 231 -1328 265
rect -1386 197 -1328 231
rect -1386 163 -1374 197
rect -1340 163 -1328 197
rect -1386 118 -1328 163
rect -1268 673 -1210 718
rect -1268 639 -1256 673
rect -1222 639 -1210 673
rect -1268 605 -1210 639
rect -1268 571 -1256 605
rect -1222 571 -1210 605
rect -1268 537 -1210 571
rect -1268 503 -1256 537
rect -1222 503 -1210 537
rect -1268 469 -1210 503
rect -1268 435 -1256 469
rect -1222 435 -1210 469
rect -1268 401 -1210 435
rect -1268 367 -1256 401
rect -1222 367 -1210 401
rect -1268 333 -1210 367
rect -1268 299 -1256 333
rect -1222 299 -1210 333
rect -1268 265 -1210 299
rect -1268 231 -1256 265
rect -1222 231 -1210 265
rect -1268 197 -1210 231
rect -1268 163 -1256 197
rect -1222 163 -1210 197
rect -1268 118 -1210 163
rect -1150 673 -1092 718
rect -1150 639 -1138 673
rect -1104 639 -1092 673
rect -1150 605 -1092 639
rect -1150 571 -1138 605
rect -1104 571 -1092 605
rect -1150 537 -1092 571
rect -1150 503 -1138 537
rect -1104 503 -1092 537
rect -1150 469 -1092 503
rect -1150 435 -1138 469
rect -1104 435 -1092 469
rect -1150 401 -1092 435
rect -1150 367 -1138 401
rect -1104 367 -1092 401
rect -1150 333 -1092 367
rect -1150 299 -1138 333
rect -1104 299 -1092 333
rect -1150 265 -1092 299
rect -1150 231 -1138 265
rect -1104 231 -1092 265
rect -1150 197 -1092 231
rect -1150 163 -1138 197
rect -1104 163 -1092 197
rect -1150 118 -1092 163
rect -1032 673 -974 718
rect -1032 639 -1020 673
rect -986 639 -974 673
rect -1032 605 -974 639
rect -1032 571 -1020 605
rect -986 571 -974 605
rect -1032 537 -974 571
rect -1032 503 -1020 537
rect -986 503 -974 537
rect -1032 469 -974 503
rect -1032 435 -1020 469
rect -986 435 -974 469
rect -1032 401 -974 435
rect -1032 367 -1020 401
rect -986 367 -974 401
rect -1032 333 -974 367
rect -1032 299 -1020 333
rect -986 299 -974 333
rect -1032 265 -974 299
rect -1032 231 -1020 265
rect -986 231 -974 265
rect -1032 197 -974 231
rect -1032 163 -1020 197
rect -986 163 -974 197
rect -1032 118 -974 163
rect -914 673 -856 718
rect -914 639 -902 673
rect -868 639 -856 673
rect -914 605 -856 639
rect -914 571 -902 605
rect -868 571 -856 605
rect -914 537 -856 571
rect -914 503 -902 537
rect -868 503 -856 537
rect -914 469 -856 503
rect -914 435 -902 469
rect -868 435 -856 469
rect -914 401 -856 435
rect -914 367 -902 401
rect -868 367 -856 401
rect -914 333 -856 367
rect -914 299 -902 333
rect -868 299 -856 333
rect -914 265 -856 299
rect -914 231 -902 265
rect -868 231 -856 265
rect -914 197 -856 231
rect -914 163 -902 197
rect -868 163 -856 197
rect -914 118 -856 163
rect -796 673 -738 718
rect -796 639 -784 673
rect -750 639 -738 673
rect -796 605 -738 639
rect -796 571 -784 605
rect -750 571 -738 605
rect -796 537 -738 571
rect -796 503 -784 537
rect -750 503 -738 537
rect -796 469 -738 503
rect -796 435 -784 469
rect -750 435 -738 469
rect -796 401 -738 435
rect -796 367 -784 401
rect -750 367 -738 401
rect -796 333 -738 367
rect -796 299 -784 333
rect -750 299 -738 333
rect -796 265 -738 299
rect -796 231 -784 265
rect -750 231 -738 265
rect -796 197 -738 231
rect -796 163 -784 197
rect -750 163 -738 197
rect -796 118 -738 163
rect -678 673 -620 718
rect -678 639 -666 673
rect -632 639 -620 673
rect -678 605 -620 639
rect -678 571 -666 605
rect -632 571 -620 605
rect -678 537 -620 571
rect -678 503 -666 537
rect -632 503 -620 537
rect -678 469 -620 503
rect -678 435 -666 469
rect -632 435 -620 469
rect -678 401 -620 435
rect -678 367 -666 401
rect -632 367 -620 401
rect -678 333 -620 367
rect -678 299 -666 333
rect -632 299 -620 333
rect -678 265 -620 299
rect -678 231 -666 265
rect -632 231 -620 265
rect -678 197 -620 231
rect -678 163 -666 197
rect -632 163 -620 197
rect -678 118 -620 163
rect -560 673 -502 718
rect -560 639 -548 673
rect -514 639 -502 673
rect -560 605 -502 639
rect -560 571 -548 605
rect -514 571 -502 605
rect -560 537 -502 571
rect -560 503 -548 537
rect -514 503 -502 537
rect -560 469 -502 503
rect -560 435 -548 469
rect -514 435 -502 469
rect -560 401 -502 435
rect -560 367 -548 401
rect -514 367 -502 401
rect -560 333 -502 367
rect -560 299 -548 333
rect -514 299 -502 333
rect -560 265 -502 299
rect -560 231 -548 265
rect -514 231 -502 265
rect -560 197 -502 231
rect -560 163 -548 197
rect -514 163 -502 197
rect -560 118 -502 163
rect -442 673 -384 718
rect -442 639 -430 673
rect -396 639 -384 673
rect -442 605 -384 639
rect -442 571 -430 605
rect -396 571 -384 605
rect -442 537 -384 571
rect -442 503 -430 537
rect -396 503 -384 537
rect -442 469 -384 503
rect -442 435 -430 469
rect -396 435 -384 469
rect -442 401 -384 435
rect -442 367 -430 401
rect -396 367 -384 401
rect -442 333 -384 367
rect -442 299 -430 333
rect -396 299 -384 333
rect -442 265 -384 299
rect -442 231 -430 265
rect -396 231 -384 265
rect -442 197 -384 231
rect -442 163 -430 197
rect -396 163 -384 197
rect -442 118 -384 163
rect -324 673 -266 718
rect -324 639 -312 673
rect -278 639 -266 673
rect -324 605 -266 639
rect -324 571 -312 605
rect -278 571 -266 605
rect -324 537 -266 571
rect -324 503 -312 537
rect -278 503 -266 537
rect -324 469 -266 503
rect -324 435 -312 469
rect -278 435 -266 469
rect -324 401 -266 435
rect -324 367 -312 401
rect -278 367 -266 401
rect -324 333 -266 367
rect -324 299 -312 333
rect -278 299 -266 333
rect -324 265 -266 299
rect -324 231 -312 265
rect -278 231 -266 265
rect -324 197 -266 231
rect -324 163 -312 197
rect -278 163 -266 197
rect -324 118 -266 163
rect -206 673 -148 718
rect -206 639 -194 673
rect -160 639 -148 673
rect -206 605 -148 639
rect -206 571 -194 605
rect -160 571 -148 605
rect -206 537 -148 571
rect -206 503 -194 537
rect -160 503 -148 537
rect -206 469 -148 503
rect -206 435 -194 469
rect -160 435 -148 469
rect -206 401 -148 435
rect -206 367 -194 401
rect -160 367 -148 401
rect -206 333 -148 367
rect -206 299 -194 333
rect -160 299 -148 333
rect -206 265 -148 299
rect -206 231 -194 265
rect -160 231 -148 265
rect -206 197 -148 231
rect -206 163 -194 197
rect -160 163 -148 197
rect -206 118 -148 163
rect -88 673 -30 718
rect -88 639 -76 673
rect -42 639 -30 673
rect -88 605 -30 639
rect -88 571 -76 605
rect -42 571 -30 605
rect -88 537 -30 571
rect -88 503 -76 537
rect -42 503 -30 537
rect -88 469 -30 503
rect -88 435 -76 469
rect -42 435 -30 469
rect -88 401 -30 435
rect -88 367 -76 401
rect -42 367 -30 401
rect -88 333 -30 367
rect -88 299 -76 333
rect -42 299 -30 333
rect -88 265 -30 299
rect -88 231 -76 265
rect -42 231 -30 265
rect -88 197 -30 231
rect -88 163 -76 197
rect -42 163 -30 197
rect -88 118 -30 163
rect 30 673 88 718
rect 30 639 42 673
rect 76 639 88 673
rect 30 605 88 639
rect 30 571 42 605
rect 76 571 88 605
rect 30 537 88 571
rect 30 503 42 537
rect 76 503 88 537
rect 30 469 88 503
rect 30 435 42 469
rect 76 435 88 469
rect 30 401 88 435
rect 30 367 42 401
rect 76 367 88 401
rect 30 333 88 367
rect 30 299 42 333
rect 76 299 88 333
rect 30 265 88 299
rect 30 231 42 265
rect 76 231 88 265
rect 30 197 88 231
rect 30 163 42 197
rect 76 163 88 197
rect 30 118 88 163
rect 148 673 206 718
rect 148 639 160 673
rect 194 639 206 673
rect 148 605 206 639
rect 148 571 160 605
rect 194 571 206 605
rect 148 537 206 571
rect 148 503 160 537
rect 194 503 206 537
rect 148 469 206 503
rect 148 435 160 469
rect 194 435 206 469
rect 148 401 206 435
rect 148 367 160 401
rect 194 367 206 401
rect 148 333 206 367
rect 148 299 160 333
rect 194 299 206 333
rect 148 265 206 299
rect 148 231 160 265
rect 194 231 206 265
rect 148 197 206 231
rect 148 163 160 197
rect 194 163 206 197
rect 148 118 206 163
rect 266 673 324 718
rect 266 639 278 673
rect 312 639 324 673
rect 266 605 324 639
rect 266 571 278 605
rect 312 571 324 605
rect 266 537 324 571
rect 266 503 278 537
rect 312 503 324 537
rect 266 469 324 503
rect 266 435 278 469
rect 312 435 324 469
rect 266 401 324 435
rect 266 367 278 401
rect 312 367 324 401
rect 266 333 324 367
rect 266 299 278 333
rect 312 299 324 333
rect 266 265 324 299
rect 266 231 278 265
rect 312 231 324 265
rect 266 197 324 231
rect 266 163 278 197
rect 312 163 324 197
rect 266 118 324 163
rect 384 673 442 718
rect 384 639 396 673
rect 430 639 442 673
rect 384 605 442 639
rect 384 571 396 605
rect 430 571 442 605
rect 384 537 442 571
rect 384 503 396 537
rect 430 503 442 537
rect 384 469 442 503
rect 384 435 396 469
rect 430 435 442 469
rect 384 401 442 435
rect 384 367 396 401
rect 430 367 442 401
rect 384 333 442 367
rect 384 299 396 333
rect 430 299 442 333
rect 384 265 442 299
rect 384 231 396 265
rect 430 231 442 265
rect 384 197 442 231
rect 384 163 396 197
rect 430 163 442 197
rect 384 118 442 163
rect 502 673 560 718
rect 502 639 514 673
rect 548 639 560 673
rect 502 605 560 639
rect 502 571 514 605
rect 548 571 560 605
rect 502 537 560 571
rect 502 503 514 537
rect 548 503 560 537
rect 502 469 560 503
rect 502 435 514 469
rect 548 435 560 469
rect 502 401 560 435
rect 502 367 514 401
rect 548 367 560 401
rect 502 333 560 367
rect 502 299 514 333
rect 548 299 560 333
rect 502 265 560 299
rect 502 231 514 265
rect 548 231 560 265
rect 502 197 560 231
rect 502 163 514 197
rect 548 163 560 197
rect 502 118 560 163
rect 620 673 678 718
rect 620 639 632 673
rect 666 639 678 673
rect 620 605 678 639
rect 620 571 632 605
rect 666 571 678 605
rect 620 537 678 571
rect 620 503 632 537
rect 666 503 678 537
rect 620 469 678 503
rect 620 435 632 469
rect 666 435 678 469
rect 620 401 678 435
rect 620 367 632 401
rect 666 367 678 401
rect 620 333 678 367
rect 620 299 632 333
rect 666 299 678 333
rect 620 265 678 299
rect 620 231 632 265
rect 666 231 678 265
rect 620 197 678 231
rect 620 163 632 197
rect 666 163 678 197
rect 620 118 678 163
rect 738 673 796 718
rect 738 639 750 673
rect 784 639 796 673
rect 738 605 796 639
rect 738 571 750 605
rect 784 571 796 605
rect 738 537 796 571
rect 738 503 750 537
rect 784 503 796 537
rect 738 469 796 503
rect 738 435 750 469
rect 784 435 796 469
rect 738 401 796 435
rect 738 367 750 401
rect 784 367 796 401
rect 738 333 796 367
rect 738 299 750 333
rect 784 299 796 333
rect 738 265 796 299
rect 738 231 750 265
rect 784 231 796 265
rect 738 197 796 231
rect 738 163 750 197
rect 784 163 796 197
rect 738 118 796 163
rect 856 673 914 718
rect 856 639 868 673
rect 902 639 914 673
rect 856 605 914 639
rect 856 571 868 605
rect 902 571 914 605
rect 856 537 914 571
rect 856 503 868 537
rect 902 503 914 537
rect 856 469 914 503
rect 856 435 868 469
rect 902 435 914 469
rect 856 401 914 435
rect 856 367 868 401
rect 902 367 914 401
rect 856 333 914 367
rect 856 299 868 333
rect 902 299 914 333
rect 856 265 914 299
rect 856 231 868 265
rect 902 231 914 265
rect 856 197 914 231
rect 856 163 868 197
rect 902 163 914 197
rect 856 118 914 163
rect 974 673 1032 718
rect 974 639 986 673
rect 1020 639 1032 673
rect 974 605 1032 639
rect 974 571 986 605
rect 1020 571 1032 605
rect 974 537 1032 571
rect 974 503 986 537
rect 1020 503 1032 537
rect 974 469 1032 503
rect 974 435 986 469
rect 1020 435 1032 469
rect 974 401 1032 435
rect 974 367 986 401
rect 1020 367 1032 401
rect 974 333 1032 367
rect 974 299 986 333
rect 1020 299 1032 333
rect 974 265 1032 299
rect 974 231 986 265
rect 1020 231 1032 265
rect 974 197 1032 231
rect 974 163 986 197
rect 1020 163 1032 197
rect 974 118 1032 163
rect 1092 673 1150 718
rect 1092 639 1104 673
rect 1138 639 1150 673
rect 1092 605 1150 639
rect 1092 571 1104 605
rect 1138 571 1150 605
rect 1092 537 1150 571
rect 1092 503 1104 537
rect 1138 503 1150 537
rect 1092 469 1150 503
rect 1092 435 1104 469
rect 1138 435 1150 469
rect 1092 401 1150 435
rect 1092 367 1104 401
rect 1138 367 1150 401
rect 1092 333 1150 367
rect 1092 299 1104 333
rect 1138 299 1150 333
rect 1092 265 1150 299
rect 1092 231 1104 265
rect 1138 231 1150 265
rect 1092 197 1150 231
rect 1092 163 1104 197
rect 1138 163 1150 197
rect 1092 118 1150 163
rect 1210 673 1268 718
rect 1210 639 1222 673
rect 1256 639 1268 673
rect 1210 605 1268 639
rect 1210 571 1222 605
rect 1256 571 1268 605
rect 1210 537 1268 571
rect 1210 503 1222 537
rect 1256 503 1268 537
rect 1210 469 1268 503
rect 1210 435 1222 469
rect 1256 435 1268 469
rect 1210 401 1268 435
rect 1210 367 1222 401
rect 1256 367 1268 401
rect 1210 333 1268 367
rect 1210 299 1222 333
rect 1256 299 1268 333
rect 1210 265 1268 299
rect 1210 231 1222 265
rect 1256 231 1268 265
rect 1210 197 1268 231
rect 1210 163 1222 197
rect 1256 163 1268 197
rect 1210 118 1268 163
rect 1328 673 1386 718
rect 1328 639 1340 673
rect 1374 639 1386 673
rect 1328 605 1386 639
rect 1328 571 1340 605
rect 1374 571 1386 605
rect 1328 537 1386 571
rect 1328 503 1340 537
rect 1374 503 1386 537
rect 1328 469 1386 503
rect 1328 435 1340 469
rect 1374 435 1386 469
rect 1328 401 1386 435
rect 1328 367 1340 401
rect 1374 367 1386 401
rect 1328 333 1386 367
rect 1328 299 1340 333
rect 1374 299 1386 333
rect 1328 265 1386 299
rect 1328 231 1340 265
rect 1374 231 1386 265
rect 1328 197 1386 231
rect 1328 163 1340 197
rect 1374 163 1386 197
rect 1328 118 1386 163
rect 1446 673 1504 718
rect 1446 639 1458 673
rect 1492 639 1504 673
rect 1446 605 1504 639
rect 1446 571 1458 605
rect 1492 571 1504 605
rect 1446 537 1504 571
rect 1446 503 1458 537
rect 1492 503 1504 537
rect 1446 469 1504 503
rect 1446 435 1458 469
rect 1492 435 1504 469
rect 1446 401 1504 435
rect 1446 367 1458 401
rect 1492 367 1504 401
rect 1446 333 1504 367
rect 1446 299 1458 333
rect 1492 299 1504 333
rect 1446 265 1504 299
rect 1446 231 1458 265
rect 1492 231 1504 265
rect 1446 197 1504 231
rect 1446 163 1458 197
rect 1492 163 1504 197
rect 1446 118 1504 163
rect -1504 -163 -1446 -118
rect -1504 -197 -1492 -163
rect -1458 -197 -1446 -163
rect -1504 -231 -1446 -197
rect -1504 -265 -1492 -231
rect -1458 -265 -1446 -231
rect -1504 -299 -1446 -265
rect -1504 -333 -1492 -299
rect -1458 -333 -1446 -299
rect -1504 -367 -1446 -333
rect -1504 -401 -1492 -367
rect -1458 -401 -1446 -367
rect -1504 -435 -1446 -401
rect -1504 -469 -1492 -435
rect -1458 -469 -1446 -435
rect -1504 -503 -1446 -469
rect -1504 -537 -1492 -503
rect -1458 -537 -1446 -503
rect -1504 -571 -1446 -537
rect -1504 -605 -1492 -571
rect -1458 -605 -1446 -571
rect -1504 -639 -1446 -605
rect -1504 -673 -1492 -639
rect -1458 -673 -1446 -639
rect -1504 -718 -1446 -673
rect -1386 -163 -1328 -118
rect -1386 -197 -1374 -163
rect -1340 -197 -1328 -163
rect -1386 -231 -1328 -197
rect -1386 -265 -1374 -231
rect -1340 -265 -1328 -231
rect -1386 -299 -1328 -265
rect -1386 -333 -1374 -299
rect -1340 -333 -1328 -299
rect -1386 -367 -1328 -333
rect -1386 -401 -1374 -367
rect -1340 -401 -1328 -367
rect -1386 -435 -1328 -401
rect -1386 -469 -1374 -435
rect -1340 -469 -1328 -435
rect -1386 -503 -1328 -469
rect -1386 -537 -1374 -503
rect -1340 -537 -1328 -503
rect -1386 -571 -1328 -537
rect -1386 -605 -1374 -571
rect -1340 -605 -1328 -571
rect -1386 -639 -1328 -605
rect -1386 -673 -1374 -639
rect -1340 -673 -1328 -639
rect -1386 -718 -1328 -673
rect -1268 -163 -1210 -118
rect -1268 -197 -1256 -163
rect -1222 -197 -1210 -163
rect -1268 -231 -1210 -197
rect -1268 -265 -1256 -231
rect -1222 -265 -1210 -231
rect -1268 -299 -1210 -265
rect -1268 -333 -1256 -299
rect -1222 -333 -1210 -299
rect -1268 -367 -1210 -333
rect -1268 -401 -1256 -367
rect -1222 -401 -1210 -367
rect -1268 -435 -1210 -401
rect -1268 -469 -1256 -435
rect -1222 -469 -1210 -435
rect -1268 -503 -1210 -469
rect -1268 -537 -1256 -503
rect -1222 -537 -1210 -503
rect -1268 -571 -1210 -537
rect -1268 -605 -1256 -571
rect -1222 -605 -1210 -571
rect -1268 -639 -1210 -605
rect -1268 -673 -1256 -639
rect -1222 -673 -1210 -639
rect -1268 -718 -1210 -673
rect -1150 -163 -1092 -118
rect -1150 -197 -1138 -163
rect -1104 -197 -1092 -163
rect -1150 -231 -1092 -197
rect -1150 -265 -1138 -231
rect -1104 -265 -1092 -231
rect -1150 -299 -1092 -265
rect -1150 -333 -1138 -299
rect -1104 -333 -1092 -299
rect -1150 -367 -1092 -333
rect -1150 -401 -1138 -367
rect -1104 -401 -1092 -367
rect -1150 -435 -1092 -401
rect -1150 -469 -1138 -435
rect -1104 -469 -1092 -435
rect -1150 -503 -1092 -469
rect -1150 -537 -1138 -503
rect -1104 -537 -1092 -503
rect -1150 -571 -1092 -537
rect -1150 -605 -1138 -571
rect -1104 -605 -1092 -571
rect -1150 -639 -1092 -605
rect -1150 -673 -1138 -639
rect -1104 -673 -1092 -639
rect -1150 -718 -1092 -673
rect -1032 -163 -974 -118
rect -1032 -197 -1020 -163
rect -986 -197 -974 -163
rect -1032 -231 -974 -197
rect -1032 -265 -1020 -231
rect -986 -265 -974 -231
rect -1032 -299 -974 -265
rect -1032 -333 -1020 -299
rect -986 -333 -974 -299
rect -1032 -367 -974 -333
rect -1032 -401 -1020 -367
rect -986 -401 -974 -367
rect -1032 -435 -974 -401
rect -1032 -469 -1020 -435
rect -986 -469 -974 -435
rect -1032 -503 -974 -469
rect -1032 -537 -1020 -503
rect -986 -537 -974 -503
rect -1032 -571 -974 -537
rect -1032 -605 -1020 -571
rect -986 -605 -974 -571
rect -1032 -639 -974 -605
rect -1032 -673 -1020 -639
rect -986 -673 -974 -639
rect -1032 -718 -974 -673
rect -914 -163 -856 -118
rect -914 -197 -902 -163
rect -868 -197 -856 -163
rect -914 -231 -856 -197
rect -914 -265 -902 -231
rect -868 -265 -856 -231
rect -914 -299 -856 -265
rect -914 -333 -902 -299
rect -868 -333 -856 -299
rect -914 -367 -856 -333
rect -914 -401 -902 -367
rect -868 -401 -856 -367
rect -914 -435 -856 -401
rect -914 -469 -902 -435
rect -868 -469 -856 -435
rect -914 -503 -856 -469
rect -914 -537 -902 -503
rect -868 -537 -856 -503
rect -914 -571 -856 -537
rect -914 -605 -902 -571
rect -868 -605 -856 -571
rect -914 -639 -856 -605
rect -914 -673 -902 -639
rect -868 -673 -856 -639
rect -914 -718 -856 -673
rect -796 -163 -738 -118
rect -796 -197 -784 -163
rect -750 -197 -738 -163
rect -796 -231 -738 -197
rect -796 -265 -784 -231
rect -750 -265 -738 -231
rect -796 -299 -738 -265
rect -796 -333 -784 -299
rect -750 -333 -738 -299
rect -796 -367 -738 -333
rect -796 -401 -784 -367
rect -750 -401 -738 -367
rect -796 -435 -738 -401
rect -796 -469 -784 -435
rect -750 -469 -738 -435
rect -796 -503 -738 -469
rect -796 -537 -784 -503
rect -750 -537 -738 -503
rect -796 -571 -738 -537
rect -796 -605 -784 -571
rect -750 -605 -738 -571
rect -796 -639 -738 -605
rect -796 -673 -784 -639
rect -750 -673 -738 -639
rect -796 -718 -738 -673
rect -678 -163 -620 -118
rect -678 -197 -666 -163
rect -632 -197 -620 -163
rect -678 -231 -620 -197
rect -678 -265 -666 -231
rect -632 -265 -620 -231
rect -678 -299 -620 -265
rect -678 -333 -666 -299
rect -632 -333 -620 -299
rect -678 -367 -620 -333
rect -678 -401 -666 -367
rect -632 -401 -620 -367
rect -678 -435 -620 -401
rect -678 -469 -666 -435
rect -632 -469 -620 -435
rect -678 -503 -620 -469
rect -678 -537 -666 -503
rect -632 -537 -620 -503
rect -678 -571 -620 -537
rect -678 -605 -666 -571
rect -632 -605 -620 -571
rect -678 -639 -620 -605
rect -678 -673 -666 -639
rect -632 -673 -620 -639
rect -678 -718 -620 -673
rect -560 -163 -502 -118
rect -560 -197 -548 -163
rect -514 -197 -502 -163
rect -560 -231 -502 -197
rect -560 -265 -548 -231
rect -514 -265 -502 -231
rect -560 -299 -502 -265
rect -560 -333 -548 -299
rect -514 -333 -502 -299
rect -560 -367 -502 -333
rect -560 -401 -548 -367
rect -514 -401 -502 -367
rect -560 -435 -502 -401
rect -560 -469 -548 -435
rect -514 -469 -502 -435
rect -560 -503 -502 -469
rect -560 -537 -548 -503
rect -514 -537 -502 -503
rect -560 -571 -502 -537
rect -560 -605 -548 -571
rect -514 -605 -502 -571
rect -560 -639 -502 -605
rect -560 -673 -548 -639
rect -514 -673 -502 -639
rect -560 -718 -502 -673
rect -442 -163 -384 -118
rect -442 -197 -430 -163
rect -396 -197 -384 -163
rect -442 -231 -384 -197
rect -442 -265 -430 -231
rect -396 -265 -384 -231
rect -442 -299 -384 -265
rect -442 -333 -430 -299
rect -396 -333 -384 -299
rect -442 -367 -384 -333
rect -442 -401 -430 -367
rect -396 -401 -384 -367
rect -442 -435 -384 -401
rect -442 -469 -430 -435
rect -396 -469 -384 -435
rect -442 -503 -384 -469
rect -442 -537 -430 -503
rect -396 -537 -384 -503
rect -442 -571 -384 -537
rect -442 -605 -430 -571
rect -396 -605 -384 -571
rect -442 -639 -384 -605
rect -442 -673 -430 -639
rect -396 -673 -384 -639
rect -442 -718 -384 -673
rect -324 -163 -266 -118
rect -324 -197 -312 -163
rect -278 -197 -266 -163
rect -324 -231 -266 -197
rect -324 -265 -312 -231
rect -278 -265 -266 -231
rect -324 -299 -266 -265
rect -324 -333 -312 -299
rect -278 -333 -266 -299
rect -324 -367 -266 -333
rect -324 -401 -312 -367
rect -278 -401 -266 -367
rect -324 -435 -266 -401
rect -324 -469 -312 -435
rect -278 -469 -266 -435
rect -324 -503 -266 -469
rect -324 -537 -312 -503
rect -278 -537 -266 -503
rect -324 -571 -266 -537
rect -324 -605 -312 -571
rect -278 -605 -266 -571
rect -324 -639 -266 -605
rect -324 -673 -312 -639
rect -278 -673 -266 -639
rect -324 -718 -266 -673
rect -206 -163 -148 -118
rect -206 -197 -194 -163
rect -160 -197 -148 -163
rect -206 -231 -148 -197
rect -206 -265 -194 -231
rect -160 -265 -148 -231
rect -206 -299 -148 -265
rect -206 -333 -194 -299
rect -160 -333 -148 -299
rect -206 -367 -148 -333
rect -206 -401 -194 -367
rect -160 -401 -148 -367
rect -206 -435 -148 -401
rect -206 -469 -194 -435
rect -160 -469 -148 -435
rect -206 -503 -148 -469
rect -206 -537 -194 -503
rect -160 -537 -148 -503
rect -206 -571 -148 -537
rect -206 -605 -194 -571
rect -160 -605 -148 -571
rect -206 -639 -148 -605
rect -206 -673 -194 -639
rect -160 -673 -148 -639
rect -206 -718 -148 -673
rect -88 -163 -30 -118
rect -88 -197 -76 -163
rect -42 -197 -30 -163
rect -88 -231 -30 -197
rect -88 -265 -76 -231
rect -42 -265 -30 -231
rect -88 -299 -30 -265
rect -88 -333 -76 -299
rect -42 -333 -30 -299
rect -88 -367 -30 -333
rect -88 -401 -76 -367
rect -42 -401 -30 -367
rect -88 -435 -30 -401
rect -88 -469 -76 -435
rect -42 -469 -30 -435
rect -88 -503 -30 -469
rect -88 -537 -76 -503
rect -42 -537 -30 -503
rect -88 -571 -30 -537
rect -88 -605 -76 -571
rect -42 -605 -30 -571
rect -88 -639 -30 -605
rect -88 -673 -76 -639
rect -42 -673 -30 -639
rect -88 -718 -30 -673
rect 30 -163 88 -118
rect 30 -197 42 -163
rect 76 -197 88 -163
rect 30 -231 88 -197
rect 30 -265 42 -231
rect 76 -265 88 -231
rect 30 -299 88 -265
rect 30 -333 42 -299
rect 76 -333 88 -299
rect 30 -367 88 -333
rect 30 -401 42 -367
rect 76 -401 88 -367
rect 30 -435 88 -401
rect 30 -469 42 -435
rect 76 -469 88 -435
rect 30 -503 88 -469
rect 30 -537 42 -503
rect 76 -537 88 -503
rect 30 -571 88 -537
rect 30 -605 42 -571
rect 76 -605 88 -571
rect 30 -639 88 -605
rect 30 -673 42 -639
rect 76 -673 88 -639
rect 30 -718 88 -673
rect 148 -163 206 -118
rect 148 -197 160 -163
rect 194 -197 206 -163
rect 148 -231 206 -197
rect 148 -265 160 -231
rect 194 -265 206 -231
rect 148 -299 206 -265
rect 148 -333 160 -299
rect 194 -333 206 -299
rect 148 -367 206 -333
rect 148 -401 160 -367
rect 194 -401 206 -367
rect 148 -435 206 -401
rect 148 -469 160 -435
rect 194 -469 206 -435
rect 148 -503 206 -469
rect 148 -537 160 -503
rect 194 -537 206 -503
rect 148 -571 206 -537
rect 148 -605 160 -571
rect 194 -605 206 -571
rect 148 -639 206 -605
rect 148 -673 160 -639
rect 194 -673 206 -639
rect 148 -718 206 -673
rect 266 -163 324 -118
rect 266 -197 278 -163
rect 312 -197 324 -163
rect 266 -231 324 -197
rect 266 -265 278 -231
rect 312 -265 324 -231
rect 266 -299 324 -265
rect 266 -333 278 -299
rect 312 -333 324 -299
rect 266 -367 324 -333
rect 266 -401 278 -367
rect 312 -401 324 -367
rect 266 -435 324 -401
rect 266 -469 278 -435
rect 312 -469 324 -435
rect 266 -503 324 -469
rect 266 -537 278 -503
rect 312 -537 324 -503
rect 266 -571 324 -537
rect 266 -605 278 -571
rect 312 -605 324 -571
rect 266 -639 324 -605
rect 266 -673 278 -639
rect 312 -673 324 -639
rect 266 -718 324 -673
rect 384 -163 442 -118
rect 384 -197 396 -163
rect 430 -197 442 -163
rect 384 -231 442 -197
rect 384 -265 396 -231
rect 430 -265 442 -231
rect 384 -299 442 -265
rect 384 -333 396 -299
rect 430 -333 442 -299
rect 384 -367 442 -333
rect 384 -401 396 -367
rect 430 -401 442 -367
rect 384 -435 442 -401
rect 384 -469 396 -435
rect 430 -469 442 -435
rect 384 -503 442 -469
rect 384 -537 396 -503
rect 430 -537 442 -503
rect 384 -571 442 -537
rect 384 -605 396 -571
rect 430 -605 442 -571
rect 384 -639 442 -605
rect 384 -673 396 -639
rect 430 -673 442 -639
rect 384 -718 442 -673
rect 502 -163 560 -118
rect 502 -197 514 -163
rect 548 -197 560 -163
rect 502 -231 560 -197
rect 502 -265 514 -231
rect 548 -265 560 -231
rect 502 -299 560 -265
rect 502 -333 514 -299
rect 548 -333 560 -299
rect 502 -367 560 -333
rect 502 -401 514 -367
rect 548 -401 560 -367
rect 502 -435 560 -401
rect 502 -469 514 -435
rect 548 -469 560 -435
rect 502 -503 560 -469
rect 502 -537 514 -503
rect 548 -537 560 -503
rect 502 -571 560 -537
rect 502 -605 514 -571
rect 548 -605 560 -571
rect 502 -639 560 -605
rect 502 -673 514 -639
rect 548 -673 560 -639
rect 502 -718 560 -673
rect 620 -163 678 -118
rect 620 -197 632 -163
rect 666 -197 678 -163
rect 620 -231 678 -197
rect 620 -265 632 -231
rect 666 -265 678 -231
rect 620 -299 678 -265
rect 620 -333 632 -299
rect 666 -333 678 -299
rect 620 -367 678 -333
rect 620 -401 632 -367
rect 666 -401 678 -367
rect 620 -435 678 -401
rect 620 -469 632 -435
rect 666 -469 678 -435
rect 620 -503 678 -469
rect 620 -537 632 -503
rect 666 -537 678 -503
rect 620 -571 678 -537
rect 620 -605 632 -571
rect 666 -605 678 -571
rect 620 -639 678 -605
rect 620 -673 632 -639
rect 666 -673 678 -639
rect 620 -718 678 -673
rect 738 -163 796 -118
rect 738 -197 750 -163
rect 784 -197 796 -163
rect 738 -231 796 -197
rect 738 -265 750 -231
rect 784 -265 796 -231
rect 738 -299 796 -265
rect 738 -333 750 -299
rect 784 -333 796 -299
rect 738 -367 796 -333
rect 738 -401 750 -367
rect 784 -401 796 -367
rect 738 -435 796 -401
rect 738 -469 750 -435
rect 784 -469 796 -435
rect 738 -503 796 -469
rect 738 -537 750 -503
rect 784 -537 796 -503
rect 738 -571 796 -537
rect 738 -605 750 -571
rect 784 -605 796 -571
rect 738 -639 796 -605
rect 738 -673 750 -639
rect 784 -673 796 -639
rect 738 -718 796 -673
rect 856 -163 914 -118
rect 856 -197 868 -163
rect 902 -197 914 -163
rect 856 -231 914 -197
rect 856 -265 868 -231
rect 902 -265 914 -231
rect 856 -299 914 -265
rect 856 -333 868 -299
rect 902 -333 914 -299
rect 856 -367 914 -333
rect 856 -401 868 -367
rect 902 -401 914 -367
rect 856 -435 914 -401
rect 856 -469 868 -435
rect 902 -469 914 -435
rect 856 -503 914 -469
rect 856 -537 868 -503
rect 902 -537 914 -503
rect 856 -571 914 -537
rect 856 -605 868 -571
rect 902 -605 914 -571
rect 856 -639 914 -605
rect 856 -673 868 -639
rect 902 -673 914 -639
rect 856 -718 914 -673
rect 974 -163 1032 -118
rect 974 -197 986 -163
rect 1020 -197 1032 -163
rect 974 -231 1032 -197
rect 974 -265 986 -231
rect 1020 -265 1032 -231
rect 974 -299 1032 -265
rect 974 -333 986 -299
rect 1020 -333 1032 -299
rect 974 -367 1032 -333
rect 974 -401 986 -367
rect 1020 -401 1032 -367
rect 974 -435 1032 -401
rect 974 -469 986 -435
rect 1020 -469 1032 -435
rect 974 -503 1032 -469
rect 974 -537 986 -503
rect 1020 -537 1032 -503
rect 974 -571 1032 -537
rect 974 -605 986 -571
rect 1020 -605 1032 -571
rect 974 -639 1032 -605
rect 974 -673 986 -639
rect 1020 -673 1032 -639
rect 974 -718 1032 -673
rect 1092 -163 1150 -118
rect 1092 -197 1104 -163
rect 1138 -197 1150 -163
rect 1092 -231 1150 -197
rect 1092 -265 1104 -231
rect 1138 -265 1150 -231
rect 1092 -299 1150 -265
rect 1092 -333 1104 -299
rect 1138 -333 1150 -299
rect 1092 -367 1150 -333
rect 1092 -401 1104 -367
rect 1138 -401 1150 -367
rect 1092 -435 1150 -401
rect 1092 -469 1104 -435
rect 1138 -469 1150 -435
rect 1092 -503 1150 -469
rect 1092 -537 1104 -503
rect 1138 -537 1150 -503
rect 1092 -571 1150 -537
rect 1092 -605 1104 -571
rect 1138 -605 1150 -571
rect 1092 -639 1150 -605
rect 1092 -673 1104 -639
rect 1138 -673 1150 -639
rect 1092 -718 1150 -673
rect 1210 -163 1268 -118
rect 1210 -197 1222 -163
rect 1256 -197 1268 -163
rect 1210 -231 1268 -197
rect 1210 -265 1222 -231
rect 1256 -265 1268 -231
rect 1210 -299 1268 -265
rect 1210 -333 1222 -299
rect 1256 -333 1268 -299
rect 1210 -367 1268 -333
rect 1210 -401 1222 -367
rect 1256 -401 1268 -367
rect 1210 -435 1268 -401
rect 1210 -469 1222 -435
rect 1256 -469 1268 -435
rect 1210 -503 1268 -469
rect 1210 -537 1222 -503
rect 1256 -537 1268 -503
rect 1210 -571 1268 -537
rect 1210 -605 1222 -571
rect 1256 -605 1268 -571
rect 1210 -639 1268 -605
rect 1210 -673 1222 -639
rect 1256 -673 1268 -639
rect 1210 -718 1268 -673
rect 1328 -163 1386 -118
rect 1328 -197 1340 -163
rect 1374 -197 1386 -163
rect 1328 -231 1386 -197
rect 1328 -265 1340 -231
rect 1374 -265 1386 -231
rect 1328 -299 1386 -265
rect 1328 -333 1340 -299
rect 1374 -333 1386 -299
rect 1328 -367 1386 -333
rect 1328 -401 1340 -367
rect 1374 -401 1386 -367
rect 1328 -435 1386 -401
rect 1328 -469 1340 -435
rect 1374 -469 1386 -435
rect 1328 -503 1386 -469
rect 1328 -537 1340 -503
rect 1374 -537 1386 -503
rect 1328 -571 1386 -537
rect 1328 -605 1340 -571
rect 1374 -605 1386 -571
rect 1328 -639 1386 -605
rect 1328 -673 1340 -639
rect 1374 -673 1386 -639
rect 1328 -718 1386 -673
rect 1446 -163 1504 -118
rect 1446 -197 1458 -163
rect 1492 -197 1504 -163
rect 1446 -231 1504 -197
rect 1446 -265 1458 -231
rect 1492 -265 1504 -231
rect 1446 -299 1504 -265
rect 1446 -333 1458 -299
rect 1492 -333 1504 -299
rect 1446 -367 1504 -333
rect 1446 -401 1458 -367
rect 1492 -401 1504 -367
rect 1446 -435 1504 -401
rect 1446 -469 1458 -435
rect 1492 -469 1504 -435
rect 1446 -503 1504 -469
rect 1446 -537 1458 -503
rect 1492 -537 1504 -503
rect 1446 -571 1504 -537
rect 1446 -605 1458 -571
rect 1492 -605 1504 -571
rect 1446 -639 1504 -605
rect 1446 -673 1458 -639
rect 1492 -673 1504 -639
rect 1446 -718 1504 -673
<< pdiffc >>
rect -1492 639 -1458 673
rect -1492 571 -1458 605
rect -1492 503 -1458 537
rect -1492 435 -1458 469
rect -1492 367 -1458 401
rect -1492 299 -1458 333
rect -1492 231 -1458 265
rect -1492 163 -1458 197
rect -1374 639 -1340 673
rect -1374 571 -1340 605
rect -1374 503 -1340 537
rect -1374 435 -1340 469
rect -1374 367 -1340 401
rect -1374 299 -1340 333
rect -1374 231 -1340 265
rect -1374 163 -1340 197
rect -1256 639 -1222 673
rect -1256 571 -1222 605
rect -1256 503 -1222 537
rect -1256 435 -1222 469
rect -1256 367 -1222 401
rect -1256 299 -1222 333
rect -1256 231 -1222 265
rect -1256 163 -1222 197
rect -1138 639 -1104 673
rect -1138 571 -1104 605
rect -1138 503 -1104 537
rect -1138 435 -1104 469
rect -1138 367 -1104 401
rect -1138 299 -1104 333
rect -1138 231 -1104 265
rect -1138 163 -1104 197
rect -1020 639 -986 673
rect -1020 571 -986 605
rect -1020 503 -986 537
rect -1020 435 -986 469
rect -1020 367 -986 401
rect -1020 299 -986 333
rect -1020 231 -986 265
rect -1020 163 -986 197
rect -902 639 -868 673
rect -902 571 -868 605
rect -902 503 -868 537
rect -902 435 -868 469
rect -902 367 -868 401
rect -902 299 -868 333
rect -902 231 -868 265
rect -902 163 -868 197
rect -784 639 -750 673
rect -784 571 -750 605
rect -784 503 -750 537
rect -784 435 -750 469
rect -784 367 -750 401
rect -784 299 -750 333
rect -784 231 -750 265
rect -784 163 -750 197
rect -666 639 -632 673
rect -666 571 -632 605
rect -666 503 -632 537
rect -666 435 -632 469
rect -666 367 -632 401
rect -666 299 -632 333
rect -666 231 -632 265
rect -666 163 -632 197
rect -548 639 -514 673
rect -548 571 -514 605
rect -548 503 -514 537
rect -548 435 -514 469
rect -548 367 -514 401
rect -548 299 -514 333
rect -548 231 -514 265
rect -548 163 -514 197
rect -430 639 -396 673
rect -430 571 -396 605
rect -430 503 -396 537
rect -430 435 -396 469
rect -430 367 -396 401
rect -430 299 -396 333
rect -430 231 -396 265
rect -430 163 -396 197
rect -312 639 -278 673
rect -312 571 -278 605
rect -312 503 -278 537
rect -312 435 -278 469
rect -312 367 -278 401
rect -312 299 -278 333
rect -312 231 -278 265
rect -312 163 -278 197
rect -194 639 -160 673
rect -194 571 -160 605
rect -194 503 -160 537
rect -194 435 -160 469
rect -194 367 -160 401
rect -194 299 -160 333
rect -194 231 -160 265
rect -194 163 -160 197
rect -76 639 -42 673
rect -76 571 -42 605
rect -76 503 -42 537
rect -76 435 -42 469
rect -76 367 -42 401
rect -76 299 -42 333
rect -76 231 -42 265
rect -76 163 -42 197
rect 42 639 76 673
rect 42 571 76 605
rect 42 503 76 537
rect 42 435 76 469
rect 42 367 76 401
rect 42 299 76 333
rect 42 231 76 265
rect 42 163 76 197
rect 160 639 194 673
rect 160 571 194 605
rect 160 503 194 537
rect 160 435 194 469
rect 160 367 194 401
rect 160 299 194 333
rect 160 231 194 265
rect 160 163 194 197
rect 278 639 312 673
rect 278 571 312 605
rect 278 503 312 537
rect 278 435 312 469
rect 278 367 312 401
rect 278 299 312 333
rect 278 231 312 265
rect 278 163 312 197
rect 396 639 430 673
rect 396 571 430 605
rect 396 503 430 537
rect 396 435 430 469
rect 396 367 430 401
rect 396 299 430 333
rect 396 231 430 265
rect 396 163 430 197
rect 514 639 548 673
rect 514 571 548 605
rect 514 503 548 537
rect 514 435 548 469
rect 514 367 548 401
rect 514 299 548 333
rect 514 231 548 265
rect 514 163 548 197
rect 632 639 666 673
rect 632 571 666 605
rect 632 503 666 537
rect 632 435 666 469
rect 632 367 666 401
rect 632 299 666 333
rect 632 231 666 265
rect 632 163 666 197
rect 750 639 784 673
rect 750 571 784 605
rect 750 503 784 537
rect 750 435 784 469
rect 750 367 784 401
rect 750 299 784 333
rect 750 231 784 265
rect 750 163 784 197
rect 868 639 902 673
rect 868 571 902 605
rect 868 503 902 537
rect 868 435 902 469
rect 868 367 902 401
rect 868 299 902 333
rect 868 231 902 265
rect 868 163 902 197
rect 986 639 1020 673
rect 986 571 1020 605
rect 986 503 1020 537
rect 986 435 1020 469
rect 986 367 1020 401
rect 986 299 1020 333
rect 986 231 1020 265
rect 986 163 1020 197
rect 1104 639 1138 673
rect 1104 571 1138 605
rect 1104 503 1138 537
rect 1104 435 1138 469
rect 1104 367 1138 401
rect 1104 299 1138 333
rect 1104 231 1138 265
rect 1104 163 1138 197
rect 1222 639 1256 673
rect 1222 571 1256 605
rect 1222 503 1256 537
rect 1222 435 1256 469
rect 1222 367 1256 401
rect 1222 299 1256 333
rect 1222 231 1256 265
rect 1222 163 1256 197
rect 1340 639 1374 673
rect 1340 571 1374 605
rect 1340 503 1374 537
rect 1340 435 1374 469
rect 1340 367 1374 401
rect 1340 299 1374 333
rect 1340 231 1374 265
rect 1340 163 1374 197
rect 1458 639 1492 673
rect 1458 571 1492 605
rect 1458 503 1492 537
rect 1458 435 1492 469
rect 1458 367 1492 401
rect 1458 299 1492 333
rect 1458 231 1492 265
rect 1458 163 1492 197
rect -1492 -197 -1458 -163
rect -1492 -265 -1458 -231
rect -1492 -333 -1458 -299
rect -1492 -401 -1458 -367
rect -1492 -469 -1458 -435
rect -1492 -537 -1458 -503
rect -1492 -605 -1458 -571
rect -1492 -673 -1458 -639
rect -1374 -197 -1340 -163
rect -1374 -265 -1340 -231
rect -1374 -333 -1340 -299
rect -1374 -401 -1340 -367
rect -1374 -469 -1340 -435
rect -1374 -537 -1340 -503
rect -1374 -605 -1340 -571
rect -1374 -673 -1340 -639
rect -1256 -197 -1222 -163
rect -1256 -265 -1222 -231
rect -1256 -333 -1222 -299
rect -1256 -401 -1222 -367
rect -1256 -469 -1222 -435
rect -1256 -537 -1222 -503
rect -1256 -605 -1222 -571
rect -1256 -673 -1222 -639
rect -1138 -197 -1104 -163
rect -1138 -265 -1104 -231
rect -1138 -333 -1104 -299
rect -1138 -401 -1104 -367
rect -1138 -469 -1104 -435
rect -1138 -537 -1104 -503
rect -1138 -605 -1104 -571
rect -1138 -673 -1104 -639
rect -1020 -197 -986 -163
rect -1020 -265 -986 -231
rect -1020 -333 -986 -299
rect -1020 -401 -986 -367
rect -1020 -469 -986 -435
rect -1020 -537 -986 -503
rect -1020 -605 -986 -571
rect -1020 -673 -986 -639
rect -902 -197 -868 -163
rect -902 -265 -868 -231
rect -902 -333 -868 -299
rect -902 -401 -868 -367
rect -902 -469 -868 -435
rect -902 -537 -868 -503
rect -902 -605 -868 -571
rect -902 -673 -868 -639
rect -784 -197 -750 -163
rect -784 -265 -750 -231
rect -784 -333 -750 -299
rect -784 -401 -750 -367
rect -784 -469 -750 -435
rect -784 -537 -750 -503
rect -784 -605 -750 -571
rect -784 -673 -750 -639
rect -666 -197 -632 -163
rect -666 -265 -632 -231
rect -666 -333 -632 -299
rect -666 -401 -632 -367
rect -666 -469 -632 -435
rect -666 -537 -632 -503
rect -666 -605 -632 -571
rect -666 -673 -632 -639
rect -548 -197 -514 -163
rect -548 -265 -514 -231
rect -548 -333 -514 -299
rect -548 -401 -514 -367
rect -548 -469 -514 -435
rect -548 -537 -514 -503
rect -548 -605 -514 -571
rect -548 -673 -514 -639
rect -430 -197 -396 -163
rect -430 -265 -396 -231
rect -430 -333 -396 -299
rect -430 -401 -396 -367
rect -430 -469 -396 -435
rect -430 -537 -396 -503
rect -430 -605 -396 -571
rect -430 -673 -396 -639
rect -312 -197 -278 -163
rect -312 -265 -278 -231
rect -312 -333 -278 -299
rect -312 -401 -278 -367
rect -312 -469 -278 -435
rect -312 -537 -278 -503
rect -312 -605 -278 -571
rect -312 -673 -278 -639
rect -194 -197 -160 -163
rect -194 -265 -160 -231
rect -194 -333 -160 -299
rect -194 -401 -160 -367
rect -194 -469 -160 -435
rect -194 -537 -160 -503
rect -194 -605 -160 -571
rect -194 -673 -160 -639
rect -76 -197 -42 -163
rect -76 -265 -42 -231
rect -76 -333 -42 -299
rect -76 -401 -42 -367
rect -76 -469 -42 -435
rect -76 -537 -42 -503
rect -76 -605 -42 -571
rect -76 -673 -42 -639
rect 42 -197 76 -163
rect 42 -265 76 -231
rect 42 -333 76 -299
rect 42 -401 76 -367
rect 42 -469 76 -435
rect 42 -537 76 -503
rect 42 -605 76 -571
rect 42 -673 76 -639
rect 160 -197 194 -163
rect 160 -265 194 -231
rect 160 -333 194 -299
rect 160 -401 194 -367
rect 160 -469 194 -435
rect 160 -537 194 -503
rect 160 -605 194 -571
rect 160 -673 194 -639
rect 278 -197 312 -163
rect 278 -265 312 -231
rect 278 -333 312 -299
rect 278 -401 312 -367
rect 278 -469 312 -435
rect 278 -537 312 -503
rect 278 -605 312 -571
rect 278 -673 312 -639
rect 396 -197 430 -163
rect 396 -265 430 -231
rect 396 -333 430 -299
rect 396 -401 430 -367
rect 396 -469 430 -435
rect 396 -537 430 -503
rect 396 -605 430 -571
rect 396 -673 430 -639
rect 514 -197 548 -163
rect 514 -265 548 -231
rect 514 -333 548 -299
rect 514 -401 548 -367
rect 514 -469 548 -435
rect 514 -537 548 -503
rect 514 -605 548 -571
rect 514 -673 548 -639
rect 632 -197 666 -163
rect 632 -265 666 -231
rect 632 -333 666 -299
rect 632 -401 666 -367
rect 632 -469 666 -435
rect 632 -537 666 -503
rect 632 -605 666 -571
rect 632 -673 666 -639
rect 750 -197 784 -163
rect 750 -265 784 -231
rect 750 -333 784 -299
rect 750 -401 784 -367
rect 750 -469 784 -435
rect 750 -537 784 -503
rect 750 -605 784 -571
rect 750 -673 784 -639
rect 868 -197 902 -163
rect 868 -265 902 -231
rect 868 -333 902 -299
rect 868 -401 902 -367
rect 868 -469 902 -435
rect 868 -537 902 -503
rect 868 -605 902 -571
rect 868 -673 902 -639
rect 986 -197 1020 -163
rect 986 -265 1020 -231
rect 986 -333 1020 -299
rect 986 -401 1020 -367
rect 986 -469 1020 -435
rect 986 -537 1020 -503
rect 986 -605 1020 -571
rect 986 -673 1020 -639
rect 1104 -197 1138 -163
rect 1104 -265 1138 -231
rect 1104 -333 1138 -299
rect 1104 -401 1138 -367
rect 1104 -469 1138 -435
rect 1104 -537 1138 -503
rect 1104 -605 1138 -571
rect 1104 -673 1138 -639
rect 1222 -197 1256 -163
rect 1222 -265 1256 -231
rect 1222 -333 1256 -299
rect 1222 -401 1256 -367
rect 1222 -469 1256 -435
rect 1222 -537 1256 -503
rect 1222 -605 1256 -571
rect 1222 -673 1256 -639
rect 1340 -197 1374 -163
rect 1340 -265 1374 -231
rect 1340 -333 1374 -299
rect 1340 -401 1374 -367
rect 1340 -469 1374 -435
rect 1340 -537 1374 -503
rect 1340 -605 1374 -571
rect 1340 -673 1374 -639
rect 1458 -197 1492 -163
rect 1458 -265 1492 -231
rect 1458 -333 1492 -299
rect 1458 -401 1492 -367
rect 1458 -469 1492 -435
rect 1458 -537 1492 -503
rect 1458 -605 1492 -571
rect 1458 -673 1492 -639
<< nsubdiff >>
rect -1606 867 -1479 901
rect -1445 867 -1411 901
rect -1377 867 -1343 901
rect -1309 867 -1275 901
rect -1241 867 -1207 901
rect -1173 867 -1139 901
rect -1105 867 -1071 901
rect -1037 867 -1003 901
rect -969 867 -935 901
rect -901 867 -867 901
rect -833 867 -799 901
rect -765 867 -731 901
rect -697 867 -663 901
rect -629 867 -595 901
rect -561 867 -527 901
rect -493 867 -459 901
rect -425 867 -391 901
rect -357 867 -323 901
rect -289 867 -255 901
rect -221 867 -187 901
rect -153 867 -119 901
rect -85 867 -51 901
rect -17 867 17 901
rect 51 867 85 901
rect 119 867 153 901
rect 187 867 221 901
rect 255 867 289 901
rect 323 867 357 901
rect 391 867 425 901
rect 459 867 493 901
rect 527 867 561 901
rect 595 867 629 901
rect 663 867 697 901
rect 731 867 765 901
rect 799 867 833 901
rect 867 867 901 901
rect 935 867 969 901
rect 1003 867 1037 901
rect 1071 867 1105 901
rect 1139 867 1173 901
rect 1207 867 1241 901
rect 1275 867 1309 901
rect 1343 867 1377 901
rect 1411 867 1445 901
rect 1479 867 1606 901
rect -1606 799 -1572 867
rect -1606 731 -1572 765
rect 1572 799 1606 867
rect 1572 731 1606 765
rect -1606 663 -1572 697
rect -1606 595 -1572 629
rect -1606 527 -1572 561
rect -1606 459 -1572 493
rect -1606 391 -1572 425
rect -1606 323 -1572 357
rect -1606 255 -1572 289
rect -1606 187 -1572 221
rect -1606 119 -1572 153
rect 1572 663 1606 697
rect 1572 595 1606 629
rect 1572 527 1606 561
rect 1572 459 1606 493
rect 1572 391 1606 425
rect 1572 323 1606 357
rect 1572 255 1606 289
rect 1572 187 1606 221
rect 1572 119 1606 153
rect -1606 51 -1572 85
rect 1572 51 1606 85
rect -1606 -17 -1572 17
rect 1572 -17 1606 17
rect -1606 -85 -1572 -51
rect 1572 -85 1606 -51
rect -1606 -153 -1572 -119
rect -1606 -221 -1572 -187
rect -1606 -289 -1572 -255
rect -1606 -357 -1572 -323
rect -1606 -425 -1572 -391
rect -1606 -493 -1572 -459
rect -1606 -561 -1572 -527
rect -1606 -629 -1572 -595
rect -1606 -697 -1572 -663
rect 1572 -153 1606 -119
rect 1572 -221 1606 -187
rect 1572 -289 1606 -255
rect 1572 -357 1606 -323
rect 1572 -425 1606 -391
rect 1572 -493 1606 -459
rect 1572 -561 1606 -527
rect 1572 -629 1606 -595
rect 1572 -697 1606 -663
rect -1606 -765 -1572 -731
rect -1606 -867 -1572 -799
rect 1572 -765 1606 -731
rect 1572 -867 1606 -799
rect -1606 -901 -1479 -867
rect -1445 -901 -1411 -867
rect -1377 -901 -1343 -867
rect -1309 -901 -1275 -867
rect -1241 -901 -1207 -867
rect -1173 -901 -1139 -867
rect -1105 -901 -1071 -867
rect -1037 -901 -1003 -867
rect -969 -901 -935 -867
rect -901 -901 -867 -867
rect -833 -901 -799 -867
rect -765 -901 -731 -867
rect -697 -901 -663 -867
rect -629 -901 -595 -867
rect -561 -901 -527 -867
rect -493 -901 -459 -867
rect -425 -901 -391 -867
rect -357 -901 -323 -867
rect -289 -901 -255 -867
rect -221 -901 -187 -867
rect -153 -901 -119 -867
rect -85 -901 -51 -867
rect -17 -901 17 -867
rect 51 -901 85 -867
rect 119 -901 153 -867
rect 187 -901 221 -867
rect 255 -901 289 -867
rect 323 -901 357 -867
rect 391 -901 425 -867
rect 459 -901 493 -867
rect 527 -901 561 -867
rect 595 -901 629 -867
rect 663 -901 697 -867
rect 731 -901 765 -867
rect 799 -901 833 -867
rect 867 -901 901 -867
rect 935 -901 969 -867
rect 1003 -901 1037 -867
rect 1071 -901 1105 -867
rect 1139 -901 1173 -867
rect 1207 -901 1241 -867
rect 1275 -901 1309 -867
rect 1343 -901 1377 -867
rect 1411 -901 1445 -867
rect 1479 -901 1606 -867
<< nsubdiffcont >>
rect -1479 867 -1445 901
rect -1411 867 -1377 901
rect -1343 867 -1309 901
rect -1275 867 -1241 901
rect -1207 867 -1173 901
rect -1139 867 -1105 901
rect -1071 867 -1037 901
rect -1003 867 -969 901
rect -935 867 -901 901
rect -867 867 -833 901
rect -799 867 -765 901
rect -731 867 -697 901
rect -663 867 -629 901
rect -595 867 -561 901
rect -527 867 -493 901
rect -459 867 -425 901
rect -391 867 -357 901
rect -323 867 -289 901
rect -255 867 -221 901
rect -187 867 -153 901
rect -119 867 -85 901
rect -51 867 -17 901
rect 17 867 51 901
rect 85 867 119 901
rect 153 867 187 901
rect 221 867 255 901
rect 289 867 323 901
rect 357 867 391 901
rect 425 867 459 901
rect 493 867 527 901
rect 561 867 595 901
rect 629 867 663 901
rect 697 867 731 901
rect 765 867 799 901
rect 833 867 867 901
rect 901 867 935 901
rect 969 867 1003 901
rect 1037 867 1071 901
rect 1105 867 1139 901
rect 1173 867 1207 901
rect 1241 867 1275 901
rect 1309 867 1343 901
rect 1377 867 1411 901
rect 1445 867 1479 901
rect -1606 765 -1572 799
rect 1572 765 1606 799
rect -1606 697 -1572 731
rect -1606 629 -1572 663
rect -1606 561 -1572 595
rect -1606 493 -1572 527
rect -1606 425 -1572 459
rect -1606 357 -1572 391
rect -1606 289 -1572 323
rect -1606 221 -1572 255
rect -1606 153 -1572 187
rect -1606 85 -1572 119
rect 1572 697 1606 731
rect 1572 629 1606 663
rect 1572 561 1606 595
rect 1572 493 1606 527
rect 1572 425 1606 459
rect 1572 357 1606 391
rect 1572 289 1606 323
rect 1572 221 1606 255
rect 1572 153 1606 187
rect -1606 17 -1572 51
rect 1572 85 1606 119
rect -1606 -51 -1572 -17
rect 1572 17 1606 51
rect -1606 -119 -1572 -85
rect 1572 -51 1606 -17
rect -1606 -187 -1572 -153
rect -1606 -255 -1572 -221
rect -1606 -323 -1572 -289
rect -1606 -391 -1572 -357
rect -1606 -459 -1572 -425
rect -1606 -527 -1572 -493
rect -1606 -595 -1572 -561
rect -1606 -663 -1572 -629
rect -1606 -731 -1572 -697
rect 1572 -119 1606 -85
rect 1572 -187 1606 -153
rect 1572 -255 1606 -221
rect 1572 -323 1606 -289
rect 1572 -391 1606 -357
rect 1572 -459 1606 -425
rect 1572 -527 1606 -493
rect 1572 -595 1606 -561
rect 1572 -663 1606 -629
rect 1572 -731 1606 -697
rect -1606 -799 -1572 -765
rect 1572 -799 1606 -765
rect -1479 -901 -1445 -867
rect -1411 -901 -1377 -867
rect -1343 -901 -1309 -867
rect -1275 -901 -1241 -867
rect -1207 -901 -1173 -867
rect -1139 -901 -1105 -867
rect -1071 -901 -1037 -867
rect -1003 -901 -969 -867
rect -935 -901 -901 -867
rect -867 -901 -833 -867
rect -799 -901 -765 -867
rect -731 -901 -697 -867
rect -663 -901 -629 -867
rect -595 -901 -561 -867
rect -527 -901 -493 -867
rect -459 -901 -425 -867
rect -391 -901 -357 -867
rect -323 -901 -289 -867
rect -255 -901 -221 -867
rect -187 -901 -153 -867
rect -119 -901 -85 -867
rect -51 -901 -17 -867
rect 17 -901 51 -867
rect 85 -901 119 -867
rect 153 -901 187 -867
rect 221 -901 255 -867
rect 289 -901 323 -867
rect 357 -901 391 -867
rect 425 -901 459 -867
rect 493 -901 527 -867
rect 561 -901 595 -867
rect 629 -901 663 -867
rect 697 -901 731 -867
rect 765 -901 799 -867
rect 833 -901 867 -867
rect 901 -901 935 -867
rect 969 -901 1003 -867
rect 1037 -901 1071 -867
rect 1105 -901 1139 -867
rect 1173 -901 1207 -867
rect 1241 -901 1275 -867
rect 1309 -901 1343 -867
rect 1377 -901 1411 -867
rect 1445 -901 1479 -867
<< poly >>
rect -1449 749 -1383 815
rect -1331 749 -1265 815
rect -1213 749 -1147 815
rect -1095 749 -1029 815
rect -977 749 -911 815
rect -859 749 -793 815
rect -741 749 -675 815
rect -623 749 -557 815
rect -505 749 -439 815
rect -387 749 -321 815
rect -269 749 -203 815
rect -151 749 -85 815
rect -33 749 33 815
rect 85 749 151 815
rect 203 749 269 815
rect 321 749 387 815
rect 439 749 505 815
rect 557 749 623 815
rect 675 749 741 815
rect 793 749 859 815
rect 911 749 977 815
rect 1029 749 1095 815
rect 1147 749 1213 815
rect 1265 749 1331 815
rect 1383 749 1449 815
rect -1446 718 -1386 749
rect -1328 718 -1268 749
rect -1210 718 -1150 749
rect -1092 718 -1032 749
rect -974 718 -914 749
rect -856 718 -796 749
rect -738 718 -678 749
rect -620 718 -560 749
rect -502 718 -442 749
rect -384 718 -324 749
rect -266 718 -206 749
rect -148 718 -88 749
rect -30 718 30 749
rect 88 718 148 749
rect 206 718 266 749
rect 324 718 384 749
rect 442 718 502 749
rect 560 718 620 749
rect 678 718 738 749
rect 796 718 856 749
rect 914 718 974 749
rect 1032 718 1092 749
rect 1150 718 1210 749
rect 1268 718 1328 749
rect 1386 718 1446 749
rect -1446 87 -1386 118
rect -1328 87 -1268 118
rect -1210 87 -1150 118
rect -1092 87 -1032 118
rect -974 87 -914 118
rect -856 87 -796 118
rect -738 87 -678 118
rect -620 87 -560 118
rect -502 87 -442 118
rect -384 87 -324 118
rect -266 87 -206 118
rect -148 87 -88 118
rect -30 87 30 118
rect 88 87 148 118
rect 206 87 266 118
rect 324 87 384 118
rect 442 87 502 118
rect 560 87 620 118
rect 678 87 738 118
rect 796 87 856 118
rect 914 87 974 118
rect 1032 87 1092 118
rect 1150 87 1210 118
rect 1268 87 1328 118
rect 1386 87 1446 118
rect -1449 71 -1383 87
rect -1449 37 -1433 71
rect -1399 37 -1383 71
rect -1449 21 -1383 37
rect -1331 71 -1265 87
rect -1331 37 -1315 71
rect -1281 37 -1265 71
rect -1331 21 -1265 37
rect -1213 71 -1147 87
rect -1213 37 -1197 71
rect -1163 37 -1147 71
rect -1213 21 -1147 37
rect -1095 71 -1029 87
rect -1095 37 -1079 71
rect -1045 37 -1029 71
rect -1095 21 -1029 37
rect -977 71 -911 87
rect -977 37 -961 71
rect -927 37 -911 71
rect -977 21 -911 37
rect -859 71 -793 87
rect -859 37 -843 71
rect -809 37 -793 71
rect -859 21 -793 37
rect -741 71 -675 87
rect -741 37 -725 71
rect -691 37 -675 71
rect -741 21 -675 37
rect -623 71 -557 87
rect -623 37 -607 71
rect -573 37 -557 71
rect -623 21 -557 37
rect -505 71 -439 87
rect -505 37 -489 71
rect -455 37 -439 71
rect -505 21 -439 37
rect -387 71 -321 87
rect -387 37 -371 71
rect -337 37 -321 71
rect -387 21 -321 37
rect -269 71 -203 87
rect -269 37 -253 71
rect -219 37 -203 71
rect -269 21 -203 37
rect -151 71 -85 87
rect -151 37 -135 71
rect -101 37 -85 71
rect -151 21 -85 37
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect 85 71 151 87
rect 85 37 101 71
rect 135 37 151 71
rect 85 21 151 37
rect 203 71 269 87
rect 203 37 219 71
rect 253 37 269 71
rect 203 21 269 37
rect 321 71 387 87
rect 321 37 337 71
rect 371 37 387 71
rect 321 21 387 37
rect 439 71 505 87
rect 439 37 455 71
rect 489 37 505 71
rect 439 21 505 37
rect 557 71 623 87
rect 557 37 573 71
rect 607 37 623 71
rect 557 21 623 37
rect 675 71 741 87
rect 675 37 691 71
rect 725 37 741 71
rect 675 21 741 37
rect 793 71 859 87
rect 793 37 809 71
rect 843 37 859 71
rect 793 21 859 37
rect 911 71 977 87
rect 911 37 927 71
rect 961 37 977 71
rect 911 21 977 37
rect 1029 71 1095 87
rect 1029 37 1045 71
rect 1079 37 1095 71
rect 1029 21 1095 37
rect 1147 71 1213 87
rect 1147 37 1163 71
rect 1197 37 1213 71
rect 1147 21 1213 37
rect 1265 71 1331 87
rect 1265 37 1281 71
rect 1315 37 1331 71
rect 1265 21 1331 37
rect 1383 71 1449 87
rect 1383 37 1399 71
rect 1433 37 1449 71
rect 1383 21 1449 37
rect -1449 -37 -1383 -21
rect -1449 -71 -1433 -37
rect -1399 -71 -1383 -37
rect -1449 -87 -1383 -71
rect -1331 -37 -1265 -21
rect -1331 -71 -1315 -37
rect -1281 -71 -1265 -37
rect -1331 -87 -1265 -71
rect -1213 -37 -1147 -21
rect -1213 -71 -1197 -37
rect -1163 -71 -1147 -37
rect -1213 -87 -1147 -71
rect -1095 -37 -1029 -21
rect -1095 -71 -1079 -37
rect -1045 -71 -1029 -37
rect -1095 -87 -1029 -71
rect -977 -37 -911 -21
rect -977 -71 -961 -37
rect -927 -71 -911 -37
rect -977 -87 -911 -71
rect -859 -37 -793 -21
rect -859 -71 -843 -37
rect -809 -71 -793 -37
rect -859 -87 -793 -71
rect -741 -37 -675 -21
rect -741 -71 -725 -37
rect -691 -71 -675 -37
rect -741 -87 -675 -71
rect -623 -37 -557 -21
rect -623 -71 -607 -37
rect -573 -71 -557 -37
rect -623 -87 -557 -71
rect -505 -37 -439 -21
rect -505 -71 -489 -37
rect -455 -71 -439 -37
rect -505 -87 -439 -71
rect -387 -37 -321 -21
rect -387 -71 -371 -37
rect -337 -71 -321 -37
rect -387 -87 -321 -71
rect -269 -37 -203 -21
rect -269 -71 -253 -37
rect -219 -71 -203 -37
rect -269 -87 -203 -71
rect -151 -37 -85 -21
rect -151 -71 -135 -37
rect -101 -71 -85 -37
rect -151 -87 -85 -71
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect 85 -37 151 -21
rect 85 -71 101 -37
rect 135 -71 151 -37
rect 85 -87 151 -71
rect 203 -37 269 -21
rect 203 -71 219 -37
rect 253 -71 269 -37
rect 203 -87 269 -71
rect 321 -37 387 -21
rect 321 -71 337 -37
rect 371 -71 387 -37
rect 321 -87 387 -71
rect 439 -37 505 -21
rect 439 -71 455 -37
rect 489 -71 505 -37
rect 439 -87 505 -71
rect 557 -37 623 -21
rect 557 -71 573 -37
rect 607 -71 623 -37
rect 557 -87 623 -71
rect 675 -37 741 -21
rect 675 -71 691 -37
rect 725 -71 741 -37
rect 675 -87 741 -71
rect 793 -37 859 -21
rect 793 -71 809 -37
rect 843 -71 859 -37
rect 793 -87 859 -71
rect 911 -37 977 -21
rect 911 -71 927 -37
rect 961 -71 977 -37
rect 911 -87 977 -71
rect 1029 -37 1095 -21
rect 1029 -71 1045 -37
rect 1079 -71 1095 -37
rect 1029 -87 1095 -71
rect 1147 -37 1213 -21
rect 1147 -71 1163 -37
rect 1197 -71 1213 -37
rect 1147 -87 1213 -71
rect 1265 -37 1331 -21
rect 1265 -71 1281 -37
rect 1315 -71 1331 -37
rect 1265 -87 1331 -71
rect 1383 -37 1449 -21
rect 1383 -71 1399 -37
rect 1433 -71 1449 -37
rect 1383 -87 1449 -71
rect -1446 -118 -1386 -87
rect -1328 -118 -1268 -87
rect -1210 -118 -1150 -87
rect -1092 -118 -1032 -87
rect -974 -118 -914 -87
rect -856 -118 -796 -87
rect -738 -118 -678 -87
rect -620 -118 -560 -87
rect -502 -118 -442 -87
rect -384 -118 -324 -87
rect -266 -118 -206 -87
rect -148 -118 -88 -87
rect -30 -118 30 -87
rect 88 -118 148 -87
rect 206 -118 266 -87
rect 324 -118 384 -87
rect 442 -118 502 -87
rect 560 -118 620 -87
rect 678 -118 738 -87
rect 796 -118 856 -87
rect 914 -118 974 -87
rect 1032 -118 1092 -87
rect 1150 -118 1210 -87
rect 1268 -118 1328 -87
rect 1386 -118 1446 -87
rect -1446 -749 -1386 -718
rect -1328 -749 -1268 -718
rect -1210 -749 -1150 -718
rect -1092 -749 -1032 -718
rect -974 -749 -914 -718
rect -856 -749 -796 -718
rect -738 -749 -678 -718
rect -620 -749 -560 -718
rect -502 -749 -442 -718
rect -384 -749 -324 -718
rect -266 -749 -206 -718
rect -148 -749 -88 -718
rect -30 -749 30 -718
rect 88 -749 148 -718
rect 206 -749 266 -718
rect 324 -749 384 -718
rect 442 -749 502 -718
rect 560 -749 620 -718
rect 678 -749 738 -718
rect 796 -749 856 -718
rect 914 -749 974 -718
rect 1032 -749 1092 -718
rect 1150 -749 1210 -718
rect 1268 -749 1328 -718
rect 1386 -749 1446 -718
rect -1449 -815 -1383 -749
rect -1331 -815 -1265 -749
rect -1213 -815 -1147 -749
rect -1095 -815 -1029 -749
rect -977 -815 -911 -749
rect -859 -815 -793 -749
rect -741 -815 -675 -749
rect -623 -815 -557 -749
rect -505 -815 -439 -749
rect -387 -815 -321 -749
rect -269 -815 -203 -749
rect -151 -815 -85 -749
rect -33 -815 33 -749
rect 85 -815 151 -749
rect 203 -815 269 -749
rect 321 -815 387 -749
rect 439 -815 505 -749
rect 557 -815 623 -749
rect 675 -815 741 -749
rect 793 -815 859 -749
rect 911 -815 977 -749
rect 1029 -815 1095 -749
rect 1147 -815 1213 -749
rect 1265 -815 1331 -749
rect 1383 -815 1449 -749
<< polycont >>
rect -1433 37 -1399 71
rect -1315 37 -1281 71
rect -1197 37 -1163 71
rect -1079 37 -1045 71
rect -961 37 -927 71
rect -843 37 -809 71
rect -725 37 -691 71
rect -607 37 -573 71
rect -489 37 -455 71
rect -371 37 -337 71
rect -253 37 -219 71
rect -135 37 -101 71
rect -17 37 17 71
rect 101 37 135 71
rect 219 37 253 71
rect 337 37 371 71
rect 455 37 489 71
rect 573 37 607 71
rect 691 37 725 71
rect 809 37 843 71
rect 927 37 961 71
rect 1045 37 1079 71
rect 1163 37 1197 71
rect 1281 37 1315 71
rect 1399 37 1433 71
rect -1433 -71 -1399 -37
rect -1315 -71 -1281 -37
rect -1197 -71 -1163 -37
rect -1079 -71 -1045 -37
rect -961 -71 -927 -37
rect -843 -71 -809 -37
rect -725 -71 -691 -37
rect -607 -71 -573 -37
rect -489 -71 -455 -37
rect -371 -71 -337 -37
rect -253 -71 -219 -37
rect -135 -71 -101 -37
rect -17 -71 17 -37
rect 101 -71 135 -37
rect 219 -71 253 -37
rect 337 -71 371 -37
rect 455 -71 489 -37
rect 573 -71 607 -37
rect 691 -71 725 -37
rect 809 -71 843 -37
rect 927 -71 961 -37
rect 1045 -71 1079 -37
rect 1163 -71 1197 -37
rect 1281 -71 1315 -37
rect 1399 -71 1433 -37
<< locali >>
rect -1606 867 -1479 901
rect -1445 867 -1411 901
rect -1377 867 -1343 901
rect -1309 867 -1275 901
rect -1241 867 -1207 901
rect -1173 867 -1139 901
rect -1105 867 -1071 901
rect -1037 867 -1003 901
rect -969 867 -935 901
rect -901 867 -867 901
rect -833 867 -799 901
rect -765 867 -731 901
rect -697 867 -663 901
rect -629 867 -595 901
rect -561 867 -527 901
rect -493 867 -459 901
rect -425 867 -391 901
rect -357 867 -323 901
rect -289 867 -255 901
rect -221 867 -187 901
rect -153 867 -119 901
rect -85 867 -51 901
rect -17 867 17 901
rect 51 867 85 901
rect 119 867 153 901
rect 187 867 221 901
rect 255 867 289 901
rect 323 867 357 901
rect 391 867 425 901
rect 459 867 493 901
rect 527 867 561 901
rect 595 867 629 901
rect 663 867 697 901
rect 731 867 765 901
rect 799 867 833 901
rect 867 867 901 901
rect 935 867 969 901
rect 1003 867 1037 901
rect 1071 867 1105 901
rect 1139 867 1173 901
rect 1207 867 1241 901
rect 1275 867 1309 901
rect 1343 867 1377 901
rect 1411 867 1445 901
rect 1479 867 1606 901
rect -1606 799 -1572 867
rect -1606 731 -1572 765
rect 1572 799 1606 867
rect 1572 731 1606 765
rect -1606 663 -1572 697
rect -1606 595 -1572 629
rect -1606 527 -1572 561
rect -1606 459 -1572 493
rect -1606 391 -1572 425
rect -1606 323 -1572 357
rect -1606 255 -1572 289
rect -1606 187 -1572 221
rect -1606 119 -1572 153
rect -1492 687 -1458 722
rect -1492 615 -1458 639
rect -1492 543 -1458 571
rect -1492 471 -1458 503
rect -1492 401 -1458 435
rect -1492 333 -1458 365
rect -1492 265 -1458 293
rect -1492 197 -1458 221
rect -1492 114 -1458 149
rect -1374 687 -1340 722
rect -1374 615 -1340 639
rect -1374 543 -1340 571
rect -1374 471 -1340 503
rect -1374 401 -1340 435
rect -1374 333 -1340 365
rect -1374 265 -1340 293
rect -1374 197 -1340 221
rect -1374 114 -1340 149
rect -1256 687 -1222 722
rect -1256 615 -1222 639
rect -1256 543 -1222 571
rect -1256 471 -1222 503
rect -1256 401 -1222 435
rect -1256 333 -1222 365
rect -1256 265 -1222 293
rect -1256 197 -1222 221
rect -1256 114 -1222 149
rect -1138 687 -1104 722
rect -1138 615 -1104 639
rect -1138 543 -1104 571
rect -1138 471 -1104 503
rect -1138 401 -1104 435
rect -1138 333 -1104 365
rect -1138 265 -1104 293
rect -1138 197 -1104 221
rect -1138 114 -1104 149
rect -1020 687 -986 722
rect -1020 615 -986 639
rect -1020 543 -986 571
rect -1020 471 -986 503
rect -1020 401 -986 435
rect -1020 333 -986 365
rect -1020 265 -986 293
rect -1020 197 -986 221
rect -1020 114 -986 149
rect -902 687 -868 722
rect -902 615 -868 639
rect -902 543 -868 571
rect -902 471 -868 503
rect -902 401 -868 435
rect -902 333 -868 365
rect -902 265 -868 293
rect -902 197 -868 221
rect -902 114 -868 149
rect -784 687 -750 722
rect -784 615 -750 639
rect -784 543 -750 571
rect -784 471 -750 503
rect -784 401 -750 435
rect -784 333 -750 365
rect -784 265 -750 293
rect -784 197 -750 221
rect -784 114 -750 149
rect -666 687 -632 722
rect -666 615 -632 639
rect -666 543 -632 571
rect -666 471 -632 503
rect -666 401 -632 435
rect -666 333 -632 365
rect -666 265 -632 293
rect -666 197 -632 221
rect -666 114 -632 149
rect -548 687 -514 722
rect -548 615 -514 639
rect -548 543 -514 571
rect -548 471 -514 503
rect -548 401 -514 435
rect -548 333 -514 365
rect -548 265 -514 293
rect -548 197 -514 221
rect -548 114 -514 149
rect -430 687 -396 722
rect -430 615 -396 639
rect -430 543 -396 571
rect -430 471 -396 503
rect -430 401 -396 435
rect -430 333 -396 365
rect -430 265 -396 293
rect -430 197 -396 221
rect -430 114 -396 149
rect -312 687 -278 722
rect -312 615 -278 639
rect -312 543 -278 571
rect -312 471 -278 503
rect -312 401 -278 435
rect -312 333 -278 365
rect -312 265 -278 293
rect -312 197 -278 221
rect -312 114 -278 149
rect -194 687 -160 722
rect -194 615 -160 639
rect -194 543 -160 571
rect -194 471 -160 503
rect -194 401 -160 435
rect -194 333 -160 365
rect -194 265 -160 293
rect -194 197 -160 221
rect -194 114 -160 149
rect -76 687 -42 722
rect -76 615 -42 639
rect -76 543 -42 571
rect -76 471 -42 503
rect -76 401 -42 435
rect -76 333 -42 365
rect -76 265 -42 293
rect -76 197 -42 221
rect -76 114 -42 149
rect 42 687 76 722
rect 42 615 76 639
rect 42 543 76 571
rect 42 471 76 503
rect 42 401 76 435
rect 42 333 76 365
rect 42 265 76 293
rect 42 197 76 221
rect 42 114 76 149
rect 160 687 194 722
rect 160 615 194 639
rect 160 543 194 571
rect 160 471 194 503
rect 160 401 194 435
rect 160 333 194 365
rect 160 265 194 293
rect 160 197 194 221
rect 160 114 194 149
rect 278 687 312 722
rect 278 615 312 639
rect 278 543 312 571
rect 278 471 312 503
rect 278 401 312 435
rect 278 333 312 365
rect 278 265 312 293
rect 278 197 312 221
rect 278 114 312 149
rect 396 687 430 722
rect 396 615 430 639
rect 396 543 430 571
rect 396 471 430 503
rect 396 401 430 435
rect 396 333 430 365
rect 396 265 430 293
rect 396 197 430 221
rect 396 114 430 149
rect 514 687 548 722
rect 514 615 548 639
rect 514 543 548 571
rect 514 471 548 503
rect 514 401 548 435
rect 514 333 548 365
rect 514 265 548 293
rect 514 197 548 221
rect 514 114 548 149
rect 632 687 666 722
rect 632 615 666 639
rect 632 543 666 571
rect 632 471 666 503
rect 632 401 666 435
rect 632 333 666 365
rect 632 265 666 293
rect 632 197 666 221
rect 632 114 666 149
rect 750 687 784 722
rect 750 615 784 639
rect 750 543 784 571
rect 750 471 784 503
rect 750 401 784 435
rect 750 333 784 365
rect 750 265 784 293
rect 750 197 784 221
rect 750 114 784 149
rect 868 687 902 722
rect 868 615 902 639
rect 868 543 902 571
rect 868 471 902 503
rect 868 401 902 435
rect 868 333 902 365
rect 868 265 902 293
rect 868 197 902 221
rect 868 114 902 149
rect 986 687 1020 722
rect 986 615 1020 639
rect 986 543 1020 571
rect 986 471 1020 503
rect 986 401 1020 435
rect 986 333 1020 365
rect 986 265 1020 293
rect 986 197 1020 221
rect 986 114 1020 149
rect 1104 687 1138 722
rect 1104 615 1138 639
rect 1104 543 1138 571
rect 1104 471 1138 503
rect 1104 401 1138 435
rect 1104 333 1138 365
rect 1104 265 1138 293
rect 1104 197 1138 221
rect 1104 114 1138 149
rect 1222 687 1256 722
rect 1222 615 1256 639
rect 1222 543 1256 571
rect 1222 471 1256 503
rect 1222 401 1256 435
rect 1222 333 1256 365
rect 1222 265 1256 293
rect 1222 197 1256 221
rect 1222 114 1256 149
rect 1340 687 1374 722
rect 1340 615 1374 639
rect 1340 543 1374 571
rect 1340 471 1374 503
rect 1340 401 1374 435
rect 1340 333 1374 365
rect 1340 265 1374 293
rect 1340 197 1374 221
rect 1340 114 1374 149
rect 1458 687 1492 722
rect 1458 615 1492 639
rect 1458 543 1492 571
rect 1458 471 1492 503
rect 1458 401 1492 435
rect 1458 333 1492 365
rect 1458 265 1492 293
rect 1458 197 1492 221
rect 1458 114 1492 149
rect 1572 663 1606 697
rect 1572 595 1606 629
rect 1572 527 1606 561
rect 1572 459 1606 493
rect 1572 391 1606 425
rect 1572 323 1606 357
rect 1572 255 1606 289
rect 1572 187 1606 221
rect 1572 119 1606 153
rect -1606 51 -1572 85
rect -1449 37 -1433 71
rect -1399 37 -1383 71
rect -1331 37 -1315 71
rect -1281 37 -1265 71
rect -1213 37 -1197 71
rect -1163 37 -1147 71
rect -1095 37 -1079 71
rect -1045 37 -1029 71
rect -977 37 -961 71
rect -927 37 -911 71
rect -859 37 -843 71
rect -809 37 -793 71
rect -741 37 -725 71
rect -691 37 -675 71
rect -623 37 -607 71
rect -573 37 -557 71
rect -505 37 -489 71
rect -455 37 -439 71
rect -387 37 -371 71
rect -337 37 -321 71
rect -269 37 -253 71
rect -219 37 -203 71
rect -151 37 -135 71
rect -101 37 -85 71
rect -33 37 -17 71
rect 17 37 33 71
rect 85 37 101 71
rect 135 37 151 71
rect 203 37 219 71
rect 253 37 269 71
rect 321 37 337 71
rect 371 37 387 71
rect 439 37 455 71
rect 489 37 505 71
rect 557 37 573 71
rect 607 37 623 71
rect 675 37 691 71
rect 725 37 741 71
rect 793 37 809 71
rect 843 37 859 71
rect 911 37 927 71
rect 961 37 977 71
rect 1029 37 1045 71
rect 1079 37 1095 71
rect 1147 37 1163 71
rect 1197 37 1213 71
rect 1265 37 1281 71
rect 1315 37 1331 71
rect 1383 37 1399 71
rect 1433 37 1449 71
rect 1572 51 1606 85
rect -1606 -17 -1572 17
rect 1572 -17 1606 17
rect -1606 -85 -1572 -51
rect -1449 -71 -1433 -37
rect -1399 -71 -1383 -37
rect -1331 -71 -1315 -37
rect -1281 -71 -1265 -37
rect -1213 -71 -1197 -37
rect -1163 -71 -1147 -37
rect -1095 -71 -1079 -37
rect -1045 -71 -1029 -37
rect -977 -71 -961 -37
rect -927 -71 -911 -37
rect -859 -71 -843 -37
rect -809 -71 -793 -37
rect -741 -71 -725 -37
rect -691 -71 -675 -37
rect -623 -71 -607 -37
rect -573 -71 -557 -37
rect -505 -71 -489 -37
rect -455 -71 -439 -37
rect -387 -71 -371 -37
rect -337 -71 -321 -37
rect -269 -71 -253 -37
rect -219 -71 -203 -37
rect -151 -71 -135 -37
rect -101 -71 -85 -37
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect 85 -71 101 -37
rect 135 -71 151 -37
rect 203 -71 219 -37
rect 253 -71 269 -37
rect 321 -71 337 -37
rect 371 -71 387 -37
rect 439 -71 455 -37
rect 489 -71 505 -37
rect 557 -71 573 -37
rect 607 -71 623 -37
rect 675 -71 691 -37
rect 725 -71 741 -37
rect 793 -71 809 -37
rect 843 -71 859 -37
rect 911 -71 927 -37
rect 961 -71 977 -37
rect 1029 -71 1045 -37
rect 1079 -71 1095 -37
rect 1147 -71 1163 -37
rect 1197 -71 1213 -37
rect 1265 -71 1281 -37
rect 1315 -71 1331 -37
rect 1383 -71 1399 -37
rect 1433 -71 1449 -37
rect 1572 -85 1606 -51
rect -1606 -153 -1572 -119
rect -1606 -221 -1572 -187
rect -1606 -289 -1572 -255
rect -1606 -357 -1572 -323
rect -1606 -425 -1572 -391
rect -1606 -493 -1572 -459
rect -1606 -561 -1572 -527
rect -1606 -629 -1572 -595
rect -1606 -697 -1572 -663
rect -1492 -149 -1458 -114
rect -1492 -221 -1458 -197
rect -1492 -293 -1458 -265
rect -1492 -365 -1458 -333
rect -1492 -435 -1458 -401
rect -1492 -503 -1458 -471
rect -1492 -571 -1458 -543
rect -1492 -639 -1458 -615
rect -1492 -722 -1458 -687
rect -1374 -149 -1340 -114
rect -1374 -221 -1340 -197
rect -1374 -293 -1340 -265
rect -1374 -365 -1340 -333
rect -1374 -435 -1340 -401
rect -1374 -503 -1340 -471
rect -1374 -571 -1340 -543
rect -1374 -639 -1340 -615
rect -1374 -722 -1340 -687
rect -1256 -149 -1222 -114
rect -1256 -221 -1222 -197
rect -1256 -293 -1222 -265
rect -1256 -365 -1222 -333
rect -1256 -435 -1222 -401
rect -1256 -503 -1222 -471
rect -1256 -571 -1222 -543
rect -1256 -639 -1222 -615
rect -1256 -722 -1222 -687
rect -1138 -149 -1104 -114
rect -1138 -221 -1104 -197
rect -1138 -293 -1104 -265
rect -1138 -365 -1104 -333
rect -1138 -435 -1104 -401
rect -1138 -503 -1104 -471
rect -1138 -571 -1104 -543
rect -1138 -639 -1104 -615
rect -1138 -722 -1104 -687
rect -1020 -149 -986 -114
rect -1020 -221 -986 -197
rect -1020 -293 -986 -265
rect -1020 -365 -986 -333
rect -1020 -435 -986 -401
rect -1020 -503 -986 -471
rect -1020 -571 -986 -543
rect -1020 -639 -986 -615
rect -1020 -722 -986 -687
rect -902 -149 -868 -114
rect -902 -221 -868 -197
rect -902 -293 -868 -265
rect -902 -365 -868 -333
rect -902 -435 -868 -401
rect -902 -503 -868 -471
rect -902 -571 -868 -543
rect -902 -639 -868 -615
rect -902 -722 -868 -687
rect -784 -149 -750 -114
rect -784 -221 -750 -197
rect -784 -293 -750 -265
rect -784 -365 -750 -333
rect -784 -435 -750 -401
rect -784 -503 -750 -471
rect -784 -571 -750 -543
rect -784 -639 -750 -615
rect -784 -722 -750 -687
rect -666 -149 -632 -114
rect -666 -221 -632 -197
rect -666 -293 -632 -265
rect -666 -365 -632 -333
rect -666 -435 -632 -401
rect -666 -503 -632 -471
rect -666 -571 -632 -543
rect -666 -639 -632 -615
rect -666 -722 -632 -687
rect -548 -149 -514 -114
rect -548 -221 -514 -197
rect -548 -293 -514 -265
rect -548 -365 -514 -333
rect -548 -435 -514 -401
rect -548 -503 -514 -471
rect -548 -571 -514 -543
rect -548 -639 -514 -615
rect -548 -722 -514 -687
rect -430 -149 -396 -114
rect -430 -221 -396 -197
rect -430 -293 -396 -265
rect -430 -365 -396 -333
rect -430 -435 -396 -401
rect -430 -503 -396 -471
rect -430 -571 -396 -543
rect -430 -639 -396 -615
rect -430 -722 -396 -687
rect -312 -149 -278 -114
rect -312 -221 -278 -197
rect -312 -293 -278 -265
rect -312 -365 -278 -333
rect -312 -435 -278 -401
rect -312 -503 -278 -471
rect -312 -571 -278 -543
rect -312 -639 -278 -615
rect -312 -722 -278 -687
rect -194 -149 -160 -114
rect -194 -221 -160 -197
rect -194 -293 -160 -265
rect -194 -365 -160 -333
rect -194 -435 -160 -401
rect -194 -503 -160 -471
rect -194 -571 -160 -543
rect -194 -639 -160 -615
rect -194 -722 -160 -687
rect -76 -149 -42 -114
rect -76 -221 -42 -197
rect -76 -293 -42 -265
rect -76 -365 -42 -333
rect -76 -435 -42 -401
rect -76 -503 -42 -471
rect -76 -571 -42 -543
rect -76 -639 -42 -615
rect -76 -722 -42 -687
rect 42 -149 76 -114
rect 42 -221 76 -197
rect 42 -293 76 -265
rect 42 -365 76 -333
rect 42 -435 76 -401
rect 42 -503 76 -471
rect 42 -571 76 -543
rect 42 -639 76 -615
rect 42 -722 76 -687
rect 160 -149 194 -114
rect 160 -221 194 -197
rect 160 -293 194 -265
rect 160 -365 194 -333
rect 160 -435 194 -401
rect 160 -503 194 -471
rect 160 -571 194 -543
rect 160 -639 194 -615
rect 160 -722 194 -687
rect 278 -149 312 -114
rect 278 -221 312 -197
rect 278 -293 312 -265
rect 278 -365 312 -333
rect 278 -435 312 -401
rect 278 -503 312 -471
rect 278 -571 312 -543
rect 278 -639 312 -615
rect 278 -722 312 -687
rect 396 -149 430 -114
rect 396 -221 430 -197
rect 396 -293 430 -265
rect 396 -365 430 -333
rect 396 -435 430 -401
rect 396 -503 430 -471
rect 396 -571 430 -543
rect 396 -639 430 -615
rect 396 -722 430 -687
rect 514 -149 548 -114
rect 514 -221 548 -197
rect 514 -293 548 -265
rect 514 -365 548 -333
rect 514 -435 548 -401
rect 514 -503 548 -471
rect 514 -571 548 -543
rect 514 -639 548 -615
rect 514 -722 548 -687
rect 632 -149 666 -114
rect 632 -221 666 -197
rect 632 -293 666 -265
rect 632 -365 666 -333
rect 632 -435 666 -401
rect 632 -503 666 -471
rect 632 -571 666 -543
rect 632 -639 666 -615
rect 632 -722 666 -687
rect 750 -149 784 -114
rect 750 -221 784 -197
rect 750 -293 784 -265
rect 750 -365 784 -333
rect 750 -435 784 -401
rect 750 -503 784 -471
rect 750 -571 784 -543
rect 750 -639 784 -615
rect 750 -722 784 -687
rect 868 -149 902 -114
rect 868 -221 902 -197
rect 868 -293 902 -265
rect 868 -365 902 -333
rect 868 -435 902 -401
rect 868 -503 902 -471
rect 868 -571 902 -543
rect 868 -639 902 -615
rect 868 -722 902 -687
rect 986 -149 1020 -114
rect 986 -221 1020 -197
rect 986 -293 1020 -265
rect 986 -365 1020 -333
rect 986 -435 1020 -401
rect 986 -503 1020 -471
rect 986 -571 1020 -543
rect 986 -639 1020 -615
rect 986 -722 1020 -687
rect 1104 -149 1138 -114
rect 1104 -221 1138 -197
rect 1104 -293 1138 -265
rect 1104 -365 1138 -333
rect 1104 -435 1138 -401
rect 1104 -503 1138 -471
rect 1104 -571 1138 -543
rect 1104 -639 1138 -615
rect 1104 -722 1138 -687
rect 1222 -149 1256 -114
rect 1222 -221 1256 -197
rect 1222 -293 1256 -265
rect 1222 -365 1256 -333
rect 1222 -435 1256 -401
rect 1222 -503 1256 -471
rect 1222 -571 1256 -543
rect 1222 -639 1256 -615
rect 1222 -722 1256 -687
rect 1340 -149 1374 -114
rect 1340 -221 1374 -197
rect 1340 -293 1374 -265
rect 1340 -365 1374 -333
rect 1340 -435 1374 -401
rect 1340 -503 1374 -471
rect 1340 -571 1374 -543
rect 1340 -639 1374 -615
rect 1340 -722 1374 -687
rect 1458 -149 1492 -114
rect 1458 -221 1492 -197
rect 1458 -293 1492 -265
rect 1458 -365 1492 -333
rect 1458 -435 1492 -401
rect 1458 -503 1492 -471
rect 1458 -571 1492 -543
rect 1458 -639 1492 -615
rect 1458 -722 1492 -687
rect 1572 -153 1606 -119
rect 1572 -221 1606 -187
rect 1572 -289 1606 -255
rect 1572 -357 1606 -323
rect 1572 -425 1606 -391
rect 1572 -493 1606 -459
rect 1572 -561 1606 -527
rect 1572 -629 1606 -595
rect 1572 -697 1606 -663
rect -1606 -765 -1572 -731
rect -1606 -867 -1572 -799
rect 1572 -765 1606 -731
rect 1572 -867 1606 -799
rect -1606 -901 -1479 -867
rect -1445 -901 -1411 -867
rect -1377 -901 -1343 -867
rect -1309 -901 -1275 -867
rect -1241 -901 -1207 -867
rect -1173 -901 -1139 -867
rect -1105 -901 -1071 -867
rect -1037 -901 -1003 -867
rect -969 -901 -935 -867
rect -901 -901 -867 -867
rect -833 -901 -799 -867
rect -765 -901 -731 -867
rect -697 -901 -663 -867
rect -629 -901 -595 -867
rect -561 -901 -527 -867
rect -493 -901 -459 -867
rect -425 -901 -391 -867
rect -357 -901 -323 -867
rect -289 -901 -255 -867
rect -221 -901 -187 -867
rect -153 -901 -119 -867
rect -85 -901 -51 -867
rect -17 -901 17 -867
rect 51 -901 85 -867
rect 119 -901 153 -867
rect 187 -901 221 -867
rect 255 -901 289 -867
rect 323 -901 357 -867
rect 391 -901 425 -867
rect 459 -901 493 -867
rect 527 -901 561 -867
rect 595 -901 629 -867
rect 663 -901 697 -867
rect 731 -901 765 -867
rect 799 -901 833 -867
rect 867 -901 901 -867
rect 935 -901 969 -867
rect 1003 -901 1037 -867
rect 1071 -901 1105 -867
rect 1139 -901 1173 -867
rect 1207 -901 1241 -867
rect 1275 -901 1309 -867
rect 1343 -901 1377 -867
rect 1411 -901 1445 -867
rect 1479 -901 1606 -867
<< viali >>
rect -1492 673 -1458 687
rect -1492 653 -1458 673
rect -1492 605 -1458 615
rect -1492 581 -1458 605
rect -1492 537 -1458 543
rect -1492 509 -1458 537
rect -1492 469 -1458 471
rect -1492 437 -1458 469
rect -1492 367 -1458 399
rect -1492 365 -1458 367
rect -1492 299 -1458 327
rect -1492 293 -1458 299
rect -1492 231 -1458 255
rect -1492 221 -1458 231
rect -1492 163 -1458 183
rect -1492 149 -1458 163
rect -1374 673 -1340 687
rect -1374 653 -1340 673
rect -1374 605 -1340 615
rect -1374 581 -1340 605
rect -1374 537 -1340 543
rect -1374 509 -1340 537
rect -1374 469 -1340 471
rect -1374 437 -1340 469
rect -1374 367 -1340 399
rect -1374 365 -1340 367
rect -1374 299 -1340 327
rect -1374 293 -1340 299
rect -1374 231 -1340 255
rect -1374 221 -1340 231
rect -1374 163 -1340 183
rect -1374 149 -1340 163
rect -1256 673 -1222 687
rect -1256 653 -1222 673
rect -1256 605 -1222 615
rect -1256 581 -1222 605
rect -1256 537 -1222 543
rect -1256 509 -1222 537
rect -1256 469 -1222 471
rect -1256 437 -1222 469
rect -1256 367 -1222 399
rect -1256 365 -1222 367
rect -1256 299 -1222 327
rect -1256 293 -1222 299
rect -1256 231 -1222 255
rect -1256 221 -1222 231
rect -1256 163 -1222 183
rect -1256 149 -1222 163
rect -1138 673 -1104 687
rect -1138 653 -1104 673
rect -1138 605 -1104 615
rect -1138 581 -1104 605
rect -1138 537 -1104 543
rect -1138 509 -1104 537
rect -1138 469 -1104 471
rect -1138 437 -1104 469
rect -1138 367 -1104 399
rect -1138 365 -1104 367
rect -1138 299 -1104 327
rect -1138 293 -1104 299
rect -1138 231 -1104 255
rect -1138 221 -1104 231
rect -1138 163 -1104 183
rect -1138 149 -1104 163
rect -1020 673 -986 687
rect -1020 653 -986 673
rect -1020 605 -986 615
rect -1020 581 -986 605
rect -1020 537 -986 543
rect -1020 509 -986 537
rect -1020 469 -986 471
rect -1020 437 -986 469
rect -1020 367 -986 399
rect -1020 365 -986 367
rect -1020 299 -986 327
rect -1020 293 -986 299
rect -1020 231 -986 255
rect -1020 221 -986 231
rect -1020 163 -986 183
rect -1020 149 -986 163
rect -902 673 -868 687
rect -902 653 -868 673
rect -902 605 -868 615
rect -902 581 -868 605
rect -902 537 -868 543
rect -902 509 -868 537
rect -902 469 -868 471
rect -902 437 -868 469
rect -902 367 -868 399
rect -902 365 -868 367
rect -902 299 -868 327
rect -902 293 -868 299
rect -902 231 -868 255
rect -902 221 -868 231
rect -902 163 -868 183
rect -902 149 -868 163
rect -784 673 -750 687
rect -784 653 -750 673
rect -784 605 -750 615
rect -784 581 -750 605
rect -784 537 -750 543
rect -784 509 -750 537
rect -784 469 -750 471
rect -784 437 -750 469
rect -784 367 -750 399
rect -784 365 -750 367
rect -784 299 -750 327
rect -784 293 -750 299
rect -784 231 -750 255
rect -784 221 -750 231
rect -784 163 -750 183
rect -784 149 -750 163
rect -666 673 -632 687
rect -666 653 -632 673
rect -666 605 -632 615
rect -666 581 -632 605
rect -666 537 -632 543
rect -666 509 -632 537
rect -666 469 -632 471
rect -666 437 -632 469
rect -666 367 -632 399
rect -666 365 -632 367
rect -666 299 -632 327
rect -666 293 -632 299
rect -666 231 -632 255
rect -666 221 -632 231
rect -666 163 -632 183
rect -666 149 -632 163
rect -548 673 -514 687
rect -548 653 -514 673
rect -548 605 -514 615
rect -548 581 -514 605
rect -548 537 -514 543
rect -548 509 -514 537
rect -548 469 -514 471
rect -548 437 -514 469
rect -548 367 -514 399
rect -548 365 -514 367
rect -548 299 -514 327
rect -548 293 -514 299
rect -548 231 -514 255
rect -548 221 -514 231
rect -548 163 -514 183
rect -548 149 -514 163
rect -430 673 -396 687
rect -430 653 -396 673
rect -430 605 -396 615
rect -430 581 -396 605
rect -430 537 -396 543
rect -430 509 -396 537
rect -430 469 -396 471
rect -430 437 -396 469
rect -430 367 -396 399
rect -430 365 -396 367
rect -430 299 -396 327
rect -430 293 -396 299
rect -430 231 -396 255
rect -430 221 -396 231
rect -430 163 -396 183
rect -430 149 -396 163
rect -312 673 -278 687
rect -312 653 -278 673
rect -312 605 -278 615
rect -312 581 -278 605
rect -312 537 -278 543
rect -312 509 -278 537
rect -312 469 -278 471
rect -312 437 -278 469
rect -312 367 -278 399
rect -312 365 -278 367
rect -312 299 -278 327
rect -312 293 -278 299
rect -312 231 -278 255
rect -312 221 -278 231
rect -312 163 -278 183
rect -312 149 -278 163
rect -194 673 -160 687
rect -194 653 -160 673
rect -194 605 -160 615
rect -194 581 -160 605
rect -194 537 -160 543
rect -194 509 -160 537
rect -194 469 -160 471
rect -194 437 -160 469
rect -194 367 -160 399
rect -194 365 -160 367
rect -194 299 -160 327
rect -194 293 -160 299
rect -194 231 -160 255
rect -194 221 -160 231
rect -194 163 -160 183
rect -194 149 -160 163
rect -76 673 -42 687
rect -76 653 -42 673
rect -76 605 -42 615
rect -76 581 -42 605
rect -76 537 -42 543
rect -76 509 -42 537
rect -76 469 -42 471
rect -76 437 -42 469
rect -76 367 -42 399
rect -76 365 -42 367
rect -76 299 -42 327
rect -76 293 -42 299
rect -76 231 -42 255
rect -76 221 -42 231
rect -76 163 -42 183
rect -76 149 -42 163
rect 42 673 76 687
rect 42 653 76 673
rect 42 605 76 615
rect 42 581 76 605
rect 42 537 76 543
rect 42 509 76 537
rect 42 469 76 471
rect 42 437 76 469
rect 42 367 76 399
rect 42 365 76 367
rect 42 299 76 327
rect 42 293 76 299
rect 42 231 76 255
rect 42 221 76 231
rect 42 163 76 183
rect 42 149 76 163
rect 160 673 194 687
rect 160 653 194 673
rect 160 605 194 615
rect 160 581 194 605
rect 160 537 194 543
rect 160 509 194 537
rect 160 469 194 471
rect 160 437 194 469
rect 160 367 194 399
rect 160 365 194 367
rect 160 299 194 327
rect 160 293 194 299
rect 160 231 194 255
rect 160 221 194 231
rect 160 163 194 183
rect 160 149 194 163
rect 278 673 312 687
rect 278 653 312 673
rect 278 605 312 615
rect 278 581 312 605
rect 278 537 312 543
rect 278 509 312 537
rect 278 469 312 471
rect 278 437 312 469
rect 278 367 312 399
rect 278 365 312 367
rect 278 299 312 327
rect 278 293 312 299
rect 278 231 312 255
rect 278 221 312 231
rect 278 163 312 183
rect 278 149 312 163
rect 396 673 430 687
rect 396 653 430 673
rect 396 605 430 615
rect 396 581 430 605
rect 396 537 430 543
rect 396 509 430 537
rect 396 469 430 471
rect 396 437 430 469
rect 396 367 430 399
rect 396 365 430 367
rect 396 299 430 327
rect 396 293 430 299
rect 396 231 430 255
rect 396 221 430 231
rect 396 163 430 183
rect 396 149 430 163
rect 514 673 548 687
rect 514 653 548 673
rect 514 605 548 615
rect 514 581 548 605
rect 514 537 548 543
rect 514 509 548 537
rect 514 469 548 471
rect 514 437 548 469
rect 514 367 548 399
rect 514 365 548 367
rect 514 299 548 327
rect 514 293 548 299
rect 514 231 548 255
rect 514 221 548 231
rect 514 163 548 183
rect 514 149 548 163
rect 632 673 666 687
rect 632 653 666 673
rect 632 605 666 615
rect 632 581 666 605
rect 632 537 666 543
rect 632 509 666 537
rect 632 469 666 471
rect 632 437 666 469
rect 632 367 666 399
rect 632 365 666 367
rect 632 299 666 327
rect 632 293 666 299
rect 632 231 666 255
rect 632 221 666 231
rect 632 163 666 183
rect 632 149 666 163
rect 750 673 784 687
rect 750 653 784 673
rect 750 605 784 615
rect 750 581 784 605
rect 750 537 784 543
rect 750 509 784 537
rect 750 469 784 471
rect 750 437 784 469
rect 750 367 784 399
rect 750 365 784 367
rect 750 299 784 327
rect 750 293 784 299
rect 750 231 784 255
rect 750 221 784 231
rect 750 163 784 183
rect 750 149 784 163
rect 868 673 902 687
rect 868 653 902 673
rect 868 605 902 615
rect 868 581 902 605
rect 868 537 902 543
rect 868 509 902 537
rect 868 469 902 471
rect 868 437 902 469
rect 868 367 902 399
rect 868 365 902 367
rect 868 299 902 327
rect 868 293 902 299
rect 868 231 902 255
rect 868 221 902 231
rect 868 163 902 183
rect 868 149 902 163
rect 986 673 1020 687
rect 986 653 1020 673
rect 986 605 1020 615
rect 986 581 1020 605
rect 986 537 1020 543
rect 986 509 1020 537
rect 986 469 1020 471
rect 986 437 1020 469
rect 986 367 1020 399
rect 986 365 1020 367
rect 986 299 1020 327
rect 986 293 1020 299
rect 986 231 1020 255
rect 986 221 1020 231
rect 986 163 1020 183
rect 986 149 1020 163
rect 1104 673 1138 687
rect 1104 653 1138 673
rect 1104 605 1138 615
rect 1104 581 1138 605
rect 1104 537 1138 543
rect 1104 509 1138 537
rect 1104 469 1138 471
rect 1104 437 1138 469
rect 1104 367 1138 399
rect 1104 365 1138 367
rect 1104 299 1138 327
rect 1104 293 1138 299
rect 1104 231 1138 255
rect 1104 221 1138 231
rect 1104 163 1138 183
rect 1104 149 1138 163
rect 1222 673 1256 687
rect 1222 653 1256 673
rect 1222 605 1256 615
rect 1222 581 1256 605
rect 1222 537 1256 543
rect 1222 509 1256 537
rect 1222 469 1256 471
rect 1222 437 1256 469
rect 1222 367 1256 399
rect 1222 365 1256 367
rect 1222 299 1256 327
rect 1222 293 1256 299
rect 1222 231 1256 255
rect 1222 221 1256 231
rect 1222 163 1256 183
rect 1222 149 1256 163
rect 1340 673 1374 687
rect 1340 653 1374 673
rect 1340 605 1374 615
rect 1340 581 1374 605
rect 1340 537 1374 543
rect 1340 509 1374 537
rect 1340 469 1374 471
rect 1340 437 1374 469
rect 1340 367 1374 399
rect 1340 365 1374 367
rect 1340 299 1374 327
rect 1340 293 1374 299
rect 1340 231 1374 255
rect 1340 221 1374 231
rect 1340 163 1374 183
rect 1340 149 1374 163
rect 1458 673 1492 687
rect 1458 653 1492 673
rect 1458 605 1492 615
rect 1458 581 1492 605
rect 1458 537 1492 543
rect 1458 509 1492 537
rect 1458 469 1492 471
rect 1458 437 1492 469
rect 1458 367 1492 399
rect 1458 365 1492 367
rect 1458 299 1492 327
rect 1458 293 1492 299
rect 1458 231 1492 255
rect 1458 221 1492 231
rect 1458 163 1492 183
rect 1458 149 1492 163
rect -1433 37 -1399 71
rect -1315 37 -1281 71
rect -1197 37 -1163 71
rect -1079 37 -1045 71
rect -961 37 -927 71
rect -843 37 -809 71
rect -725 37 -691 71
rect -607 37 -573 71
rect -489 37 -455 71
rect -371 37 -337 71
rect -253 37 -219 71
rect -135 37 -101 71
rect -17 37 17 71
rect 101 37 135 71
rect 219 37 253 71
rect 337 37 371 71
rect 455 37 489 71
rect 573 37 607 71
rect 691 37 725 71
rect 809 37 843 71
rect 927 37 961 71
rect 1045 37 1079 71
rect 1163 37 1197 71
rect 1281 37 1315 71
rect 1399 37 1433 71
rect -1433 -71 -1399 -37
rect -1315 -71 -1281 -37
rect -1197 -71 -1163 -37
rect -1079 -71 -1045 -37
rect -961 -71 -927 -37
rect -843 -71 -809 -37
rect -725 -71 -691 -37
rect -607 -71 -573 -37
rect -489 -71 -455 -37
rect -371 -71 -337 -37
rect -253 -71 -219 -37
rect -135 -71 -101 -37
rect -17 -71 17 -37
rect 101 -71 135 -37
rect 219 -71 253 -37
rect 337 -71 371 -37
rect 455 -71 489 -37
rect 573 -71 607 -37
rect 691 -71 725 -37
rect 809 -71 843 -37
rect 927 -71 961 -37
rect 1045 -71 1079 -37
rect 1163 -71 1197 -37
rect 1281 -71 1315 -37
rect 1399 -71 1433 -37
rect -1492 -163 -1458 -149
rect -1492 -183 -1458 -163
rect -1492 -231 -1458 -221
rect -1492 -255 -1458 -231
rect -1492 -299 -1458 -293
rect -1492 -327 -1458 -299
rect -1492 -367 -1458 -365
rect -1492 -399 -1458 -367
rect -1492 -469 -1458 -437
rect -1492 -471 -1458 -469
rect -1492 -537 -1458 -509
rect -1492 -543 -1458 -537
rect -1492 -605 -1458 -581
rect -1492 -615 -1458 -605
rect -1492 -673 -1458 -653
rect -1492 -687 -1458 -673
rect -1374 -163 -1340 -149
rect -1374 -183 -1340 -163
rect -1374 -231 -1340 -221
rect -1374 -255 -1340 -231
rect -1374 -299 -1340 -293
rect -1374 -327 -1340 -299
rect -1374 -367 -1340 -365
rect -1374 -399 -1340 -367
rect -1374 -469 -1340 -437
rect -1374 -471 -1340 -469
rect -1374 -537 -1340 -509
rect -1374 -543 -1340 -537
rect -1374 -605 -1340 -581
rect -1374 -615 -1340 -605
rect -1374 -673 -1340 -653
rect -1374 -687 -1340 -673
rect -1256 -163 -1222 -149
rect -1256 -183 -1222 -163
rect -1256 -231 -1222 -221
rect -1256 -255 -1222 -231
rect -1256 -299 -1222 -293
rect -1256 -327 -1222 -299
rect -1256 -367 -1222 -365
rect -1256 -399 -1222 -367
rect -1256 -469 -1222 -437
rect -1256 -471 -1222 -469
rect -1256 -537 -1222 -509
rect -1256 -543 -1222 -537
rect -1256 -605 -1222 -581
rect -1256 -615 -1222 -605
rect -1256 -673 -1222 -653
rect -1256 -687 -1222 -673
rect -1138 -163 -1104 -149
rect -1138 -183 -1104 -163
rect -1138 -231 -1104 -221
rect -1138 -255 -1104 -231
rect -1138 -299 -1104 -293
rect -1138 -327 -1104 -299
rect -1138 -367 -1104 -365
rect -1138 -399 -1104 -367
rect -1138 -469 -1104 -437
rect -1138 -471 -1104 -469
rect -1138 -537 -1104 -509
rect -1138 -543 -1104 -537
rect -1138 -605 -1104 -581
rect -1138 -615 -1104 -605
rect -1138 -673 -1104 -653
rect -1138 -687 -1104 -673
rect -1020 -163 -986 -149
rect -1020 -183 -986 -163
rect -1020 -231 -986 -221
rect -1020 -255 -986 -231
rect -1020 -299 -986 -293
rect -1020 -327 -986 -299
rect -1020 -367 -986 -365
rect -1020 -399 -986 -367
rect -1020 -469 -986 -437
rect -1020 -471 -986 -469
rect -1020 -537 -986 -509
rect -1020 -543 -986 -537
rect -1020 -605 -986 -581
rect -1020 -615 -986 -605
rect -1020 -673 -986 -653
rect -1020 -687 -986 -673
rect -902 -163 -868 -149
rect -902 -183 -868 -163
rect -902 -231 -868 -221
rect -902 -255 -868 -231
rect -902 -299 -868 -293
rect -902 -327 -868 -299
rect -902 -367 -868 -365
rect -902 -399 -868 -367
rect -902 -469 -868 -437
rect -902 -471 -868 -469
rect -902 -537 -868 -509
rect -902 -543 -868 -537
rect -902 -605 -868 -581
rect -902 -615 -868 -605
rect -902 -673 -868 -653
rect -902 -687 -868 -673
rect -784 -163 -750 -149
rect -784 -183 -750 -163
rect -784 -231 -750 -221
rect -784 -255 -750 -231
rect -784 -299 -750 -293
rect -784 -327 -750 -299
rect -784 -367 -750 -365
rect -784 -399 -750 -367
rect -784 -469 -750 -437
rect -784 -471 -750 -469
rect -784 -537 -750 -509
rect -784 -543 -750 -537
rect -784 -605 -750 -581
rect -784 -615 -750 -605
rect -784 -673 -750 -653
rect -784 -687 -750 -673
rect -666 -163 -632 -149
rect -666 -183 -632 -163
rect -666 -231 -632 -221
rect -666 -255 -632 -231
rect -666 -299 -632 -293
rect -666 -327 -632 -299
rect -666 -367 -632 -365
rect -666 -399 -632 -367
rect -666 -469 -632 -437
rect -666 -471 -632 -469
rect -666 -537 -632 -509
rect -666 -543 -632 -537
rect -666 -605 -632 -581
rect -666 -615 -632 -605
rect -666 -673 -632 -653
rect -666 -687 -632 -673
rect -548 -163 -514 -149
rect -548 -183 -514 -163
rect -548 -231 -514 -221
rect -548 -255 -514 -231
rect -548 -299 -514 -293
rect -548 -327 -514 -299
rect -548 -367 -514 -365
rect -548 -399 -514 -367
rect -548 -469 -514 -437
rect -548 -471 -514 -469
rect -548 -537 -514 -509
rect -548 -543 -514 -537
rect -548 -605 -514 -581
rect -548 -615 -514 -605
rect -548 -673 -514 -653
rect -548 -687 -514 -673
rect -430 -163 -396 -149
rect -430 -183 -396 -163
rect -430 -231 -396 -221
rect -430 -255 -396 -231
rect -430 -299 -396 -293
rect -430 -327 -396 -299
rect -430 -367 -396 -365
rect -430 -399 -396 -367
rect -430 -469 -396 -437
rect -430 -471 -396 -469
rect -430 -537 -396 -509
rect -430 -543 -396 -537
rect -430 -605 -396 -581
rect -430 -615 -396 -605
rect -430 -673 -396 -653
rect -430 -687 -396 -673
rect -312 -163 -278 -149
rect -312 -183 -278 -163
rect -312 -231 -278 -221
rect -312 -255 -278 -231
rect -312 -299 -278 -293
rect -312 -327 -278 -299
rect -312 -367 -278 -365
rect -312 -399 -278 -367
rect -312 -469 -278 -437
rect -312 -471 -278 -469
rect -312 -537 -278 -509
rect -312 -543 -278 -537
rect -312 -605 -278 -581
rect -312 -615 -278 -605
rect -312 -673 -278 -653
rect -312 -687 -278 -673
rect -194 -163 -160 -149
rect -194 -183 -160 -163
rect -194 -231 -160 -221
rect -194 -255 -160 -231
rect -194 -299 -160 -293
rect -194 -327 -160 -299
rect -194 -367 -160 -365
rect -194 -399 -160 -367
rect -194 -469 -160 -437
rect -194 -471 -160 -469
rect -194 -537 -160 -509
rect -194 -543 -160 -537
rect -194 -605 -160 -581
rect -194 -615 -160 -605
rect -194 -673 -160 -653
rect -194 -687 -160 -673
rect -76 -163 -42 -149
rect -76 -183 -42 -163
rect -76 -231 -42 -221
rect -76 -255 -42 -231
rect -76 -299 -42 -293
rect -76 -327 -42 -299
rect -76 -367 -42 -365
rect -76 -399 -42 -367
rect -76 -469 -42 -437
rect -76 -471 -42 -469
rect -76 -537 -42 -509
rect -76 -543 -42 -537
rect -76 -605 -42 -581
rect -76 -615 -42 -605
rect -76 -673 -42 -653
rect -76 -687 -42 -673
rect 42 -163 76 -149
rect 42 -183 76 -163
rect 42 -231 76 -221
rect 42 -255 76 -231
rect 42 -299 76 -293
rect 42 -327 76 -299
rect 42 -367 76 -365
rect 42 -399 76 -367
rect 42 -469 76 -437
rect 42 -471 76 -469
rect 42 -537 76 -509
rect 42 -543 76 -537
rect 42 -605 76 -581
rect 42 -615 76 -605
rect 42 -673 76 -653
rect 42 -687 76 -673
rect 160 -163 194 -149
rect 160 -183 194 -163
rect 160 -231 194 -221
rect 160 -255 194 -231
rect 160 -299 194 -293
rect 160 -327 194 -299
rect 160 -367 194 -365
rect 160 -399 194 -367
rect 160 -469 194 -437
rect 160 -471 194 -469
rect 160 -537 194 -509
rect 160 -543 194 -537
rect 160 -605 194 -581
rect 160 -615 194 -605
rect 160 -673 194 -653
rect 160 -687 194 -673
rect 278 -163 312 -149
rect 278 -183 312 -163
rect 278 -231 312 -221
rect 278 -255 312 -231
rect 278 -299 312 -293
rect 278 -327 312 -299
rect 278 -367 312 -365
rect 278 -399 312 -367
rect 278 -469 312 -437
rect 278 -471 312 -469
rect 278 -537 312 -509
rect 278 -543 312 -537
rect 278 -605 312 -581
rect 278 -615 312 -605
rect 278 -673 312 -653
rect 278 -687 312 -673
rect 396 -163 430 -149
rect 396 -183 430 -163
rect 396 -231 430 -221
rect 396 -255 430 -231
rect 396 -299 430 -293
rect 396 -327 430 -299
rect 396 -367 430 -365
rect 396 -399 430 -367
rect 396 -469 430 -437
rect 396 -471 430 -469
rect 396 -537 430 -509
rect 396 -543 430 -537
rect 396 -605 430 -581
rect 396 -615 430 -605
rect 396 -673 430 -653
rect 396 -687 430 -673
rect 514 -163 548 -149
rect 514 -183 548 -163
rect 514 -231 548 -221
rect 514 -255 548 -231
rect 514 -299 548 -293
rect 514 -327 548 -299
rect 514 -367 548 -365
rect 514 -399 548 -367
rect 514 -469 548 -437
rect 514 -471 548 -469
rect 514 -537 548 -509
rect 514 -543 548 -537
rect 514 -605 548 -581
rect 514 -615 548 -605
rect 514 -673 548 -653
rect 514 -687 548 -673
rect 632 -163 666 -149
rect 632 -183 666 -163
rect 632 -231 666 -221
rect 632 -255 666 -231
rect 632 -299 666 -293
rect 632 -327 666 -299
rect 632 -367 666 -365
rect 632 -399 666 -367
rect 632 -469 666 -437
rect 632 -471 666 -469
rect 632 -537 666 -509
rect 632 -543 666 -537
rect 632 -605 666 -581
rect 632 -615 666 -605
rect 632 -673 666 -653
rect 632 -687 666 -673
rect 750 -163 784 -149
rect 750 -183 784 -163
rect 750 -231 784 -221
rect 750 -255 784 -231
rect 750 -299 784 -293
rect 750 -327 784 -299
rect 750 -367 784 -365
rect 750 -399 784 -367
rect 750 -469 784 -437
rect 750 -471 784 -469
rect 750 -537 784 -509
rect 750 -543 784 -537
rect 750 -605 784 -581
rect 750 -615 784 -605
rect 750 -673 784 -653
rect 750 -687 784 -673
rect 868 -163 902 -149
rect 868 -183 902 -163
rect 868 -231 902 -221
rect 868 -255 902 -231
rect 868 -299 902 -293
rect 868 -327 902 -299
rect 868 -367 902 -365
rect 868 -399 902 -367
rect 868 -469 902 -437
rect 868 -471 902 -469
rect 868 -537 902 -509
rect 868 -543 902 -537
rect 868 -605 902 -581
rect 868 -615 902 -605
rect 868 -673 902 -653
rect 868 -687 902 -673
rect 986 -163 1020 -149
rect 986 -183 1020 -163
rect 986 -231 1020 -221
rect 986 -255 1020 -231
rect 986 -299 1020 -293
rect 986 -327 1020 -299
rect 986 -367 1020 -365
rect 986 -399 1020 -367
rect 986 -469 1020 -437
rect 986 -471 1020 -469
rect 986 -537 1020 -509
rect 986 -543 1020 -537
rect 986 -605 1020 -581
rect 986 -615 1020 -605
rect 986 -673 1020 -653
rect 986 -687 1020 -673
rect 1104 -163 1138 -149
rect 1104 -183 1138 -163
rect 1104 -231 1138 -221
rect 1104 -255 1138 -231
rect 1104 -299 1138 -293
rect 1104 -327 1138 -299
rect 1104 -367 1138 -365
rect 1104 -399 1138 -367
rect 1104 -469 1138 -437
rect 1104 -471 1138 -469
rect 1104 -537 1138 -509
rect 1104 -543 1138 -537
rect 1104 -605 1138 -581
rect 1104 -615 1138 -605
rect 1104 -673 1138 -653
rect 1104 -687 1138 -673
rect 1222 -163 1256 -149
rect 1222 -183 1256 -163
rect 1222 -231 1256 -221
rect 1222 -255 1256 -231
rect 1222 -299 1256 -293
rect 1222 -327 1256 -299
rect 1222 -367 1256 -365
rect 1222 -399 1256 -367
rect 1222 -469 1256 -437
rect 1222 -471 1256 -469
rect 1222 -537 1256 -509
rect 1222 -543 1256 -537
rect 1222 -605 1256 -581
rect 1222 -615 1256 -605
rect 1222 -673 1256 -653
rect 1222 -687 1256 -673
rect 1340 -163 1374 -149
rect 1340 -183 1374 -163
rect 1340 -231 1374 -221
rect 1340 -255 1374 -231
rect 1340 -299 1374 -293
rect 1340 -327 1374 -299
rect 1340 -367 1374 -365
rect 1340 -399 1374 -367
rect 1340 -469 1374 -437
rect 1340 -471 1374 -469
rect 1340 -537 1374 -509
rect 1340 -543 1374 -537
rect 1340 -605 1374 -581
rect 1340 -615 1374 -605
rect 1340 -673 1374 -653
rect 1340 -687 1374 -673
rect 1458 -163 1492 -149
rect 1458 -183 1492 -163
rect 1458 -231 1492 -221
rect 1458 -255 1492 -231
rect 1458 -299 1492 -293
rect 1458 -327 1492 -299
rect 1458 -367 1492 -365
rect 1458 -399 1492 -367
rect 1458 -469 1492 -437
rect 1458 -471 1492 -469
rect 1458 -537 1492 -509
rect 1458 -543 1492 -537
rect 1458 -605 1492 -581
rect 1458 -615 1492 -605
rect 1458 -673 1492 -653
rect 1458 -687 1492 -673
<< metal1 >>
rect -1498 687 -1452 718
rect -1498 653 -1492 687
rect -1458 653 -1452 687
rect -1498 615 -1452 653
rect -1498 581 -1492 615
rect -1458 581 -1452 615
rect -1498 543 -1452 581
rect -1498 509 -1492 543
rect -1458 509 -1452 543
rect -1498 471 -1452 509
rect -1498 437 -1492 471
rect -1458 437 -1452 471
rect -1498 399 -1452 437
rect -1498 365 -1492 399
rect -1458 365 -1452 399
rect -1498 327 -1452 365
rect -1498 293 -1492 327
rect -1458 293 -1452 327
rect -1498 255 -1452 293
rect -1498 221 -1492 255
rect -1458 221 -1452 255
rect -1498 183 -1452 221
rect -1498 149 -1492 183
rect -1458 149 -1452 183
rect -1498 118 -1452 149
rect -1380 687 -1334 718
rect -1380 653 -1374 687
rect -1340 653 -1334 687
rect -1380 615 -1334 653
rect -1380 581 -1374 615
rect -1340 581 -1334 615
rect -1380 543 -1334 581
rect -1380 509 -1374 543
rect -1340 509 -1334 543
rect -1380 471 -1334 509
rect -1380 437 -1374 471
rect -1340 437 -1334 471
rect -1380 399 -1334 437
rect -1380 365 -1374 399
rect -1340 365 -1334 399
rect -1380 327 -1334 365
rect -1380 293 -1374 327
rect -1340 293 -1334 327
rect -1380 255 -1334 293
rect -1380 221 -1374 255
rect -1340 221 -1334 255
rect -1380 183 -1334 221
rect -1380 149 -1374 183
rect -1340 149 -1334 183
rect -1380 118 -1334 149
rect -1262 687 -1216 718
rect -1262 653 -1256 687
rect -1222 653 -1216 687
rect -1262 615 -1216 653
rect -1262 581 -1256 615
rect -1222 581 -1216 615
rect -1262 543 -1216 581
rect -1262 509 -1256 543
rect -1222 509 -1216 543
rect -1262 471 -1216 509
rect -1262 437 -1256 471
rect -1222 437 -1216 471
rect -1262 399 -1216 437
rect -1262 365 -1256 399
rect -1222 365 -1216 399
rect -1262 327 -1216 365
rect -1262 293 -1256 327
rect -1222 293 -1216 327
rect -1262 255 -1216 293
rect -1262 221 -1256 255
rect -1222 221 -1216 255
rect -1262 183 -1216 221
rect -1262 149 -1256 183
rect -1222 149 -1216 183
rect -1262 118 -1216 149
rect -1144 687 -1098 718
rect -1144 653 -1138 687
rect -1104 653 -1098 687
rect -1144 615 -1098 653
rect -1144 581 -1138 615
rect -1104 581 -1098 615
rect -1144 543 -1098 581
rect -1144 509 -1138 543
rect -1104 509 -1098 543
rect -1144 471 -1098 509
rect -1144 437 -1138 471
rect -1104 437 -1098 471
rect -1144 399 -1098 437
rect -1144 365 -1138 399
rect -1104 365 -1098 399
rect -1144 327 -1098 365
rect -1144 293 -1138 327
rect -1104 293 -1098 327
rect -1144 255 -1098 293
rect -1144 221 -1138 255
rect -1104 221 -1098 255
rect -1144 183 -1098 221
rect -1144 149 -1138 183
rect -1104 149 -1098 183
rect -1144 118 -1098 149
rect -1026 687 -980 718
rect -1026 653 -1020 687
rect -986 653 -980 687
rect -1026 615 -980 653
rect -1026 581 -1020 615
rect -986 581 -980 615
rect -1026 543 -980 581
rect -1026 509 -1020 543
rect -986 509 -980 543
rect -1026 471 -980 509
rect -1026 437 -1020 471
rect -986 437 -980 471
rect -1026 399 -980 437
rect -1026 365 -1020 399
rect -986 365 -980 399
rect -1026 327 -980 365
rect -1026 293 -1020 327
rect -986 293 -980 327
rect -1026 255 -980 293
rect -1026 221 -1020 255
rect -986 221 -980 255
rect -1026 183 -980 221
rect -1026 149 -1020 183
rect -986 149 -980 183
rect -1026 118 -980 149
rect -908 687 -862 718
rect -908 653 -902 687
rect -868 653 -862 687
rect -908 615 -862 653
rect -908 581 -902 615
rect -868 581 -862 615
rect -908 543 -862 581
rect -908 509 -902 543
rect -868 509 -862 543
rect -908 471 -862 509
rect -908 437 -902 471
rect -868 437 -862 471
rect -908 399 -862 437
rect -908 365 -902 399
rect -868 365 -862 399
rect -908 327 -862 365
rect -908 293 -902 327
rect -868 293 -862 327
rect -908 255 -862 293
rect -908 221 -902 255
rect -868 221 -862 255
rect -908 183 -862 221
rect -908 149 -902 183
rect -868 149 -862 183
rect -908 118 -862 149
rect -790 687 -744 718
rect -790 653 -784 687
rect -750 653 -744 687
rect -790 615 -744 653
rect -790 581 -784 615
rect -750 581 -744 615
rect -790 543 -744 581
rect -790 509 -784 543
rect -750 509 -744 543
rect -790 471 -744 509
rect -790 437 -784 471
rect -750 437 -744 471
rect -790 399 -744 437
rect -790 365 -784 399
rect -750 365 -744 399
rect -790 327 -744 365
rect -790 293 -784 327
rect -750 293 -744 327
rect -790 255 -744 293
rect -790 221 -784 255
rect -750 221 -744 255
rect -790 183 -744 221
rect -790 149 -784 183
rect -750 149 -744 183
rect -790 118 -744 149
rect -672 687 -626 718
rect -672 653 -666 687
rect -632 653 -626 687
rect -672 615 -626 653
rect -672 581 -666 615
rect -632 581 -626 615
rect -672 543 -626 581
rect -672 509 -666 543
rect -632 509 -626 543
rect -672 471 -626 509
rect -672 437 -666 471
rect -632 437 -626 471
rect -672 399 -626 437
rect -672 365 -666 399
rect -632 365 -626 399
rect -672 327 -626 365
rect -672 293 -666 327
rect -632 293 -626 327
rect -672 255 -626 293
rect -672 221 -666 255
rect -632 221 -626 255
rect -672 183 -626 221
rect -672 149 -666 183
rect -632 149 -626 183
rect -672 118 -626 149
rect -554 687 -508 718
rect -554 653 -548 687
rect -514 653 -508 687
rect -554 615 -508 653
rect -554 581 -548 615
rect -514 581 -508 615
rect -554 543 -508 581
rect -554 509 -548 543
rect -514 509 -508 543
rect -554 471 -508 509
rect -554 437 -548 471
rect -514 437 -508 471
rect -554 399 -508 437
rect -554 365 -548 399
rect -514 365 -508 399
rect -554 327 -508 365
rect -554 293 -548 327
rect -514 293 -508 327
rect -554 255 -508 293
rect -554 221 -548 255
rect -514 221 -508 255
rect -554 183 -508 221
rect -554 149 -548 183
rect -514 149 -508 183
rect -554 118 -508 149
rect -436 687 -390 718
rect -436 653 -430 687
rect -396 653 -390 687
rect -436 615 -390 653
rect -436 581 -430 615
rect -396 581 -390 615
rect -436 543 -390 581
rect -436 509 -430 543
rect -396 509 -390 543
rect -436 471 -390 509
rect -436 437 -430 471
rect -396 437 -390 471
rect -436 399 -390 437
rect -436 365 -430 399
rect -396 365 -390 399
rect -436 327 -390 365
rect -436 293 -430 327
rect -396 293 -390 327
rect -436 255 -390 293
rect -436 221 -430 255
rect -396 221 -390 255
rect -436 183 -390 221
rect -436 149 -430 183
rect -396 149 -390 183
rect -436 118 -390 149
rect -318 687 -272 718
rect -318 653 -312 687
rect -278 653 -272 687
rect -318 615 -272 653
rect -318 581 -312 615
rect -278 581 -272 615
rect -318 543 -272 581
rect -318 509 -312 543
rect -278 509 -272 543
rect -318 471 -272 509
rect -318 437 -312 471
rect -278 437 -272 471
rect -318 399 -272 437
rect -318 365 -312 399
rect -278 365 -272 399
rect -318 327 -272 365
rect -318 293 -312 327
rect -278 293 -272 327
rect -318 255 -272 293
rect -318 221 -312 255
rect -278 221 -272 255
rect -318 183 -272 221
rect -318 149 -312 183
rect -278 149 -272 183
rect -318 118 -272 149
rect -200 687 -154 718
rect -200 653 -194 687
rect -160 653 -154 687
rect -200 615 -154 653
rect -200 581 -194 615
rect -160 581 -154 615
rect -200 543 -154 581
rect -200 509 -194 543
rect -160 509 -154 543
rect -200 471 -154 509
rect -200 437 -194 471
rect -160 437 -154 471
rect -200 399 -154 437
rect -200 365 -194 399
rect -160 365 -154 399
rect -200 327 -154 365
rect -200 293 -194 327
rect -160 293 -154 327
rect -200 255 -154 293
rect -200 221 -194 255
rect -160 221 -154 255
rect -200 183 -154 221
rect -200 149 -194 183
rect -160 149 -154 183
rect -200 118 -154 149
rect -82 687 -36 718
rect -82 653 -76 687
rect -42 653 -36 687
rect -82 615 -36 653
rect -82 581 -76 615
rect -42 581 -36 615
rect -82 543 -36 581
rect -82 509 -76 543
rect -42 509 -36 543
rect -82 471 -36 509
rect -82 437 -76 471
rect -42 437 -36 471
rect -82 399 -36 437
rect -82 365 -76 399
rect -42 365 -36 399
rect -82 327 -36 365
rect -82 293 -76 327
rect -42 293 -36 327
rect -82 255 -36 293
rect -82 221 -76 255
rect -42 221 -36 255
rect -82 183 -36 221
rect -82 149 -76 183
rect -42 149 -36 183
rect -82 118 -36 149
rect 36 687 82 718
rect 36 653 42 687
rect 76 653 82 687
rect 36 615 82 653
rect 36 581 42 615
rect 76 581 82 615
rect 36 543 82 581
rect 36 509 42 543
rect 76 509 82 543
rect 36 471 82 509
rect 36 437 42 471
rect 76 437 82 471
rect 36 399 82 437
rect 36 365 42 399
rect 76 365 82 399
rect 36 327 82 365
rect 36 293 42 327
rect 76 293 82 327
rect 36 255 82 293
rect 36 221 42 255
rect 76 221 82 255
rect 36 183 82 221
rect 36 149 42 183
rect 76 149 82 183
rect 36 118 82 149
rect 154 687 200 718
rect 154 653 160 687
rect 194 653 200 687
rect 154 615 200 653
rect 154 581 160 615
rect 194 581 200 615
rect 154 543 200 581
rect 154 509 160 543
rect 194 509 200 543
rect 154 471 200 509
rect 154 437 160 471
rect 194 437 200 471
rect 154 399 200 437
rect 154 365 160 399
rect 194 365 200 399
rect 154 327 200 365
rect 154 293 160 327
rect 194 293 200 327
rect 154 255 200 293
rect 154 221 160 255
rect 194 221 200 255
rect 154 183 200 221
rect 154 149 160 183
rect 194 149 200 183
rect 154 118 200 149
rect 272 687 318 718
rect 272 653 278 687
rect 312 653 318 687
rect 272 615 318 653
rect 272 581 278 615
rect 312 581 318 615
rect 272 543 318 581
rect 272 509 278 543
rect 312 509 318 543
rect 272 471 318 509
rect 272 437 278 471
rect 312 437 318 471
rect 272 399 318 437
rect 272 365 278 399
rect 312 365 318 399
rect 272 327 318 365
rect 272 293 278 327
rect 312 293 318 327
rect 272 255 318 293
rect 272 221 278 255
rect 312 221 318 255
rect 272 183 318 221
rect 272 149 278 183
rect 312 149 318 183
rect 272 118 318 149
rect 390 687 436 718
rect 390 653 396 687
rect 430 653 436 687
rect 390 615 436 653
rect 390 581 396 615
rect 430 581 436 615
rect 390 543 436 581
rect 390 509 396 543
rect 430 509 436 543
rect 390 471 436 509
rect 390 437 396 471
rect 430 437 436 471
rect 390 399 436 437
rect 390 365 396 399
rect 430 365 436 399
rect 390 327 436 365
rect 390 293 396 327
rect 430 293 436 327
rect 390 255 436 293
rect 390 221 396 255
rect 430 221 436 255
rect 390 183 436 221
rect 390 149 396 183
rect 430 149 436 183
rect 390 118 436 149
rect 508 687 554 718
rect 508 653 514 687
rect 548 653 554 687
rect 508 615 554 653
rect 508 581 514 615
rect 548 581 554 615
rect 508 543 554 581
rect 508 509 514 543
rect 548 509 554 543
rect 508 471 554 509
rect 508 437 514 471
rect 548 437 554 471
rect 508 399 554 437
rect 508 365 514 399
rect 548 365 554 399
rect 508 327 554 365
rect 508 293 514 327
rect 548 293 554 327
rect 508 255 554 293
rect 508 221 514 255
rect 548 221 554 255
rect 508 183 554 221
rect 508 149 514 183
rect 548 149 554 183
rect 508 118 554 149
rect 626 687 672 718
rect 626 653 632 687
rect 666 653 672 687
rect 626 615 672 653
rect 626 581 632 615
rect 666 581 672 615
rect 626 543 672 581
rect 626 509 632 543
rect 666 509 672 543
rect 626 471 672 509
rect 626 437 632 471
rect 666 437 672 471
rect 626 399 672 437
rect 626 365 632 399
rect 666 365 672 399
rect 626 327 672 365
rect 626 293 632 327
rect 666 293 672 327
rect 626 255 672 293
rect 626 221 632 255
rect 666 221 672 255
rect 626 183 672 221
rect 626 149 632 183
rect 666 149 672 183
rect 626 118 672 149
rect 744 687 790 718
rect 744 653 750 687
rect 784 653 790 687
rect 744 615 790 653
rect 744 581 750 615
rect 784 581 790 615
rect 744 543 790 581
rect 744 509 750 543
rect 784 509 790 543
rect 744 471 790 509
rect 744 437 750 471
rect 784 437 790 471
rect 744 399 790 437
rect 744 365 750 399
rect 784 365 790 399
rect 744 327 790 365
rect 744 293 750 327
rect 784 293 790 327
rect 744 255 790 293
rect 744 221 750 255
rect 784 221 790 255
rect 744 183 790 221
rect 744 149 750 183
rect 784 149 790 183
rect 744 118 790 149
rect 862 687 908 718
rect 862 653 868 687
rect 902 653 908 687
rect 862 615 908 653
rect 862 581 868 615
rect 902 581 908 615
rect 862 543 908 581
rect 862 509 868 543
rect 902 509 908 543
rect 862 471 908 509
rect 862 437 868 471
rect 902 437 908 471
rect 862 399 908 437
rect 862 365 868 399
rect 902 365 908 399
rect 862 327 908 365
rect 862 293 868 327
rect 902 293 908 327
rect 862 255 908 293
rect 862 221 868 255
rect 902 221 908 255
rect 862 183 908 221
rect 862 149 868 183
rect 902 149 908 183
rect 862 118 908 149
rect 980 687 1026 718
rect 980 653 986 687
rect 1020 653 1026 687
rect 980 615 1026 653
rect 980 581 986 615
rect 1020 581 1026 615
rect 980 543 1026 581
rect 980 509 986 543
rect 1020 509 1026 543
rect 980 471 1026 509
rect 980 437 986 471
rect 1020 437 1026 471
rect 980 399 1026 437
rect 980 365 986 399
rect 1020 365 1026 399
rect 980 327 1026 365
rect 980 293 986 327
rect 1020 293 1026 327
rect 980 255 1026 293
rect 980 221 986 255
rect 1020 221 1026 255
rect 980 183 1026 221
rect 980 149 986 183
rect 1020 149 1026 183
rect 980 118 1026 149
rect 1098 687 1144 718
rect 1098 653 1104 687
rect 1138 653 1144 687
rect 1098 615 1144 653
rect 1098 581 1104 615
rect 1138 581 1144 615
rect 1098 543 1144 581
rect 1098 509 1104 543
rect 1138 509 1144 543
rect 1098 471 1144 509
rect 1098 437 1104 471
rect 1138 437 1144 471
rect 1098 399 1144 437
rect 1098 365 1104 399
rect 1138 365 1144 399
rect 1098 327 1144 365
rect 1098 293 1104 327
rect 1138 293 1144 327
rect 1098 255 1144 293
rect 1098 221 1104 255
rect 1138 221 1144 255
rect 1098 183 1144 221
rect 1098 149 1104 183
rect 1138 149 1144 183
rect 1098 118 1144 149
rect 1216 687 1262 718
rect 1216 653 1222 687
rect 1256 653 1262 687
rect 1216 615 1262 653
rect 1216 581 1222 615
rect 1256 581 1262 615
rect 1216 543 1262 581
rect 1216 509 1222 543
rect 1256 509 1262 543
rect 1216 471 1262 509
rect 1216 437 1222 471
rect 1256 437 1262 471
rect 1216 399 1262 437
rect 1216 365 1222 399
rect 1256 365 1262 399
rect 1216 327 1262 365
rect 1216 293 1222 327
rect 1256 293 1262 327
rect 1216 255 1262 293
rect 1216 221 1222 255
rect 1256 221 1262 255
rect 1216 183 1262 221
rect 1216 149 1222 183
rect 1256 149 1262 183
rect 1216 118 1262 149
rect 1334 687 1380 718
rect 1334 653 1340 687
rect 1374 653 1380 687
rect 1334 615 1380 653
rect 1334 581 1340 615
rect 1374 581 1380 615
rect 1334 543 1380 581
rect 1334 509 1340 543
rect 1374 509 1380 543
rect 1334 471 1380 509
rect 1334 437 1340 471
rect 1374 437 1380 471
rect 1334 399 1380 437
rect 1334 365 1340 399
rect 1374 365 1380 399
rect 1334 327 1380 365
rect 1334 293 1340 327
rect 1374 293 1380 327
rect 1334 255 1380 293
rect 1334 221 1340 255
rect 1374 221 1380 255
rect 1334 183 1380 221
rect 1334 149 1340 183
rect 1374 149 1380 183
rect 1334 118 1380 149
rect 1452 687 1498 718
rect 1452 653 1458 687
rect 1492 653 1498 687
rect 1452 615 1498 653
rect 1452 581 1458 615
rect 1492 581 1498 615
rect 1452 543 1498 581
rect 1452 509 1458 543
rect 1492 509 1498 543
rect 1452 471 1498 509
rect 1452 437 1458 471
rect 1492 437 1498 471
rect 1452 399 1498 437
rect 1452 365 1458 399
rect 1492 365 1498 399
rect 1452 327 1498 365
rect 1452 293 1458 327
rect 1492 293 1498 327
rect 1452 255 1498 293
rect 1452 221 1458 255
rect 1492 221 1498 255
rect 1452 183 1498 221
rect 1452 149 1458 183
rect 1492 149 1498 183
rect 1452 118 1498 149
rect -1445 71 -1387 77
rect -1445 37 -1433 71
rect -1399 37 -1387 71
rect -1445 31 -1387 37
rect -1327 71 -1269 77
rect -1327 37 -1315 71
rect -1281 37 -1269 71
rect -1327 31 -1269 37
rect -1209 71 -1151 77
rect -1209 37 -1197 71
rect -1163 37 -1151 71
rect -1209 31 -1151 37
rect -1091 71 -1033 77
rect -1091 37 -1079 71
rect -1045 37 -1033 71
rect -1091 31 -1033 37
rect -973 71 -915 77
rect -973 37 -961 71
rect -927 37 -915 71
rect -973 31 -915 37
rect -855 71 -797 77
rect -855 37 -843 71
rect -809 37 -797 71
rect -855 31 -797 37
rect -737 71 -679 77
rect -737 37 -725 71
rect -691 37 -679 71
rect -737 31 -679 37
rect -619 71 -561 77
rect -619 37 -607 71
rect -573 37 -561 71
rect -619 31 -561 37
rect -501 71 -443 77
rect -501 37 -489 71
rect -455 37 -443 71
rect -501 31 -443 37
rect -383 71 -325 77
rect -383 37 -371 71
rect -337 37 -325 71
rect -383 31 -325 37
rect -265 71 -207 77
rect -265 37 -253 71
rect -219 37 -207 71
rect -265 31 -207 37
rect -147 71 -89 77
rect -147 37 -135 71
rect -101 37 -89 71
rect -147 31 -89 37
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect 89 71 147 77
rect 89 37 101 71
rect 135 37 147 71
rect 89 31 147 37
rect 207 71 265 77
rect 207 37 219 71
rect 253 37 265 71
rect 207 31 265 37
rect 325 71 383 77
rect 325 37 337 71
rect 371 37 383 71
rect 325 31 383 37
rect 443 71 501 77
rect 443 37 455 71
rect 489 37 501 71
rect 443 31 501 37
rect 561 71 619 77
rect 561 37 573 71
rect 607 37 619 71
rect 561 31 619 37
rect 679 71 737 77
rect 679 37 691 71
rect 725 37 737 71
rect 679 31 737 37
rect 797 71 855 77
rect 797 37 809 71
rect 843 37 855 71
rect 797 31 855 37
rect 915 71 973 77
rect 915 37 927 71
rect 961 37 973 71
rect 915 31 973 37
rect 1033 71 1091 77
rect 1033 37 1045 71
rect 1079 37 1091 71
rect 1033 31 1091 37
rect 1151 71 1209 77
rect 1151 37 1163 71
rect 1197 37 1209 71
rect 1151 31 1209 37
rect 1269 71 1327 77
rect 1269 37 1281 71
rect 1315 37 1327 71
rect 1269 31 1327 37
rect 1387 71 1445 77
rect 1387 37 1399 71
rect 1433 37 1445 71
rect 1387 31 1445 37
rect -1445 -37 -1387 -31
rect -1445 -71 -1433 -37
rect -1399 -71 -1387 -37
rect -1445 -77 -1387 -71
rect -1327 -37 -1269 -31
rect -1327 -71 -1315 -37
rect -1281 -71 -1269 -37
rect -1327 -77 -1269 -71
rect -1209 -37 -1151 -31
rect -1209 -71 -1197 -37
rect -1163 -71 -1151 -37
rect -1209 -77 -1151 -71
rect -1091 -37 -1033 -31
rect -1091 -71 -1079 -37
rect -1045 -71 -1033 -37
rect -1091 -77 -1033 -71
rect -973 -37 -915 -31
rect -973 -71 -961 -37
rect -927 -71 -915 -37
rect -973 -77 -915 -71
rect -855 -37 -797 -31
rect -855 -71 -843 -37
rect -809 -71 -797 -37
rect -855 -77 -797 -71
rect -737 -37 -679 -31
rect -737 -71 -725 -37
rect -691 -71 -679 -37
rect -737 -77 -679 -71
rect -619 -37 -561 -31
rect -619 -71 -607 -37
rect -573 -71 -561 -37
rect -619 -77 -561 -71
rect -501 -37 -443 -31
rect -501 -71 -489 -37
rect -455 -71 -443 -37
rect -501 -77 -443 -71
rect -383 -37 -325 -31
rect -383 -71 -371 -37
rect -337 -71 -325 -37
rect -383 -77 -325 -71
rect -265 -37 -207 -31
rect -265 -71 -253 -37
rect -219 -71 -207 -37
rect -265 -77 -207 -71
rect -147 -37 -89 -31
rect -147 -71 -135 -37
rect -101 -71 -89 -37
rect -147 -77 -89 -71
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect 89 -37 147 -31
rect 89 -71 101 -37
rect 135 -71 147 -37
rect 89 -77 147 -71
rect 207 -37 265 -31
rect 207 -71 219 -37
rect 253 -71 265 -37
rect 207 -77 265 -71
rect 325 -37 383 -31
rect 325 -71 337 -37
rect 371 -71 383 -37
rect 325 -77 383 -71
rect 443 -37 501 -31
rect 443 -71 455 -37
rect 489 -71 501 -37
rect 443 -77 501 -71
rect 561 -37 619 -31
rect 561 -71 573 -37
rect 607 -71 619 -37
rect 561 -77 619 -71
rect 679 -37 737 -31
rect 679 -71 691 -37
rect 725 -71 737 -37
rect 679 -77 737 -71
rect 797 -37 855 -31
rect 797 -71 809 -37
rect 843 -71 855 -37
rect 797 -77 855 -71
rect 915 -37 973 -31
rect 915 -71 927 -37
rect 961 -71 973 -37
rect 915 -77 973 -71
rect 1033 -37 1091 -31
rect 1033 -71 1045 -37
rect 1079 -71 1091 -37
rect 1033 -77 1091 -71
rect 1151 -37 1209 -31
rect 1151 -71 1163 -37
rect 1197 -71 1209 -37
rect 1151 -77 1209 -71
rect 1269 -37 1327 -31
rect 1269 -71 1281 -37
rect 1315 -71 1327 -37
rect 1269 -77 1327 -71
rect 1387 -37 1445 -31
rect 1387 -71 1399 -37
rect 1433 -71 1445 -37
rect 1387 -77 1445 -71
rect -1498 -149 -1452 -118
rect -1498 -183 -1492 -149
rect -1458 -183 -1452 -149
rect -1498 -221 -1452 -183
rect -1498 -255 -1492 -221
rect -1458 -255 -1452 -221
rect -1498 -293 -1452 -255
rect -1498 -327 -1492 -293
rect -1458 -327 -1452 -293
rect -1498 -365 -1452 -327
rect -1498 -399 -1492 -365
rect -1458 -399 -1452 -365
rect -1498 -437 -1452 -399
rect -1498 -471 -1492 -437
rect -1458 -471 -1452 -437
rect -1498 -509 -1452 -471
rect -1498 -543 -1492 -509
rect -1458 -543 -1452 -509
rect -1498 -581 -1452 -543
rect -1498 -615 -1492 -581
rect -1458 -615 -1452 -581
rect -1498 -653 -1452 -615
rect -1498 -687 -1492 -653
rect -1458 -687 -1452 -653
rect -1498 -718 -1452 -687
rect -1380 -149 -1334 -118
rect -1380 -183 -1374 -149
rect -1340 -183 -1334 -149
rect -1380 -221 -1334 -183
rect -1380 -255 -1374 -221
rect -1340 -255 -1334 -221
rect -1380 -293 -1334 -255
rect -1380 -327 -1374 -293
rect -1340 -327 -1334 -293
rect -1380 -365 -1334 -327
rect -1380 -399 -1374 -365
rect -1340 -399 -1334 -365
rect -1380 -437 -1334 -399
rect -1380 -471 -1374 -437
rect -1340 -471 -1334 -437
rect -1380 -509 -1334 -471
rect -1380 -543 -1374 -509
rect -1340 -543 -1334 -509
rect -1380 -581 -1334 -543
rect -1380 -615 -1374 -581
rect -1340 -615 -1334 -581
rect -1380 -653 -1334 -615
rect -1380 -687 -1374 -653
rect -1340 -687 -1334 -653
rect -1380 -718 -1334 -687
rect -1262 -149 -1216 -118
rect -1262 -183 -1256 -149
rect -1222 -183 -1216 -149
rect -1262 -221 -1216 -183
rect -1262 -255 -1256 -221
rect -1222 -255 -1216 -221
rect -1262 -293 -1216 -255
rect -1262 -327 -1256 -293
rect -1222 -327 -1216 -293
rect -1262 -365 -1216 -327
rect -1262 -399 -1256 -365
rect -1222 -399 -1216 -365
rect -1262 -437 -1216 -399
rect -1262 -471 -1256 -437
rect -1222 -471 -1216 -437
rect -1262 -509 -1216 -471
rect -1262 -543 -1256 -509
rect -1222 -543 -1216 -509
rect -1262 -581 -1216 -543
rect -1262 -615 -1256 -581
rect -1222 -615 -1216 -581
rect -1262 -653 -1216 -615
rect -1262 -687 -1256 -653
rect -1222 -687 -1216 -653
rect -1262 -718 -1216 -687
rect -1144 -149 -1098 -118
rect -1144 -183 -1138 -149
rect -1104 -183 -1098 -149
rect -1144 -221 -1098 -183
rect -1144 -255 -1138 -221
rect -1104 -255 -1098 -221
rect -1144 -293 -1098 -255
rect -1144 -327 -1138 -293
rect -1104 -327 -1098 -293
rect -1144 -365 -1098 -327
rect -1144 -399 -1138 -365
rect -1104 -399 -1098 -365
rect -1144 -437 -1098 -399
rect -1144 -471 -1138 -437
rect -1104 -471 -1098 -437
rect -1144 -509 -1098 -471
rect -1144 -543 -1138 -509
rect -1104 -543 -1098 -509
rect -1144 -581 -1098 -543
rect -1144 -615 -1138 -581
rect -1104 -615 -1098 -581
rect -1144 -653 -1098 -615
rect -1144 -687 -1138 -653
rect -1104 -687 -1098 -653
rect -1144 -718 -1098 -687
rect -1026 -149 -980 -118
rect -1026 -183 -1020 -149
rect -986 -183 -980 -149
rect -1026 -221 -980 -183
rect -1026 -255 -1020 -221
rect -986 -255 -980 -221
rect -1026 -293 -980 -255
rect -1026 -327 -1020 -293
rect -986 -327 -980 -293
rect -1026 -365 -980 -327
rect -1026 -399 -1020 -365
rect -986 -399 -980 -365
rect -1026 -437 -980 -399
rect -1026 -471 -1020 -437
rect -986 -471 -980 -437
rect -1026 -509 -980 -471
rect -1026 -543 -1020 -509
rect -986 -543 -980 -509
rect -1026 -581 -980 -543
rect -1026 -615 -1020 -581
rect -986 -615 -980 -581
rect -1026 -653 -980 -615
rect -1026 -687 -1020 -653
rect -986 -687 -980 -653
rect -1026 -718 -980 -687
rect -908 -149 -862 -118
rect -908 -183 -902 -149
rect -868 -183 -862 -149
rect -908 -221 -862 -183
rect -908 -255 -902 -221
rect -868 -255 -862 -221
rect -908 -293 -862 -255
rect -908 -327 -902 -293
rect -868 -327 -862 -293
rect -908 -365 -862 -327
rect -908 -399 -902 -365
rect -868 -399 -862 -365
rect -908 -437 -862 -399
rect -908 -471 -902 -437
rect -868 -471 -862 -437
rect -908 -509 -862 -471
rect -908 -543 -902 -509
rect -868 -543 -862 -509
rect -908 -581 -862 -543
rect -908 -615 -902 -581
rect -868 -615 -862 -581
rect -908 -653 -862 -615
rect -908 -687 -902 -653
rect -868 -687 -862 -653
rect -908 -718 -862 -687
rect -790 -149 -744 -118
rect -790 -183 -784 -149
rect -750 -183 -744 -149
rect -790 -221 -744 -183
rect -790 -255 -784 -221
rect -750 -255 -744 -221
rect -790 -293 -744 -255
rect -790 -327 -784 -293
rect -750 -327 -744 -293
rect -790 -365 -744 -327
rect -790 -399 -784 -365
rect -750 -399 -744 -365
rect -790 -437 -744 -399
rect -790 -471 -784 -437
rect -750 -471 -744 -437
rect -790 -509 -744 -471
rect -790 -543 -784 -509
rect -750 -543 -744 -509
rect -790 -581 -744 -543
rect -790 -615 -784 -581
rect -750 -615 -744 -581
rect -790 -653 -744 -615
rect -790 -687 -784 -653
rect -750 -687 -744 -653
rect -790 -718 -744 -687
rect -672 -149 -626 -118
rect -672 -183 -666 -149
rect -632 -183 -626 -149
rect -672 -221 -626 -183
rect -672 -255 -666 -221
rect -632 -255 -626 -221
rect -672 -293 -626 -255
rect -672 -327 -666 -293
rect -632 -327 -626 -293
rect -672 -365 -626 -327
rect -672 -399 -666 -365
rect -632 -399 -626 -365
rect -672 -437 -626 -399
rect -672 -471 -666 -437
rect -632 -471 -626 -437
rect -672 -509 -626 -471
rect -672 -543 -666 -509
rect -632 -543 -626 -509
rect -672 -581 -626 -543
rect -672 -615 -666 -581
rect -632 -615 -626 -581
rect -672 -653 -626 -615
rect -672 -687 -666 -653
rect -632 -687 -626 -653
rect -672 -718 -626 -687
rect -554 -149 -508 -118
rect -554 -183 -548 -149
rect -514 -183 -508 -149
rect -554 -221 -508 -183
rect -554 -255 -548 -221
rect -514 -255 -508 -221
rect -554 -293 -508 -255
rect -554 -327 -548 -293
rect -514 -327 -508 -293
rect -554 -365 -508 -327
rect -554 -399 -548 -365
rect -514 -399 -508 -365
rect -554 -437 -508 -399
rect -554 -471 -548 -437
rect -514 -471 -508 -437
rect -554 -509 -508 -471
rect -554 -543 -548 -509
rect -514 -543 -508 -509
rect -554 -581 -508 -543
rect -554 -615 -548 -581
rect -514 -615 -508 -581
rect -554 -653 -508 -615
rect -554 -687 -548 -653
rect -514 -687 -508 -653
rect -554 -718 -508 -687
rect -436 -149 -390 -118
rect -436 -183 -430 -149
rect -396 -183 -390 -149
rect -436 -221 -390 -183
rect -436 -255 -430 -221
rect -396 -255 -390 -221
rect -436 -293 -390 -255
rect -436 -327 -430 -293
rect -396 -327 -390 -293
rect -436 -365 -390 -327
rect -436 -399 -430 -365
rect -396 -399 -390 -365
rect -436 -437 -390 -399
rect -436 -471 -430 -437
rect -396 -471 -390 -437
rect -436 -509 -390 -471
rect -436 -543 -430 -509
rect -396 -543 -390 -509
rect -436 -581 -390 -543
rect -436 -615 -430 -581
rect -396 -615 -390 -581
rect -436 -653 -390 -615
rect -436 -687 -430 -653
rect -396 -687 -390 -653
rect -436 -718 -390 -687
rect -318 -149 -272 -118
rect -318 -183 -312 -149
rect -278 -183 -272 -149
rect -318 -221 -272 -183
rect -318 -255 -312 -221
rect -278 -255 -272 -221
rect -318 -293 -272 -255
rect -318 -327 -312 -293
rect -278 -327 -272 -293
rect -318 -365 -272 -327
rect -318 -399 -312 -365
rect -278 -399 -272 -365
rect -318 -437 -272 -399
rect -318 -471 -312 -437
rect -278 -471 -272 -437
rect -318 -509 -272 -471
rect -318 -543 -312 -509
rect -278 -543 -272 -509
rect -318 -581 -272 -543
rect -318 -615 -312 -581
rect -278 -615 -272 -581
rect -318 -653 -272 -615
rect -318 -687 -312 -653
rect -278 -687 -272 -653
rect -318 -718 -272 -687
rect -200 -149 -154 -118
rect -200 -183 -194 -149
rect -160 -183 -154 -149
rect -200 -221 -154 -183
rect -200 -255 -194 -221
rect -160 -255 -154 -221
rect -200 -293 -154 -255
rect -200 -327 -194 -293
rect -160 -327 -154 -293
rect -200 -365 -154 -327
rect -200 -399 -194 -365
rect -160 -399 -154 -365
rect -200 -437 -154 -399
rect -200 -471 -194 -437
rect -160 -471 -154 -437
rect -200 -509 -154 -471
rect -200 -543 -194 -509
rect -160 -543 -154 -509
rect -200 -581 -154 -543
rect -200 -615 -194 -581
rect -160 -615 -154 -581
rect -200 -653 -154 -615
rect -200 -687 -194 -653
rect -160 -687 -154 -653
rect -200 -718 -154 -687
rect -82 -149 -36 -118
rect -82 -183 -76 -149
rect -42 -183 -36 -149
rect -82 -221 -36 -183
rect -82 -255 -76 -221
rect -42 -255 -36 -221
rect -82 -293 -36 -255
rect -82 -327 -76 -293
rect -42 -327 -36 -293
rect -82 -365 -36 -327
rect -82 -399 -76 -365
rect -42 -399 -36 -365
rect -82 -437 -36 -399
rect -82 -471 -76 -437
rect -42 -471 -36 -437
rect -82 -509 -36 -471
rect -82 -543 -76 -509
rect -42 -543 -36 -509
rect -82 -581 -36 -543
rect -82 -615 -76 -581
rect -42 -615 -36 -581
rect -82 -653 -36 -615
rect -82 -687 -76 -653
rect -42 -687 -36 -653
rect -82 -718 -36 -687
rect 36 -149 82 -118
rect 36 -183 42 -149
rect 76 -183 82 -149
rect 36 -221 82 -183
rect 36 -255 42 -221
rect 76 -255 82 -221
rect 36 -293 82 -255
rect 36 -327 42 -293
rect 76 -327 82 -293
rect 36 -365 82 -327
rect 36 -399 42 -365
rect 76 -399 82 -365
rect 36 -437 82 -399
rect 36 -471 42 -437
rect 76 -471 82 -437
rect 36 -509 82 -471
rect 36 -543 42 -509
rect 76 -543 82 -509
rect 36 -581 82 -543
rect 36 -615 42 -581
rect 76 -615 82 -581
rect 36 -653 82 -615
rect 36 -687 42 -653
rect 76 -687 82 -653
rect 36 -718 82 -687
rect 154 -149 200 -118
rect 154 -183 160 -149
rect 194 -183 200 -149
rect 154 -221 200 -183
rect 154 -255 160 -221
rect 194 -255 200 -221
rect 154 -293 200 -255
rect 154 -327 160 -293
rect 194 -327 200 -293
rect 154 -365 200 -327
rect 154 -399 160 -365
rect 194 -399 200 -365
rect 154 -437 200 -399
rect 154 -471 160 -437
rect 194 -471 200 -437
rect 154 -509 200 -471
rect 154 -543 160 -509
rect 194 -543 200 -509
rect 154 -581 200 -543
rect 154 -615 160 -581
rect 194 -615 200 -581
rect 154 -653 200 -615
rect 154 -687 160 -653
rect 194 -687 200 -653
rect 154 -718 200 -687
rect 272 -149 318 -118
rect 272 -183 278 -149
rect 312 -183 318 -149
rect 272 -221 318 -183
rect 272 -255 278 -221
rect 312 -255 318 -221
rect 272 -293 318 -255
rect 272 -327 278 -293
rect 312 -327 318 -293
rect 272 -365 318 -327
rect 272 -399 278 -365
rect 312 -399 318 -365
rect 272 -437 318 -399
rect 272 -471 278 -437
rect 312 -471 318 -437
rect 272 -509 318 -471
rect 272 -543 278 -509
rect 312 -543 318 -509
rect 272 -581 318 -543
rect 272 -615 278 -581
rect 312 -615 318 -581
rect 272 -653 318 -615
rect 272 -687 278 -653
rect 312 -687 318 -653
rect 272 -718 318 -687
rect 390 -149 436 -118
rect 390 -183 396 -149
rect 430 -183 436 -149
rect 390 -221 436 -183
rect 390 -255 396 -221
rect 430 -255 436 -221
rect 390 -293 436 -255
rect 390 -327 396 -293
rect 430 -327 436 -293
rect 390 -365 436 -327
rect 390 -399 396 -365
rect 430 -399 436 -365
rect 390 -437 436 -399
rect 390 -471 396 -437
rect 430 -471 436 -437
rect 390 -509 436 -471
rect 390 -543 396 -509
rect 430 -543 436 -509
rect 390 -581 436 -543
rect 390 -615 396 -581
rect 430 -615 436 -581
rect 390 -653 436 -615
rect 390 -687 396 -653
rect 430 -687 436 -653
rect 390 -718 436 -687
rect 508 -149 554 -118
rect 508 -183 514 -149
rect 548 -183 554 -149
rect 508 -221 554 -183
rect 508 -255 514 -221
rect 548 -255 554 -221
rect 508 -293 554 -255
rect 508 -327 514 -293
rect 548 -327 554 -293
rect 508 -365 554 -327
rect 508 -399 514 -365
rect 548 -399 554 -365
rect 508 -437 554 -399
rect 508 -471 514 -437
rect 548 -471 554 -437
rect 508 -509 554 -471
rect 508 -543 514 -509
rect 548 -543 554 -509
rect 508 -581 554 -543
rect 508 -615 514 -581
rect 548 -615 554 -581
rect 508 -653 554 -615
rect 508 -687 514 -653
rect 548 -687 554 -653
rect 508 -718 554 -687
rect 626 -149 672 -118
rect 626 -183 632 -149
rect 666 -183 672 -149
rect 626 -221 672 -183
rect 626 -255 632 -221
rect 666 -255 672 -221
rect 626 -293 672 -255
rect 626 -327 632 -293
rect 666 -327 672 -293
rect 626 -365 672 -327
rect 626 -399 632 -365
rect 666 -399 672 -365
rect 626 -437 672 -399
rect 626 -471 632 -437
rect 666 -471 672 -437
rect 626 -509 672 -471
rect 626 -543 632 -509
rect 666 -543 672 -509
rect 626 -581 672 -543
rect 626 -615 632 -581
rect 666 -615 672 -581
rect 626 -653 672 -615
rect 626 -687 632 -653
rect 666 -687 672 -653
rect 626 -718 672 -687
rect 744 -149 790 -118
rect 744 -183 750 -149
rect 784 -183 790 -149
rect 744 -221 790 -183
rect 744 -255 750 -221
rect 784 -255 790 -221
rect 744 -293 790 -255
rect 744 -327 750 -293
rect 784 -327 790 -293
rect 744 -365 790 -327
rect 744 -399 750 -365
rect 784 -399 790 -365
rect 744 -437 790 -399
rect 744 -471 750 -437
rect 784 -471 790 -437
rect 744 -509 790 -471
rect 744 -543 750 -509
rect 784 -543 790 -509
rect 744 -581 790 -543
rect 744 -615 750 -581
rect 784 -615 790 -581
rect 744 -653 790 -615
rect 744 -687 750 -653
rect 784 -687 790 -653
rect 744 -718 790 -687
rect 862 -149 908 -118
rect 862 -183 868 -149
rect 902 -183 908 -149
rect 862 -221 908 -183
rect 862 -255 868 -221
rect 902 -255 908 -221
rect 862 -293 908 -255
rect 862 -327 868 -293
rect 902 -327 908 -293
rect 862 -365 908 -327
rect 862 -399 868 -365
rect 902 -399 908 -365
rect 862 -437 908 -399
rect 862 -471 868 -437
rect 902 -471 908 -437
rect 862 -509 908 -471
rect 862 -543 868 -509
rect 902 -543 908 -509
rect 862 -581 908 -543
rect 862 -615 868 -581
rect 902 -615 908 -581
rect 862 -653 908 -615
rect 862 -687 868 -653
rect 902 -687 908 -653
rect 862 -718 908 -687
rect 980 -149 1026 -118
rect 980 -183 986 -149
rect 1020 -183 1026 -149
rect 980 -221 1026 -183
rect 980 -255 986 -221
rect 1020 -255 1026 -221
rect 980 -293 1026 -255
rect 980 -327 986 -293
rect 1020 -327 1026 -293
rect 980 -365 1026 -327
rect 980 -399 986 -365
rect 1020 -399 1026 -365
rect 980 -437 1026 -399
rect 980 -471 986 -437
rect 1020 -471 1026 -437
rect 980 -509 1026 -471
rect 980 -543 986 -509
rect 1020 -543 1026 -509
rect 980 -581 1026 -543
rect 980 -615 986 -581
rect 1020 -615 1026 -581
rect 980 -653 1026 -615
rect 980 -687 986 -653
rect 1020 -687 1026 -653
rect 980 -718 1026 -687
rect 1098 -149 1144 -118
rect 1098 -183 1104 -149
rect 1138 -183 1144 -149
rect 1098 -221 1144 -183
rect 1098 -255 1104 -221
rect 1138 -255 1144 -221
rect 1098 -293 1144 -255
rect 1098 -327 1104 -293
rect 1138 -327 1144 -293
rect 1098 -365 1144 -327
rect 1098 -399 1104 -365
rect 1138 -399 1144 -365
rect 1098 -437 1144 -399
rect 1098 -471 1104 -437
rect 1138 -471 1144 -437
rect 1098 -509 1144 -471
rect 1098 -543 1104 -509
rect 1138 -543 1144 -509
rect 1098 -581 1144 -543
rect 1098 -615 1104 -581
rect 1138 -615 1144 -581
rect 1098 -653 1144 -615
rect 1098 -687 1104 -653
rect 1138 -687 1144 -653
rect 1098 -718 1144 -687
rect 1216 -149 1262 -118
rect 1216 -183 1222 -149
rect 1256 -183 1262 -149
rect 1216 -221 1262 -183
rect 1216 -255 1222 -221
rect 1256 -255 1262 -221
rect 1216 -293 1262 -255
rect 1216 -327 1222 -293
rect 1256 -327 1262 -293
rect 1216 -365 1262 -327
rect 1216 -399 1222 -365
rect 1256 -399 1262 -365
rect 1216 -437 1262 -399
rect 1216 -471 1222 -437
rect 1256 -471 1262 -437
rect 1216 -509 1262 -471
rect 1216 -543 1222 -509
rect 1256 -543 1262 -509
rect 1216 -581 1262 -543
rect 1216 -615 1222 -581
rect 1256 -615 1262 -581
rect 1216 -653 1262 -615
rect 1216 -687 1222 -653
rect 1256 -687 1262 -653
rect 1216 -718 1262 -687
rect 1334 -149 1380 -118
rect 1334 -183 1340 -149
rect 1374 -183 1380 -149
rect 1334 -221 1380 -183
rect 1334 -255 1340 -221
rect 1374 -255 1380 -221
rect 1334 -293 1380 -255
rect 1334 -327 1340 -293
rect 1374 -327 1380 -293
rect 1334 -365 1380 -327
rect 1334 -399 1340 -365
rect 1374 -399 1380 -365
rect 1334 -437 1380 -399
rect 1334 -471 1340 -437
rect 1374 -471 1380 -437
rect 1334 -509 1380 -471
rect 1334 -543 1340 -509
rect 1374 -543 1380 -509
rect 1334 -581 1380 -543
rect 1334 -615 1340 -581
rect 1374 -615 1380 -581
rect 1334 -653 1380 -615
rect 1334 -687 1340 -653
rect 1374 -687 1380 -653
rect 1334 -718 1380 -687
rect 1452 -149 1498 -118
rect 1452 -183 1458 -149
rect 1492 -183 1498 -149
rect 1452 -221 1498 -183
rect 1452 -255 1458 -221
rect 1492 -255 1498 -221
rect 1452 -293 1498 -255
rect 1452 -327 1458 -293
rect 1492 -327 1498 -293
rect 1452 -365 1498 -327
rect 1452 -399 1458 -365
rect 1492 -399 1498 -365
rect 1452 -437 1498 -399
rect 1452 -471 1458 -437
rect 1492 -471 1498 -437
rect 1452 -509 1498 -471
rect 1452 -543 1458 -509
rect 1492 -543 1498 -509
rect 1452 -581 1498 -543
rect 1452 -615 1458 -581
rect 1492 -615 1498 -581
rect 1452 -653 1498 -615
rect 1452 -687 1458 -653
rect 1492 -687 1498 -653
rect 1452 -718 1498 -687
<< properties >>
string FIXED_BBOX -1589 -884 1589 884
<< end >>
