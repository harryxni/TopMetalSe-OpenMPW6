magic
tech sky130A
magscale 1 2
timestamp 1655248036
<< nmoslvt >>
rect 540 -6800 2140 -6400
rect 3540 -6800 5140 -6400
rect 6540 -6800 8140 -6400
<< ndiff >>
rect 540 -6320 2140 -6300
rect 540 -6380 560 -6320
rect 2120 -6380 2140 -6320
rect 540 -6400 2140 -6380
rect 3540 -6320 5140 -6300
rect 3540 -6380 3560 -6320
rect 5120 -6380 5140 -6320
rect 3540 -6400 5140 -6380
rect 6540 -6320 8140 -6300
rect 6540 -6380 6560 -6320
rect 8120 -6380 8140 -6320
rect 6540 -6400 8140 -6380
rect 540 -6830 2140 -6800
rect 540 -6870 560 -6830
rect 2120 -6870 2140 -6830
rect 540 -6880 2140 -6870
rect 3540 -6830 5140 -6800
rect 3540 -6870 3560 -6830
rect 5120 -6870 5140 -6830
rect 3540 -6880 5140 -6870
rect 6540 -6830 8140 -6800
rect 6540 -6870 6560 -6830
rect 8120 -6870 8140 -6830
rect 6540 -6880 8140 -6870
<< ndiffc >>
rect 560 -6380 2120 -6320
rect 3560 -6380 5120 -6320
rect 6560 -6380 8120 -6320
rect 560 -6870 2120 -6830
rect 3560 -6870 5120 -6830
rect 6560 -6870 8120 -6830
<< poly >>
rect 510 -6490 540 -6400
rect 220 -6500 540 -6490
rect 220 -6700 240 -6500
rect 420 -6700 540 -6500
rect 220 -6710 540 -6700
rect 510 -6800 540 -6710
rect 2140 -6800 2170 -6400
rect 3510 -6490 3540 -6400
rect 3220 -6500 3540 -6490
rect 3220 -6700 3240 -6500
rect 3420 -6700 3540 -6500
rect 3220 -6710 3540 -6700
rect 3510 -6800 3540 -6710
rect 5140 -6800 5170 -6400
rect 6510 -6490 6540 -6400
rect 6220 -6500 6540 -6490
rect 6220 -6700 6240 -6500
rect 6420 -6700 6540 -6500
rect 6220 -6710 6540 -6700
rect 6510 -6800 6540 -6710
rect 8140 -6800 8170 -6400
<< polycont >>
rect 240 -6700 420 -6500
rect 3240 -6700 3420 -6500
rect 6240 -6700 6420 -6500
<< locali >>
rect 540 -6290 560 -6230
rect 2120 -6290 2140 -6230
rect 540 -6320 2140 -6290
rect 540 -6380 560 -6320
rect 2120 -6380 2140 -6320
rect 3540 -6290 3560 -6230
rect 5120 -6290 5140 -6230
rect 3540 -6320 5140 -6290
rect 3540 -6380 3560 -6320
rect 5120 -6380 5140 -6320
rect 6540 -6290 6560 -6230
rect 8120 -6290 8140 -6230
rect 6540 -6320 8140 -6290
rect 6540 -6380 6560 -6320
rect 8120 -6380 8140 -6320
rect 220 -6500 440 -6490
rect 220 -6700 240 -6500
rect 420 -6700 440 -6500
rect 220 -6710 440 -6700
rect 3220 -6500 3440 -6490
rect 3220 -6700 3240 -6500
rect 3420 -6700 3440 -6500
rect 3220 -6710 3440 -6700
rect 6220 -6500 6440 -6490
rect 6220 -6700 6240 -6500
rect 6420 -6700 6440 -6500
rect 6220 -6710 6440 -6700
rect 540 -6830 2140 -6800
rect 540 -6870 560 -6830
rect 2120 -6870 2140 -6830
rect 540 -6920 2140 -6870
rect 540 -6980 560 -6920
rect 2120 -6980 2140 -6920
rect 540 -7000 2140 -6980
rect 3540 -6830 5140 -6800
rect 3540 -6870 3560 -6830
rect 5120 -6870 5140 -6830
rect 3540 -6920 5140 -6870
rect 3540 -6980 3560 -6920
rect 5120 -6980 5140 -6920
rect 3540 -7000 5140 -6980
rect 6540 -6830 8140 -6800
rect 6540 -6870 6560 -6830
rect 8120 -6870 8140 -6830
rect 6540 -6920 8140 -6870
rect 6540 -6980 6560 -6920
rect 8120 -6980 8140 -6920
rect 6540 -7000 8140 -6980
<< viali >>
rect 9426 -604 9734 -296
rect 560 -6290 2120 -6230
rect 3560 -6290 5120 -6230
rect 6560 -6290 8120 -6230
rect 240 -6700 420 -6500
rect 3240 -6700 3420 -6500
rect 6240 -6700 6420 -6500
rect 560 -6980 2120 -6920
rect 3560 -6980 5120 -6920
rect 6560 -6980 8120 -6920
<< metal1 >>
rect -1770 3450 8000 3460
rect -900 3360 50 3450
rect 140 3360 3050 3450
rect 3140 3360 6050 3450
rect 6140 3360 8000 3450
rect -1770 3350 8000 3360
rect -2000 2970 -1800 2990
rect -2000 2880 40 2970
rect -2000 2820 0 2880
rect -2000 2170 -1800 2820
rect 9400 2580 9600 2710
rect 10610 2580 10930 2586
rect 9400 2260 10610 2580
rect -2006 1970 -2000 2170
rect -1800 1970 -1794 2170
rect -2000 -20 -1800 1970
rect -1600 1560 0 1570
rect -1600 1490 -1580 1560
rect -1180 1490 -540 1560
rect -260 1490 0 1560
rect -1600 1480 0 1490
rect 9400 180 9600 2260
rect 10610 2254 10930 2260
rect 9000 30 9600 180
rect -2006 -220 -2000 -20
rect -1800 -30 -1794 -20
rect -1800 -120 40 -30
rect -1800 -180 0 -120
rect -1800 -220 -1794 -180
rect -2000 -3030 -1800 -220
rect 9400 -284 9600 30
rect 9400 -290 9740 -284
rect 9400 -610 9420 -290
rect 9740 -610 9746 -290
rect 9400 -616 9740 -610
rect -1600 -1440 0 -1430
rect -1600 -1510 -1580 -1440
rect -1180 -1510 -540 -1440
rect -260 -1510 0 -1440
rect -1600 -1520 0 -1510
rect 9400 -2820 9600 -616
rect 9000 -2970 9600 -2820
rect -2000 -3040 40 -3030
rect -2006 -3240 -2000 -3040
rect -1800 -3120 40 -3040
rect -1800 -3180 0 -3120
rect -1800 -3240 -1794 -3180
rect -2000 -5800 -1800 -3240
rect 9400 -3884 9600 -2970
rect 9400 -3890 9720 -3884
rect 9400 -4216 9720 -4210
rect -1600 -4440 0 -4430
rect -1600 -4510 -1580 -4440
rect -1180 -4510 -540 -4440
rect -260 -4510 0 -4440
rect -1600 -4520 0 -4510
rect -2006 -6000 -2000 -5800
rect -1800 -6000 -1794 -5800
rect 9400 -5820 9600 -4216
rect 2860 -5910 3000 -5830
rect 9000 -5970 9600 -5820
rect 540 -6200 560 -6130
rect 2120 -6200 2140 -6130
rect 540 -6230 2140 -6200
rect 540 -6290 560 -6230
rect 2120 -6290 2140 -6230
rect 540 -6300 2140 -6290
rect 3540 -6200 3560 -6130
rect 5120 -6200 5140 -6130
rect 3540 -6230 5140 -6200
rect 3540 -6290 3560 -6230
rect 5120 -6290 5140 -6230
rect 3540 -6300 5140 -6290
rect 6540 -6200 6560 -6130
rect 8120 -6200 8140 -6130
rect 6540 -6230 8140 -6200
rect 6540 -6290 6560 -6230
rect 8120 -6290 8140 -6230
rect 6540 -6300 8140 -6290
rect 220 -6500 440 -6490
rect 220 -6700 240 -6500
rect 420 -6700 440 -6500
rect 220 -6710 440 -6700
rect 3220 -6500 3440 -6490
rect 3220 -6700 3240 -6500
rect 3420 -6700 3440 -6500
rect 3220 -6710 3440 -6700
rect 6220 -6500 6440 -6490
rect 6220 -6700 6240 -6500
rect 6420 -6700 6440 -6500
rect 6220 -6710 6440 -6700
rect 540 -6920 9740 -6900
rect 540 -7080 560 -6920
rect 540 -7100 9740 -7080
<< via1 >>
rect -1770 3360 -900 3450
rect 50 3360 140 3450
rect 3050 3360 3140 3450
rect 6050 3360 6140 3450
rect 10610 2260 10930 2580
rect -2000 1970 -1800 2170
rect -1580 1490 -1180 1560
rect -540 1490 -260 1560
rect -2000 -220 -1800 -20
rect 9420 -296 9740 -290
rect 9420 -604 9426 -296
rect 9426 -604 9734 -296
rect 9734 -604 9740 -296
rect 9420 -610 9740 -604
rect -1580 -1510 -1180 -1440
rect -540 -1510 -260 -1440
rect -2000 -3240 -1800 -3040
rect 9400 -4210 9720 -3890
rect -1580 -4510 -1180 -4440
rect -540 -4510 -260 -4440
rect -2000 -6000 -1800 -5800
rect 560 -6200 2120 -6130
rect 3560 -6200 5120 -6130
rect 6560 -6200 8120 -6130
rect 240 -6700 420 -6500
rect 3240 -6700 3420 -6500
rect 6240 -6700 6420 -6500
rect 560 -6980 2120 -6920
rect 2120 -6980 3560 -6920
rect 3560 -6980 5120 -6920
rect 5120 -6980 6560 -6920
rect 6560 -6980 8120 -6920
rect 8120 -6980 9740 -6920
rect 560 -7080 9740 -6980
<< metal2 >>
rect 0 4040 9000 4150
rect -3000 3450 -890 3460
rect -3000 3360 -1770 3450
rect -900 3360 -890 3450
rect -3000 3350 -890 3360
rect -2000 2170 -1800 2176
rect -2009 1970 -2000 2170
rect -1800 1970 -1791 2170
rect -2000 1964 -1800 1970
rect -3000 1560 -1000 1570
rect -3000 1490 -1580 1560
rect -1180 1490 -1000 1560
rect -3000 1480 -1000 1490
rect -750 230 -640 4000
rect 480 3650 590 3660
rect 60 3460 130 3600
rect 480 3560 490 3650
rect 580 3560 590 3650
rect 480 3550 590 3560
rect 40 3450 150 3460
rect 40 3360 50 3450
rect 140 3360 150 3450
rect 40 3350 150 3360
rect 60 3000 130 3350
rect 500 3000 570 3550
rect 1020 3000 1090 4040
rect 3480 3650 3590 3660
rect 3060 3460 3130 3600
rect 3480 3560 3490 3650
rect 3580 3560 3590 3650
rect 3480 3550 3590 3560
rect 3040 3450 3150 3460
rect 3040 3360 3050 3450
rect 3140 3360 3150 3450
rect 3040 3350 3150 3360
rect 3060 3000 3130 3350
rect 3500 3000 3570 3550
rect 4020 3000 4090 4040
rect 6480 3650 6590 3660
rect 6060 3460 6130 3600
rect 6480 3560 6490 3650
rect 6580 3560 6590 3650
rect 6480 3550 6590 3560
rect 6040 3450 6150 3460
rect 6040 3360 6050 3450
rect 6140 3360 6150 3450
rect 6040 3350 6150 3360
rect 6060 3000 6130 3350
rect 6500 3000 6570 3550
rect 7020 3000 7090 4040
rect 10615 2580 10925 2584
rect 10604 2260 10610 2580
rect 10930 2260 10936 2580
rect 10615 2256 10925 2260
rect -560 1560 -260 1570
rect -560 1490 -540 1560
rect -560 1480 -260 1490
rect -750 160 -740 230
rect -650 160 -640 230
rect -2000 -20 -1800 -14
rect -2009 -220 -2000 -20
rect -1800 -220 -1791 -20
rect -2000 -226 -1800 -220
rect -3000 -1440 -1000 -1430
rect -3000 -1510 -1580 -1440
rect -1180 -1510 -1000 -1440
rect -3000 -1520 -1000 -1510
rect -750 -2770 -640 160
rect 9425 -290 9735 -286
rect 9414 -610 9420 -290
rect 9740 -610 9746 -290
rect 9425 -614 9735 -610
rect -560 -1440 -260 -1430
rect -560 -1510 -540 -1440
rect -560 -1520 -260 -1510
rect -750 -2840 -740 -2770
rect -650 -2840 -640 -2770
rect -2000 -3040 -1800 -3034
rect -2009 -3240 -2000 -3040
rect -1800 -3240 -1791 -3040
rect -2000 -3246 -1800 -3240
rect -3000 -4440 -1000 -4430
rect -3000 -4510 -1580 -4440
rect -1180 -4510 -1000 -4440
rect -3000 -4520 -1000 -4510
rect -750 -5770 -640 -2840
rect 10615 -3890 10925 -3886
rect 9394 -4210 9400 -3890
rect 9720 -3895 10930 -3890
rect 9720 -4205 10615 -3895
rect 10925 -4205 10930 -3895
rect 9720 -4210 10930 -4205
rect 10615 -4214 10925 -4210
rect -560 -4440 -260 -4430
rect -560 -4510 -540 -4440
rect -560 -4520 -260 -4510
rect -2000 -5800 -1800 -5794
rect -2009 -6000 -2000 -5800
rect -1800 -6000 -1791 -5800
rect -750 -5840 -740 -5770
rect -650 -5840 -640 -5770
rect -750 -6000 -640 -5840
rect -2000 -6006 -1800 -6000
rect 540 -6080 2780 -6060
rect 540 -6200 560 -6080
rect 2760 -6180 2780 -6080
rect 2120 -6200 2780 -6180
rect 3540 -6080 5780 -6060
rect 3540 -6200 3560 -6080
rect 5760 -6180 5780 -6080
rect 5120 -6200 5780 -6180
rect 6540 -6080 8780 -6060
rect 6540 -6200 6560 -6080
rect 8760 -6180 8780 -6080
rect 8120 -6200 8780 -6180
rect 220 -6500 440 -6490
rect 220 -6700 240 -6500
rect 420 -6700 440 -6500
rect 220 -6710 440 -6700
rect 3220 -6500 3440 -6490
rect 3220 -6700 3240 -6500
rect 3420 -6700 3440 -6500
rect 3220 -6710 3440 -6700
rect 6220 -6500 6440 -6490
rect 6220 -6700 6240 -6500
rect 6420 -6700 6440 -6500
rect 6220 -6710 6440 -6700
rect 540 -6920 9740 -6900
rect 540 -7080 560 -6920
rect 540 -7100 9740 -7080
<< via2 >>
rect -2000 1970 -1800 2170
rect 490 3560 580 3650
rect 3490 3560 3580 3650
rect 6490 3560 6580 3650
rect 10615 2265 10925 2575
rect -540 1490 -260 1560
rect -740 160 -650 230
rect -2000 -220 -1800 -20
rect 9425 -605 9735 -295
rect -540 -1510 -260 -1440
rect -740 -2840 -650 -2770
rect -2000 -3240 -1800 -3040
rect 10615 -4205 10925 -3895
rect -540 -4510 -260 -4440
rect -2000 -6000 -1800 -5800
rect -740 -5840 -650 -5770
rect 560 -6130 2760 -6080
rect 560 -6180 2120 -6130
rect 2120 -6180 2760 -6130
rect 3560 -6130 5760 -6080
rect 3560 -6180 5120 -6130
rect 5120 -6180 5760 -6130
rect 6560 -6130 8760 -6080
rect 6560 -6180 8120 -6130
rect 8120 -6180 8760 -6130
rect 240 -6700 420 -6500
rect 3240 -6700 3420 -6500
rect 6240 -6700 6420 -6500
<< metal3 >>
rect -1200 2840 -1110 5000
rect 480 3650 590 3660
rect 480 3560 490 3650
rect 580 3560 590 3650
rect 480 3550 590 3560
rect 3480 3650 3590 3660
rect 3480 3560 3490 3650
rect 3580 3560 3590 3650
rect 3480 3550 3590 3560
rect 6480 3650 6590 3660
rect 6480 3560 6490 3650
rect 6580 3560 6590 3650
rect 6480 3550 6590 3560
rect -1200 2750 200 2840
rect -2011 1965 -2005 2175
rect -1805 2170 -1795 2175
rect -1800 1970 -1795 2170
rect -1805 1965 -1795 1970
rect -2011 -225 -2005 -15
rect -1805 -20 -1795 -15
rect -1800 -220 -1795 -20
rect -1805 -225 -1795 -220
rect -1200 -160 -1110 2750
rect 10611 2580 10929 2585
rect 10610 2579 10930 2580
rect -480 2550 -370 2560
rect -560 2540 520 2550
rect -560 2470 -470 2540
rect -380 2470 520 2540
rect -560 2460 520 2470
rect -480 2450 -370 2460
rect 10610 2261 10611 2579
rect 10929 2261 10930 2579
rect 10610 2260 10930 2261
rect 10611 2255 10929 2260
rect -560 1560 440 1570
rect -560 1490 -540 1560
rect -260 1490 440 1560
rect -560 1480 440 1490
rect -760 230 40 250
rect -760 160 -740 230
rect -650 160 40 230
rect -750 140 -640 160
rect -1200 -250 200 -160
rect -2011 -3245 -2005 -3035
rect -1805 -3040 -1795 -3035
rect -1800 -3240 -1795 -3040
rect -1805 -3245 -1795 -3240
rect -1200 -3160 -1110 -250
rect 10611 -290 10929 -285
rect 9420 -291 10930 -290
rect 9420 -295 10611 -291
rect -480 -450 -370 -440
rect -560 -460 520 -450
rect -560 -530 -470 -460
rect -380 -530 520 -460
rect -560 -540 520 -530
rect -480 -550 -370 -540
rect 9420 -605 9425 -295
rect 9735 -605 10611 -295
rect 9420 -609 10611 -605
rect 10929 -609 10930 -291
rect 9420 -610 10930 -609
rect 10611 -615 10929 -610
rect -560 -1440 440 -1430
rect -560 -1510 -540 -1440
rect -260 -1510 440 -1440
rect -560 -1520 440 -1510
rect -760 -2770 40 -2750
rect -760 -2840 -740 -2770
rect -650 -2840 40 -2770
rect -750 -2860 -640 -2840
rect -1200 -3250 200 -3160
rect -1200 -4000 -1110 -3250
rect -480 -3450 -370 -3440
rect -560 -3460 520 -3450
rect -560 -3530 -470 -3460
rect -380 -3530 520 -3460
rect -560 -3540 520 -3530
rect -480 -3550 -370 -3540
rect 10611 -3890 10929 -3885
rect 10610 -3891 10930 -3890
rect 10610 -4209 10611 -3891
rect 10929 -4209 10930 -3891
rect 10610 -4210 10930 -4209
rect 10611 -4215 10929 -4210
rect -560 -4440 440 -4430
rect -560 -4510 -540 -4440
rect -260 -4510 440 -4440
rect -560 -4520 440 -4510
rect -760 -5770 40 -5750
rect -2005 -5800 -1795 -5795
rect -2446 -6000 -2440 -5800
rect -2240 -6000 -2000 -5800
rect -1800 -6000 -1795 -5800
rect -760 -5840 -740 -5770
rect -650 -5840 40 -5770
rect -750 -5860 -640 -5840
rect -2005 -6005 -1795 -6000
rect 540 -6080 2780 -6060
rect 540 -6180 560 -6080
rect 2760 -6180 2780 -6080
rect 540 -6200 2780 -6180
rect 3540 -6080 5780 -6060
rect 3540 -6180 3560 -6080
rect 5760 -6180 5780 -6080
rect 3540 -6200 5780 -6180
rect 6540 -6080 8780 -6060
rect 6540 -6180 6560 -6080
rect 8760 -6180 8780 -6080
rect 6540 -6200 8780 -6180
rect 220 -6500 440 -6490
rect 220 -6700 240 -6500
rect 420 -6700 440 -6500
rect 220 -6710 440 -6700
rect 3220 -6500 3440 -6490
rect 3220 -6700 3240 -6500
rect 3420 -6700 3440 -6500
rect 3220 -6710 3440 -6700
rect 6220 -6500 6440 -6490
rect 6220 -6700 6240 -6500
rect 6420 -6700 6440 -6500
rect 6220 -6710 6440 -6700
<< via3 >>
rect 490 3560 580 3650
rect 3490 3560 3580 3650
rect 6490 3560 6580 3650
rect -2005 2170 -1805 2175
rect -2005 1970 -2000 2170
rect -2000 1970 -1805 2170
rect -2005 1965 -1805 1970
rect -2005 -20 -1805 -15
rect -2005 -220 -2000 -20
rect -2000 -220 -1805 -20
rect -2005 -225 -1805 -220
rect -470 2470 -380 2540
rect 10611 2575 10929 2579
rect 10611 2265 10615 2575
rect 10615 2265 10925 2575
rect 10925 2265 10929 2575
rect 10611 2261 10929 2265
rect -2005 -3040 -1805 -3035
rect -2005 -3240 -2000 -3040
rect -2000 -3240 -1805 -3040
rect -2005 -3245 -1805 -3240
rect -470 -530 -380 -460
rect 10611 -609 10929 -291
rect -470 -3530 -380 -3460
rect 10611 -3895 10929 -3891
rect 10611 -4205 10615 -3895
rect 10615 -4205 10925 -3895
rect 10925 -4205 10929 -3895
rect 10611 -4209 10929 -4205
rect -2440 -6000 -2240 -5800
rect 560 -6180 2760 -6080
rect 3560 -6180 5760 -6080
rect 6560 -6180 8760 -6080
rect 240 -6700 420 -6500
rect 3240 -6700 3420 -6500
rect 6240 -6700 6420 -6500
<< metal4 >>
rect -3000 3650 8200 3660
rect -3000 3560 490 3650
rect 580 3560 3490 3650
rect 3580 3560 6490 3650
rect 6580 3560 8200 3650
rect -3000 3550 8200 3560
rect -480 2540 -370 2600
rect -480 2470 -470 2540
rect -380 2470 -370 2540
rect -480 -460 -370 2470
rect 10610 2579 10930 2580
rect 10610 2261 10611 2579
rect 10929 2261 10930 2579
rect 10610 2260 10930 2261
rect -480 -530 -470 -460
rect -380 -530 -370 -460
rect -480 -3460 -370 -530
rect 10610 -291 10930 -290
rect 10610 -609 10611 -291
rect 10929 -609 10930 -291
rect 10610 -610 10930 -609
rect -480 -3530 -470 -3460
rect -380 -3530 -370 -3460
rect -2441 -5800 -2239 -5799
rect -2530 -6000 -2440 -5800
rect -2240 -6000 -2239 -5800
rect -2441 -6001 -2239 -6000
rect -480 -7600 -370 -3530
rect 10610 -3891 10930 -3890
rect 10610 -4209 10611 -3891
rect 10929 -4209 10930 -3891
rect 10610 -4210 10930 -4209
rect 2630 -6060 2780 -6000
rect 5630 -6060 5780 -6000
rect 8630 -6060 8780 -6000
rect 540 -6080 2780 -6060
rect 540 -6180 560 -6080
rect 2760 -6180 2780 -6080
rect 540 -6200 2780 -6180
rect 3540 -6080 5780 -6060
rect 3540 -6180 3560 -6080
rect 5760 -6180 5780 -6080
rect 3540 -6200 5780 -6180
rect 6540 -6080 8780 -6060
rect 6540 -6180 6560 -6080
rect 8760 -6180 8780 -6080
rect 6540 -6200 8780 -6180
rect 220 -6500 440 -6490
rect 220 -6700 240 -6500
rect 420 -6700 440 -6500
rect 220 -7100 440 -6700
rect 3220 -6500 3440 -6490
rect 3220 -6700 3240 -6500
rect 3420 -6700 3440 -6500
rect 3220 -7100 3440 -6700
rect 6220 -6500 6440 -6490
rect 6220 -6700 6240 -6500
rect 6420 -6700 6440 -6500
rect 6220 -7100 6440 -6700
<< via4 >>
rect -2065 2175 -1745 2230
rect -2065 1965 -2005 2175
rect -2005 1965 -1805 2175
rect -1805 1965 -1745 2175
rect -2065 1910 -1745 1965
rect -2065 -15 -1745 40
rect -2065 -225 -2005 -15
rect -2005 -225 -1805 -15
rect -1805 -225 -1745 -15
rect -2065 -280 -1745 -225
rect 10634 2284 10906 2556
rect -2065 -3035 -1745 -2980
rect -2065 -3245 -2005 -3035
rect -2005 -3245 -1805 -3035
rect -1805 -3245 -1745 -3035
rect -2065 -3300 -1745 -3245
rect 10634 -586 10906 -314
rect -2850 -6060 -2530 -5740
rect 10634 -4186 10906 -3914
<< metal5 >>
rect -3720 5500 11230 5820
rect -3720 -8280 -3400 5500
rect -2850 3990 9900 4310
rect -2850 2230 -2530 3990
rect -2000 2840 0 3160
rect -2089 2230 -1721 2254
rect -2850 1910 -2065 2230
rect -1745 1910 -1721 2230
rect -2850 40 -2530 1910
rect -2089 1886 -1721 1910
rect 1040 1040 1240 1240
rect 4040 1040 4240 1240
rect 7040 1040 7240 1240
rect -2089 40 -1721 64
rect -2860 -280 -2065 40
rect -1745 -280 -1721 40
rect -2850 -2980 -2530 -280
rect -2089 -304 -1721 -280
rect 1040 -1960 1240 -1760
rect 4040 -1960 4240 -1760
rect 7040 -1960 7240 -1760
rect -2089 -2980 -1721 -2956
rect -2850 -3300 -2065 -2980
rect -1745 -3300 -1721 -2980
rect -2850 -5716 -2530 -3300
rect -2089 -3324 -1721 -3300
rect 1040 -4960 1240 -4760
rect 4040 -4960 4240 -4760
rect 7040 -4960 7240 -4760
rect -2874 -5740 -2506 -5716
rect -2874 -6060 -2850 -5740
rect -2530 -6060 -2506 -5740
rect -2874 -6084 -2506 -6060
rect -2850 -7250 -2530 -6084
rect 9580 -7250 9900 3990
rect 10610 3060 10930 5500
rect 10560 2740 10930 3060
rect -2850 -7560 9900 -7250
rect -2820 -7570 9900 -7560
rect 10610 2556 10930 2740
rect 10610 2284 10634 2556
rect 10906 2284 10930 2556
rect 10610 -314 10930 2284
rect 10610 -586 10634 -314
rect 10906 -586 10930 -314
rect 10610 -3914 10930 -586
rect 10610 -4186 10634 -3914
rect 10906 -4186 10930 -3914
rect 10610 -8280 10930 -4186
rect -3720 -8600 10930 -8280
use pixel  pixel_0
timestamp 1655248036
transform 1 0 -3800 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_1
timestamp 1655248036
transform 1 0 -800 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_2
timestamp 1655248036
transform 1 0 2200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_3
timestamp 1655248036
transform 1 0 -3800 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_4
timestamp 1655248036
transform 1 0 -800 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_5
timestamp 1655248036
transform 1 0 2200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_6
timestamp 1655248036
transform 1 0 -3800 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_7
timestamp 1655248036
transform 1 0 -800 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_8
timestamp 1655248036
transform 1 0 2200 0 1 -3300
box 3640 -2860 6960 460
<< labels >>
rlabel metal2 500 3000 570 3600 1 VBIAS
port 202 n
rlabel metal2 60 3000 130 3600 1 VREF
port 203 n
rlabel metal2 1020 3000 1090 3600 1 NB2
port 204 n
rlabel metal3 -560 2750 40 2840 1 SF_IB
port 206 n
rlabel metal3 -560 2460 40 2550 1 CSA_VREF
port 207 n
rlabel metal3 -560 160 40 250 1 NB1
port 208 n
rlabel metal3 -560 1480 40 1570 1 ROW_SEL0
port 209 n
rlabel metal2 3500 3000 3570 3600 1 VBIAS
rlabel metal2 3060 3000 3130 3600 1 VREF
rlabel metal2 4020 3000 4090 3600 1 NB2
rlabel metal2 6500 3000 6570 3600 1 VBIAS
rlabel metal2 6060 3000 6130 3600 1 VREF
rlabel metal2 7020 3000 7090 3600 1 NB2
rlabel metal1 9000 30 9600 120 1 GND
port 212 n
rlabel metal1 -560 -120 40 -30 1 VDD
rlabel metal3 -560 -250 40 -160 1 SF_IB
rlabel metal3 -560 -540 40 -450 1 CSA_VREF
rlabel metal3 -560 -2840 40 -2750 1 NB1
rlabel metal3 -560 -1520 40 -1430 1 ROW_SEL1
port 214 n
rlabel metal1 9000 -2970 9600 -2880 1 GND
rlabel metal1 -560 -3120 40 -3030 1 VDD
rlabel metal3 -560 -3250 40 -3160 1 SF_IB
rlabel metal3 -560 -3540 40 -3450 1 CSA_VREF
rlabel metal3 -560 -5840 40 -5750 1 NB1
rlabel metal3 -560 -4520 40 -4430 1 ROW_SEL2
port 220 n
rlabel metal1 9000 -5970 9600 -5880 1 GND
rlabel metal4 -1000 3550 -1000 3550 1 VBIAS
port 202 n
rlabel metal1 -1000 3350 -1000 3350 3 VREF
port 203 e
rlabel metal2 -3000 1480 -3000 1480 3 ROW_SEL0
port 209 e
rlabel metal2 -3000 -1520 -3000 -1520 3 ROW_SEL1
port 214 e
rlabel metal2 -3000 -4520 -3000 -4520 3 ROW_SEL2
port 220 e
rlabel metal5 1040 1040 1240 1240 1 PIX0_IN
port 244 n
rlabel metal4 -3000 3550 -3000 3660 1 VBIAS
port 202 n
rlabel metal2 -3000 3350 -3000 3450 3 VREF
port 203 e
rlabel metal2 0 4040 0 4040 1 NB2
port 204 n
rlabel metal1 -2000 0 -2000 0 1 VDD
port 205 n
rlabel metal2 -740 3560 -740 3560 1 NB1
port 208 n
rlabel metal2 -3000 1480 -3000 1570 3 ROW_SEL0
port 209 e
rlabel metal5 -2000 2840 -2000 2840 1 GRING
port 245 n
rlabel metal5 4040 1040 4240 1240 1 PIX1_IN
port 246 n
rlabel metal5 7040 1040 7240 1240 1 PIX2_IN
port 247 n
rlabel metal1 9400 30 9400 30 1 GND
port 212 n
rlabel metal5 1040 -1960 1240 -1760 1 PIX3_IN
port 248 n
rlabel metal2 -3000 -1520 -3000 -1430 3 ROW_SEL1
port 214 e
rlabel metal5 4040 -1960 4240 -1760 1 PIX4_IN
port 249 n
rlabel metal5 7040 -1960 7240 -1760 1 PIX5_IN
port 250 n
rlabel metal5 1040 -4960 1240 -4760 1 PIX6_IN
port 251 n
rlabel metal4 2630 -6200 2780 -6000 1 PIX_OUT0
port 252 n
rlabel metal4 -480 -7600 -480 -7600 1 CSA_VREF
port 207 n
rlabel metal2 -3000 -4520 -3000 -4430 3 ROW_SEL2
port 220 e
rlabel metal5 4040 -4960 4240 -4760 1 PIX7_IN
port 254 n
rlabel metal4 5630 -6200 5780 -6000 1 PIX_OUT1
port 255 n
rlabel metal5 7040 -4960 7240 -4760 1 PIX8_IN
port 257 n
rlabel metal4 8630 -6200 8780 -6000 1 PIX_OUT2
port 258 n
rlabel metal2 8940 -7100 8940 -7100 1 ARRAY_OUT
port 259 n
rlabel metal1 -560 2880 40 2970 1 VDD
port 205 n
rlabel metal4 283 -6958 283 -6958 1 COL_SEL0
port 260 n
rlabel metal4 3346 -6841 3346 -6841 1 COL_SEl1
port 261 n
rlabel metal4 6337 -6795 6337 -6795 1 COL_SEL2
port 262 n
<< end >>
