magic
tech sky130A
timestamp 1654709086
<< nmoslvt >>
rect 270 -118900 1070 -118700
rect 1770 -118900 2570 -118700
rect 3270 -118900 4070 -118700
rect 4770 -118900 5570 -118700
rect 6270 -118900 7070 -118700
rect 7770 -118900 8570 -118700
rect 9270 -118900 10070 -118700
rect 10770 -118900 11570 -118700
rect 12270 -118900 13070 -118700
rect 13770 -118900 14570 -118700
rect 15270 -118900 16070 -118700
rect 16770 -118900 17570 -118700
rect 18270 -118900 19070 -118700
rect 19770 -118900 20570 -118700
rect 21270 -118900 22070 -118700
rect 22770 -118900 23570 -118700
rect 24270 -118900 25070 -118700
rect 25770 -118900 26570 -118700
rect 27270 -118900 28070 -118700
rect 28770 -118900 29570 -118700
rect 30270 -118900 31070 -118700
rect 31770 -118900 32570 -118700
rect 33270 -118900 34070 -118700
rect 34770 -118900 35570 -118700
rect 36270 -118900 37070 -118700
rect 37770 -118900 38570 -118700
rect 39270 -118900 40070 -118700
rect 40770 -118900 41570 -118700
rect 42270 -118900 43070 -118700
rect 43770 -118900 44570 -118700
rect 45270 -118900 46070 -118700
rect 46770 -118900 47570 -118700
rect 48270 -118900 49070 -118700
rect 49770 -118900 50570 -118700
rect 51270 -118900 52070 -118700
rect 52770 -118900 53570 -118700
rect 54270 -118900 55070 -118700
rect 55770 -118900 56570 -118700
rect 57270 -118900 58070 -118700
rect 58770 -118900 59570 -118700
rect 60270 -118900 61070 -118700
rect 61770 -118900 62570 -118700
rect 63270 -118900 64070 -118700
rect 64770 -118900 65570 -118700
rect 66270 -118900 67070 -118700
rect 67770 -118900 68570 -118700
rect 69270 -118900 70070 -118700
rect 70770 -118900 71570 -118700
rect 72270 -118900 73070 -118700
rect 73770 -118900 74570 -118700
rect 75270 -118900 76070 -118700
rect 76770 -118900 77570 -118700
rect 78270 -118900 79070 -118700
rect 79770 -118900 80570 -118700
rect 81270 -118900 82070 -118700
rect 82770 -118900 83570 -118700
rect 84270 -118900 85070 -118700
rect 85770 -118900 86570 -118700
rect 87270 -118900 88070 -118700
rect 88770 -118900 89570 -118700
rect 90270 -118900 91070 -118700
rect 91770 -118900 92570 -118700
rect 93270 -118900 94070 -118700
rect 94770 -118900 95570 -118700
rect 96270 -118900 97070 -118700
rect 97770 -118900 98570 -118700
rect 99270 -118900 100070 -118700
rect 100770 -118900 101570 -118700
rect 102270 -118900 103070 -118700
rect 103770 -118900 104570 -118700
rect 105270 -118900 106070 -118700
rect 106770 -118900 107570 -118700
rect 108270 -118900 109070 -118700
rect 109770 -118900 110570 -118700
rect 111270 -118900 112070 -118700
rect 112770 -118900 113570 -118700
rect 114270 -118900 115070 -118700
rect 115770 -118900 116570 -118700
rect 117270 -118900 118070 -118700
rect 118770 -118900 119570 -118700
<< ndiff >>
rect 270 -118660 1070 -118650
rect 270 -118690 280 -118660
rect 1060 -118690 1070 -118660
rect 270 -118700 1070 -118690
rect 1770 -118660 2570 -118650
rect 1770 -118690 1780 -118660
rect 2560 -118690 2570 -118660
rect 1770 -118700 2570 -118690
rect 3270 -118660 4070 -118650
rect 3270 -118690 3280 -118660
rect 4060 -118690 4070 -118660
rect 3270 -118700 4070 -118690
rect 4770 -118660 5570 -118650
rect 4770 -118690 4780 -118660
rect 5560 -118690 5570 -118660
rect 4770 -118700 5570 -118690
rect 6270 -118660 7070 -118650
rect 6270 -118690 6280 -118660
rect 7060 -118690 7070 -118660
rect 6270 -118700 7070 -118690
rect 7770 -118660 8570 -118650
rect 7770 -118690 7780 -118660
rect 8560 -118690 8570 -118660
rect 7770 -118700 8570 -118690
rect 9270 -118660 10070 -118650
rect 9270 -118690 9280 -118660
rect 10060 -118690 10070 -118660
rect 9270 -118700 10070 -118690
rect 10770 -118660 11570 -118650
rect 10770 -118690 10780 -118660
rect 11560 -118690 11570 -118660
rect 10770 -118700 11570 -118690
rect 12270 -118660 13070 -118650
rect 12270 -118690 12280 -118660
rect 13060 -118690 13070 -118660
rect 12270 -118700 13070 -118690
rect 13770 -118660 14570 -118650
rect 13770 -118690 13780 -118660
rect 14560 -118690 14570 -118660
rect 13770 -118700 14570 -118690
rect 15270 -118660 16070 -118650
rect 15270 -118690 15280 -118660
rect 16060 -118690 16070 -118660
rect 15270 -118700 16070 -118690
rect 16770 -118660 17570 -118650
rect 16770 -118690 16780 -118660
rect 17560 -118690 17570 -118660
rect 16770 -118700 17570 -118690
rect 18270 -118660 19070 -118650
rect 18270 -118690 18280 -118660
rect 19060 -118690 19070 -118660
rect 18270 -118700 19070 -118690
rect 19770 -118660 20570 -118650
rect 19770 -118690 19780 -118660
rect 20560 -118690 20570 -118660
rect 19770 -118700 20570 -118690
rect 21270 -118660 22070 -118650
rect 21270 -118690 21280 -118660
rect 22060 -118690 22070 -118660
rect 21270 -118700 22070 -118690
rect 22770 -118660 23570 -118650
rect 22770 -118690 22780 -118660
rect 23560 -118690 23570 -118660
rect 22770 -118700 23570 -118690
rect 24270 -118660 25070 -118650
rect 24270 -118690 24280 -118660
rect 25060 -118690 25070 -118660
rect 24270 -118700 25070 -118690
rect 25770 -118660 26570 -118650
rect 25770 -118690 25780 -118660
rect 26560 -118690 26570 -118660
rect 25770 -118700 26570 -118690
rect 27270 -118660 28070 -118650
rect 27270 -118690 27280 -118660
rect 28060 -118690 28070 -118660
rect 27270 -118700 28070 -118690
rect 28770 -118660 29570 -118650
rect 28770 -118690 28780 -118660
rect 29560 -118690 29570 -118660
rect 28770 -118700 29570 -118690
rect 30270 -118660 31070 -118650
rect 30270 -118690 30280 -118660
rect 31060 -118690 31070 -118660
rect 30270 -118700 31070 -118690
rect 31770 -118660 32570 -118650
rect 31770 -118690 31780 -118660
rect 32560 -118690 32570 -118660
rect 31770 -118700 32570 -118690
rect 33270 -118660 34070 -118650
rect 33270 -118690 33280 -118660
rect 34060 -118690 34070 -118660
rect 33270 -118700 34070 -118690
rect 34770 -118660 35570 -118650
rect 34770 -118690 34780 -118660
rect 35560 -118690 35570 -118660
rect 34770 -118700 35570 -118690
rect 36270 -118660 37070 -118650
rect 36270 -118690 36280 -118660
rect 37060 -118690 37070 -118660
rect 36270 -118700 37070 -118690
rect 37770 -118660 38570 -118650
rect 37770 -118690 37780 -118660
rect 38560 -118690 38570 -118660
rect 37770 -118700 38570 -118690
rect 39270 -118660 40070 -118650
rect 39270 -118690 39280 -118660
rect 40060 -118690 40070 -118660
rect 39270 -118700 40070 -118690
rect 40770 -118660 41570 -118650
rect 40770 -118690 40780 -118660
rect 41560 -118690 41570 -118660
rect 40770 -118700 41570 -118690
rect 42270 -118660 43070 -118650
rect 42270 -118690 42280 -118660
rect 43060 -118690 43070 -118660
rect 42270 -118700 43070 -118690
rect 43770 -118660 44570 -118650
rect 43770 -118690 43780 -118660
rect 44560 -118690 44570 -118660
rect 43770 -118700 44570 -118690
rect 45270 -118660 46070 -118650
rect 45270 -118690 45280 -118660
rect 46060 -118690 46070 -118660
rect 45270 -118700 46070 -118690
rect 46770 -118660 47570 -118650
rect 46770 -118690 46780 -118660
rect 47560 -118690 47570 -118660
rect 46770 -118700 47570 -118690
rect 48270 -118660 49070 -118650
rect 48270 -118690 48280 -118660
rect 49060 -118690 49070 -118660
rect 48270 -118700 49070 -118690
rect 49770 -118660 50570 -118650
rect 49770 -118690 49780 -118660
rect 50560 -118690 50570 -118660
rect 49770 -118700 50570 -118690
rect 51270 -118660 52070 -118650
rect 51270 -118690 51280 -118660
rect 52060 -118690 52070 -118660
rect 51270 -118700 52070 -118690
rect 52770 -118660 53570 -118650
rect 52770 -118690 52780 -118660
rect 53560 -118690 53570 -118660
rect 52770 -118700 53570 -118690
rect 54270 -118660 55070 -118650
rect 54270 -118690 54280 -118660
rect 55060 -118690 55070 -118660
rect 54270 -118700 55070 -118690
rect 55770 -118660 56570 -118650
rect 55770 -118690 55780 -118660
rect 56560 -118690 56570 -118660
rect 55770 -118700 56570 -118690
rect 57270 -118660 58070 -118650
rect 57270 -118690 57280 -118660
rect 58060 -118690 58070 -118660
rect 57270 -118700 58070 -118690
rect 58770 -118660 59570 -118650
rect 58770 -118690 58780 -118660
rect 59560 -118690 59570 -118660
rect 58770 -118700 59570 -118690
rect 60270 -118660 61070 -118650
rect 60270 -118690 60280 -118660
rect 61060 -118690 61070 -118660
rect 60270 -118700 61070 -118690
rect 61770 -118660 62570 -118650
rect 61770 -118690 61780 -118660
rect 62560 -118690 62570 -118660
rect 61770 -118700 62570 -118690
rect 63270 -118660 64070 -118650
rect 63270 -118690 63280 -118660
rect 64060 -118690 64070 -118660
rect 63270 -118700 64070 -118690
rect 64770 -118660 65570 -118650
rect 64770 -118690 64780 -118660
rect 65560 -118690 65570 -118660
rect 64770 -118700 65570 -118690
rect 66270 -118660 67070 -118650
rect 66270 -118690 66280 -118660
rect 67060 -118690 67070 -118660
rect 66270 -118700 67070 -118690
rect 67770 -118660 68570 -118650
rect 67770 -118690 67780 -118660
rect 68560 -118690 68570 -118660
rect 67770 -118700 68570 -118690
rect 69270 -118660 70070 -118650
rect 69270 -118690 69280 -118660
rect 70060 -118690 70070 -118660
rect 69270 -118700 70070 -118690
rect 70770 -118660 71570 -118650
rect 70770 -118690 70780 -118660
rect 71560 -118690 71570 -118660
rect 70770 -118700 71570 -118690
rect 72270 -118660 73070 -118650
rect 72270 -118690 72280 -118660
rect 73060 -118690 73070 -118660
rect 72270 -118700 73070 -118690
rect 73770 -118660 74570 -118650
rect 73770 -118690 73780 -118660
rect 74560 -118690 74570 -118660
rect 73770 -118700 74570 -118690
rect 75270 -118660 76070 -118650
rect 75270 -118690 75280 -118660
rect 76060 -118690 76070 -118660
rect 75270 -118700 76070 -118690
rect 76770 -118660 77570 -118650
rect 76770 -118690 76780 -118660
rect 77560 -118690 77570 -118660
rect 76770 -118700 77570 -118690
rect 78270 -118660 79070 -118650
rect 78270 -118690 78280 -118660
rect 79060 -118690 79070 -118660
rect 78270 -118700 79070 -118690
rect 79770 -118660 80570 -118650
rect 79770 -118690 79780 -118660
rect 80560 -118690 80570 -118660
rect 79770 -118700 80570 -118690
rect 81270 -118660 82070 -118650
rect 81270 -118690 81280 -118660
rect 82060 -118690 82070 -118660
rect 81270 -118700 82070 -118690
rect 82770 -118660 83570 -118650
rect 82770 -118690 82780 -118660
rect 83560 -118690 83570 -118660
rect 82770 -118700 83570 -118690
rect 84270 -118660 85070 -118650
rect 84270 -118690 84280 -118660
rect 85060 -118690 85070 -118660
rect 84270 -118700 85070 -118690
rect 85770 -118660 86570 -118650
rect 85770 -118690 85780 -118660
rect 86560 -118690 86570 -118660
rect 85770 -118700 86570 -118690
rect 87270 -118660 88070 -118650
rect 87270 -118690 87280 -118660
rect 88060 -118690 88070 -118660
rect 87270 -118700 88070 -118690
rect 88770 -118660 89570 -118650
rect 88770 -118690 88780 -118660
rect 89560 -118690 89570 -118660
rect 88770 -118700 89570 -118690
rect 90270 -118660 91070 -118650
rect 90270 -118690 90280 -118660
rect 91060 -118690 91070 -118660
rect 90270 -118700 91070 -118690
rect 91770 -118660 92570 -118650
rect 91770 -118690 91780 -118660
rect 92560 -118690 92570 -118660
rect 91770 -118700 92570 -118690
rect 93270 -118660 94070 -118650
rect 93270 -118690 93280 -118660
rect 94060 -118690 94070 -118660
rect 93270 -118700 94070 -118690
rect 94770 -118660 95570 -118650
rect 94770 -118690 94780 -118660
rect 95560 -118690 95570 -118660
rect 94770 -118700 95570 -118690
rect 96270 -118660 97070 -118650
rect 96270 -118690 96280 -118660
rect 97060 -118690 97070 -118660
rect 96270 -118700 97070 -118690
rect 97770 -118660 98570 -118650
rect 97770 -118690 97780 -118660
rect 98560 -118690 98570 -118660
rect 97770 -118700 98570 -118690
rect 99270 -118660 100070 -118650
rect 99270 -118690 99280 -118660
rect 100060 -118690 100070 -118660
rect 99270 -118700 100070 -118690
rect 100770 -118660 101570 -118650
rect 100770 -118690 100780 -118660
rect 101560 -118690 101570 -118660
rect 100770 -118700 101570 -118690
rect 102270 -118660 103070 -118650
rect 102270 -118690 102280 -118660
rect 103060 -118690 103070 -118660
rect 102270 -118700 103070 -118690
rect 103770 -118660 104570 -118650
rect 103770 -118690 103780 -118660
rect 104560 -118690 104570 -118660
rect 103770 -118700 104570 -118690
rect 105270 -118660 106070 -118650
rect 105270 -118690 105280 -118660
rect 106060 -118690 106070 -118660
rect 105270 -118700 106070 -118690
rect 106770 -118660 107570 -118650
rect 106770 -118690 106780 -118660
rect 107560 -118690 107570 -118660
rect 106770 -118700 107570 -118690
rect 108270 -118660 109070 -118650
rect 108270 -118690 108280 -118660
rect 109060 -118690 109070 -118660
rect 108270 -118700 109070 -118690
rect 109770 -118660 110570 -118650
rect 109770 -118690 109780 -118660
rect 110560 -118690 110570 -118660
rect 109770 -118700 110570 -118690
rect 111270 -118660 112070 -118650
rect 111270 -118690 111280 -118660
rect 112060 -118690 112070 -118660
rect 111270 -118700 112070 -118690
rect 112770 -118660 113570 -118650
rect 112770 -118690 112780 -118660
rect 113560 -118690 113570 -118660
rect 112770 -118700 113570 -118690
rect 114270 -118660 115070 -118650
rect 114270 -118690 114280 -118660
rect 115060 -118690 115070 -118660
rect 114270 -118700 115070 -118690
rect 115770 -118660 116570 -118650
rect 115770 -118690 115780 -118660
rect 116560 -118690 116570 -118660
rect 115770 -118700 116570 -118690
rect 117270 -118660 118070 -118650
rect 117270 -118690 117280 -118660
rect 118060 -118690 118070 -118660
rect 117270 -118700 118070 -118690
rect 118770 -118660 119570 -118650
rect 118770 -118690 118780 -118660
rect 119560 -118690 119570 -118660
rect 118770 -118700 119570 -118690
rect 270 -118915 1070 -118900
rect 270 -118935 280 -118915
rect 1060 -118935 1070 -118915
rect 270 -118940 1070 -118935
rect 1770 -118915 2570 -118900
rect 1770 -118935 1780 -118915
rect 2560 -118935 2570 -118915
rect 1770 -118940 2570 -118935
rect 3270 -118915 4070 -118900
rect 3270 -118935 3280 -118915
rect 4060 -118935 4070 -118915
rect 3270 -118940 4070 -118935
rect 4770 -118915 5570 -118900
rect 4770 -118935 4780 -118915
rect 5560 -118935 5570 -118915
rect 4770 -118940 5570 -118935
rect 6270 -118915 7070 -118900
rect 6270 -118935 6280 -118915
rect 7060 -118935 7070 -118915
rect 6270 -118940 7070 -118935
rect 7770 -118915 8570 -118900
rect 7770 -118935 7780 -118915
rect 8560 -118935 8570 -118915
rect 7770 -118940 8570 -118935
rect 9270 -118915 10070 -118900
rect 9270 -118935 9280 -118915
rect 10060 -118935 10070 -118915
rect 9270 -118940 10070 -118935
rect 10770 -118915 11570 -118900
rect 10770 -118935 10780 -118915
rect 11560 -118935 11570 -118915
rect 10770 -118940 11570 -118935
rect 12270 -118915 13070 -118900
rect 12270 -118935 12280 -118915
rect 13060 -118935 13070 -118915
rect 12270 -118940 13070 -118935
rect 13770 -118915 14570 -118900
rect 13770 -118935 13780 -118915
rect 14560 -118935 14570 -118915
rect 13770 -118940 14570 -118935
rect 15270 -118915 16070 -118900
rect 15270 -118935 15280 -118915
rect 16060 -118935 16070 -118915
rect 15270 -118940 16070 -118935
rect 16770 -118915 17570 -118900
rect 16770 -118935 16780 -118915
rect 17560 -118935 17570 -118915
rect 16770 -118940 17570 -118935
rect 18270 -118915 19070 -118900
rect 18270 -118935 18280 -118915
rect 19060 -118935 19070 -118915
rect 18270 -118940 19070 -118935
rect 19770 -118915 20570 -118900
rect 19770 -118935 19780 -118915
rect 20560 -118935 20570 -118915
rect 19770 -118940 20570 -118935
rect 21270 -118915 22070 -118900
rect 21270 -118935 21280 -118915
rect 22060 -118935 22070 -118915
rect 21270 -118940 22070 -118935
rect 22770 -118915 23570 -118900
rect 22770 -118935 22780 -118915
rect 23560 -118935 23570 -118915
rect 22770 -118940 23570 -118935
rect 24270 -118915 25070 -118900
rect 24270 -118935 24280 -118915
rect 25060 -118935 25070 -118915
rect 24270 -118940 25070 -118935
rect 25770 -118915 26570 -118900
rect 25770 -118935 25780 -118915
rect 26560 -118935 26570 -118915
rect 25770 -118940 26570 -118935
rect 27270 -118915 28070 -118900
rect 27270 -118935 27280 -118915
rect 28060 -118935 28070 -118915
rect 27270 -118940 28070 -118935
rect 28770 -118915 29570 -118900
rect 28770 -118935 28780 -118915
rect 29560 -118935 29570 -118915
rect 28770 -118940 29570 -118935
rect 30270 -118915 31070 -118900
rect 30270 -118935 30280 -118915
rect 31060 -118935 31070 -118915
rect 30270 -118940 31070 -118935
rect 31770 -118915 32570 -118900
rect 31770 -118935 31780 -118915
rect 32560 -118935 32570 -118915
rect 31770 -118940 32570 -118935
rect 33270 -118915 34070 -118900
rect 33270 -118935 33280 -118915
rect 34060 -118935 34070 -118915
rect 33270 -118940 34070 -118935
rect 34770 -118915 35570 -118900
rect 34770 -118935 34780 -118915
rect 35560 -118935 35570 -118915
rect 34770 -118940 35570 -118935
rect 36270 -118915 37070 -118900
rect 36270 -118935 36280 -118915
rect 37060 -118935 37070 -118915
rect 36270 -118940 37070 -118935
rect 37770 -118915 38570 -118900
rect 37770 -118935 37780 -118915
rect 38560 -118935 38570 -118915
rect 37770 -118940 38570 -118935
rect 39270 -118915 40070 -118900
rect 39270 -118935 39280 -118915
rect 40060 -118935 40070 -118915
rect 39270 -118940 40070 -118935
rect 40770 -118915 41570 -118900
rect 40770 -118935 40780 -118915
rect 41560 -118935 41570 -118915
rect 40770 -118940 41570 -118935
rect 42270 -118915 43070 -118900
rect 42270 -118935 42280 -118915
rect 43060 -118935 43070 -118915
rect 42270 -118940 43070 -118935
rect 43770 -118915 44570 -118900
rect 43770 -118935 43780 -118915
rect 44560 -118935 44570 -118915
rect 43770 -118940 44570 -118935
rect 45270 -118915 46070 -118900
rect 45270 -118935 45280 -118915
rect 46060 -118935 46070 -118915
rect 45270 -118940 46070 -118935
rect 46770 -118915 47570 -118900
rect 46770 -118935 46780 -118915
rect 47560 -118935 47570 -118915
rect 46770 -118940 47570 -118935
rect 48270 -118915 49070 -118900
rect 48270 -118935 48280 -118915
rect 49060 -118935 49070 -118915
rect 48270 -118940 49070 -118935
rect 49770 -118915 50570 -118900
rect 49770 -118935 49780 -118915
rect 50560 -118935 50570 -118915
rect 49770 -118940 50570 -118935
rect 51270 -118915 52070 -118900
rect 51270 -118935 51280 -118915
rect 52060 -118935 52070 -118915
rect 51270 -118940 52070 -118935
rect 52770 -118915 53570 -118900
rect 52770 -118935 52780 -118915
rect 53560 -118935 53570 -118915
rect 52770 -118940 53570 -118935
rect 54270 -118915 55070 -118900
rect 54270 -118935 54280 -118915
rect 55060 -118935 55070 -118915
rect 54270 -118940 55070 -118935
rect 55770 -118915 56570 -118900
rect 55770 -118935 55780 -118915
rect 56560 -118935 56570 -118915
rect 55770 -118940 56570 -118935
rect 57270 -118915 58070 -118900
rect 57270 -118935 57280 -118915
rect 58060 -118935 58070 -118915
rect 57270 -118940 58070 -118935
rect 58770 -118915 59570 -118900
rect 58770 -118935 58780 -118915
rect 59560 -118935 59570 -118915
rect 58770 -118940 59570 -118935
rect 60270 -118915 61070 -118900
rect 60270 -118935 60280 -118915
rect 61060 -118935 61070 -118915
rect 60270 -118940 61070 -118935
rect 61770 -118915 62570 -118900
rect 61770 -118935 61780 -118915
rect 62560 -118935 62570 -118915
rect 61770 -118940 62570 -118935
rect 63270 -118915 64070 -118900
rect 63270 -118935 63280 -118915
rect 64060 -118935 64070 -118915
rect 63270 -118940 64070 -118935
rect 64770 -118915 65570 -118900
rect 64770 -118935 64780 -118915
rect 65560 -118935 65570 -118915
rect 64770 -118940 65570 -118935
rect 66270 -118915 67070 -118900
rect 66270 -118935 66280 -118915
rect 67060 -118935 67070 -118915
rect 66270 -118940 67070 -118935
rect 67770 -118915 68570 -118900
rect 67770 -118935 67780 -118915
rect 68560 -118935 68570 -118915
rect 67770 -118940 68570 -118935
rect 69270 -118915 70070 -118900
rect 69270 -118935 69280 -118915
rect 70060 -118935 70070 -118915
rect 69270 -118940 70070 -118935
rect 70770 -118915 71570 -118900
rect 70770 -118935 70780 -118915
rect 71560 -118935 71570 -118915
rect 70770 -118940 71570 -118935
rect 72270 -118915 73070 -118900
rect 72270 -118935 72280 -118915
rect 73060 -118935 73070 -118915
rect 72270 -118940 73070 -118935
rect 73770 -118915 74570 -118900
rect 73770 -118935 73780 -118915
rect 74560 -118935 74570 -118915
rect 73770 -118940 74570 -118935
rect 75270 -118915 76070 -118900
rect 75270 -118935 75280 -118915
rect 76060 -118935 76070 -118915
rect 75270 -118940 76070 -118935
rect 76770 -118915 77570 -118900
rect 76770 -118935 76780 -118915
rect 77560 -118935 77570 -118915
rect 76770 -118940 77570 -118935
rect 78270 -118915 79070 -118900
rect 78270 -118935 78280 -118915
rect 79060 -118935 79070 -118915
rect 78270 -118940 79070 -118935
rect 79770 -118915 80570 -118900
rect 79770 -118935 79780 -118915
rect 80560 -118935 80570 -118915
rect 79770 -118940 80570 -118935
rect 81270 -118915 82070 -118900
rect 81270 -118935 81280 -118915
rect 82060 -118935 82070 -118915
rect 81270 -118940 82070 -118935
rect 82770 -118915 83570 -118900
rect 82770 -118935 82780 -118915
rect 83560 -118935 83570 -118915
rect 82770 -118940 83570 -118935
rect 84270 -118915 85070 -118900
rect 84270 -118935 84280 -118915
rect 85060 -118935 85070 -118915
rect 84270 -118940 85070 -118935
rect 85770 -118915 86570 -118900
rect 85770 -118935 85780 -118915
rect 86560 -118935 86570 -118915
rect 85770 -118940 86570 -118935
rect 87270 -118915 88070 -118900
rect 87270 -118935 87280 -118915
rect 88060 -118935 88070 -118915
rect 87270 -118940 88070 -118935
rect 88770 -118915 89570 -118900
rect 88770 -118935 88780 -118915
rect 89560 -118935 89570 -118915
rect 88770 -118940 89570 -118935
rect 90270 -118915 91070 -118900
rect 90270 -118935 90280 -118915
rect 91060 -118935 91070 -118915
rect 90270 -118940 91070 -118935
rect 91770 -118915 92570 -118900
rect 91770 -118935 91780 -118915
rect 92560 -118935 92570 -118915
rect 91770 -118940 92570 -118935
rect 93270 -118915 94070 -118900
rect 93270 -118935 93280 -118915
rect 94060 -118935 94070 -118915
rect 93270 -118940 94070 -118935
rect 94770 -118915 95570 -118900
rect 94770 -118935 94780 -118915
rect 95560 -118935 95570 -118915
rect 94770 -118940 95570 -118935
rect 96270 -118915 97070 -118900
rect 96270 -118935 96280 -118915
rect 97060 -118935 97070 -118915
rect 96270 -118940 97070 -118935
rect 97770 -118915 98570 -118900
rect 97770 -118935 97780 -118915
rect 98560 -118935 98570 -118915
rect 97770 -118940 98570 -118935
rect 99270 -118915 100070 -118900
rect 99270 -118935 99280 -118915
rect 100060 -118935 100070 -118915
rect 99270 -118940 100070 -118935
rect 100770 -118915 101570 -118900
rect 100770 -118935 100780 -118915
rect 101560 -118935 101570 -118915
rect 100770 -118940 101570 -118935
rect 102270 -118915 103070 -118900
rect 102270 -118935 102280 -118915
rect 103060 -118935 103070 -118915
rect 102270 -118940 103070 -118935
rect 103770 -118915 104570 -118900
rect 103770 -118935 103780 -118915
rect 104560 -118935 104570 -118915
rect 103770 -118940 104570 -118935
rect 105270 -118915 106070 -118900
rect 105270 -118935 105280 -118915
rect 106060 -118935 106070 -118915
rect 105270 -118940 106070 -118935
rect 106770 -118915 107570 -118900
rect 106770 -118935 106780 -118915
rect 107560 -118935 107570 -118915
rect 106770 -118940 107570 -118935
rect 108270 -118915 109070 -118900
rect 108270 -118935 108280 -118915
rect 109060 -118935 109070 -118915
rect 108270 -118940 109070 -118935
rect 109770 -118915 110570 -118900
rect 109770 -118935 109780 -118915
rect 110560 -118935 110570 -118915
rect 109770 -118940 110570 -118935
rect 111270 -118915 112070 -118900
rect 111270 -118935 111280 -118915
rect 112060 -118935 112070 -118915
rect 111270 -118940 112070 -118935
rect 112770 -118915 113570 -118900
rect 112770 -118935 112780 -118915
rect 113560 -118935 113570 -118915
rect 112770 -118940 113570 -118935
rect 114270 -118915 115070 -118900
rect 114270 -118935 114280 -118915
rect 115060 -118935 115070 -118915
rect 114270 -118940 115070 -118935
rect 115770 -118915 116570 -118900
rect 115770 -118935 115780 -118915
rect 116560 -118935 116570 -118915
rect 115770 -118940 116570 -118935
rect 117270 -118915 118070 -118900
rect 117270 -118935 117280 -118915
rect 118060 -118935 118070 -118915
rect 117270 -118940 118070 -118935
rect 118770 -118915 119570 -118900
rect 118770 -118935 118780 -118915
rect 119560 -118935 119570 -118915
rect 118770 -118940 119570 -118935
<< ndiffc >>
rect 280 -118690 1060 -118660
rect 1780 -118690 2560 -118660
rect 3280 -118690 4060 -118660
rect 4780 -118690 5560 -118660
rect 6280 -118690 7060 -118660
rect 7780 -118690 8560 -118660
rect 9280 -118690 10060 -118660
rect 10780 -118690 11560 -118660
rect 12280 -118690 13060 -118660
rect 13780 -118690 14560 -118660
rect 15280 -118690 16060 -118660
rect 16780 -118690 17560 -118660
rect 18280 -118690 19060 -118660
rect 19780 -118690 20560 -118660
rect 21280 -118690 22060 -118660
rect 22780 -118690 23560 -118660
rect 24280 -118690 25060 -118660
rect 25780 -118690 26560 -118660
rect 27280 -118690 28060 -118660
rect 28780 -118690 29560 -118660
rect 30280 -118690 31060 -118660
rect 31780 -118690 32560 -118660
rect 33280 -118690 34060 -118660
rect 34780 -118690 35560 -118660
rect 36280 -118690 37060 -118660
rect 37780 -118690 38560 -118660
rect 39280 -118690 40060 -118660
rect 40780 -118690 41560 -118660
rect 42280 -118690 43060 -118660
rect 43780 -118690 44560 -118660
rect 45280 -118690 46060 -118660
rect 46780 -118690 47560 -118660
rect 48280 -118690 49060 -118660
rect 49780 -118690 50560 -118660
rect 51280 -118690 52060 -118660
rect 52780 -118690 53560 -118660
rect 54280 -118690 55060 -118660
rect 55780 -118690 56560 -118660
rect 57280 -118690 58060 -118660
rect 58780 -118690 59560 -118660
rect 60280 -118690 61060 -118660
rect 61780 -118690 62560 -118660
rect 63280 -118690 64060 -118660
rect 64780 -118690 65560 -118660
rect 66280 -118690 67060 -118660
rect 67780 -118690 68560 -118660
rect 69280 -118690 70060 -118660
rect 70780 -118690 71560 -118660
rect 72280 -118690 73060 -118660
rect 73780 -118690 74560 -118660
rect 75280 -118690 76060 -118660
rect 76780 -118690 77560 -118660
rect 78280 -118690 79060 -118660
rect 79780 -118690 80560 -118660
rect 81280 -118690 82060 -118660
rect 82780 -118690 83560 -118660
rect 84280 -118690 85060 -118660
rect 85780 -118690 86560 -118660
rect 87280 -118690 88060 -118660
rect 88780 -118690 89560 -118660
rect 90280 -118690 91060 -118660
rect 91780 -118690 92560 -118660
rect 93280 -118690 94060 -118660
rect 94780 -118690 95560 -118660
rect 96280 -118690 97060 -118660
rect 97780 -118690 98560 -118660
rect 99280 -118690 100060 -118660
rect 100780 -118690 101560 -118660
rect 102280 -118690 103060 -118660
rect 103780 -118690 104560 -118660
rect 105280 -118690 106060 -118660
rect 106780 -118690 107560 -118660
rect 108280 -118690 109060 -118660
rect 109780 -118690 110560 -118660
rect 111280 -118690 112060 -118660
rect 112780 -118690 113560 -118660
rect 114280 -118690 115060 -118660
rect 115780 -118690 116560 -118660
rect 117280 -118690 118060 -118660
rect 118780 -118690 119560 -118660
rect 280 -118935 1060 -118915
rect 1780 -118935 2560 -118915
rect 3280 -118935 4060 -118915
rect 4780 -118935 5560 -118915
rect 6280 -118935 7060 -118915
rect 7780 -118935 8560 -118915
rect 9280 -118935 10060 -118915
rect 10780 -118935 11560 -118915
rect 12280 -118935 13060 -118915
rect 13780 -118935 14560 -118915
rect 15280 -118935 16060 -118915
rect 16780 -118935 17560 -118915
rect 18280 -118935 19060 -118915
rect 19780 -118935 20560 -118915
rect 21280 -118935 22060 -118915
rect 22780 -118935 23560 -118915
rect 24280 -118935 25060 -118915
rect 25780 -118935 26560 -118915
rect 27280 -118935 28060 -118915
rect 28780 -118935 29560 -118915
rect 30280 -118935 31060 -118915
rect 31780 -118935 32560 -118915
rect 33280 -118935 34060 -118915
rect 34780 -118935 35560 -118915
rect 36280 -118935 37060 -118915
rect 37780 -118935 38560 -118915
rect 39280 -118935 40060 -118915
rect 40780 -118935 41560 -118915
rect 42280 -118935 43060 -118915
rect 43780 -118935 44560 -118915
rect 45280 -118935 46060 -118915
rect 46780 -118935 47560 -118915
rect 48280 -118935 49060 -118915
rect 49780 -118935 50560 -118915
rect 51280 -118935 52060 -118915
rect 52780 -118935 53560 -118915
rect 54280 -118935 55060 -118915
rect 55780 -118935 56560 -118915
rect 57280 -118935 58060 -118915
rect 58780 -118935 59560 -118915
rect 60280 -118935 61060 -118915
rect 61780 -118935 62560 -118915
rect 63280 -118935 64060 -118915
rect 64780 -118935 65560 -118915
rect 66280 -118935 67060 -118915
rect 67780 -118935 68560 -118915
rect 69280 -118935 70060 -118915
rect 70780 -118935 71560 -118915
rect 72280 -118935 73060 -118915
rect 73780 -118935 74560 -118915
rect 75280 -118935 76060 -118915
rect 76780 -118935 77560 -118915
rect 78280 -118935 79060 -118915
rect 79780 -118935 80560 -118915
rect 81280 -118935 82060 -118915
rect 82780 -118935 83560 -118915
rect 84280 -118935 85060 -118915
rect 85780 -118935 86560 -118915
rect 87280 -118935 88060 -118915
rect 88780 -118935 89560 -118915
rect 90280 -118935 91060 -118915
rect 91780 -118935 92560 -118915
rect 93280 -118935 94060 -118915
rect 94780 -118935 95560 -118915
rect 96280 -118935 97060 -118915
rect 97780 -118935 98560 -118915
rect 99280 -118935 100060 -118915
rect 100780 -118935 101560 -118915
rect 102280 -118935 103060 -118915
rect 103780 -118935 104560 -118915
rect 105280 -118935 106060 -118915
rect 106780 -118935 107560 -118915
rect 108280 -118935 109060 -118915
rect 109780 -118935 110560 -118915
rect 111280 -118935 112060 -118915
rect 112780 -118935 113560 -118915
rect 114280 -118935 115060 -118915
rect 115780 -118935 116560 -118915
rect 117280 -118935 118060 -118915
rect 118780 -118935 119560 -118915
<< poly >>
rect 255 -118745 270 -118700
rect 110 -118750 270 -118745
rect 110 -118850 120 -118750
rect 210 -118850 270 -118750
rect 110 -118855 270 -118850
rect 255 -118900 270 -118855
rect 1070 -118900 1085 -118700
rect 1755 -118745 1770 -118700
rect 1610 -118750 1770 -118745
rect 1610 -118850 1620 -118750
rect 1710 -118850 1770 -118750
rect 1610 -118855 1770 -118850
rect 1755 -118900 1770 -118855
rect 2570 -118900 2585 -118700
rect 3255 -118745 3270 -118700
rect 3110 -118750 3270 -118745
rect 3110 -118850 3120 -118750
rect 3210 -118850 3270 -118750
rect 3110 -118855 3270 -118850
rect 3255 -118900 3270 -118855
rect 4070 -118900 4085 -118700
rect 4755 -118745 4770 -118700
rect 4610 -118750 4770 -118745
rect 4610 -118850 4620 -118750
rect 4710 -118850 4770 -118750
rect 4610 -118855 4770 -118850
rect 4755 -118900 4770 -118855
rect 5570 -118900 5585 -118700
rect 6255 -118745 6270 -118700
rect 6110 -118750 6270 -118745
rect 6110 -118850 6120 -118750
rect 6210 -118850 6270 -118750
rect 6110 -118855 6270 -118850
rect 6255 -118900 6270 -118855
rect 7070 -118900 7085 -118700
rect 7755 -118745 7770 -118700
rect 7610 -118750 7770 -118745
rect 7610 -118850 7620 -118750
rect 7710 -118850 7770 -118750
rect 7610 -118855 7770 -118850
rect 7755 -118900 7770 -118855
rect 8570 -118900 8585 -118700
rect 9255 -118745 9270 -118700
rect 9110 -118750 9270 -118745
rect 9110 -118850 9120 -118750
rect 9210 -118850 9270 -118750
rect 9110 -118855 9270 -118850
rect 9255 -118900 9270 -118855
rect 10070 -118900 10085 -118700
rect 10755 -118745 10770 -118700
rect 10610 -118750 10770 -118745
rect 10610 -118850 10620 -118750
rect 10710 -118850 10770 -118750
rect 10610 -118855 10770 -118850
rect 10755 -118900 10770 -118855
rect 11570 -118900 11585 -118700
rect 12255 -118745 12270 -118700
rect 12110 -118750 12270 -118745
rect 12110 -118850 12120 -118750
rect 12210 -118850 12270 -118750
rect 12110 -118855 12270 -118850
rect 12255 -118900 12270 -118855
rect 13070 -118900 13085 -118700
rect 13755 -118745 13770 -118700
rect 13610 -118750 13770 -118745
rect 13610 -118850 13620 -118750
rect 13710 -118850 13770 -118750
rect 13610 -118855 13770 -118850
rect 13755 -118900 13770 -118855
rect 14570 -118900 14585 -118700
rect 15255 -118745 15270 -118700
rect 15110 -118750 15270 -118745
rect 15110 -118850 15120 -118750
rect 15210 -118850 15270 -118750
rect 15110 -118855 15270 -118850
rect 15255 -118900 15270 -118855
rect 16070 -118900 16085 -118700
rect 16755 -118745 16770 -118700
rect 16610 -118750 16770 -118745
rect 16610 -118850 16620 -118750
rect 16710 -118850 16770 -118750
rect 16610 -118855 16770 -118850
rect 16755 -118900 16770 -118855
rect 17570 -118900 17585 -118700
rect 18255 -118745 18270 -118700
rect 18110 -118750 18270 -118745
rect 18110 -118850 18120 -118750
rect 18210 -118850 18270 -118750
rect 18110 -118855 18270 -118850
rect 18255 -118900 18270 -118855
rect 19070 -118900 19085 -118700
rect 19755 -118745 19770 -118700
rect 19610 -118750 19770 -118745
rect 19610 -118850 19620 -118750
rect 19710 -118850 19770 -118750
rect 19610 -118855 19770 -118850
rect 19755 -118900 19770 -118855
rect 20570 -118900 20585 -118700
rect 21255 -118745 21270 -118700
rect 21110 -118750 21270 -118745
rect 21110 -118850 21120 -118750
rect 21210 -118850 21270 -118750
rect 21110 -118855 21270 -118850
rect 21255 -118900 21270 -118855
rect 22070 -118900 22085 -118700
rect 22755 -118745 22770 -118700
rect 22610 -118750 22770 -118745
rect 22610 -118850 22620 -118750
rect 22710 -118850 22770 -118750
rect 22610 -118855 22770 -118850
rect 22755 -118900 22770 -118855
rect 23570 -118900 23585 -118700
rect 24255 -118745 24270 -118700
rect 24110 -118750 24270 -118745
rect 24110 -118850 24120 -118750
rect 24210 -118850 24270 -118750
rect 24110 -118855 24270 -118850
rect 24255 -118900 24270 -118855
rect 25070 -118900 25085 -118700
rect 25755 -118745 25770 -118700
rect 25610 -118750 25770 -118745
rect 25610 -118850 25620 -118750
rect 25710 -118850 25770 -118750
rect 25610 -118855 25770 -118850
rect 25755 -118900 25770 -118855
rect 26570 -118900 26585 -118700
rect 27255 -118745 27270 -118700
rect 27110 -118750 27270 -118745
rect 27110 -118850 27120 -118750
rect 27210 -118850 27270 -118750
rect 27110 -118855 27270 -118850
rect 27255 -118900 27270 -118855
rect 28070 -118900 28085 -118700
rect 28755 -118745 28770 -118700
rect 28610 -118750 28770 -118745
rect 28610 -118850 28620 -118750
rect 28710 -118850 28770 -118750
rect 28610 -118855 28770 -118850
rect 28755 -118900 28770 -118855
rect 29570 -118900 29585 -118700
rect 30255 -118745 30270 -118700
rect 30110 -118750 30270 -118745
rect 30110 -118850 30120 -118750
rect 30210 -118850 30270 -118750
rect 30110 -118855 30270 -118850
rect 30255 -118900 30270 -118855
rect 31070 -118900 31085 -118700
rect 31755 -118745 31770 -118700
rect 31610 -118750 31770 -118745
rect 31610 -118850 31620 -118750
rect 31710 -118850 31770 -118750
rect 31610 -118855 31770 -118850
rect 31755 -118900 31770 -118855
rect 32570 -118900 32585 -118700
rect 33255 -118745 33270 -118700
rect 33110 -118750 33270 -118745
rect 33110 -118850 33120 -118750
rect 33210 -118850 33270 -118750
rect 33110 -118855 33270 -118850
rect 33255 -118900 33270 -118855
rect 34070 -118900 34085 -118700
rect 34755 -118745 34770 -118700
rect 34610 -118750 34770 -118745
rect 34610 -118850 34620 -118750
rect 34710 -118850 34770 -118750
rect 34610 -118855 34770 -118850
rect 34755 -118900 34770 -118855
rect 35570 -118900 35585 -118700
rect 36255 -118745 36270 -118700
rect 36110 -118750 36270 -118745
rect 36110 -118850 36120 -118750
rect 36210 -118850 36270 -118750
rect 36110 -118855 36270 -118850
rect 36255 -118900 36270 -118855
rect 37070 -118900 37085 -118700
rect 37755 -118745 37770 -118700
rect 37610 -118750 37770 -118745
rect 37610 -118850 37620 -118750
rect 37710 -118850 37770 -118750
rect 37610 -118855 37770 -118850
rect 37755 -118900 37770 -118855
rect 38570 -118900 38585 -118700
rect 39255 -118745 39270 -118700
rect 39110 -118750 39270 -118745
rect 39110 -118850 39120 -118750
rect 39210 -118850 39270 -118750
rect 39110 -118855 39270 -118850
rect 39255 -118900 39270 -118855
rect 40070 -118900 40085 -118700
rect 40755 -118745 40770 -118700
rect 40610 -118750 40770 -118745
rect 40610 -118850 40620 -118750
rect 40710 -118850 40770 -118750
rect 40610 -118855 40770 -118850
rect 40755 -118900 40770 -118855
rect 41570 -118900 41585 -118700
rect 42255 -118745 42270 -118700
rect 42110 -118750 42270 -118745
rect 42110 -118850 42120 -118750
rect 42210 -118850 42270 -118750
rect 42110 -118855 42270 -118850
rect 42255 -118900 42270 -118855
rect 43070 -118900 43085 -118700
rect 43755 -118745 43770 -118700
rect 43610 -118750 43770 -118745
rect 43610 -118850 43620 -118750
rect 43710 -118850 43770 -118750
rect 43610 -118855 43770 -118850
rect 43755 -118900 43770 -118855
rect 44570 -118900 44585 -118700
rect 45255 -118745 45270 -118700
rect 45110 -118750 45270 -118745
rect 45110 -118850 45120 -118750
rect 45210 -118850 45270 -118750
rect 45110 -118855 45270 -118850
rect 45255 -118900 45270 -118855
rect 46070 -118900 46085 -118700
rect 46755 -118745 46770 -118700
rect 46610 -118750 46770 -118745
rect 46610 -118850 46620 -118750
rect 46710 -118850 46770 -118750
rect 46610 -118855 46770 -118850
rect 46755 -118900 46770 -118855
rect 47570 -118900 47585 -118700
rect 48255 -118745 48270 -118700
rect 48110 -118750 48270 -118745
rect 48110 -118850 48120 -118750
rect 48210 -118850 48270 -118750
rect 48110 -118855 48270 -118850
rect 48255 -118900 48270 -118855
rect 49070 -118900 49085 -118700
rect 49755 -118745 49770 -118700
rect 49610 -118750 49770 -118745
rect 49610 -118850 49620 -118750
rect 49710 -118850 49770 -118750
rect 49610 -118855 49770 -118850
rect 49755 -118900 49770 -118855
rect 50570 -118900 50585 -118700
rect 51255 -118745 51270 -118700
rect 51110 -118750 51270 -118745
rect 51110 -118850 51120 -118750
rect 51210 -118850 51270 -118750
rect 51110 -118855 51270 -118850
rect 51255 -118900 51270 -118855
rect 52070 -118900 52085 -118700
rect 52755 -118745 52770 -118700
rect 52610 -118750 52770 -118745
rect 52610 -118850 52620 -118750
rect 52710 -118850 52770 -118750
rect 52610 -118855 52770 -118850
rect 52755 -118900 52770 -118855
rect 53570 -118900 53585 -118700
rect 54255 -118745 54270 -118700
rect 54110 -118750 54270 -118745
rect 54110 -118850 54120 -118750
rect 54210 -118850 54270 -118750
rect 54110 -118855 54270 -118850
rect 54255 -118900 54270 -118855
rect 55070 -118900 55085 -118700
rect 55755 -118745 55770 -118700
rect 55610 -118750 55770 -118745
rect 55610 -118850 55620 -118750
rect 55710 -118850 55770 -118750
rect 55610 -118855 55770 -118850
rect 55755 -118900 55770 -118855
rect 56570 -118900 56585 -118700
rect 57255 -118745 57270 -118700
rect 57110 -118750 57270 -118745
rect 57110 -118850 57120 -118750
rect 57210 -118850 57270 -118750
rect 57110 -118855 57270 -118850
rect 57255 -118900 57270 -118855
rect 58070 -118900 58085 -118700
rect 58755 -118745 58770 -118700
rect 58610 -118750 58770 -118745
rect 58610 -118850 58620 -118750
rect 58710 -118850 58770 -118750
rect 58610 -118855 58770 -118850
rect 58755 -118900 58770 -118855
rect 59570 -118900 59585 -118700
rect 60255 -118745 60270 -118700
rect 60110 -118750 60270 -118745
rect 60110 -118850 60120 -118750
rect 60210 -118850 60270 -118750
rect 60110 -118855 60270 -118850
rect 60255 -118900 60270 -118855
rect 61070 -118900 61085 -118700
rect 61755 -118745 61770 -118700
rect 61610 -118750 61770 -118745
rect 61610 -118850 61620 -118750
rect 61710 -118850 61770 -118750
rect 61610 -118855 61770 -118850
rect 61755 -118900 61770 -118855
rect 62570 -118900 62585 -118700
rect 63255 -118745 63270 -118700
rect 63110 -118750 63270 -118745
rect 63110 -118850 63120 -118750
rect 63210 -118850 63270 -118750
rect 63110 -118855 63270 -118850
rect 63255 -118900 63270 -118855
rect 64070 -118900 64085 -118700
rect 64755 -118745 64770 -118700
rect 64610 -118750 64770 -118745
rect 64610 -118850 64620 -118750
rect 64710 -118850 64770 -118750
rect 64610 -118855 64770 -118850
rect 64755 -118900 64770 -118855
rect 65570 -118900 65585 -118700
rect 66255 -118745 66270 -118700
rect 66110 -118750 66270 -118745
rect 66110 -118850 66120 -118750
rect 66210 -118850 66270 -118750
rect 66110 -118855 66270 -118850
rect 66255 -118900 66270 -118855
rect 67070 -118900 67085 -118700
rect 67755 -118745 67770 -118700
rect 67610 -118750 67770 -118745
rect 67610 -118850 67620 -118750
rect 67710 -118850 67770 -118750
rect 67610 -118855 67770 -118850
rect 67755 -118900 67770 -118855
rect 68570 -118900 68585 -118700
rect 69255 -118745 69270 -118700
rect 69110 -118750 69270 -118745
rect 69110 -118850 69120 -118750
rect 69210 -118850 69270 -118750
rect 69110 -118855 69270 -118850
rect 69255 -118900 69270 -118855
rect 70070 -118900 70085 -118700
rect 70755 -118745 70770 -118700
rect 70610 -118750 70770 -118745
rect 70610 -118850 70620 -118750
rect 70710 -118850 70770 -118750
rect 70610 -118855 70770 -118850
rect 70755 -118900 70770 -118855
rect 71570 -118900 71585 -118700
rect 72255 -118745 72270 -118700
rect 72110 -118750 72270 -118745
rect 72110 -118850 72120 -118750
rect 72210 -118850 72270 -118750
rect 72110 -118855 72270 -118850
rect 72255 -118900 72270 -118855
rect 73070 -118900 73085 -118700
rect 73755 -118745 73770 -118700
rect 73610 -118750 73770 -118745
rect 73610 -118850 73620 -118750
rect 73710 -118850 73770 -118750
rect 73610 -118855 73770 -118850
rect 73755 -118900 73770 -118855
rect 74570 -118900 74585 -118700
rect 75255 -118745 75270 -118700
rect 75110 -118750 75270 -118745
rect 75110 -118850 75120 -118750
rect 75210 -118850 75270 -118750
rect 75110 -118855 75270 -118850
rect 75255 -118900 75270 -118855
rect 76070 -118900 76085 -118700
rect 76755 -118745 76770 -118700
rect 76610 -118750 76770 -118745
rect 76610 -118850 76620 -118750
rect 76710 -118850 76770 -118750
rect 76610 -118855 76770 -118850
rect 76755 -118900 76770 -118855
rect 77570 -118900 77585 -118700
rect 78255 -118745 78270 -118700
rect 78110 -118750 78270 -118745
rect 78110 -118850 78120 -118750
rect 78210 -118850 78270 -118750
rect 78110 -118855 78270 -118850
rect 78255 -118900 78270 -118855
rect 79070 -118900 79085 -118700
rect 79755 -118745 79770 -118700
rect 79610 -118750 79770 -118745
rect 79610 -118850 79620 -118750
rect 79710 -118850 79770 -118750
rect 79610 -118855 79770 -118850
rect 79755 -118900 79770 -118855
rect 80570 -118900 80585 -118700
rect 81255 -118745 81270 -118700
rect 81110 -118750 81270 -118745
rect 81110 -118850 81120 -118750
rect 81210 -118850 81270 -118750
rect 81110 -118855 81270 -118850
rect 81255 -118900 81270 -118855
rect 82070 -118900 82085 -118700
rect 82755 -118745 82770 -118700
rect 82610 -118750 82770 -118745
rect 82610 -118850 82620 -118750
rect 82710 -118850 82770 -118750
rect 82610 -118855 82770 -118850
rect 82755 -118900 82770 -118855
rect 83570 -118900 83585 -118700
rect 84255 -118745 84270 -118700
rect 84110 -118750 84270 -118745
rect 84110 -118850 84120 -118750
rect 84210 -118850 84270 -118750
rect 84110 -118855 84270 -118850
rect 84255 -118900 84270 -118855
rect 85070 -118900 85085 -118700
rect 85755 -118745 85770 -118700
rect 85610 -118750 85770 -118745
rect 85610 -118850 85620 -118750
rect 85710 -118850 85770 -118750
rect 85610 -118855 85770 -118850
rect 85755 -118900 85770 -118855
rect 86570 -118900 86585 -118700
rect 87255 -118745 87270 -118700
rect 87110 -118750 87270 -118745
rect 87110 -118850 87120 -118750
rect 87210 -118850 87270 -118750
rect 87110 -118855 87270 -118850
rect 87255 -118900 87270 -118855
rect 88070 -118900 88085 -118700
rect 88755 -118745 88770 -118700
rect 88610 -118750 88770 -118745
rect 88610 -118850 88620 -118750
rect 88710 -118850 88770 -118750
rect 88610 -118855 88770 -118850
rect 88755 -118900 88770 -118855
rect 89570 -118900 89585 -118700
rect 90255 -118745 90270 -118700
rect 90110 -118750 90270 -118745
rect 90110 -118850 90120 -118750
rect 90210 -118850 90270 -118750
rect 90110 -118855 90270 -118850
rect 90255 -118900 90270 -118855
rect 91070 -118900 91085 -118700
rect 91755 -118745 91770 -118700
rect 91610 -118750 91770 -118745
rect 91610 -118850 91620 -118750
rect 91710 -118850 91770 -118750
rect 91610 -118855 91770 -118850
rect 91755 -118900 91770 -118855
rect 92570 -118900 92585 -118700
rect 93255 -118745 93270 -118700
rect 93110 -118750 93270 -118745
rect 93110 -118850 93120 -118750
rect 93210 -118850 93270 -118750
rect 93110 -118855 93270 -118850
rect 93255 -118900 93270 -118855
rect 94070 -118900 94085 -118700
rect 94755 -118745 94770 -118700
rect 94610 -118750 94770 -118745
rect 94610 -118850 94620 -118750
rect 94710 -118850 94770 -118750
rect 94610 -118855 94770 -118850
rect 94755 -118900 94770 -118855
rect 95570 -118900 95585 -118700
rect 96255 -118745 96270 -118700
rect 96110 -118750 96270 -118745
rect 96110 -118850 96120 -118750
rect 96210 -118850 96270 -118750
rect 96110 -118855 96270 -118850
rect 96255 -118900 96270 -118855
rect 97070 -118900 97085 -118700
rect 97755 -118745 97770 -118700
rect 97610 -118750 97770 -118745
rect 97610 -118850 97620 -118750
rect 97710 -118850 97770 -118750
rect 97610 -118855 97770 -118850
rect 97755 -118900 97770 -118855
rect 98570 -118900 98585 -118700
rect 99255 -118745 99270 -118700
rect 99110 -118750 99270 -118745
rect 99110 -118850 99120 -118750
rect 99210 -118850 99270 -118750
rect 99110 -118855 99270 -118850
rect 99255 -118900 99270 -118855
rect 100070 -118900 100085 -118700
rect 100755 -118745 100770 -118700
rect 100610 -118750 100770 -118745
rect 100610 -118850 100620 -118750
rect 100710 -118850 100770 -118750
rect 100610 -118855 100770 -118850
rect 100755 -118900 100770 -118855
rect 101570 -118900 101585 -118700
rect 102255 -118745 102270 -118700
rect 102110 -118750 102270 -118745
rect 102110 -118850 102120 -118750
rect 102210 -118850 102270 -118750
rect 102110 -118855 102270 -118850
rect 102255 -118900 102270 -118855
rect 103070 -118900 103085 -118700
rect 103755 -118745 103770 -118700
rect 103610 -118750 103770 -118745
rect 103610 -118850 103620 -118750
rect 103710 -118850 103770 -118750
rect 103610 -118855 103770 -118850
rect 103755 -118900 103770 -118855
rect 104570 -118900 104585 -118700
rect 105255 -118745 105270 -118700
rect 105110 -118750 105270 -118745
rect 105110 -118850 105120 -118750
rect 105210 -118850 105270 -118750
rect 105110 -118855 105270 -118850
rect 105255 -118900 105270 -118855
rect 106070 -118900 106085 -118700
rect 106755 -118745 106770 -118700
rect 106610 -118750 106770 -118745
rect 106610 -118850 106620 -118750
rect 106710 -118850 106770 -118750
rect 106610 -118855 106770 -118850
rect 106755 -118900 106770 -118855
rect 107570 -118900 107585 -118700
rect 108255 -118745 108270 -118700
rect 108110 -118750 108270 -118745
rect 108110 -118850 108120 -118750
rect 108210 -118850 108270 -118750
rect 108110 -118855 108270 -118850
rect 108255 -118900 108270 -118855
rect 109070 -118900 109085 -118700
rect 109755 -118745 109770 -118700
rect 109610 -118750 109770 -118745
rect 109610 -118850 109620 -118750
rect 109710 -118850 109770 -118750
rect 109610 -118855 109770 -118850
rect 109755 -118900 109770 -118855
rect 110570 -118900 110585 -118700
rect 111255 -118745 111270 -118700
rect 111110 -118750 111270 -118745
rect 111110 -118850 111120 -118750
rect 111210 -118850 111270 -118750
rect 111110 -118855 111270 -118850
rect 111255 -118900 111270 -118855
rect 112070 -118900 112085 -118700
rect 112755 -118745 112770 -118700
rect 112610 -118750 112770 -118745
rect 112610 -118850 112620 -118750
rect 112710 -118850 112770 -118750
rect 112610 -118855 112770 -118850
rect 112755 -118900 112770 -118855
rect 113570 -118900 113585 -118700
rect 114255 -118745 114270 -118700
rect 114110 -118750 114270 -118745
rect 114110 -118850 114120 -118750
rect 114210 -118850 114270 -118750
rect 114110 -118855 114270 -118850
rect 114255 -118900 114270 -118855
rect 115070 -118900 115085 -118700
rect 115755 -118745 115770 -118700
rect 115610 -118750 115770 -118745
rect 115610 -118850 115620 -118750
rect 115710 -118850 115770 -118750
rect 115610 -118855 115770 -118850
rect 115755 -118900 115770 -118855
rect 116570 -118900 116585 -118700
rect 117255 -118745 117270 -118700
rect 117110 -118750 117270 -118745
rect 117110 -118850 117120 -118750
rect 117210 -118850 117270 -118750
rect 117110 -118855 117270 -118850
rect 117255 -118900 117270 -118855
rect 118070 -118900 118085 -118700
rect 118755 -118745 118770 -118700
rect 118610 -118750 118770 -118745
rect 118610 -118850 118620 -118750
rect 118710 -118850 118770 -118750
rect 118610 -118855 118770 -118850
rect 118755 -118900 118770 -118855
rect 119570 -118900 119585 -118700
<< polycont >>
rect 120 -118850 210 -118750
rect 1620 -118850 1710 -118750
rect 3120 -118850 3210 -118750
rect 4620 -118850 4710 -118750
rect 6120 -118850 6210 -118750
rect 7620 -118850 7710 -118750
rect 9120 -118850 9210 -118750
rect 10620 -118850 10710 -118750
rect 12120 -118850 12210 -118750
rect 13620 -118850 13710 -118750
rect 15120 -118850 15210 -118750
rect 16620 -118850 16710 -118750
rect 18120 -118850 18210 -118750
rect 19620 -118850 19710 -118750
rect 21120 -118850 21210 -118750
rect 22620 -118850 22710 -118750
rect 24120 -118850 24210 -118750
rect 25620 -118850 25710 -118750
rect 27120 -118850 27210 -118750
rect 28620 -118850 28710 -118750
rect 30120 -118850 30210 -118750
rect 31620 -118850 31710 -118750
rect 33120 -118850 33210 -118750
rect 34620 -118850 34710 -118750
rect 36120 -118850 36210 -118750
rect 37620 -118850 37710 -118750
rect 39120 -118850 39210 -118750
rect 40620 -118850 40710 -118750
rect 42120 -118850 42210 -118750
rect 43620 -118850 43710 -118750
rect 45120 -118850 45210 -118750
rect 46620 -118850 46710 -118750
rect 48120 -118850 48210 -118750
rect 49620 -118850 49710 -118750
rect 51120 -118850 51210 -118750
rect 52620 -118850 52710 -118750
rect 54120 -118850 54210 -118750
rect 55620 -118850 55710 -118750
rect 57120 -118850 57210 -118750
rect 58620 -118850 58710 -118750
rect 60120 -118850 60210 -118750
rect 61620 -118850 61710 -118750
rect 63120 -118850 63210 -118750
rect 64620 -118850 64710 -118750
rect 66120 -118850 66210 -118750
rect 67620 -118850 67710 -118750
rect 69120 -118850 69210 -118750
rect 70620 -118850 70710 -118750
rect 72120 -118850 72210 -118750
rect 73620 -118850 73710 -118750
rect 75120 -118850 75210 -118750
rect 76620 -118850 76710 -118750
rect 78120 -118850 78210 -118750
rect 79620 -118850 79710 -118750
rect 81120 -118850 81210 -118750
rect 82620 -118850 82710 -118750
rect 84120 -118850 84210 -118750
rect 85620 -118850 85710 -118750
rect 87120 -118850 87210 -118750
rect 88620 -118850 88710 -118750
rect 90120 -118850 90210 -118750
rect 91620 -118850 91710 -118750
rect 93120 -118850 93210 -118750
rect 94620 -118850 94710 -118750
rect 96120 -118850 96210 -118750
rect 97620 -118850 97710 -118750
rect 99120 -118850 99210 -118750
rect 100620 -118850 100710 -118750
rect 102120 -118850 102210 -118750
rect 103620 -118850 103710 -118750
rect 105120 -118850 105210 -118750
rect 106620 -118850 106710 -118750
rect 108120 -118850 108210 -118750
rect 109620 -118850 109710 -118750
rect 111120 -118850 111210 -118750
rect 112620 -118850 112710 -118750
rect 114120 -118850 114210 -118750
rect 115620 -118850 115710 -118750
rect 117120 -118850 117210 -118750
rect 118620 -118850 118710 -118750
<< locali >>
rect 270 -118645 280 -118615
rect 1060 -118645 1070 -118615
rect 270 -118660 1070 -118645
rect 270 -118690 280 -118660
rect 1060 -118690 1070 -118660
rect 1770 -118645 1780 -118615
rect 2560 -118645 2570 -118615
rect 1770 -118660 2570 -118645
rect 1770 -118690 1780 -118660
rect 2560 -118690 2570 -118660
rect 3270 -118645 3280 -118615
rect 4060 -118645 4070 -118615
rect 3270 -118660 4070 -118645
rect 3270 -118690 3280 -118660
rect 4060 -118690 4070 -118660
rect 4770 -118645 4780 -118615
rect 5560 -118645 5570 -118615
rect 4770 -118660 5570 -118645
rect 4770 -118690 4780 -118660
rect 5560 -118690 5570 -118660
rect 6270 -118645 6280 -118615
rect 7060 -118645 7070 -118615
rect 6270 -118660 7070 -118645
rect 6270 -118690 6280 -118660
rect 7060 -118690 7070 -118660
rect 7770 -118645 7780 -118615
rect 8560 -118645 8570 -118615
rect 7770 -118660 8570 -118645
rect 7770 -118690 7780 -118660
rect 8560 -118690 8570 -118660
rect 9270 -118645 9280 -118615
rect 10060 -118645 10070 -118615
rect 9270 -118660 10070 -118645
rect 9270 -118690 9280 -118660
rect 10060 -118690 10070 -118660
rect 10770 -118645 10780 -118615
rect 11560 -118645 11570 -118615
rect 10770 -118660 11570 -118645
rect 10770 -118690 10780 -118660
rect 11560 -118690 11570 -118660
rect 12270 -118645 12280 -118615
rect 13060 -118645 13070 -118615
rect 12270 -118660 13070 -118645
rect 12270 -118690 12280 -118660
rect 13060 -118690 13070 -118660
rect 13770 -118645 13780 -118615
rect 14560 -118645 14570 -118615
rect 13770 -118660 14570 -118645
rect 13770 -118690 13780 -118660
rect 14560 -118690 14570 -118660
rect 15270 -118645 15280 -118615
rect 16060 -118645 16070 -118615
rect 15270 -118660 16070 -118645
rect 15270 -118690 15280 -118660
rect 16060 -118690 16070 -118660
rect 16770 -118645 16780 -118615
rect 17560 -118645 17570 -118615
rect 16770 -118660 17570 -118645
rect 16770 -118690 16780 -118660
rect 17560 -118690 17570 -118660
rect 18270 -118645 18280 -118615
rect 19060 -118645 19070 -118615
rect 18270 -118660 19070 -118645
rect 18270 -118690 18280 -118660
rect 19060 -118690 19070 -118660
rect 19770 -118645 19780 -118615
rect 20560 -118645 20570 -118615
rect 19770 -118660 20570 -118645
rect 19770 -118690 19780 -118660
rect 20560 -118690 20570 -118660
rect 21270 -118645 21280 -118615
rect 22060 -118645 22070 -118615
rect 21270 -118660 22070 -118645
rect 21270 -118690 21280 -118660
rect 22060 -118690 22070 -118660
rect 22770 -118645 22780 -118615
rect 23560 -118645 23570 -118615
rect 22770 -118660 23570 -118645
rect 22770 -118690 22780 -118660
rect 23560 -118690 23570 -118660
rect 24270 -118645 24280 -118615
rect 25060 -118645 25070 -118615
rect 24270 -118660 25070 -118645
rect 24270 -118690 24280 -118660
rect 25060 -118690 25070 -118660
rect 25770 -118645 25780 -118615
rect 26560 -118645 26570 -118615
rect 25770 -118660 26570 -118645
rect 25770 -118690 25780 -118660
rect 26560 -118690 26570 -118660
rect 27270 -118645 27280 -118615
rect 28060 -118645 28070 -118615
rect 27270 -118660 28070 -118645
rect 27270 -118690 27280 -118660
rect 28060 -118690 28070 -118660
rect 28770 -118645 28780 -118615
rect 29560 -118645 29570 -118615
rect 28770 -118660 29570 -118645
rect 28770 -118690 28780 -118660
rect 29560 -118690 29570 -118660
rect 30270 -118645 30280 -118615
rect 31060 -118645 31070 -118615
rect 30270 -118660 31070 -118645
rect 30270 -118690 30280 -118660
rect 31060 -118690 31070 -118660
rect 31770 -118645 31780 -118615
rect 32560 -118645 32570 -118615
rect 31770 -118660 32570 -118645
rect 31770 -118690 31780 -118660
rect 32560 -118690 32570 -118660
rect 33270 -118645 33280 -118615
rect 34060 -118645 34070 -118615
rect 33270 -118660 34070 -118645
rect 33270 -118690 33280 -118660
rect 34060 -118690 34070 -118660
rect 34770 -118645 34780 -118615
rect 35560 -118645 35570 -118615
rect 34770 -118660 35570 -118645
rect 34770 -118690 34780 -118660
rect 35560 -118690 35570 -118660
rect 36270 -118645 36280 -118615
rect 37060 -118645 37070 -118615
rect 36270 -118660 37070 -118645
rect 36270 -118690 36280 -118660
rect 37060 -118690 37070 -118660
rect 37770 -118645 37780 -118615
rect 38560 -118645 38570 -118615
rect 37770 -118660 38570 -118645
rect 37770 -118690 37780 -118660
rect 38560 -118690 38570 -118660
rect 39270 -118645 39280 -118615
rect 40060 -118645 40070 -118615
rect 39270 -118660 40070 -118645
rect 39270 -118690 39280 -118660
rect 40060 -118690 40070 -118660
rect 40770 -118645 40780 -118615
rect 41560 -118645 41570 -118615
rect 40770 -118660 41570 -118645
rect 40770 -118690 40780 -118660
rect 41560 -118690 41570 -118660
rect 42270 -118645 42280 -118615
rect 43060 -118645 43070 -118615
rect 42270 -118660 43070 -118645
rect 42270 -118690 42280 -118660
rect 43060 -118690 43070 -118660
rect 43770 -118645 43780 -118615
rect 44560 -118645 44570 -118615
rect 43770 -118660 44570 -118645
rect 43770 -118690 43780 -118660
rect 44560 -118690 44570 -118660
rect 45270 -118645 45280 -118615
rect 46060 -118645 46070 -118615
rect 45270 -118660 46070 -118645
rect 45270 -118690 45280 -118660
rect 46060 -118690 46070 -118660
rect 46770 -118645 46780 -118615
rect 47560 -118645 47570 -118615
rect 46770 -118660 47570 -118645
rect 46770 -118690 46780 -118660
rect 47560 -118690 47570 -118660
rect 48270 -118645 48280 -118615
rect 49060 -118645 49070 -118615
rect 48270 -118660 49070 -118645
rect 48270 -118690 48280 -118660
rect 49060 -118690 49070 -118660
rect 49770 -118645 49780 -118615
rect 50560 -118645 50570 -118615
rect 49770 -118660 50570 -118645
rect 49770 -118690 49780 -118660
rect 50560 -118690 50570 -118660
rect 51270 -118645 51280 -118615
rect 52060 -118645 52070 -118615
rect 51270 -118660 52070 -118645
rect 51270 -118690 51280 -118660
rect 52060 -118690 52070 -118660
rect 52770 -118645 52780 -118615
rect 53560 -118645 53570 -118615
rect 52770 -118660 53570 -118645
rect 52770 -118690 52780 -118660
rect 53560 -118690 53570 -118660
rect 54270 -118645 54280 -118615
rect 55060 -118645 55070 -118615
rect 54270 -118660 55070 -118645
rect 54270 -118690 54280 -118660
rect 55060 -118690 55070 -118660
rect 55770 -118645 55780 -118615
rect 56560 -118645 56570 -118615
rect 55770 -118660 56570 -118645
rect 55770 -118690 55780 -118660
rect 56560 -118690 56570 -118660
rect 57270 -118645 57280 -118615
rect 58060 -118645 58070 -118615
rect 57270 -118660 58070 -118645
rect 57270 -118690 57280 -118660
rect 58060 -118690 58070 -118660
rect 58770 -118645 58780 -118615
rect 59560 -118645 59570 -118615
rect 58770 -118660 59570 -118645
rect 58770 -118690 58780 -118660
rect 59560 -118690 59570 -118660
rect 60270 -118645 60280 -118615
rect 61060 -118645 61070 -118615
rect 60270 -118660 61070 -118645
rect 60270 -118690 60280 -118660
rect 61060 -118690 61070 -118660
rect 61770 -118645 61780 -118615
rect 62560 -118645 62570 -118615
rect 61770 -118660 62570 -118645
rect 61770 -118690 61780 -118660
rect 62560 -118690 62570 -118660
rect 63270 -118645 63280 -118615
rect 64060 -118645 64070 -118615
rect 63270 -118660 64070 -118645
rect 63270 -118690 63280 -118660
rect 64060 -118690 64070 -118660
rect 64770 -118645 64780 -118615
rect 65560 -118645 65570 -118615
rect 64770 -118660 65570 -118645
rect 64770 -118690 64780 -118660
rect 65560 -118690 65570 -118660
rect 66270 -118645 66280 -118615
rect 67060 -118645 67070 -118615
rect 66270 -118660 67070 -118645
rect 66270 -118690 66280 -118660
rect 67060 -118690 67070 -118660
rect 67770 -118645 67780 -118615
rect 68560 -118645 68570 -118615
rect 67770 -118660 68570 -118645
rect 67770 -118690 67780 -118660
rect 68560 -118690 68570 -118660
rect 69270 -118645 69280 -118615
rect 70060 -118645 70070 -118615
rect 69270 -118660 70070 -118645
rect 69270 -118690 69280 -118660
rect 70060 -118690 70070 -118660
rect 70770 -118645 70780 -118615
rect 71560 -118645 71570 -118615
rect 70770 -118660 71570 -118645
rect 70770 -118690 70780 -118660
rect 71560 -118690 71570 -118660
rect 72270 -118645 72280 -118615
rect 73060 -118645 73070 -118615
rect 72270 -118660 73070 -118645
rect 72270 -118690 72280 -118660
rect 73060 -118690 73070 -118660
rect 73770 -118645 73780 -118615
rect 74560 -118645 74570 -118615
rect 73770 -118660 74570 -118645
rect 73770 -118690 73780 -118660
rect 74560 -118690 74570 -118660
rect 75270 -118645 75280 -118615
rect 76060 -118645 76070 -118615
rect 75270 -118660 76070 -118645
rect 75270 -118690 75280 -118660
rect 76060 -118690 76070 -118660
rect 76770 -118645 76780 -118615
rect 77560 -118645 77570 -118615
rect 76770 -118660 77570 -118645
rect 76770 -118690 76780 -118660
rect 77560 -118690 77570 -118660
rect 78270 -118645 78280 -118615
rect 79060 -118645 79070 -118615
rect 78270 -118660 79070 -118645
rect 78270 -118690 78280 -118660
rect 79060 -118690 79070 -118660
rect 79770 -118645 79780 -118615
rect 80560 -118645 80570 -118615
rect 79770 -118660 80570 -118645
rect 79770 -118690 79780 -118660
rect 80560 -118690 80570 -118660
rect 81270 -118645 81280 -118615
rect 82060 -118645 82070 -118615
rect 81270 -118660 82070 -118645
rect 81270 -118690 81280 -118660
rect 82060 -118690 82070 -118660
rect 82770 -118645 82780 -118615
rect 83560 -118645 83570 -118615
rect 82770 -118660 83570 -118645
rect 82770 -118690 82780 -118660
rect 83560 -118690 83570 -118660
rect 84270 -118645 84280 -118615
rect 85060 -118645 85070 -118615
rect 84270 -118660 85070 -118645
rect 84270 -118690 84280 -118660
rect 85060 -118690 85070 -118660
rect 85770 -118645 85780 -118615
rect 86560 -118645 86570 -118615
rect 85770 -118660 86570 -118645
rect 85770 -118690 85780 -118660
rect 86560 -118690 86570 -118660
rect 87270 -118645 87280 -118615
rect 88060 -118645 88070 -118615
rect 87270 -118660 88070 -118645
rect 87270 -118690 87280 -118660
rect 88060 -118690 88070 -118660
rect 88770 -118645 88780 -118615
rect 89560 -118645 89570 -118615
rect 88770 -118660 89570 -118645
rect 88770 -118690 88780 -118660
rect 89560 -118690 89570 -118660
rect 90270 -118645 90280 -118615
rect 91060 -118645 91070 -118615
rect 90270 -118660 91070 -118645
rect 90270 -118690 90280 -118660
rect 91060 -118690 91070 -118660
rect 91770 -118645 91780 -118615
rect 92560 -118645 92570 -118615
rect 91770 -118660 92570 -118645
rect 91770 -118690 91780 -118660
rect 92560 -118690 92570 -118660
rect 93270 -118645 93280 -118615
rect 94060 -118645 94070 -118615
rect 93270 -118660 94070 -118645
rect 93270 -118690 93280 -118660
rect 94060 -118690 94070 -118660
rect 94770 -118645 94780 -118615
rect 95560 -118645 95570 -118615
rect 94770 -118660 95570 -118645
rect 94770 -118690 94780 -118660
rect 95560 -118690 95570 -118660
rect 96270 -118645 96280 -118615
rect 97060 -118645 97070 -118615
rect 96270 -118660 97070 -118645
rect 96270 -118690 96280 -118660
rect 97060 -118690 97070 -118660
rect 97770 -118645 97780 -118615
rect 98560 -118645 98570 -118615
rect 97770 -118660 98570 -118645
rect 97770 -118690 97780 -118660
rect 98560 -118690 98570 -118660
rect 99270 -118645 99280 -118615
rect 100060 -118645 100070 -118615
rect 99270 -118660 100070 -118645
rect 99270 -118690 99280 -118660
rect 100060 -118690 100070 -118660
rect 100770 -118645 100780 -118615
rect 101560 -118645 101570 -118615
rect 100770 -118660 101570 -118645
rect 100770 -118690 100780 -118660
rect 101560 -118690 101570 -118660
rect 102270 -118645 102280 -118615
rect 103060 -118645 103070 -118615
rect 102270 -118660 103070 -118645
rect 102270 -118690 102280 -118660
rect 103060 -118690 103070 -118660
rect 103770 -118645 103780 -118615
rect 104560 -118645 104570 -118615
rect 103770 -118660 104570 -118645
rect 103770 -118690 103780 -118660
rect 104560 -118690 104570 -118660
rect 105270 -118645 105280 -118615
rect 106060 -118645 106070 -118615
rect 105270 -118660 106070 -118645
rect 105270 -118690 105280 -118660
rect 106060 -118690 106070 -118660
rect 106770 -118645 106780 -118615
rect 107560 -118645 107570 -118615
rect 106770 -118660 107570 -118645
rect 106770 -118690 106780 -118660
rect 107560 -118690 107570 -118660
rect 108270 -118645 108280 -118615
rect 109060 -118645 109070 -118615
rect 108270 -118660 109070 -118645
rect 108270 -118690 108280 -118660
rect 109060 -118690 109070 -118660
rect 109770 -118645 109780 -118615
rect 110560 -118645 110570 -118615
rect 109770 -118660 110570 -118645
rect 109770 -118690 109780 -118660
rect 110560 -118690 110570 -118660
rect 111270 -118645 111280 -118615
rect 112060 -118645 112070 -118615
rect 111270 -118660 112070 -118645
rect 111270 -118690 111280 -118660
rect 112060 -118690 112070 -118660
rect 112770 -118645 112780 -118615
rect 113560 -118645 113570 -118615
rect 112770 -118660 113570 -118645
rect 112770 -118690 112780 -118660
rect 113560 -118690 113570 -118660
rect 114270 -118645 114280 -118615
rect 115060 -118645 115070 -118615
rect 114270 -118660 115070 -118645
rect 114270 -118690 114280 -118660
rect 115060 -118690 115070 -118660
rect 115770 -118645 115780 -118615
rect 116560 -118645 116570 -118615
rect 115770 -118660 116570 -118645
rect 115770 -118690 115780 -118660
rect 116560 -118690 116570 -118660
rect 117270 -118645 117280 -118615
rect 118060 -118645 118070 -118615
rect 117270 -118660 118070 -118645
rect 117270 -118690 117280 -118660
rect 118060 -118690 118070 -118660
rect 118770 -118645 118780 -118615
rect 119560 -118645 119570 -118615
rect 118770 -118660 119570 -118645
rect 118770 -118690 118780 -118660
rect 119560 -118690 119570 -118660
rect 110 -118750 220 -118745
rect 110 -118850 120 -118750
rect 210 -118850 220 -118750
rect 110 -118855 220 -118850
rect 1610 -118750 1720 -118745
rect 1610 -118850 1620 -118750
rect 1710 -118850 1720 -118750
rect 1610 -118855 1720 -118850
rect 3110 -118750 3220 -118745
rect 3110 -118850 3120 -118750
rect 3210 -118850 3220 -118750
rect 3110 -118855 3220 -118850
rect 4610 -118750 4720 -118745
rect 4610 -118850 4620 -118750
rect 4710 -118850 4720 -118750
rect 4610 -118855 4720 -118850
rect 6110 -118750 6220 -118745
rect 6110 -118850 6120 -118750
rect 6210 -118850 6220 -118750
rect 6110 -118855 6220 -118850
rect 7610 -118750 7720 -118745
rect 7610 -118850 7620 -118750
rect 7710 -118850 7720 -118750
rect 7610 -118855 7720 -118850
rect 9110 -118750 9220 -118745
rect 9110 -118850 9120 -118750
rect 9210 -118850 9220 -118750
rect 9110 -118855 9220 -118850
rect 10610 -118750 10720 -118745
rect 10610 -118850 10620 -118750
rect 10710 -118850 10720 -118750
rect 10610 -118855 10720 -118850
rect 12110 -118750 12220 -118745
rect 12110 -118850 12120 -118750
rect 12210 -118850 12220 -118750
rect 12110 -118855 12220 -118850
rect 13610 -118750 13720 -118745
rect 13610 -118850 13620 -118750
rect 13710 -118850 13720 -118750
rect 13610 -118855 13720 -118850
rect 15110 -118750 15220 -118745
rect 15110 -118850 15120 -118750
rect 15210 -118850 15220 -118750
rect 15110 -118855 15220 -118850
rect 16610 -118750 16720 -118745
rect 16610 -118850 16620 -118750
rect 16710 -118850 16720 -118750
rect 16610 -118855 16720 -118850
rect 18110 -118750 18220 -118745
rect 18110 -118850 18120 -118750
rect 18210 -118850 18220 -118750
rect 18110 -118855 18220 -118850
rect 19610 -118750 19720 -118745
rect 19610 -118850 19620 -118750
rect 19710 -118850 19720 -118750
rect 19610 -118855 19720 -118850
rect 21110 -118750 21220 -118745
rect 21110 -118850 21120 -118750
rect 21210 -118850 21220 -118750
rect 21110 -118855 21220 -118850
rect 22610 -118750 22720 -118745
rect 22610 -118850 22620 -118750
rect 22710 -118850 22720 -118750
rect 22610 -118855 22720 -118850
rect 24110 -118750 24220 -118745
rect 24110 -118850 24120 -118750
rect 24210 -118850 24220 -118750
rect 24110 -118855 24220 -118850
rect 25610 -118750 25720 -118745
rect 25610 -118850 25620 -118750
rect 25710 -118850 25720 -118750
rect 25610 -118855 25720 -118850
rect 27110 -118750 27220 -118745
rect 27110 -118850 27120 -118750
rect 27210 -118850 27220 -118750
rect 27110 -118855 27220 -118850
rect 28610 -118750 28720 -118745
rect 28610 -118850 28620 -118750
rect 28710 -118850 28720 -118750
rect 28610 -118855 28720 -118850
rect 30110 -118750 30220 -118745
rect 30110 -118850 30120 -118750
rect 30210 -118850 30220 -118750
rect 30110 -118855 30220 -118850
rect 31610 -118750 31720 -118745
rect 31610 -118850 31620 -118750
rect 31710 -118850 31720 -118750
rect 31610 -118855 31720 -118850
rect 33110 -118750 33220 -118745
rect 33110 -118850 33120 -118750
rect 33210 -118850 33220 -118750
rect 33110 -118855 33220 -118850
rect 34610 -118750 34720 -118745
rect 34610 -118850 34620 -118750
rect 34710 -118850 34720 -118750
rect 34610 -118855 34720 -118850
rect 36110 -118750 36220 -118745
rect 36110 -118850 36120 -118750
rect 36210 -118850 36220 -118750
rect 36110 -118855 36220 -118850
rect 37610 -118750 37720 -118745
rect 37610 -118850 37620 -118750
rect 37710 -118850 37720 -118750
rect 37610 -118855 37720 -118850
rect 39110 -118750 39220 -118745
rect 39110 -118850 39120 -118750
rect 39210 -118850 39220 -118750
rect 39110 -118855 39220 -118850
rect 40610 -118750 40720 -118745
rect 40610 -118850 40620 -118750
rect 40710 -118850 40720 -118750
rect 40610 -118855 40720 -118850
rect 42110 -118750 42220 -118745
rect 42110 -118850 42120 -118750
rect 42210 -118850 42220 -118750
rect 42110 -118855 42220 -118850
rect 43610 -118750 43720 -118745
rect 43610 -118850 43620 -118750
rect 43710 -118850 43720 -118750
rect 43610 -118855 43720 -118850
rect 45110 -118750 45220 -118745
rect 45110 -118850 45120 -118750
rect 45210 -118850 45220 -118750
rect 45110 -118855 45220 -118850
rect 46610 -118750 46720 -118745
rect 46610 -118850 46620 -118750
rect 46710 -118850 46720 -118750
rect 46610 -118855 46720 -118850
rect 48110 -118750 48220 -118745
rect 48110 -118850 48120 -118750
rect 48210 -118850 48220 -118750
rect 48110 -118855 48220 -118850
rect 49610 -118750 49720 -118745
rect 49610 -118850 49620 -118750
rect 49710 -118850 49720 -118750
rect 49610 -118855 49720 -118850
rect 51110 -118750 51220 -118745
rect 51110 -118850 51120 -118750
rect 51210 -118850 51220 -118750
rect 51110 -118855 51220 -118850
rect 52610 -118750 52720 -118745
rect 52610 -118850 52620 -118750
rect 52710 -118850 52720 -118750
rect 52610 -118855 52720 -118850
rect 54110 -118750 54220 -118745
rect 54110 -118850 54120 -118750
rect 54210 -118850 54220 -118750
rect 54110 -118855 54220 -118850
rect 55610 -118750 55720 -118745
rect 55610 -118850 55620 -118750
rect 55710 -118850 55720 -118750
rect 55610 -118855 55720 -118850
rect 57110 -118750 57220 -118745
rect 57110 -118850 57120 -118750
rect 57210 -118850 57220 -118750
rect 57110 -118855 57220 -118850
rect 58610 -118750 58720 -118745
rect 58610 -118850 58620 -118750
rect 58710 -118850 58720 -118750
rect 58610 -118855 58720 -118850
rect 60110 -118750 60220 -118745
rect 60110 -118850 60120 -118750
rect 60210 -118850 60220 -118750
rect 60110 -118855 60220 -118850
rect 61610 -118750 61720 -118745
rect 61610 -118850 61620 -118750
rect 61710 -118850 61720 -118750
rect 61610 -118855 61720 -118850
rect 63110 -118750 63220 -118745
rect 63110 -118850 63120 -118750
rect 63210 -118850 63220 -118750
rect 63110 -118855 63220 -118850
rect 64610 -118750 64720 -118745
rect 64610 -118850 64620 -118750
rect 64710 -118850 64720 -118750
rect 64610 -118855 64720 -118850
rect 66110 -118750 66220 -118745
rect 66110 -118850 66120 -118750
rect 66210 -118850 66220 -118750
rect 66110 -118855 66220 -118850
rect 67610 -118750 67720 -118745
rect 67610 -118850 67620 -118750
rect 67710 -118850 67720 -118750
rect 67610 -118855 67720 -118850
rect 69110 -118750 69220 -118745
rect 69110 -118850 69120 -118750
rect 69210 -118850 69220 -118750
rect 69110 -118855 69220 -118850
rect 70610 -118750 70720 -118745
rect 70610 -118850 70620 -118750
rect 70710 -118850 70720 -118750
rect 70610 -118855 70720 -118850
rect 72110 -118750 72220 -118745
rect 72110 -118850 72120 -118750
rect 72210 -118850 72220 -118750
rect 72110 -118855 72220 -118850
rect 73610 -118750 73720 -118745
rect 73610 -118850 73620 -118750
rect 73710 -118850 73720 -118750
rect 73610 -118855 73720 -118850
rect 75110 -118750 75220 -118745
rect 75110 -118850 75120 -118750
rect 75210 -118850 75220 -118750
rect 75110 -118855 75220 -118850
rect 76610 -118750 76720 -118745
rect 76610 -118850 76620 -118750
rect 76710 -118850 76720 -118750
rect 76610 -118855 76720 -118850
rect 78110 -118750 78220 -118745
rect 78110 -118850 78120 -118750
rect 78210 -118850 78220 -118750
rect 78110 -118855 78220 -118850
rect 79610 -118750 79720 -118745
rect 79610 -118850 79620 -118750
rect 79710 -118850 79720 -118750
rect 79610 -118855 79720 -118850
rect 81110 -118750 81220 -118745
rect 81110 -118850 81120 -118750
rect 81210 -118850 81220 -118750
rect 81110 -118855 81220 -118850
rect 82610 -118750 82720 -118745
rect 82610 -118850 82620 -118750
rect 82710 -118850 82720 -118750
rect 82610 -118855 82720 -118850
rect 84110 -118750 84220 -118745
rect 84110 -118850 84120 -118750
rect 84210 -118850 84220 -118750
rect 84110 -118855 84220 -118850
rect 85610 -118750 85720 -118745
rect 85610 -118850 85620 -118750
rect 85710 -118850 85720 -118750
rect 85610 -118855 85720 -118850
rect 87110 -118750 87220 -118745
rect 87110 -118850 87120 -118750
rect 87210 -118850 87220 -118750
rect 87110 -118855 87220 -118850
rect 88610 -118750 88720 -118745
rect 88610 -118850 88620 -118750
rect 88710 -118850 88720 -118750
rect 88610 -118855 88720 -118850
rect 90110 -118750 90220 -118745
rect 90110 -118850 90120 -118750
rect 90210 -118850 90220 -118750
rect 90110 -118855 90220 -118850
rect 91610 -118750 91720 -118745
rect 91610 -118850 91620 -118750
rect 91710 -118850 91720 -118750
rect 91610 -118855 91720 -118850
rect 93110 -118750 93220 -118745
rect 93110 -118850 93120 -118750
rect 93210 -118850 93220 -118750
rect 93110 -118855 93220 -118850
rect 94610 -118750 94720 -118745
rect 94610 -118850 94620 -118750
rect 94710 -118850 94720 -118750
rect 94610 -118855 94720 -118850
rect 96110 -118750 96220 -118745
rect 96110 -118850 96120 -118750
rect 96210 -118850 96220 -118750
rect 96110 -118855 96220 -118850
rect 97610 -118750 97720 -118745
rect 97610 -118850 97620 -118750
rect 97710 -118850 97720 -118750
rect 97610 -118855 97720 -118850
rect 99110 -118750 99220 -118745
rect 99110 -118850 99120 -118750
rect 99210 -118850 99220 -118750
rect 99110 -118855 99220 -118850
rect 100610 -118750 100720 -118745
rect 100610 -118850 100620 -118750
rect 100710 -118850 100720 -118750
rect 100610 -118855 100720 -118850
rect 102110 -118750 102220 -118745
rect 102110 -118850 102120 -118750
rect 102210 -118850 102220 -118750
rect 102110 -118855 102220 -118850
rect 103610 -118750 103720 -118745
rect 103610 -118850 103620 -118750
rect 103710 -118850 103720 -118750
rect 103610 -118855 103720 -118850
rect 105110 -118750 105220 -118745
rect 105110 -118850 105120 -118750
rect 105210 -118850 105220 -118750
rect 105110 -118855 105220 -118850
rect 106610 -118750 106720 -118745
rect 106610 -118850 106620 -118750
rect 106710 -118850 106720 -118750
rect 106610 -118855 106720 -118850
rect 108110 -118750 108220 -118745
rect 108110 -118850 108120 -118750
rect 108210 -118850 108220 -118750
rect 108110 -118855 108220 -118850
rect 109610 -118750 109720 -118745
rect 109610 -118850 109620 -118750
rect 109710 -118850 109720 -118750
rect 109610 -118855 109720 -118850
rect 111110 -118750 111220 -118745
rect 111110 -118850 111120 -118750
rect 111210 -118850 111220 -118750
rect 111110 -118855 111220 -118850
rect 112610 -118750 112720 -118745
rect 112610 -118850 112620 -118750
rect 112710 -118850 112720 -118750
rect 112610 -118855 112720 -118850
rect 114110 -118750 114220 -118745
rect 114110 -118850 114120 -118750
rect 114210 -118850 114220 -118750
rect 114110 -118855 114220 -118850
rect 115610 -118750 115720 -118745
rect 115610 -118850 115620 -118750
rect 115710 -118850 115720 -118750
rect 115610 -118855 115720 -118850
rect 117110 -118750 117220 -118745
rect 117110 -118850 117120 -118750
rect 117210 -118850 117220 -118750
rect 117110 -118855 117220 -118850
rect 118610 -118750 118720 -118745
rect 118610 -118850 118620 -118750
rect 118710 -118850 118720 -118750
rect 118610 -118855 118720 -118850
rect 270 -118915 1070 -118900
rect 270 -118935 280 -118915
rect 1060 -118935 1070 -118915
rect 270 -118960 1070 -118935
rect 270 -118990 280 -118960
rect 1060 -118990 1070 -118960
rect 270 -119000 1070 -118990
rect 1770 -118915 2570 -118900
rect 1770 -118935 1780 -118915
rect 2560 -118935 2570 -118915
rect 1770 -118960 2570 -118935
rect 1770 -118990 1780 -118960
rect 2560 -118990 2570 -118960
rect 1770 -119000 2570 -118990
rect 3270 -118915 4070 -118900
rect 3270 -118935 3280 -118915
rect 4060 -118935 4070 -118915
rect 3270 -118960 4070 -118935
rect 3270 -118990 3280 -118960
rect 4060 -118990 4070 -118960
rect 3270 -119000 4070 -118990
rect 4770 -118915 5570 -118900
rect 4770 -118935 4780 -118915
rect 5560 -118935 5570 -118915
rect 4770 -118960 5570 -118935
rect 4770 -118990 4780 -118960
rect 5560 -118990 5570 -118960
rect 4770 -119000 5570 -118990
rect 6270 -118915 7070 -118900
rect 6270 -118935 6280 -118915
rect 7060 -118935 7070 -118915
rect 6270 -118960 7070 -118935
rect 6270 -118990 6280 -118960
rect 7060 -118990 7070 -118960
rect 6270 -119000 7070 -118990
rect 7770 -118915 8570 -118900
rect 7770 -118935 7780 -118915
rect 8560 -118935 8570 -118915
rect 7770 -118960 8570 -118935
rect 7770 -118990 7780 -118960
rect 8560 -118990 8570 -118960
rect 7770 -119000 8570 -118990
rect 9270 -118915 10070 -118900
rect 9270 -118935 9280 -118915
rect 10060 -118935 10070 -118915
rect 9270 -118960 10070 -118935
rect 9270 -118990 9280 -118960
rect 10060 -118990 10070 -118960
rect 9270 -119000 10070 -118990
rect 10770 -118915 11570 -118900
rect 10770 -118935 10780 -118915
rect 11560 -118935 11570 -118915
rect 10770 -118960 11570 -118935
rect 10770 -118990 10780 -118960
rect 11560 -118990 11570 -118960
rect 10770 -119000 11570 -118990
rect 12270 -118915 13070 -118900
rect 12270 -118935 12280 -118915
rect 13060 -118935 13070 -118915
rect 12270 -118960 13070 -118935
rect 12270 -118990 12280 -118960
rect 13060 -118990 13070 -118960
rect 12270 -119000 13070 -118990
rect 13770 -118915 14570 -118900
rect 13770 -118935 13780 -118915
rect 14560 -118935 14570 -118915
rect 13770 -118960 14570 -118935
rect 13770 -118990 13780 -118960
rect 14560 -118990 14570 -118960
rect 13770 -119000 14570 -118990
rect 15270 -118915 16070 -118900
rect 15270 -118935 15280 -118915
rect 16060 -118935 16070 -118915
rect 15270 -118960 16070 -118935
rect 15270 -118990 15280 -118960
rect 16060 -118990 16070 -118960
rect 15270 -119000 16070 -118990
rect 16770 -118915 17570 -118900
rect 16770 -118935 16780 -118915
rect 17560 -118935 17570 -118915
rect 16770 -118960 17570 -118935
rect 16770 -118990 16780 -118960
rect 17560 -118990 17570 -118960
rect 16770 -119000 17570 -118990
rect 18270 -118915 19070 -118900
rect 18270 -118935 18280 -118915
rect 19060 -118935 19070 -118915
rect 18270 -118960 19070 -118935
rect 18270 -118990 18280 -118960
rect 19060 -118990 19070 -118960
rect 18270 -119000 19070 -118990
rect 19770 -118915 20570 -118900
rect 19770 -118935 19780 -118915
rect 20560 -118935 20570 -118915
rect 19770 -118960 20570 -118935
rect 19770 -118990 19780 -118960
rect 20560 -118990 20570 -118960
rect 19770 -119000 20570 -118990
rect 21270 -118915 22070 -118900
rect 21270 -118935 21280 -118915
rect 22060 -118935 22070 -118915
rect 21270 -118960 22070 -118935
rect 21270 -118990 21280 -118960
rect 22060 -118990 22070 -118960
rect 21270 -119000 22070 -118990
rect 22770 -118915 23570 -118900
rect 22770 -118935 22780 -118915
rect 23560 -118935 23570 -118915
rect 22770 -118960 23570 -118935
rect 22770 -118990 22780 -118960
rect 23560 -118990 23570 -118960
rect 22770 -119000 23570 -118990
rect 24270 -118915 25070 -118900
rect 24270 -118935 24280 -118915
rect 25060 -118935 25070 -118915
rect 24270 -118960 25070 -118935
rect 24270 -118990 24280 -118960
rect 25060 -118990 25070 -118960
rect 24270 -119000 25070 -118990
rect 25770 -118915 26570 -118900
rect 25770 -118935 25780 -118915
rect 26560 -118935 26570 -118915
rect 25770 -118960 26570 -118935
rect 25770 -118990 25780 -118960
rect 26560 -118990 26570 -118960
rect 25770 -119000 26570 -118990
rect 27270 -118915 28070 -118900
rect 27270 -118935 27280 -118915
rect 28060 -118935 28070 -118915
rect 27270 -118960 28070 -118935
rect 27270 -118990 27280 -118960
rect 28060 -118990 28070 -118960
rect 27270 -119000 28070 -118990
rect 28770 -118915 29570 -118900
rect 28770 -118935 28780 -118915
rect 29560 -118935 29570 -118915
rect 28770 -118960 29570 -118935
rect 28770 -118990 28780 -118960
rect 29560 -118990 29570 -118960
rect 28770 -119000 29570 -118990
rect 30270 -118915 31070 -118900
rect 30270 -118935 30280 -118915
rect 31060 -118935 31070 -118915
rect 30270 -118960 31070 -118935
rect 30270 -118990 30280 -118960
rect 31060 -118990 31070 -118960
rect 30270 -119000 31070 -118990
rect 31770 -118915 32570 -118900
rect 31770 -118935 31780 -118915
rect 32560 -118935 32570 -118915
rect 31770 -118960 32570 -118935
rect 31770 -118990 31780 -118960
rect 32560 -118990 32570 -118960
rect 31770 -119000 32570 -118990
rect 33270 -118915 34070 -118900
rect 33270 -118935 33280 -118915
rect 34060 -118935 34070 -118915
rect 33270 -118960 34070 -118935
rect 33270 -118990 33280 -118960
rect 34060 -118990 34070 -118960
rect 33270 -119000 34070 -118990
rect 34770 -118915 35570 -118900
rect 34770 -118935 34780 -118915
rect 35560 -118935 35570 -118915
rect 34770 -118960 35570 -118935
rect 34770 -118990 34780 -118960
rect 35560 -118990 35570 -118960
rect 34770 -119000 35570 -118990
rect 36270 -118915 37070 -118900
rect 36270 -118935 36280 -118915
rect 37060 -118935 37070 -118915
rect 36270 -118960 37070 -118935
rect 36270 -118990 36280 -118960
rect 37060 -118990 37070 -118960
rect 36270 -119000 37070 -118990
rect 37770 -118915 38570 -118900
rect 37770 -118935 37780 -118915
rect 38560 -118935 38570 -118915
rect 37770 -118960 38570 -118935
rect 37770 -118990 37780 -118960
rect 38560 -118990 38570 -118960
rect 37770 -119000 38570 -118990
rect 39270 -118915 40070 -118900
rect 39270 -118935 39280 -118915
rect 40060 -118935 40070 -118915
rect 39270 -118960 40070 -118935
rect 39270 -118990 39280 -118960
rect 40060 -118990 40070 -118960
rect 39270 -119000 40070 -118990
rect 40770 -118915 41570 -118900
rect 40770 -118935 40780 -118915
rect 41560 -118935 41570 -118915
rect 40770 -118960 41570 -118935
rect 40770 -118990 40780 -118960
rect 41560 -118990 41570 -118960
rect 40770 -119000 41570 -118990
rect 42270 -118915 43070 -118900
rect 42270 -118935 42280 -118915
rect 43060 -118935 43070 -118915
rect 42270 -118960 43070 -118935
rect 42270 -118990 42280 -118960
rect 43060 -118990 43070 -118960
rect 42270 -119000 43070 -118990
rect 43770 -118915 44570 -118900
rect 43770 -118935 43780 -118915
rect 44560 -118935 44570 -118915
rect 43770 -118960 44570 -118935
rect 43770 -118990 43780 -118960
rect 44560 -118990 44570 -118960
rect 43770 -119000 44570 -118990
rect 45270 -118915 46070 -118900
rect 45270 -118935 45280 -118915
rect 46060 -118935 46070 -118915
rect 45270 -118960 46070 -118935
rect 45270 -118990 45280 -118960
rect 46060 -118990 46070 -118960
rect 45270 -119000 46070 -118990
rect 46770 -118915 47570 -118900
rect 46770 -118935 46780 -118915
rect 47560 -118935 47570 -118915
rect 46770 -118960 47570 -118935
rect 46770 -118990 46780 -118960
rect 47560 -118990 47570 -118960
rect 46770 -119000 47570 -118990
rect 48270 -118915 49070 -118900
rect 48270 -118935 48280 -118915
rect 49060 -118935 49070 -118915
rect 48270 -118960 49070 -118935
rect 48270 -118990 48280 -118960
rect 49060 -118990 49070 -118960
rect 48270 -119000 49070 -118990
rect 49770 -118915 50570 -118900
rect 49770 -118935 49780 -118915
rect 50560 -118935 50570 -118915
rect 49770 -118960 50570 -118935
rect 49770 -118990 49780 -118960
rect 50560 -118990 50570 -118960
rect 49770 -119000 50570 -118990
rect 51270 -118915 52070 -118900
rect 51270 -118935 51280 -118915
rect 52060 -118935 52070 -118915
rect 51270 -118960 52070 -118935
rect 51270 -118990 51280 -118960
rect 52060 -118990 52070 -118960
rect 51270 -119000 52070 -118990
rect 52770 -118915 53570 -118900
rect 52770 -118935 52780 -118915
rect 53560 -118935 53570 -118915
rect 52770 -118960 53570 -118935
rect 52770 -118990 52780 -118960
rect 53560 -118990 53570 -118960
rect 52770 -119000 53570 -118990
rect 54270 -118915 55070 -118900
rect 54270 -118935 54280 -118915
rect 55060 -118935 55070 -118915
rect 54270 -118960 55070 -118935
rect 54270 -118990 54280 -118960
rect 55060 -118990 55070 -118960
rect 54270 -119000 55070 -118990
rect 55770 -118915 56570 -118900
rect 55770 -118935 55780 -118915
rect 56560 -118935 56570 -118915
rect 55770 -118960 56570 -118935
rect 55770 -118990 55780 -118960
rect 56560 -118990 56570 -118960
rect 55770 -119000 56570 -118990
rect 57270 -118915 58070 -118900
rect 57270 -118935 57280 -118915
rect 58060 -118935 58070 -118915
rect 57270 -118960 58070 -118935
rect 57270 -118990 57280 -118960
rect 58060 -118990 58070 -118960
rect 57270 -119000 58070 -118990
rect 58770 -118915 59570 -118900
rect 58770 -118935 58780 -118915
rect 59560 -118935 59570 -118915
rect 58770 -118960 59570 -118935
rect 58770 -118990 58780 -118960
rect 59560 -118990 59570 -118960
rect 58770 -119000 59570 -118990
rect 60270 -118915 61070 -118900
rect 60270 -118935 60280 -118915
rect 61060 -118935 61070 -118915
rect 60270 -118960 61070 -118935
rect 60270 -118990 60280 -118960
rect 61060 -118990 61070 -118960
rect 60270 -119000 61070 -118990
rect 61770 -118915 62570 -118900
rect 61770 -118935 61780 -118915
rect 62560 -118935 62570 -118915
rect 61770 -118960 62570 -118935
rect 61770 -118990 61780 -118960
rect 62560 -118990 62570 -118960
rect 61770 -119000 62570 -118990
rect 63270 -118915 64070 -118900
rect 63270 -118935 63280 -118915
rect 64060 -118935 64070 -118915
rect 63270 -118960 64070 -118935
rect 63270 -118990 63280 -118960
rect 64060 -118990 64070 -118960
rect 63270 -119000 64070 -118990
rect 64770 -118915 65570 -118900
rect 64770 -118935 64780 -118915
rect 65560 -118935 65570 -118915
rect 64770 -118960 65570 -118935
rect 64770 -118990 64780 -118960
rect 65560 -118990 65570 -118960
rect 64770 -119000 65570 -118990
rect 66270 -118915 67070 -118900
rect 66270 -118935 66280 -118915
rect 67060 -118935 67070 -118915
rect 66270 -118960 67070 -118935
rect 66270 -118990 66280 -118960
rect 67060 -118990 67070 -118960
rect 66270 -119000 67070 -118990
rect 67770 -118915 68570 -118900
rect 67770 -118935 67780 -118915
rect 68560 -118935 68570 -118915
rect 67770 -118960 68570 -118935
rect 67770 -118990 67780 -118960
rect 68560 -118990 68570 -118960
rect 67770 -119000 68570 -118990
rect 69270 -118915 70070 -118900
rect 69270 -118935 69280 -118915
rect 70060 -118935 70070 -118915
rect 69270 -118960 70070 -118935
rect 69270 -118990 69280 -118960
rect 70060 -118990 70070 -118960
rect 69270 -119000 70070 -118990
rect 70770 -118915 71570 -118900
rect 70770 -118935 70780 -118915
rect 71560 -118935 71570 -118915
rect 70770 -118960 71570 -118935
rect 70770 -118990 70780 -118960
rect 71560 -118990 71570 -118960
rect 70770 -119000 71570 -118990
rect 72270 -118915 73070 -118900
rect 72270 -118935 72280 -118915
rect 73060 -118935 73070 -118915
rect 72270 -118960 73070 -118935
rect 72270 -118990 72280 -118960
rect 73060 -118990 73070 -118960
rect 72270 -119000 73070 -118990
rect 73770 -118915 74570 -118900
rect 73770 -118935 73780 -118915
rect 74560 -118935 74570 -118915
rect 73770 -118960 74570 -118935
rect 73770 -118990 73780 -118960
rect 74560 -118990 74570 -118960
rect 73770 -119000 74570 -118990
rect 75270 -118915 76070 -118900
rect 75270 -118935 75280 -118915
rect 76060 -118935 76070 -118915
rect 75270 -118960 76070 -118935
rect 75270 -118990 75280 -118960
rect 76060 -118990 76070 -118960
rect 75270 -119000 76070 -118990
rect 76770 -118915 77570 -118900
rect 76770 -118935 76780 -118915
rect 77560 -118935 77570 -118915
rect 76770 -118960 77570 -118935
rect 76770 -118990 76780 -118960
rect 77560 -118990 77570 -118960
rect 76770 -119000 77570 -118990
rect 78270 -118915 79070 -118900
rect 78270 -118935 78280 -118915
rect 79060 -118935 79070 -118915
rect 78270 -118960 79070 -118935
rect 78270 -118990 78280 -118960
rect 79060 -118990 79070 -118960
rect 78270 -119000 79070 -118990
rect 79770 -118915 80570 -118900
rect 79770 -118935 79780 -118915
rect 80560 -118935 80570 -118915
rect 79770 -118960 80570 -118935
rect 79770 -118990 79780 -118960
rect 80560 -118990 80570 -118960
rect 79770 -119000 80570 -118990
rect 81270 -118915 82070 -118900
rect 81270 -118935 81280 -118915
rect 82060 -118935 82070 -118915
rect 81270 -118960 82070 -118935
rect 81270 -118990 81280 -118960
rect 82060 -118990 82070 -118960
rect 81270 -119000 82070 -118990
rect 82770 -118915 83570 -118900
rect 82770 -118935 82780 -118915
rect 83560 -118935 83570 -118915
rect 82770 -118960 83570 -118935
rect 82770 -118990 82780 -118960
rect 83560 -118990 83570 -118960
rect 82770 -119000 83570 -118990
rect 84270 -118915 85070 -118900
rect 84270 -118935 84280 -118915
rect 85060 -118935 85070 -118915
rect 84270 -118960 85070 -118935
rect 84270 -118990 84280 -118960
rect 85060 -118990 85070 -118960
rect 84270 -119000 85070 -118990
rect 85770 -118915 86570 -118900
rect 85770 -118935 85780 -118915
rect 86560 -118935 86570 -118915
rect 85770 -118960 86570 -118935
rect 85770 -118990 85780 -118960
rect 86560 -118990 86570 -118960
rect 85770 -119000 86570 -118990
rect 87270 -118915 88070 -118900
rect 87270 -118935 87280 -118915
rect 88060 -118935 88070 -118915
rect 87270 -118960 88070 -118935
rect 87270 -118990 87280 -118960
rect 88060 -118990 88070 -118960
rect 87270 -119000 88070 -118990
rect 88770 -118915 89570 -118900
rect 88770 -118935 88780 -118915
rect 89560 -118935 89570 -118915
rect 88770 -118960 89570 -118935
rect 88770 -118990 88780 -118960
rect 89560 -118990 89570 -118960
rect 88770 -119000 89570 -118990
rect 90270 -118915 91070 -118900
rect 90270 -118935 90280 -118915
rect 91060 -118935 91070 -118915
rect 90270 -118960 91070 -118935
rect 90270 -118990 90280 -118960
rect 91060 -118990 91070 -118960
rect 90270 -119000 91070 -118990
rect 91770 -118915 92570 -118900
rect 91770 -118935 91780 -118915
rect 92560 -118935 92570 -118915
rect 91770 -118960 92570 -118935
rect 91770 -118990 91780 -118960
rect 92560 -118990 92570 -118960
rect 91770 -119000 92570 -118990
rect 93270 -118915 94070 -118900
rect 93270 -118935 93280 -118915
rect 94060 -118935 94070 -118915
rect 93270 -118960 94070 -118935
rect 93270 -118990 93280 -118960
rect 94060 -118990 94070 -118960
rect 93270 -119000 94070 -118990
rect 94770 -118915 95570 -118900
rect 94770 -118935 94780 -118915
rect 95560 -118935 95570 -118915
rect 94770 -118960 95570 -118935
rect 94770 -118990 94780 -118960
rect 95560 -118990 95570 -118960
rect 94770 -119000 95570 -118990
rect 96270 -118915 97070 -118900
rect 96270 -118935 96280 -118915
rect 97060 -118935 97070 -118915
rect 96270 -118960 97070 -118935
rect 96270 -118990 96280 -118960
rect 97060 -118990 97070 -118960
rect 96270 -119000 97070 -118990
rect 97770 -118915 98570 -118900
rect 97770 -118935 97780 -118915
rect 98560 -118935 98570 -118915
rect 97770 -118960 98570 -118935
rect 97770 -118990 97780 -118960
rect 98560 -118990 98570 -118960
rect 97770 -119000 98570 -118990
rect 99270 -118915 100070 -118900
rect 99270 -118935 99280 -118915
rect 100060 -118935 100070 -118915
rect 99270 -118960 100070 -118935
rect 99270 -118990 99280 -118960
rect 100060 -118990 100070 -118960
rect 99270 -119000 100070 -118990
rect 100770 -118915 101570 -118900
rect 100770 -118935 100780 -118915
rect 101560 -118935 101570 -118915
rect 100770 -118960 101570 -118935
rect 100770 -118990 100780 -118960
rect 101560 -118990 101570 -118960
rect 100770 -119000 101570 -118990
rect 102270 -118915 103070 -118900
rect 102270 -118935 102280 -118915
rect 103060 -118935 103070 -118915
rect 102270 -118960 103070 -118935
rect 102270 -118990 102280 -118960
rect 103060 -118990 103070 -118960
rect 102270 -119000 103070 -118990
rect 103770 -118915 104570 -118900
rect 103770 -118935 103780 -118915
rect 104560 -118935 104570 -118915
rect 103770 -118960 104570 -118935
rect 103770 -118990 103780 -118960
rect 104560 -118990 104570 -118960
rect 103770 -119000 104570 -118990
rect 105270 -118915 106070 -118900
rect 105270 -118935 105280 -118915
rect 106060 -118935 106070 -118915
rect 105270 -118960 106070 -118935
rect 105270 -118990 105280 -118960
rect 106060 -118990 106070 -118960
rect 105270 -119000 106070 -118990
rect 106770 -118915 107570 -118900
rect 106770 -118935 106780 -118915
rect 107560 -118935 107570 -118915
rect 106770 -118960 107570 -118935
rect 106770 -118990 106780 -118960
rect 107560 -118990 107570 -118960
rect 106770 -119000 107570 -118990
rect 108270 -118915 109070 -118900
rect 108270 -118935 108280 -118915
rect 109060 -118935 109070 -118915
rect 108270 -118960 109070 -118935
rect 108270 -118990 108280 -118960
rect 109060 -118990 109070 -118960
rect 108270 -119000 109070 -118990
rect 109770 -118915 110570 -118900
rect 109770 -118935 109780 -118915
rect 110560 -118935 110570 -118915
rect 109770 -118960 110570 -118935
rect 109770 -118990 109780 -118960
rect 110560 -118990 110570 -118960
rect 109770 -119000 110570 -118990
rect 111270 -118915 112070 -118900
rect 111270 -118935 111280 -118915
rect 112060 -118935 112070 -118915
rect 111270 -118960 112070 -118935
rect 111270 -118990 111280 -118960
rect 112060 -118990 112070 -118960
rect 111270 -119000 112070 -118990
rect 112770 -118915 113570 -118900
rect 112770 -118935 112780 -118915
rect 113560 -118935 113570 -118915
rect 112770 -118960 113570 -118935
rect 112770 -118990 112780 -118960
rect 113560 -118990 113570 -118960
rect 112770 -119000 113570 -118990
rect 114270 -118915 115070 -118900
rect 114270 -118935 114280 -118915
rect 115060 -118935 115070 -118915
rect 114270 -118960 115070 -118935
rect 114270 -118990 114280 -118960
rect 115060 -118990 115070 -118960
rect 114270 -119000 115070 -118990
rect 115770 -118915 116570 -118900
rect 115770 -118935 115780 -118915
rect 116560 -118935 116570 -118915
rect 115770 -118960 116570 -118935
rect 115770 -118990 115780 -118960
rect 116560 -118990 116570 -118960
rect 115770 -119000 116570 -118990
rect 117270 -118915 118070 -118900
rect 117270 -118935 117280 -118915
rect 118060 -118935 118070 -118915
rect 117270 -118960 118070 -118935
rect 117270 -118990 117280 -118960
rect 118060 -118990 118070 -118960
rect 117270 -119000 118070 -118990
rect 118770 -118915 119570 -118900
rect 118770 -118935 118780 -118915
rect 119560 -118935 119570 -118915
rect 118770 -118960 119570 -118935
rect 118770 -118990 118780 -118960
rect 119560 -118990 119570 -118960
rect 118770 -119000 119570 -118990
<< viali >>
rect 280 -118645 1060 -118615
rect 1780 -118645 2560 -118615
rect 3280 -118645 4060 -118615
rect 4780 -118645 5560 -118615
rect 6280 -118645 7060 -118615
rect 7780 -118645 8560 -118615
rect 9280 -118645 10060 -118615
rect 10780 -118645 11560 -118615
rect 12280 -118645 13060 -118615
rect 13780 -118645 14560 -118615
rect 15280 -118645 16060 -118615
rect 16780 -118645 17560 -118615
rect 18280 -118645 19060 -118615
rect 19780 -118645 20560 -118615
rect 21280 -118645 22060 -118615
rect 22780 -118645 23560 -118615
rect 24280 -118645 25060 -118615
rect 25780 -118645 26560 -118615
rect 27280 -118645 28060 -118615
rect 28780 -118645 29560 -118615
rect 30280 -118645 31060 -118615
rect 31780 -118645 32560 -118615
rect 33280 -118645 34060 -118615
rect 34780 -118645 35560 -118615
rect 36280 -118645 37060 -118615
rect 37780 -118645 38560 -118615
rect 39280 -118645 40060 -118615
rect 40780 -118645 41560 -118615
rect 42280 -118645 43060 -118615
rect 43780 -118645 44560 -118615
rect 45280 -118645 46060 -118615
rect 46780 -118645 47560 -118615
rect 48280 -118645 49060 -118615
rect 49780 -118645 50560 -118615
rect 51280 -118645 52060 -118615
rect 52780 -118645 53560 -118615
rect 54280 -118645 55060 -118615
rect 55780 -118645 56560 -118615
rect 57280 -118645 58060 -118615
rect 58780 -118645 59560 -118615
rect 60280 -118645 61060 -118615
rect 61780 -118645 62560 -118615
rect 63280 -118645 64060 -118615
rect 64780 -118645 65560 -118615
rect 66280 -118645 67060 -118615
rect 67780 -118645 68560 -118615
rect 69280 -118645 70060 -118615
rect 70780 -118645 71560 -118615
rect 72280 -118645 73060 -118615
rect 73780 -118645 74560 -118615
rect 75280 -118645 76060 -118615
rect 76780 -118645 77560 -118615
rect 78280 -118645 79060 -118615
rect 79780 -118645 80560 -118615
rect 81280 -118645 82060 -118615
rect 82780 -118645 83560 -118615
rect 84280 -118645 85060 -118615
rect 85780 -118645 86560 -118615
rect 87280 -118645 88060 -118615
rect 88780 -118645 89560 -118615
rect 90280 -118645 91060 -118615
rect 91780 -118645 92560 -118615
rect 93280 -118645 94060 -118615
rect 94780 -118645 95560 -118615
rect 96280 -118645 97060 -118615
rect 97780 -118645 98560 -118615
rect 99280 -118645 100060 -118615
rect 100780 -118645 101560 -118615
rect 102280 -118645 103060 -118615
rect 103780 -118645 104560 -118615
rect 105280 -118645 106060 -118615
rect 106780 -118645 107560 -118615
rect 108280 -118645 109060 -118615
rect 109780 -118645 110560 -118615
rect 111280 -118645 112060 -118615
rect 112780 -118645 113560 -118615
rect 114280 -118645 115060 -118615
rect 115780 -118645 116560 -118615
rect 117280 -118645 118060 -118615
rect 118780 -118645 119560 -118615
rect 120 -118850 210 -118750
rect 1620 -118850 1710 -118750
rect 3120 -118850 3210 -118750
rect 4620 -118850 4710 -118750
rect 6120 -118850 6210 -118750
rect 7620 -118850 7710 -118750
rect 9120 -118850 9210 -118750
rect 10620 -118850 10710 -118750
rect 12120 -118850 12210 -118750
rect 13620 -118850 13710 -118750
rect 15120 -118850 15210 -118750
rect 16620 -118850 16710 -118750
rect 18120 -118850 18210 -118750
rect 19620 -118850 19710 -118750
rect 21120 -118850 21210 -118750
rect 22620 -118850 22710 -118750
rect 24120 -118850 24210 -118750
rect 25620 -118850 25710 -118750
rect 27120 -118850 27210 -118750
rect 28620 -118850 28710 -118750
rect 30120 -118850 30210 -118750
rect 31620 -118850 31710 -118750
rect 33120 -118850 33210 -118750
rect 34620 -118850 34710 -118750
rect 36120 -118850 36210 -118750
rect 37620 -118850 37710 -118750
rect 39120 -118850 39210 -118750
rect 40620 -118850 40710 -118750
rect 42120 -118850 42210 -118750
rect 43620 -118850 43710 -118750
rect 45120 -118850 45210 -118750
rect 46620 -118850 46710 -118750
rect 48120 -118850 48210 -118750
rect 49620 -118850 49710 -118750
rect 51120 -118850 51210 -118750
rect 52620 -118850 52710 -118750
rect 54120 -118850 54210 -118750
rect 55620 -118850 55710 -118750
rect 57120 -118850 57210 -118750
rect 58620 -118850 58710 -118750
rect 60120 -118850 60210 -118750
rect 61620 -118850 61710 -118750
rect 63120 -118850 63210 -118750
rect 64620 -118850 64710 -118750
rect 66120 -118850 66210 -118750
rect 67620 -118850 67710 -118750
rect 69120 -118850 69210 -118750
rect 70620 -118850 70710 -118750
rect 72120 -118850 72210 -118750
rect 73620 -118850 73710 -118750
rect 75120 -118850 75210 -118750
rect 76620 -118850 76710 -118750
rect 78120 -118850 78210 -118750
rect 79620 -118850 79710 -118750
rect 81120 -118850 81210 -118750
rect 82620 -118850 82710 -118750
rect 84120 -118850 84210 -118750
rect 85620 -118850 85710 -118750
rect 87120 -118850 87210 -118750
rect 88620 -118850 88710 -118750
rect 90120 -118850 90210 -118750
rect 91620 -118850 91710 -118750
rect 93120 -118850 93210 -118750
rect 94620 -118850 94710 -118750
rect 96120 -118850 96210 -118750
rect 97620 -118850 97710 -118750
rect 99120 -118850 99210 -118750
rect 100620 -118850 100710 -118750
rect 102120 -118850 102210 -118750
rect 103620 -118850 103710 -118750
rect 105120 -118850 105210 -118750
rect 106620 -118850 106710 -118750
rect 108120 -118850 108210 -118750
rect 109620 -118850 109710 -118750
rect 111120 -118850 111210 -118750
rect 112620 -118850 112710 -118750
rect 114120 -118850 114210 -118750
rect 115620 -118850 115710 -118750
rect 117120 -118850 117210 -118750
rect 118620 -118850 118710 -118750
rect 280 -118990 1060 -118960
rect 1780 -118990 2560 -118960
rect 3280 -118990 4060 -118960
rect 4780 -118990 5560 -118960
rect 6280 -118990 7060 -118960
rect 7780 -118990 8560 -118960
rect 9280 -118990 10060 -118960
rect 10780 -118990 11560 -118960
rect 12280 -118990 13060 -118960
rect 13780 -118990 14560 -118960
rect 15280 -118990 16060 -118960
rect 16780 -118990 17560 -118960
rect 18280 -118990 19060 -118960
rect 19780 -118990 20560 -118960
rect 21280 -118990 22060 -118960
rect 22780 -118990 23560 -118960
rect 24280 -118990 25060 -118960
rect 25780 -118990 26560 -118960
rect 27280 -118990 28060 -118960
rect 28780 -118990 29560 -118960
rect 30280 -118990 31060 -118960
rect 31780 -118990 32560 -118960
rect 33280 -118990 34060 -118960
rect 34780 -118990 35560 -118960
rect 36280 -118990 37060 -118960
rect 37780 -118990 38560 -118960
rect 39280 -118990 40060 -118960
rect 40780 -118990 41560 -118960
rect 42280 -118990 43060 -118960
rect 43780 -118990 44560 -118960
rect 45280 -118990 46060 -118960
rect 46780 -118990 47560 -118960
rect 48280 -118990 49060 -118960
rect 49780 -118990 50560 -118960
rect 51280 -118990 52060 -118960
rect 52780 -118990 53560 -118960
rect 54280 -118990 55060 -118960
rect 55780 -118990 56560 -118960
rect 57280 -118990 58060 -118960
rect 58780 -118990 59560 -118960
rect 60280 -118990 61060 -118960
rect 61780 -118990 62560 -118960
rect 63280 -118990 64060 -118960
rect 64780 -118990 65560 -118960
rect 66280 -118990 67060 -118960
rect 67780 -118990 68560 -118960
rect 69280 -118990 70060 -118960
rect 70780 -118990 71560 -118960
rect 72280 -118990 73060 -118960
rect 73780 -118990 74560 -118960
rect 75280 -118990 76060 -118960
rect 76780 -118990 77560 -118960
rect 78280 -118990 79060 -118960
rect 79780 -118990 80560 -118960
rect 81280 -118990 82060 -118960
rect 82780 -118990 83560 -118960
rect 84280 -118990 85060 -118960
rect 85780 -118990 86560 -118960
rect 87280 -118990 88060 -118960
rect 88780 -118990 89560 -118960
rect 90280 -118990 91060 -118960
rect 91780 -118990 92560 -118960
rect 93280 -118990 94060 -118960
rect 94780 -118990 95560 -118960
rect 96280 -118990 97060 -118960
rect 97780 -118990 98560 -118960
rect 99280 -118990 100060 -118960
rect 100780 -118990 101560 -118960
rect 102280 -118990 103060 -118960
rect 103780 -118990 104560 -118960
rect 105280 -118990 106060 -118960
rect 106780 -118990 107560 -118960
rect 108280 -118990 109060 -118960
rect 109780 -118990 110560 -118960
rect 111280 -118990 112060 -118960
rect 112780 -118990 113560 -118960
rect 114280 -118990 115060 -118960
rect 115780 -118990 116560 -118960
rect 117280 -118990 118060 -118960
rect 118780 -118990 119560 -118960
<< metal1 >>
rect -970 1725 119500 1730
rect -970 1680 -960 1725
rect -450 1680 25 1725
rect 70 1680 1525 1725
rect 1570 1680 3025 1725
rect 3070 1680 4525 1725
rect 4570 1680 6025 1725
rect 6070 1680 7525 1725
rect 7570 1680 9025 1725
rect 9070 1680 10525 1725
rect 10570 1680 12025 1725
rect 12070 1680 13525 1725
rect 13570 1680 15025 1725
rect 15070 1680 16525 1725
rect 16570 1680 18025 1725
rect 18070 1680 19525 1725
rect 19570 1680 21025 1725
rect 21070 1680 22525 1725
rect 22570 1680 24025 1725
rect 24070 1680 25525 1725
rect 25570 1680 27025 1725
rect 27070 1680 28525 1725
rect 28570 1680 30025 1725
rect 30070 1680 31525 1725
rect 31570 1680 33025 1725
rect 33070 1680 34525 1725
rect 34570 1680 36025 1725
rect 36070 1680 37525 1725
rect 37570 1680 39025 1725
rect 39070 1680 40525 1725
rect 40570 1680 42025 1725
rect 42070 1680 43525 1725
rect 43570 1680 45025 1725
rect 45070 1680 46525 1725
rect 46570 1680 48025 1725
rect 48070 1680 49525 1725
rect 49570 1680 51025 1725
rect 51070 1680 52525 1725
rect 52570 1680 54025 1725
rect 54070 1680 55525 1725
rect 55570 1680 57025 1725
rect 57070 1680 58525 1725
rect 58570 1680 60025 1725
rect 60070 1680 61525 1725
rect 61570 1680 63025 1725
rect 63070 1680 64525 1725
rect 64570 1680 66025 1725
rect 66070 1680 67525 1725
rect 67570 1680 69025 1725
rect 69070 1680 70525 1725
rect 70570 1680 72025 1725
rect 72070 1680 73525 1725
rect 73570 1680 75025 1725
rect 75070 1680 76525 1725
rect 76570 1680 78025 1725
rect 78070 1680 79525 1725
rect 79570 1680 81025 1725
rect 81070 1680 82525 1725
rect 82570 1680 84025 1725
rect 84070 1680 85525 1725
rect 85570 1680 87025 1725
rect 87070 1680 88525 1725
rect 88570 1680 90025 1725
rect 90070 1680 91525 1725
rect 91570 1680 93025 1725
rect 93070 1680 94525 1725
rect 94570 1680 96025 1725
rect 96070 1680 97525 1725
rect 97570 1680 99025 1725
rect 99070 1680 100525 1725
rect 100570 1680 102025 1725
rect 102070 1680 103525 1725
rect 103570 1680 105025 1725
rect 105070 1680 106525 1725
rect 106570 1680 108025 1725
rect 108070 1680 109525 1725
rect 109570 1680 111025 1725
rect 111070 1680 112525 1725
rect 112570 1680 114025 1725
rect 114070 1680 115525 1725
rect 115570 1680 117025 1725
rect 117070 1680 118525 1725
rect 118570 1680 119500 1725
rect -970 1675 119500 1680
rect -1000 1485 -900 1500
rect -1000 1410 0 1485
rect -1000 -15 -900 1410
rect -800 780 0 785
rect -800 745 -790 780
rect -590 745 -270 780
rect -130 745 0 780
rect -800 740 0 745
rect 120200 90 120300 1515
rect 120000 15 120300 90
rect -1000 -90 0 -15
rect -1000 -1515 -900 -90
rect -800 -720 0 -715
rect -800 -755 -790 -720
rect -590 -755 -270 -720
rect -130 -755 0 -720
rect -800 -760 0 -755
rect 120200 -1410 120300 15
rect 120000 -1485 120300 -1410
rect -1000 -1590 0 -1515
rect -1000 -3015 -900 -1590
rect -800 -2220 0 -2215
rect -800 -2255 -790 -2220
rect -590 -2255 -270 -2220
rect -130 -2255 0 -2220
rect -800 -2260 0 -2255
rect 120200 -2910 120300 -1485
rect 120000 -2985 120300 -2910
rect -1000 -3090 0 -3015
rect -1000 -4515 -900 -3090
rect -800 -3720 0 -3715
rect -800 -3755 -790 -3720
rect -590 -3755 -270 -3720
rect -130 -3755 0 -3720
rect -800 -3760 0 -3755
rect 120200 -4410 120300 -2985
rect 120000 -4485 120300 -4410
rect -1000 -4590 0 -4515
rect -1000 -6015 -900 -4590
rect -800 -5220 0 -5215
rect -800 -5255 -790 -5220
rect -590 -5255 -270 -5220
rect -130 -5255 0 -5220
rect -800 -5260 0 -5255
rect 120200 -5910 120300 -4485
rect 120000 -5985 120300 -5910
rect -1000 -6090 0 -6015
rect -1000 -7515 -900 -6090
rect -800 -6720 0 -6715
rect -800 -6755 -790 -6720
rect -590 -6755 -270 -6720
rect -130 -6755 0 -6720
rect -800 -6760 0 -6755
rect 120200 -7410 120300 -5985
rect 120000 -7485 120300 -7410
rect -1000 -7590 0 -7515
rect -1000 -9015 -900 -7590
rect -800 -8220 0 -8215
rect -800 -8255 -790 -8220
rect -590 -8255 -270 -8220
rect -130 -8255 0 -8220
rect -800 -8260 0 -8255
rect 120200 -8910 120300 -7485
rect 120000 -8985 120300 -8910
rect -1000 -9090 0 -9015
rect -1000 -10515 -900 -9090
rect -800 -9720 0 -9715
rect -800 -9755 -790 -9720
rect -590 -9755 -270 -9720
rect -130 -9755 0 -9720
rect -800 -9760 0 -9755
rect 120200 -10410 120300 -8985
rect 120000 -10485 120300 -10410
rect -1000 -10590 0 -10515
rect -1000 -12015 -900 -10590
rect -800 -11220 0 -11215
rect -800 -11255 -790 -11220
rect -590 -11255 -270 -11220
rect -130 -11255 0 -11220
rect -800 -11260 0 -11255
rect 120200 -11910 120300 -10485
rect 120000 -11985 120300 -11910
rect -1000 -12090 0 -12015
rect -1000 -13515 -900 -12090
rect -800 -12720 0 -12715
rect -800 -12755 -790 -12720
rect -590 -12755 -270 -12720
rect -130 -12755 0 -12720
rect -800 -12760 0 -12755
rect 120200 -13410 120300 -11985
rect 120000 -13485 120300 -13410
rect -1000 -13590 0 -13515
rect -1000 -15015 -900 -13590
rect -800 -14220 0 -14215
rect -800 -14255 -790 -14220
rect -590 -14255 -270 -14220
rect -130 -14255 0 -14220
rect -800 -14260 0 -14255
rect 120200 -14910 120300 -13485
rect 120000 -14985 120300 -14910
rect -1000 -15090 0 -15015
rect -1000 -16515 -900 -15090
rect -800 -15720 0 -15715
rect -800 -15755 -790 -15720
rect -590 -15755 -270 -15720
rect -130 -15755 0 -15720
rect -800 -15760 0 -15755
rect 120200 -16410 120300 -14985
rect 120000 -16485 120300 -16410
rect -1000 -16590 0 -16515
rect -1000 -18015 -900 -16590
rect -800 -17220 0 -17215
rect -800 -17255 -790 -17220
rect -590 -17255 -270 -17220
rect -130 -17255 0 -17220
rect -800 -17260 0 -17255
rect 120200 -17910 120300 -16485
rect 120000 -17985 120300 -17910
rect -1000 -18090 0 -18015
rect -1000 -19515 -900 -18090
rect -800 -18720 0 -18715
rect -800 -18755 -790 -18720
rect -590 -18755 -270 -18720
rect -130 -18755 0 -18720
rect -800 -18760 0 -18755
rect 120200 -19410 120300 -17985
rect 120000 -19485 120300 -19410
rect -1000 -19590 0 -19515
rect -1000 -21015 -900 -19590
rect -800 -20220 0 -20215
rect -800 -20255 -790 -20220
rect -590 -20255 -270 -20220
rect -130 -20255 0 -20220
rect -800 -20260 0 -20255
rect 120200 -20910 120300 -19485
rect 120000 -20985 120300 -20910
rect -1000 -21090 0 -21015
rect -1000 -22515 -900 -21090
rect -800 -21720 0 -21715
rect -800 -21755 -790 -21720
rect -590 -21755 -270 -21720
rect -130 -21755 0 -21720
rect -800 -21760 0 -21755
rect 120200 -22410 120300 -20985
rect 120000 -22485 120300 -22410
rect -1000 -22590 0 -22515
rect -1000 -24015 -900 -22590
rect -800 -23220 0 -23215
rect -800 -23255 -790 -23220
rect -590 -23255 -270 -23220
rect -130 -23255 0 -23220
rect -800 -23260 0 -23255
rect 120200 -23910 120300 -22485
rect 120000 -23985 120300 -23910
rect -1000 -24090 0 -24015
rect -1000 -25515 -900 -24090
rect -800 -24720 0 -24715
rect -800 -24755 -790 -24720
rect -590 -24755 -270 -24720
rect -130 -24755 0 -24720
rect -800 -24760 0 -24755
rect 120200 -25410 120300 -23985
rect 120000 -25485 120300 -25410
rect -1000 -25590 0 -25515
rect -1000 -27015 -900 -25590
rect -800 -26220 0 -26215
rect -800 -26255 -790 -26220
rect -590 -26255 -270 -26220
rect -130 -26255 0 -26220
rect -800 -26260 0 -26255
rect 120200 -26910 120300 -25485
rect 120000 -26985 120300 -26910
rect -1000 -27090 0 -27015
rect -1000 -28515 -900 -27090
rect -800 -27720 0 -27715
rect -800 -27755 -790 -27720
rect -590 -27755 -270 -27720
rect -130 -27755 0 -27720
rect -800 -27760 0 -27755
rect 120200 -28410 120300 -26985
rect 120000 -28485 120300 -28410
rect -1000 -28590 0 -28515
rect -1000 -30015 -900 -28590
rect -800 -29220 0 -29215
rect -800 -29255 -790 -29220
rect -590 -29255 -270 -29220
rect -130 -29255 0 -29220
rect -800 -29260 0 -29255
rect 120200 -29910 120300 -28485
rect 120000 -29985 120300 -29910
rect -1000 -30090 0 -30015
rect -1000 -31515 -900 -30090
rect -800 -30720 0 -30715
rect -800 -30755 -790 -30720
rect -590 -30755 -270 -30720
rect -130 -30755 0 -30720
rect -800 -30760 0 -30755
rect 120200 -31410 120300 -29985
rect 120000 -31485 120300 -31410
rect -1000 -31590 0 -31515
rect -1000 -33015 -900 -31590
rect -800 -32220 0 -32215
rect -800 -32255 -790 -32220
rect -590 -32255 -270 -32220
rect -130 -32255 0 -32220
rect -800 -32260 0 -32255
rect 120200 -32910 120300 -31485
rect 120000 -32985 120300 -32910
rect -1000 -33090 0 -33015
rect -1000 -34515 -900 -33090
rect -800 -33720 0 -33715
rect -800 -33755 -790 -33720
rect -590 -33755 -270 -33720
rect -130 -33755 0 -33720
rect -800 -33760 0 -33755
rect 120200 -34410 120300 -32985
rect 120000 -34485 120300 -34410
rect -1000 -34590 0 -34515
rect -1000 -36015 -900 -34590
rect -800 -35220 0 -35215
rect -800 -35255 -790 -35220
rect -590 -35255 -270 -35220
rect -130 -35255 0 -35220
rect -800 -35260 0 -35255
rect 120200 -35910 120300 -34485
rect 120000 -35985 120300 -35910
rect -1000 -36090 0 -36015
rect -1000 -37515 -900 -36090
rect -800 -36720 0 -36715
rect -800 -36755 -790 -36720
rect -590 -36755 -270 -36720
rect -130 -36755 0 -36720
rect -800 -36760 0 -36755
rect 120200 -37410 120300 -35985
rect 120000 -37485 120300 -37410
rect -1000 -37590 0 -37515
rect -1000 -39015 -900 -37590
rect -800 -38220 0 -38215
rect -800 -38255 -790 -38220
rect -590 -38255 -270 -38220
rect -130 -38255 0 -38220
rect -800 -38260 0 -38255
rect 120200 -38910 120300 -37485
rect 120000 -38985 120300 -38910
rect -1000 -39090 0 -39015
rect -1000 -40515 -900 -39090
rect -800 -39720 0 -39715
rect -800 -39755 -790 -39720
rect -590 -39755 -270 -39720
rect -130 -39755 0 -39720
rect -800 -39760 0 -39755
rect 120200 -40410 120300 -38985
rect 120000 -40485 120300 -40410
rect -1000 -40590 0 -40515
rect -1000 -42015 -900 -40590
rect -800 -41220 0 -41215
rect -800 -41255 -790 -41220
rect -590 -41255 -270 -41220
rect -130 -41255 0 -41220
rect -800 -41260 0 -41255
rect 120200 -41910 120300 -40485
rect 120000 -41985 120300 -41910
rect -1000 -42090 0 -42015
rect -1000 -43515 -900 -42090
rect -800 -42720 0 -42715
rect -800 -42755 -790 -42720
rect -590 -42755 -270 -42720
rect -130 -42755 0 -42720
rect -800 -42760 0 -42755
rect 120200 -43410 120300 -41985
rect 120000 -43485 120300 -43410
rect -1000 -43590 0 -43515
rect -1000 -45015 -900 -43590
rect -800 -44220 0 -44215
rect -800 -44255 -790 -44220
rect -590 -44255 -270 -44220
rect -130 -44255 0 -44220
rect -800 -44260 0 -44255
rect 120200 -44910 120300 -43485
rect 120000 -44985 120300 -44910
rect -1000 -45090 0 -45015
rect -1000 -46515 -900 -45090
rect -800 -45720 0 -45715
rect -800 -45755 -790 -45720
rect -590 -45755 -270 -45720
rect -130 -45755 0 -45720
rect -800 -45760 0 -45755
rect 120200 -46410 120300 -44985
rect 120000 -46485 120300 -46410
rect -1000 -46590 0 -46515
rect -1000 -48015 -900 -46590
rect -800 -47220 0 -47215
rect -800 -47255 -790 -47220
rect -590 -47255 -270 -47220
rect -130 -47255 0 -47220
rect -800 -47260 0 -47255
rect 120200 -47910 120300 -46485
rect 120000 -47985 120300 -47910
rect -1000 -48090 0 -48015
rect -1000 -49515 -900 -48090
rect -800 -48720 0 -48715
rect -800 -48755 -790 -48720
rect -590 -48755 -270 -48720
rect -130 -48755 0 -48720
rect -800 -48760 0 -48755
rect 120200 -49410 120300 -47985
rect 120000 -49485 120300 -49410
rect -1000 -49590 0 -49515
rect -1000 -51015 -900 -49590
rect -800 -50220 0 -50215
rect -800 -50255 -790 -50220
rect -590 -50255 -270 -50220
rect -130 -50255 0 -50220
rect -800 -50260 0 -50255
rect 120200 -50910 120300 -49485
rect 120000 -50985 120300 -50910
rect -1000 -51090 0 -51015
rect -1000 -52515 -900 -51090
rect -800 -51720 0 -51715
rect -800 -51755 -790 -51720
rect -590 -51755 -270 -51720
rect -130 -51755 0 -51720
rect -800 -51760 0 -51755
rect 120200 -52410 120300 -50985
rect 120000 -52485 120300 -52410
rect -1000 -52590 0 -52515
rect -1000 -54015 -900 -52590
rect -800 -53220 0 -53215
rect -800 -53255 -790 -53220
rect -590 -53255 -270 -53220
rect -130 -53255 0 -53220
rect -800 -53260 0 -53255
rect 120200 -53910 120300 -52485
rect 120000 -53985 120300 -53910
rect -1000 -54090 0 -54015
rect -1000 -55515 -900 -54090
rect -800 -54720 0 -54715
rect -800 -54755 -790 -54720
rect -590 -54755 -270 -54720
rect -130 -54755 0 -54720
rect -800 -54760 0 -54755
rect 120200 -55410 120300 -53985
rect 120000 -55485 120300 -55410
rect -1000 -55590 0 -55515
rect -1000 -57015 -900 -55590
rect -800 -56220 0 -56215
rect -800 -56255 -790 -56220
rect -590 -56255 -270 -56220
rect -130 -56255 0 -56220
rect -800 -56260 0 -56255
rect 120200 -56910 120300 -55485
rect 120000 -56985 120300 -56910
rect -1000 -57090 0 -57015
rect -1000 -58515 -900 -57090
rect -800 -57720 0 -57715
rect -800 -57755 -790 -57720
rect -590 -57755 -270 -57720
rect -130 -57755 0 -57720
rect -800 -57760 0 -57755
rect 120200 -58410 120300 -56985
rect 120000 -58485 120300 -58410
rect -1000 -58590 0 -58515
rect -1000 -60015 -900 -58590
rect -800 -59220 0 -59215
rect -800 -59255 -790 -59220
rect -590 -59255 -270 -59220
rect -130 -59255 0 -59220
rect -800 -59260 0 -59255
rect 120200 -59910 120300 -58485
rect 120000 -59985 120300 -59910
rect -1000 -60090 0 -60015
rect -1000 -61515 -900 -60090
rect -800 -60720 0 -60715
rect -800 -60755 -790 -60720
rect -590 -60755 -270 -60720
rect -130 -60755 0 -60720
rect -800 -60760 0 -60755
rect 120200 -61410 120300 -59985
rect 120000 -61485 120300 -61410
rect -1000 -61590 0 -61515
rect -1000 -63015 -900 -61590
rect -800 -62220 0 -62215
rect -800 -62255 -790 -62220
rect -590 -62255 -270 -62220
rect -130 -62255 0 -62220
rect -800 -62260 0 -62255
rect 120200 -62910 120300 -61485
rect 120000 -62985 120300 -62910
rect -1000 -63090 0 -63015
rect -1000 -64515 -900 -63090
rect -800 -63720 0 -63715
rect -800 -63755 -790 -63720
rect -590 -63755 -270 -63720
rect -130 -63755 0 -63720
rect -800 -63760 0 -63755
rect 120200 -64410 120300 -62985
rect 120000 -64485 120300 -64410
rect -1000 -64590 0 -64515
rect -1000 -66015 -900 -64590
rect -800 -65220 0 -65215
rect -800 -65255 -790 -65220
rect -590 -65255 -270 -65220
rect -130 -65255 0 -65220
rect -800 -65260 0 -65255
rect 120200 -65910 120300 -64485
rect 120000 -65985 120300 -65910
rect -1000 -66090 0 -66015
rect -1000 -67515 -900 -66090
rect -800 -66720 0 -66715
rect -800 -66755 -790 -66720
rect -590 -66755 -270 -66720
rect -130 -66755 0 -66720
rect -800 -66760 0 -66755
rect 120200 -67410 120300 -65985
rect 120000 -67485 120300 -67410
rect -1000 -67590 0 -67515
rect -1000 -69015 -900 -67590
rect -800 -68220 0 -68215
rect -800 -68255 -790 -68220
rect -590 -68255 -270 -68220
rect -130 -68255 0 -68220
rect -800 -68260 0 -68255
rect 120200 -68910 120300 -67485
rect 120000 -68985 120300 -68910
rect -1000 -69090 0 -69015
rect -1000 -70515 -900 -69090
rect -800 -69720 0 -69715
rect -800 -69755 -790 -69720
rect -590 -69755 -270 -69720
rect -130 -69755 0 -69720
rect -800 -69760 0 -69755
rect 120200 -70410 120300 -68985
rect 120000 -70485 120300 -70410
rect -1000 -70590 0 -70515
rect -1000 -72015 -900 -70590
rect -800 -71220 0 -71215
rect -800 -71255 -790 -71220
rect -590 -71255 -270 -71220
rect -130 -71255 0 -71220
rect -800 -71260 0 -71255
rect 120200 -71910 120300 -70485
rect 120000 -71985 120300 -71910
rect -1000 -72090 0 -72015
rect -1000 -73515 -900 -72090
rect -800 -72720 0 -72715
rect -800 -72755 -790 -72720
rect -590 -72755 -270 -72720
rect -130 -72755 0 -72720
rect -800 -72760 0 -72755
rect 120200 -73410 120300 -71985
rect 120000 -73485 120300 -73410
rect -1000 -73590 0 -73515
rect -1000 -75015 -900 -73590
rect -800 -74220 0 -74215
rect -800 -74255 -790 -74220
rect -590 -74255 -270 -74220
rect -130 -74255 0 -74220
rect -800 -74260 0 -74255
rect 120200 -74910 120300 -73485
rect 120000 -74985 120300 -74910
rect -1000 -75090 0 -75015
rect -1000 -76515 -900 -75090
rect -800 -75720 0 -75715
rect -800 -75755 -790 -75720
rect -590 -75755 -270 -75720
rect -130 -75755 0 -75720
rect -800 -75760 0 -75755
rect 120200 -76410 120300 -74985
rect 120000 -76485 120300 -76410
rect -1000 -76590 0 -76515
rect -1000 -78015 -900 -76590
rect -800 -77220 0 -77215
rect -800 -77255 -790 -77220
rect -590 -77255 -270 -77220
rect -130 -77255 0 -77220
rect -800 -77260 0 -77255
rect 120200 -77910 120300 -76485
rect 120000 -77985 120300 -77910
rect -1000 -78090 0 -78015
rect -1000 -79515 -900 -78090
rect -800 -78720 0 -78715
rect -800 -78755 -790 -78720
rect -590 -78755 -270 -78720
rect -130 -78755 0 -78720
rect -800 -78760 0 -78755
rect 120200 -79410 120300 -77985
rect 120000 -79485 120300 -79410
rect -1000 -79590 0 -79515
rect -1000 -81015 -900 -79590
rect -800 -80220 0 -80215
rect -800 -80255 -790 -80220
rect -590 -80255 -270 -80220
rect -130 -80255 0 -80220
rect -800 -80260 0 -80255
rect 120200 -80910 120300 -79485
rect 120000 -80985 120300 -80910
rect -1000 -81090 0 -81015
rect -1000 -82515 -900 -81090
rect -800 -81720 0 -81715
rect -800 -81755 -790 -81720
rect -590 -81755 -270 -81720
rect -130 -81755 0 -81720
rect -800 -81760 0 -81755
rect 120200 -82410 120300 -80985
rect 120000 -82485 120300 -82410
rect -1000 -82590 0 -82515
rect -1000 -84015 -900 -82590
rect -800 -83220 0 -83215
rect -800 -83255 -790 -83220
rect -590 -83255 -270 -83220
rect -130 -83255 0 -83220
rect -800 -83260 0 -83255
rect 120200 -83910 120300 -82485
rect 120000 -83985 120300 -83910
rect -1000 -84090 0 -84015
rect -1000 -85515 -900 -84090
rect -800 -84720 0 -84715
rect -800 -84755 -790 -84720
rect -590 -84755 -270 -84720
rect -130 -84755 0 -84720
rect -800 -84760 0 -84755
rect 120200 -85410 120300 -83985
rect 120000 -85485 120300 -85410
rect -1000 -85590 0 -85515
rect -1000 -87015 -900 -85590
rect -800 -86220 0 -86215
rect -800 -86255 -790 -86220
rect -590 -86255 -270 -86220
rect -130 -86255 0 -86220
rect -800 -86260 0 -86255
rect 120200 -86910 120300 -85485
rect 120000 -86985 120300 -86910
rect -1000 -87090 0 -87015
rect -1000 -88515 -900 -87090
rect -800 -87720 0 -87715
rect -800 -87755 -790 -87720
rect -590 -87755 -270 -87720
rect -130 -87755 0 -87720
rect -800 -87760 0 -87755
rect 120200 -88410 120300 -86985
rect 120000 -88485 120300 -88410
rect -1000 -88590 0 -88515
rect -1000 -90015 -900 -88590
rect -800 -89220 0 -89215
rect -800 -89255 -790 -89220
rect -590 -89255 -270 -89220
rect -130 -89255 0 -89220
rect -800 -89260 0 -89255
rect 120200 -89910 120300 -88485
rect 120000 -89985 120300 -89910
rect -1000 -90090 0 -90015
rect -1000 -91515 -900 -90090
rect -800 -90720 0 -90715
rect -800 -90755 -790 -90720
rect -590 -90755 -270 -90720
rect -130 -90755 0 -90720
rect -800 -90760 0 -90755
rect 120200 -91410 120300 -89985
rect 120000 -91485 120300 -91410
rect -1000 -91590 0 -91515
rect -1000 -93015 -900 -91590
rect -800 -92220 0 -92215
rect -800 -92255 -790 -92220
rect -590 -92255 -270 -92220
rect -130 -92255 0 -92220
rect -800 -92260 0 -92255
rect 120200 -92910 120300 -91485
rect 120000 -92985 120300 -92910
rect -1000 -93090 0 -93015
rect -1000 -94515 -900 -93090
rect -800 -93720 0 -93715
rect -800 -93755 -790 -93720
rect -590 -93755 -270 -93720
rect -130 -93755 0 -93720
rect -800 -93760 0 -93755
rect 120200 -94410 120300 -92985
rect 120000 -94485 120300 -94410
rect -1000 -94590 0 -94515
rect -1000 -96015 -900 -94590
rect -800 -95220 0 -95215
rect -800 -95255 -790 -95220
rect -590 -95255 -270 -95220
rect -130 -95255 0 -95220
rect -800 -95260 0 -95255
rect 120200 -95910 120300 -94485
rect 120000 -95985 120300 -95910
rect -1000 -96090 0 -96015
rect -1000 -97515 -900 -96090
rect -800 -96720 0 -96715
rect -800 -96755 -790 -96720
rect -590 -96755 -270 -96720
rect -130 -96755 0 -96720
rect -800 -96760 0 -96755
rect 120200 -97410 120300 -95985
rect 120000 -97485 120300 -97410
rect -1000 -97590 0 -97515
rect -1000 -99015 -900 -97590
rect -800 -98220 0 -98215
rect -800 -98255 -790 -98220
rect -590 -98255 -270 -98220
rect -130 -98255 0 -98220
rect -800 -98260 0 -98255
rect 120200 -98910 120300 -97485
rect 120000 -98985 120300 -98910
rect -1000 -99090 0 -99015
rect -1000 -100515 -900 -99090
rect -800 -99720 0 -99715
rect -800 -99755 -790 -99720
rect -590 -99755 -270 -99720
rect -130 -99755 0 -99720
rect -800 -99760 0 -99755
rect 120200 -100410 120300 -98985
rect 120000 -100485 120300 -100410
rect -1000 -100590 0 -100515
rect -1000 -102015 -900 -100590
rect -800 -101220 0 -101215
rect -800 -101255 -790 -101220
rect -590 -101255 -270 -101220
rect -130 -101255 0 -101220
rect -800 -101260 0 -101255
rect 120200 -101910 120300 -100485
rect 120000 -101985 120300 -101910
rect -1000 -102090 0 -102015
rect -1000 -103515 -900 -102090
rect -800 -102720 0 -102715
rect -800 -102755 -790 -102720
rect -590 -102755 -270 -102720
rect -130 -102755 0 -102720
rect -800 -102760 0 -102755
rect 120200 -103410 120300 -101985
rect 120000 -103485 120300 -103410
rect -1000 -103590 0 -103515
rect -1000 -105015 -900 -103590
rect -800 -104220 0 -104215
rect -800 -104255 -790 -104220
rect -590 -104255 -270 -104220
rect -130 -104255 0 -104220
rect -800 -104260 0 -104255
rect 120200 -104910 120300 -103485
rect 120000 -104985 120300 -104910
rect -1000 -105090 0 -105015
rect -1000 -106515 -900 -105090
rect -800 -105720 0 -105715
rect -800 -105755 -790 -105720
rect -590 -105755 -270 -105720
rect -130 -105755 0 -105720
rect -800 -105760 0 -105755
rect 120200 -106410 120300 -104985
rect 120000 -106485 120300 -106410
rect -1000 -106590 0 -106515
rect -1000 -108015 -900 -106590
rect -800 -107220 0 -107215
rect -800 -107255 -790 -107220
rect -590 -107255 -270 -107220
rect -130 -107255 0 -107220
rect -800 -107260 0 -107255
rect 120200 -107910 120300 -106485
rect 120000 -107985 120300 -107910
rect -1000 -108090 0 -108015
rect -1000 -109515 -900 -108090
rect -800 -108720 0 -108715
rect -800 -108755 -790 -108720
rect -590 -108755 -270 -108720
rect -130 -108755 0 -108720
rect -800 -108760 0 -108755
rect 120200 -109410 120300 -107985
rect 120000 -109485 120300 -109410
rect -1000 -109590 0 -109515
rect -1000 -111015 -900 -109590
rect -800 -110220 0 -110215
rect -800 -110255 -790 -110220
rect -590 -110255 -270 -110220
rect -130 -110255 0 -110220
rect -800 -110260 0 -110255
rect 120200 -110910 120300 -109485
rect 120000 -110985 120300 -110910
rect -1000 -111090 0 -111015
rect -1000 -112515 -900 -111090
rect -800 -111720 0 -111715
rect -800 -111755 -790 -111720
rect -590 -111755 -270 -111720
rect -130 -111755 0 -111720
rect -800 -111760 0 -111755
rect 120200 -112410 120300 -110985
rect 120000 -112485 120300 -112410
rect -1000 -112590 0 -112515
rect -1000 -114015 -900 -112590
rect -800 -113220 0 -113215
rect -800 -113255 -790 -113220
rect -590 -113255 -270 -113220
rect -130 -113255 0 -113220
rect -800 -113260 0 -113255
rect 120200 -113910 120300 -112485
rect 120000 -113985 120300 -113910
rect -1000 -114090 0 -114015
rect -1000 -115515 -900 -114090
rect -800 -114720 0 -114715
rect -800 -114755 -790 -114720
rect -590 -114755 -270 -114720
rect -130 -114755 0 -114720
rect -800 -114760 0 -114755
rect 120200 -115410 120300 -113985
rect 120000 -115485 120300 -115410
rect -1000 -115590 0 -115515
rect -1000 -117015 -900 -115590
rect -800 -116220 0 -116215
rect -800 -116255 -790 -116220
rect -590 -116255 -270 -116220
rect -130 -116255 0 -116220
rect -800 -116260 0 -116255
rect 120200 -116910 120300 -115485
rect 120000 -116985 120300 -116910
rect -1000 -117090 0 -117015
rect -1000 -118500 -900 -117090
rect -800 -117720 0 -117715
rect -800 -117755 -790 -117720
rect -590 -117755 -270 -117720
rect -130 -117755 0 -117720
rect -800 -117760 0 -117755
rect 120200 -118410 120300 -116985
rect 120000 -118485 120300 -118410
rect 270 -118600 280 -118565
rect 1060 -118600 1070 -118565
rect 270 -118615 1070 -118600
rect 270 -118645 280 -118615
rect 1060 -118645 1070 -118615
rect 270 -118650 1070 -118645
rect 1770 -118600 1780 -118565
rect 2560 -118600 2570 -118565
rect 1770 -118615 2570 -118600
rect 1770 -118645 1780 -118615
rect 2560 -118645 2570 -118615
rect 1770 -118650 2570 -118645
rect 3270 -118600 3280 -118565
rect 4060 -118600 4070 -118565
rect 3270 -118615 4070 -118600
rect 3270 -118645 3280 -118615
rect 4060 -118645 4070 -118615
rect 3270 -118650 4070 -118645
rect 4770 -118600 4780 -118565
rect 5560 -118600 5570 -118565
rect 4770 -118615 5570 -118600
rect 4770 -118645 4780 -118615
rect 5560 -118645 5570 -118615
rect 4770 -118650 5570 -118645
rect 6270 -118600 6280 -118565
rect 7060 -118600 7070 -118565
rect 6270 -118615 7070 -118600
rect 6270 -118645 6280 -118615
rect 7060 -118645 7070 -118615
rect 6270 -118650 7070 -118645
rect 7770 -118600 7780 -118565
rect 8560 -118600 8570 -118565
rect 7770 -118615 8570 -118600
rect 7770 -118645 7780 -118615
rect 8560 -118645 8570 -118615
rect 7770 -118650 8570 -118645
rect 9270 -118600 9280 -118565
rect 10060 -118600 10070 -118565
rect 9270 -118615 10070 -118600
rect 9270 -118645 9280 -118615
rect 10060 -118645 10070 -118615
rect 9270 -118650 10070 -118645
rect 10770 -118600 10780 -118565
rect 11560 -118600 11570 -118565
rect 10770 -118615 11570 -118600
rect 10770 -118645 10780 -118615
rect 11560 -118645 11570 -118615
rect 10770 -118650 11570 -118645
rect 12270 -118600 12280 -118565
rect 13060 -118600 13070 -118565
rect 12270 -118615 13070 -118600
rect 12270 -118645 12280 -118615
rect 13060 -118645 13070 -118615
rect 12270 -118650 13070 -118645
rect 13770 -118600 13780 -118565
rect 14560 -118600 14570 -118565
rect 13770 -118615 14570 -118600
rect 13770 -118645 13780 -118615
rect 14560 -118645 14570 -118615
rect 13770 -118650 14570 -118645
rect 15270 -118600 15280 -118565
rect 16060 -118600 16070 -118565
rect 15270 -118615 16070 -118600
rect 15270 -118645 15280 -118615
rect 16060 -118645 16070 -118615
rect 15270 -118650 16070 -118645
rect 16770 -118600 16780 -118565
rect 17560 -118600 17570 -118565
rect 16770 -118615 17570 -118600
rect 16770 -118645 16780 -118615
rect 17560 -118645 17570 -118615
rect 16770 -118650 17570 -118645
rect 18270 -118600 18280 -118565
rect 19060 -118600 19070 -118565
rect 18270 -118615 19070 -118600
rect 18270 -118645 18280 -118615
rect 19060 -118645 19070 -118615
rect 18270 -118650 19070 -118645
rect 19770 -118600 19780 -118565
rect 20560 -118600 20570 -118565
rect 19770 -118615 20570 -118600
rect 19770 -118645 19780 -118615
rect 20560 -118645 20570 -118615
rect 19770 -118650 20570 -118645
rect 21270 -118600 21280 -118565
rect 22060 -118600 22070 -118565
rect 21270 -118615 22070 -118600
rect 21270 -118645 21280 -118615
rect 22060 -118645 22070 -118615
rect 21270 -118650 22070 -118645
rect 22770 -118600 22780 -118565
rect 23560 -118600 23570 -118565
rect 22770 -118615 23570 -118600
rect 22770 -118645 22780 -118615
rect 23560 -118645 23570 -118615
rect 22770 -118650 23570 -118645
rect 24270 -118600 24280 -118565
rect 25060 -118600 25070 -118565
rect 24270 -118615 25070 -118600
rect 24270 -118645 24280 -118615
rect 25060 -118645 25070 -118615
rect 24270 -118650 25070 -118645
rect 25770 -118600 25780 -118565
rect 26560 -118600 26570 -118565
rect 25770 -118615 26570 -118600
rect 25770 -118645 25780 -118615
rect 26560 -118645 26570 -118615
rect 25770 -118650 26570 -118645
rect 27270 -118600 27280 -118565
rect 28060 -118600 28070 -118565
rect 27270 -118615 28070 -118600
rect 27270 -118645 27280 -118615
rect 28060 -118645 28070 -118615
rect 27270 -118650 28070 -118645
rect 28770 -118600 28780 -118565
rect 29560 -118600 29570 -118565
rect 28770 -118615 29570 -118600
rect 28770 -118645 28780 -118615
rect 29560 -118645 29570 -118615
rect 28770 -118650 29570 -118645
rect 30270 -118600 30280 -118565
rect 31060 -118600 31070 -118565
rect 30270 -118615 31070 -118600
rect 30270 -118645 30280 -118615
rect 31060 -118645 31070 -118615
rect 30270 -118650 31070 -118645
rect 31770 -118600 31780 -118565
rect 32560 -118600 32570 -118565
rect 31770 -118615 32570 -118600
rect 31770 -118645 31780 -118615
rect 32560 -118645 32570 -118615
rect 31770 -118650 32570 -118645
rect 33270 -118600 33280 -118565
rect 34060 -118600 34070 -118565
rect 33270 -118615 34070 -118600
rect 33270 -118645 33280 -118615
rect 34060 -118645 34070 -118615
rect 33270 -118650 34070 -118645
rect 34770 -118600 34780 -118565
rect 35560 -118600 35570 -118565
rect 34770 -118615 35570 -118600
rect 34770 -118645 34780 -118615
rect 35560 -118645 35570 -118615
rect 34770 -118650 35570 -118645
rect 36270 -118600 36280 -118565
rect 37060 -118600 37070 -118565
rect 36270 -118615 37070 -118600
rect 36270 -118645 36280 -118615
rect 37060 -118645 37070 -118615
rect 36270 -118650 37070 -118645
rect 37770 -118600 37780 -118565
rect 38560 -118600 38570 -118565
rect 37770 -118615 38570 -118600
rect 37770 -118645 37780 -118615
rect 38560 -118645 38570 -118615
rect 37770 -118650 38570 -118645
rect 39270 -118600 39280 -118565
rect 40060 -118600 40070 -118565
rect 39270 -118615 40070 -118600
rect 39270 -118645 39280 -118615
rect 40060 -118645 40070 -118615
rect 39270 -118650 40070 -118645
rect 40770 -118600 40780 -118565
rect 41560 -118600 41570 -118565
rect 40770 -118615 41570 -118600
rect 40770 -118645 40780 -118615
rect 41560 -118645 41570 -118615
rect 40770 -118650 41570 -118645
rect 42270 -118600 42280 -118565
rect 43060 -118600 43070 -118565
rect 42270 -118615 43070 -118600
rect 42270 -118645 42280 -118615
rect 43060 -118645 43070 -118615
rect 42270 -118650 43070 -118645
rect 43770 -118600 43780 -118565
rect 44560 -118600 44570 -118565
rect 43770 -118615 44570 -118600
rect 43770 -118645 43780 -118615
rect 44560 -118645 44570 -118615
rect 43770 -118650 44570 -118645
rect 45270 -118600 45280 -118565
rect 46060 -118600 46070 -118565
rect 45270 -118615 46070 -118600
rect 45270 -118645 45280 -118615
rect 46060 -118645 46070 -118615
rect 45270 -118650 46070 -118645
rect 46770 -118600 46780 -118565
rect 47560 -118600 47570 -118565
rect 46770 -118615 47570 -118600
rect 46770 -118645 46780 -118615
rect 47560 -118645 47570 -118615
rect 46770 -118650 47570 -118645
rect 48270 -118600 48280 -118565
rect 49060 -118600 49070 -118565
rect 48270 -118615 49070 -118600
rect 48270 -118645 48280 -118615
rect 49060 -118645 49070 -118615
rect 48270 -118650 49070 -118645
rect 49770 -118600 49780 -118565
rect 50560 -118600 50570 -118565
rect 49770 -118615 50570 -118600
rect 49770 -118645 49780 -118615
rect 50560 -118645 50570 -118615
rect 49770 -118650 50570 -118645
rect 51270 -118600 51280 -118565
rect 52060 -118600 52070 -118565
rect 51270 -118615 52070 -118600
rect 51270 -118645 51280 -118615
rect 52060 -118645 52070 -118615
rect 51270 -118650 52070 -118645
rect 52770 -118600 52780 -118565
rect 53560 -118600 53570 -118565
rect 52770 -118615 53570 -118600
rect 52770 -118645 52780 -118615
rect 53560 -118645 53570 -118615
rect 52770 -118650 53570 -118645
rect 54270 -118600 54280 -118565
rect 55060 -118600 55070 -118565
rect 54270 -118615 55070 -118600
rect 54270 -118645 54280 -118615
rect 55060 -118645 55070 -118615
rect 54270 -118650 55070 -118645
rect 55770 -118600 55780 -118565
rect 56560 -118600 56570 -118565
rect 55770 -118615 56570 -118600
rect 55770 -118645 55780 -118615
rect 56560 -118645 56570 -118615
rect 55770 -118650 56570 -118645
rect 57270 -118600 57280 -118565
rect 58060 -118600 58070 -118565
rect 57270 -118615 58070 -118600
rect 57270 -118645 57280 -118615
rect 58060 -118645 58070 -118615
rect 57270 -118650 58070 -118645
rect 58770 -118600 58780 -118565
rect 59560 -118600 59570 -118565
rect 58770 -118615 59570 -118600
rect 58770 -118645 58780 -118615
rect 59560 -118645 59570 -118615
rect 58770 -118650 59570 -118645
rect 60270 -118600 60280 -118565
rect 61060 -118600 61070 -118565
rect 60270 -118615 61070 -118600
rect 60270 -118645 60280 -118615
rect 61060 -118645 61070 -118615
rect 60270 -118650 61070 -118645
rect 61770 -118600 61780 -118565
rect 62560 -118600 62570 -118565
rect 61770 -118615 62570 -118600
rect 61770 -118645 61780 -118615
rect 62560 -118645 62570 -118615
rect 61770 -118650 62570 -118645
rect 63270 -118600 63280 -118565
rect 64060 -118600 64070 -118565
rect 63270 -118615 64070 -118600
rect 63270 -118645 63280 -118615
rect 64060 -118645 64070 -118615
rect 63270 -118650 64070 -118645
rect 64770 -118600 64780 -118565
rect 65560 -118600 65570 -118565
rect 64770 -118615 65570 -118600
rect 64770 -118645 64780 -118615
rect 65560 -118645 65570 -118615
rect 64770 -118650 65570 -118645
rect 66270 -118600 66280 -118565
rect 67060 -118600 67070 -118565
rect 66270 -118615 67070 -118600
rect 66270 -118645 66280 -118615
rect 67060 -118645 67070 -118615
rect 66270 -118650 67070 -118645
rect 67770 -118600 67780 -118565
rect 68560 -118600 68570 -118565
rect 67770 -118615 68570 -118600
rect 67770 -118645 67780 -118615
rect 68560 -118645 68570 -118615
rect 67770 -118650 68570 -118645
rect 69270 -118600 69280 -118565
rect 70060 -118600 70070 -118565
rect 69270 -118615 70070 -118600
rect 69270 -118645 69280 -118615
rect 70060 -118645 70070 -118615
rect 69270 -118650 70070 -118645
rect 70770 -118600 70780 -118565
rect 71560 -118600 71570 -118565
rect 70770 -118615 71570 -118600
rect 70770 -118645 70780 -118615
rect 71560 -118645 71570 -118615
rect 70770 -118650 71570 -118645
rect 72270 -118600 72280 -118565
rect 73060 -118600 73070 -118565
rect 72270 -118615 73070 -118600
rect 72270 -118645 72280 -118615
rect 73060 -118645 73070 -118615
rect 72270 -118650 73070 -118645
rect 73770 -118600 73780 -118565
rect 74560 -118600 74570 -118565
rect 73770 -118615 74570 -118600
rect 73770 -118645 73780 -118615
rect 74560 -118645 74570 -118615
rect 73770 -118650 74570 -118645
rect 75270 -118600 75280 -118565
rect 76060 -118600 76070 -118565
rect 75270 -118615 76070 -118600
rect 75270 -118645 75280 -118615
rect 76060 -118645 76070 -118615
rect 75270 -118650 76070 -118645
rect 76770 -118600 76780 -118565
rect 77560 -118600 77570 -118565
rect 76770 -118615 77570 -118600
rect 76770 -118645 76780 -118615
rect 77560 -118645 77570 -118615
rect 76770 -118650 77570 -118645
rect 78270 -118600 78280 -118565
rect 79060 -118600 79070 -118565
rect 78270 -118615 79070 -118600
rect 78270 -118645 78280 -118615
rect 79060 -118645 79070 -118615
rect 78270 -118650 79070 -118645
rect 79770 -118600 79780 -118565
rect 80560 -118600 80570 -118565
rect 79770 -118615 80570 -118600
rect 79770 -118645 79780 -118615
rect 80560 -118645 80570 -118615
rect 79770 -118650 80570 -118645
rect 81270 -118600 81280 -118565
rect 82060 -118600 82070 -118565
rect 81270 -118615 82070 -118600
rect 81270 -118645 81280 -118615
rect 82060 -118645 82070 -118615
rect 81270 -118650 82070 -118645
rect 82770 -118600 82780 -118565
rect 83560 -118600 83570 -118565
rect 82770 -118615 83570 -118600
rect 82770 -118645 82780 -118615
rect 83560 -118645 83570 -118615
rect 82770 -118650 83570 -118645
rect 84270 -118600 84280 -118565
rect 85060 -118600 85070 -118565
rect 84270 -118615 85070 -118600
rect 84270 -118645 84280 -118615
rect 85060 -118645 85070 -118615
rect 84270 -118650 85070 -118645
rect 85770 -118600 85780 -118565
rect 86560 -118600 86570 -118565
rect 85770 -118615 86570 -118600
rect 85770 -118645 85780 -118615
rect 86560 -118645 86570 -118615
rect 85770 -118650 86570 -118645
rect 87270 -118600 87280 -118565
rect 88060 -118600 88070 -118565
rect 87270 -118615 88070 -118600
rect 87270 -118645 87280 -118615
rect 88060 -118645 88070 -118615
rect 87270 -118650 88070 -118645
rect 88770 -118600 88780 -118565
rect 89560 -118600 89570 -118565
rect 88770 -118615 89570 -118600
rect 88770 -118645 88780 -118615
rect 89560 -118645 89570 -118615
rect 88770 -118650 89570 -118645
rect 90270 -118600 90280 -118565
rect 91060 -118600 91070 -118565
rect 90270 -118615 91070 -118600
rect 90270 -118645 90280 -118615
rect 91060 -118645 91070 -118615
rect 90270 -118650 91070 -118645
rect 91770 -118600 91780 -118565
rect 92560 -118600 92570 -118565
rect 91770 -118615 92570 -118600
rect 91770 -118645 91780 -118615
rect 92560 -118645 92570 -118615
rect 91770 -118650 92570 -118645
rect 93270 -118600 93280 -118565
rect 94060 -118600 94070 -118565
rect 93270 -118615 94070 -118600
rect 93270 -118645 93280 -118615
rect 94060 -118645 94070 -118615
rect 93270 -118650 94070 -118645
rect 94770 -118600 94780 -118565
rect 95560 -118600 95570 -118565
rect 94770 -118615 95570 -118600
rect 94770 -118645 94780 -118615
rect 95560 -118645 95570 -118615
rect 94770 -118650 95570 -118645
rect 96270 -118600 96280 -118565
rect 97060 -118600 97070 -118565
rect 96270 -118615 97070 -118600
rect 96270 -118645 96280 -118615
rect 97060 -118645 97070 -118615
rect 96270 -118650 97070 -118645
rect 97770 -118600 97780 -118565
rect 98560 -118600 98570 -118565
rect 97770 -118615 98570 -118600
rect 97770 -118645 97780 -118615
rect 98560 -118645 98570 -118615
rect 97770 -118650 98570 -118645
rect 99270 -118600 99280 -118565
rect 100060 -118600 100070 -118565
rect 99270 -118615 100070 -118600
rect 99270 -118645 99280 -118615
rect 100060 -118645 100070 -118615
rect 99270 -118650 100070 -118645
rect 100770 -118600 100780 -118565
rect 101560 -118600 101570 -118565
rect 100770 -118615 101570 -118600
rect 100770 -118645 100780 -118615
rect 101560 -118645 101570 -118615
rect 100770 -118650 101570 -118645
rect 102270 -118600 102280 -118565
rect 103060 -118600 103070 -118565
rect 102270 -118615 103070 -118600
rect 102270 -118645 102280 -118615
rect 103060 -118645 103070 -118615
rect 102270 -118650 103070 -118645
rect 103770 -118600 103780 -118565
rect 104560 -118600 104570 -118565
rect 103770 -118615 104570 -118600
rect 103770 -118645 103780 -118615
rect 104560 -118645 104570 -118615
rect 103770 -118650 104570 -118645
rect 105270 -118600 105280 -118565
rect 106060 -118600 106070 -118565
rect 105270 -118615 106070 -118600
rect 105270 -118645 105280 -118615
rect 106060 -118645 106070 -118615
rect 105270 -118650 106070 -118645
rect 106770 -118600 106780 -118565
rect 107560 -118600 107570 -118565
rect 106770 -118615 107570 -118600
rect 106770 -118645 106780 -118615
rect 107560 -118645 107570 -118615
rect 106770 -118650 107570 -118645
rect 108270 -118600 108280 -118565
rect 109060 -118600 109070 -118565
rect 108270 -118615 109070 -118600
rect 108270 -118645 108280 -118615
rect 109060 -118645 109070 -118615
rect 108270 -118650 109070 -118645
rect 109770 -118600 109780 -118565
rect 110560 -118600 110570 -118565
rect 109770 -118615 110570 -118600
rect 109770 -118645 109780 -118615
rect 110560 -118645 110570 -118615
rect 109770 -118650 110570 -118645
rect 111270 -118600 111280 -118565
rect 112060 -118600 112070 -118565
rect 111270 -118615 112070 -118600
rect 111270 -118645 111280 -118615
rect 112060 -118645 112070 -118615
rect 111270 -118650 112070 -118645
rect 112770 -118600 112780 -118565
rect 113560 -118600 113570 -118565
rect 112770 -118615 113570 -118600
rect 112770 -118645 112780 -118615
rect 113560 -118645 113570 -118615
rect 112770 -118650 113570 -118645
rect 114270 -118600 114280 -118565
rect 115060 -118600 115070 -118565
rect 114270 -118615 115070 -118600
rect 114270 -118645 114280 -118615
rect 115060 -118645 115070 -118615
rect 114270 -118650 115070 -118645
rect 115770 -118600 115780 -118565
rect 116560 -118600 116570 -118565
rect 115770 -118615 116570 -118600
rect 115770 -118645 115780 -118615
rect 116560 -118645 116570 -118615
rect 115770 -118650 116570 -118645
rect 117270 -118600 117280 -118565
rect 118060 -118600 118070 -118565
rect 117270 -118615 118070 -118600
rect 117270 -118645 117280 -118615
rect 118060 -118645 118070 -118615
rect 117270 -118650 118070 -118645
rect 118770 -118600 118780 -118565
rect 119560 -118600 119570 -118565
rect 118770 -118615 119570 -118600
rect 118770 -118645 118780 -118615
rect 119560 -118645 119570 -118615
rect 118770 -118650 119570 -118645
rect 110 -118750 220 -118745
rect 110 -118850 120 -118750
rect 210 -118850 220 -118750
rect 110 -118855 220 -118850
rect 1610 -118750 1720 -118745
rect 1610 -118850 1620 -118750
rect 1710 -118850 1720 -118750
rect 1610 -118855 1720 -118850
rect 3110 -118750 3220 -118745
rect 3110 -118850 3120 -118750
rect 3210 -118850 3220 -118750
rect 3110 -118855 3220 -118850
rect 4610 -118750 4720 -118745
rect 4610 -118850 4620 -118750
rect 4710 -118850 4720 -118750
rect 4610 -118855 4720 -118850
rect 6110 -118750 6220 -118745
rect 6110 -118850 6120 -118750
rect 6210 -118850 6220 -118750
rect 6110 -118855 6220 -118850
rect 7610 -118750 7720 -118745
rect 7610 -118850 7620 -118750
rect 7710 -118850 7720 -118750
rect 7610 -118855 7720 -118850
rect 9110 -118750 9220 -118745
rect 9110 -118850 9120 -118750
rect 9210 -118850 9220 -118750
rect 9110 -118855 9220 -118850
rect 10610 -118750 10720 -118745
rect 10610 -118850 10620 -118750
rect 10710 -118850 10720 -118750
rect 10610 -118855 10720 -118850
rect 12110 -118750 12220 -118745
rect 12110 -118850 12120 -118750
rect 12210 -118850 12220 -118750
rect 12110 -118855 12220 -118850
rect 13610 -118750 13720 -118745
rect 13610 -118850 13620 -118750
rect 13710 -118850 13720 -118750
rect 13610 -118855 13720 -118850
rect 15110 -118750 15220 -118745
rect 15110 -118850 15120 -118750
rect 15210 -118850 15220 -118750
rect 15110 -118855 15220 -118850
rect 16610 -118750 16720 -118745
rect 16610 -118850 16620 -118750
rect 16710 -118850 16720 -118750
rect 16610 -118855 16720 -118850
rect 18110 -118750 18220 -118745
rect 18110 -118850 18120 -118750
rect 18210 -118850 18220 -118750
rect 18110 -118855 18220 -118850
rect 19610 -118750 19720 -118745
rect 19610 -118850 19620 -118750
rect 19710 -118850 19720 -118750
rect 19610 -118855 19720 -118850
rect 21110 -118750 21220 -118745
rect 21110 -118850 21120 -118750
rect 21210 -118850 21220 -118750
rect 21110 -118855 21220 -118850
rect 22610 -118750 22720 -118745
rect 22610 -118850 22620 -118750
rect 22710 -118850 22720 -118750
rect 22610 -118855 22720 -118850
rect 24110 -118750 24220 -118745
rect 24110 -118850 24120 -118750
rect 24210 -118850 24220 -118750
rect 24110 -118855 24220 -118850
rect 25610 -118750 25720 -118745
rect 25610 -118850 25620 -118750
rect 25710 -118850 25720 -118750
rect 25610 -118855 25720 -118850
rect 27110 -118750 27220 -118745
rect 27110 -118850 27120 -118750
rect 27210 -118850 27220 -118750
rect 27110 -118855 27220 -118850
rect 28610 -118750 28720 -118745
rect 28610 -118850 28620 -118750
rect 28710 -118850 28720 -118750
rect 28610 -118855 28720 -118850
rect 30110 -118750 30220 -118745
rect 30110 -118850 30120 -118750
rect 30210 -118850 30220 -118750
rect 30110 -118855 30220 -118850
rect 31610 -118750 31720 -118745
rect 31610 -118850 31620 -118750
rect 31710 -118850 31720 -118750
rect 31610 -118855 31720 -118850
rect 33110 -118750 33220 -118745
rect 33110 -118850 33120 -118750
rect 33210 -118850 33220 -118750
rect 33110 -118855 33220 -118850
rect 34610 -118750 34720 -118745
rect 34610 -118850 34620 -118750
rect 34710 -118850 34720 -118750
rect 34610 -118855 34720 -118850
rect 36110 -118750 36220 -118745
rect 36110 -118850 36120 -118750
rect 36210 -118850 36220 -118750
rect 36110 -118855 36220 -118850
rect 37610 -118750 37720 -118745
rect 37610 -118850 37620 -118750
rect 37710 -118850 37720 -118750
rect 37610 -118855 37720 -118850
rect 39110 -118750 39220 -118745
rect 39110 -118850 39120 -118750
rect 39210 -118850 39220 -118750
rect 39110 -118855 39220 -118850
rect 40610 -118750 40720 -118745
rect 40610 -118850 40620 -118750
rect 40710 -118850 40720 -118750
rect 40610 -118855 40720 -118850
rect 42110 -118750 42220 -118745
rect 42110 -118850 42120 -118750
rect 42210 -118850 42220 -118750
rect 42110 -118855 42220 -118850
rect 43610 -118750 43720 -118745
rect 43610 -118850 43620 -118750
rect 43710 -118850 43720 -118750
rect 43610 -118855 43720 -118850
rect 45110 -118750 45220 -118745
rect 45110 -118850 45120 -118750
rect 45210 -118850 45220 -118750
rect 45110 -118855 45220 -118850
rect 46610 -118750 46720 -118745
rect 46610 -118850 46620 -118750
rect 46710 -118850 46720 -118750
rect 46610 -118855 46720 -118850
rect 48110 -118750 48220 -118745
rect 48110 -118850 48120 -118750
rect 48210 -118850 48220 -118750
rect 48110 -118855 48220 -118850
rect 49610 -118750 49720 -118745
rect 49610 -118850 49620 -118750
rect 49710 -118850 49720 -118750
rect 49610 -118855 49720 -118850
rect 51110 -118750 51220 -118745
rect 51110 -118850 51120 -118750
rect 51210 -118850 51220 -118750
rect 51110 -118855 51220 -118850
rect 52610 -118750 52720 -118745
rect 52610 -118850 52620 -118750
rect 52710 -118850 52720 -118750
rect 52610 -118855 52720 -118850
rect 54110 -118750 54220 -118745
rect 54110 -118850 54120 -118750
rect 54210 -118850 54220 -118750
rect 54110 -118855 54220 -118850
rect 55610 -118750 55720 -118745
rect 55610 -118850 55620 -118750
rect 55710 -118850 55720 -118750
rect 55610 -118855 55720 -118850
rect 57110 -118750 57220 -118745
rect 57110 -118850 57120 -118750
rect 57210 -118850 57220 -118750
rect 57110 -118855 57220 -118850
rect 58610 -118750 58720 -118745
rect 58610 -118850 58620 -118750
rect 58710 -118850 58720 -118750
rect 58610 -118855 58720 -118850
rect 60110 -118750 60220 -118745
rect 60110 -118850 60120 -118750
rect 60210 -118850 60220 -118750
rect 60110 -118855 60220 -118850
rect 61610 -118750 61720 -118745
rect 61610 -118850 61620 -118750
rect 61710 -118850 61720 -118750
rect 61610 -118855 61720 -118850
rect 63110 -118750 63220 -118745
rect 63110 -118850 63120 -118750
rect 63210 -118850 63220 -118750
rect 63110 -118855 63220 -118850
rect 64610 -118750 64720 -118745
rect 64610 -118850 64620 -118750
rect 64710 -118850 64720 -118750
rect 64610 -118855 64720 -118850
rect 66110 -118750 66220 -118745
rect 66110 -118850 66120 -118750
rect 66210 -118850 66220 -118750
rect 66110 -118855 66220 -118850
rect 67610 -118750 67720 -118745
rect 67610 -118850 67620 -118750
rect 67710 -118850 67720 -118750
rect 67610 -118855 67720 -118850
rect 69110 -118750 69220 -118745
rect 69110 -118850 69120 -118750
rect 69210 -118850 69220 -118750
rect 69110 -118855 69220 -118850
rect 70610 -118750 70720 -118745
rect 70610 -118850 70620 -118750
rect 70710 -118850 70720 -118750
rect 70610 -118855 70720 -118850
rect 72110 -118750 72220 -118745
rect 72110 -118850 72120 -118750
rect 72210 -118850 72220 -118750
rect 72110 -118855 72220 -118850
rect 73610 -118750 73720 -118745
rect 73610 -118850 73620 -118750
rect 73710 -118850 73720 -118750
rect 73610 -118855 73720 -118850
rect 75110 -118750 75220 -118745
rect 75110 -118850 75120 -118750
rect 75210 -118850 75220 -118750
rect 75110 -118855 75220 -118850
rect 76610 -118750 76720 -118745
rect 76610 -118850 76620 -118750
rect 76710 -118850 76720 -118750
rect 76610 -118855 76720 -118850
rect 78110 -118750 78220 -118745
rect 78110 -118850 78120 -118750
rect 78210 -118850 78220 -118750
rect 78110 -118855 78220 -118850
rect 79610 -118750 79720 -118745
rect 79610 -118850 79620 -118750
rect 79710 -118850 79720 -118750
rect 79610 -118855 79720 -118850
rect 81110 -118750 81220 -118745
rect 81110 -118850 81120 -118750
rect 81210 -118850 81220 -118750
rect 81110 -118855 81220 -118850
rect 82610 -118750 82720 -118745
rect 82610 -118850 82620 -118750
rect 82710 -118850 82720 -118750
rect 82610 -118855 82720 -118850
rect 84110 -118750 84220 -118745
rect 84110 -118850 84120 -118750
rect 84210 -118850 84220 -118750
rect 84110 -118855 84220 -118850
rect 85610 -118750 85720 -118745
rect 85610 -118850 85620 -118750
rect 85710 -118850 85720 -118750
rect 85610 -118855 85720 -118850
rect 87110 -118750 87220 -118745
rect 87110 -118850 87120 -118750
rect 87210 -118850 87220 -118750
rect 87110 -118855 87220 -118850
rect 88610 -118750 88720 -118745
rect 88610 -118850 88620 -118750
rect 88710 -118850 88720 -118750
rect 88610 -118855 88720 -118850
rect 90110 -118750 90220 -118745
rect 90110 -118850 90120 -118750
rect 90210 -118850 90220 -118750
rect 90110 -118855 90220 -118850
rect 91610 -118750 91720 -118745
rect 91610 -118850 91620 -118750
rect 91710 -118850 91720 -118750
rect 91610 -118855 91720 -118850
rect 93110 -118750 93220 -118745
rect 93110 -118850 93120 -118750
rect 93210 -118850 93220 -118750
rect 93110 -118855 93220 -118850
rect 94610 -118750 94720 -118745
rect 94610 -118850 94620 -118750
rect 94710 -118850 94720 -118750
rect 94610 -118855 94720 -118850
rect 96110 -118750 96220 -118745
rect 96110 -118850 96120 -118750
rect 96210 -118850 96220 -118750
rect 96110 -118855 96220 -118850
rect 97610 -118750 97720 -118745
rect 97610 -118850 97620 -118750
rect 97710 -118850 97720 -118750
rect 97610 -118855 97720 -118850
rect 99110 -118750 99220 -118745
rect 99110 -118850 99120 -118750
rect 99210 -118850 99220 -118750
rect 99110 -118855 99220 -118850
rect 100610 -118750 100720 -118745
rect 100610 -118850 100620 -118750
rect 100710 -118850 100720 -118750
rect 100610 -118855 100720 -118850
rect 102110 -118750 102220 -118745
rect 102110 -118850 102120 -118750
rect 102210 -118850 102220 -118750
rect 102110 -118855 102220 -118850
rect 103610 -118750 103720 -118745
rect 103610 -118850 103620 -118750
rect 103710 -118850 103720 -118750
rect 103610 -118855 103720 -118850
rect 105110 -118750 105220 -118745
rect 105110 -118850 105120 -118750
rect 105210 -118850 105220 -118750
rect 105110 -118855 105220 -118850
rect 106610 -118750 106720 -118745
rect 106610 -118850 106620 -118750
rect 106710 -118850 106720 -118750
rect 106610 -118855 106720 -118850
rect 108110 -118750 108220 -118745
rect 108110 -118850 108120 -118750
rect 108210 -118850 108220 -118750
rect 108110 -118855 108220 -118850
rect 109610 -118750 109720 -118745
rect 109610 -118850 109620 -118750
rect 109710 -118850 109720 -118750
rect 109610 -118855 109720 -118850
rect 111110 -118750 111220 -118745
rect 111110 -118850 111120 -118750
rect 111210 -118850 111220 -118750
rect 111110 -118855 111220 -118850
rect 112610 -118750 112720 -118745
rect 112610 -118850 112620 -118750
rect 112710 -118850 112720 -118750
rect 112610 -118855 112720 -118850
rect 114110 -118750 114220 -118745
rect 114110 -118850 114120 -118750
rect 114210 -118850 114220 -118750
rect 114110 -118855 114220 -118850
rect 115610 -118750 115720 -118745
rect 115610 -118850 115620 -118750
rect 115710 -118850 115720 -118750
rect 115610 -118855 115720 -118850
rect 117110 -118750 117220 -118745
rect 117110 -118850 117120 -118750
rect 117210 -118850 117220 -118750
rect 117110 -118855 117220 -118850
rect 118610 -118750 118720 -118745
rect 118610 -118850 118620 -118750
rect 118710 -118850 118720 -118750
rect 118610 -118855 118720 -118850
rect 270 -118960 120370 -118950
rect 270 -119040 280 -118960
rect 270 -119050 120370 -119040
<< via1 >>
rect -960 1680 -450 1725
rect 25 1680 70 1725
rect 1525 1680 1570 1725
rect 3025 1680 3070 1725
rect 4525 1680 4570 1725
rect 6025 1680 6070 1725
rect 7525 1680 7570 1725
rect 9025 1680 9070 1725
rect 10525 1680 10570 1725
rect 12025 1680 12070 1725
rect 13525 1680 13570 1725
rect 15025 1680 15070 1725
rect 16525 1680 16570 1725
rect 18025 1680 18070 1725
rect 19525 1680 19570 1725
rect 21025 1680 21070 1725
rect 22525 1680 22570 1725
rect 24025 1680 24070 1725
rect 25525 1680 25570 1725
rect 27025 1680 27070 1725
rect 28525 1680 28570 1725
rect 30025 1680 30070 1725
rect 31525 1680 31570 1725
rect 33025 1680 33070 1725
rect 34525 1680 34570 1725
rect 36025 1680 36070 1725
rect 37525 1680 37570 1725
rect 39025 1680 39070 1725
rect 40525 1680 40570 1725
rect 42025 1680 42070 1725
rect 43525 1680 43570 1725
rect 45025 1680 45070 1725
rect 46525 1680 46570 1725
rect 48025 1680 48070 1725
rect 49525 1680 49570 1725
rect 51025 1680 51070 1725
rect 52525 1680 52570 1725
rect 54025 1680 54070 1725
rect 55525 1680 55570 1725
rect 57025 1680 57070 1725
rect 58525 1680 58570 1725
rect 60025 1680 60070 1725
rect 61525 1680 61570 1725
rect 63025 1680 63070 1725
rect 64525 1680 64570 1725
rect 66025 1680 66070 1725
rect 67525 1680 67570 1725
rect 69025 1680 69070 1725
rect 70525 1680 70570 1725
rect 72025 1680 72070 1725
rect 73525 1680 73570 1725
rect 75025 1680 75070 1725
rect 76525 1680 76570 1725
rect 78025 1680 78070 1725
rect 79525 1680 79570 1725
rect 81025 1680 81070 1725
rect 82525 1680 82570 1725
rect 84025 1680 84070 1725
rect 85525 1680 85570 1725
rect 87025 1680 87070 1725
rect 88525 1680 88570 1725
rect 90025 1680 90070 1725
rect 91525 1680 91570 1725
rect 93025 1680 93070 1725
rect 94525 1680 94570 1725
rect 96025 1680 96070 1725
rect 97525 1680 97570 1725
rect 99025 1680 99070 1725
rect 100525 1680 100570 1725
rect 102025 1680 102070 1725
rect 103525 1680 103570 1725
rect 105025 1680 105070 1725
rect 106525 1680 106570 1725
rect 108025 1680 108070 1725
rect 109525 1680 109570 1725
rect 111025 1680 111070 1725
rect 112525 1680 112570 1725
rect 114025 1680 114070 1725
rect 115525 1680 115570 1725
rect 117025 1680 117070 1725
rect 118525 1680 118570 1725
rect -790 745 -590 780
rect -270 745 -130 780
rect -790 -755 -590 -720
rect -270 -755 -130 -720
rect -790 -2255 -590 -2220
rect -270 -2255 -130 -2220
rect -790 -3755 -590 -3720
rect -270 -3755 -130 -3720
rect -790 -5255 -590 -5220
rect -270 -5255 -130 -5220
rect -790 -6755 -590 -6720
rect -270 -6755 -130 -6720
rect -790 -8255 -590 -8220
rect -270 -8255 -130 -8220
rect -790 -9755 -590 -9720
rect -270 -9755 -130 -9720
rect -790 -11255 -590 -11220
rect -270 -11255 -130 -11220
rect -790 -12755 -590 -12720
rect -270 -12755 -130 -12720
rect -790 -14255 -590 -14220
rect -270 -14255 -130 -14220
rect -790 -15755 -590 -15720
rect -270 -15755 -130 -15720
rect -790 -17255 -590 -17220
rect -270 -17255 -130 -17220
rect -790 -18755 -590 -18720
rect -270 -18755 -130 -18720
rect -790 -20255 -590 -20220
rect -270 -20255 -130 -20220
rect -790 -21755 -590 -21720
rect -270 -21755 -130 -21720
rect -790 -23255 -590 -23220
rect -270 -23255 -130 -23220
rect -790 -24755 -590 -24720
rect -270 -24755 -130 -24720
rect -790 -26255 -590 -26220
rect -270 -26255 -130 -26220
rect -790 -27755 -590 -27720
rect -270 -27755 -130 -27720
rect -790 -29255 -590 -29220
rect -270 -29255 -130 -29220
rect -790 -30755 -590 -30720
rect -270 -30755 -130 -30720
rect -790 -32255 -590 -32220
rect -270 -32255 -130 -32220
rect -790 -33755 -590 -33720
rect -270 -33755 -130 -33720
rect -790 -35255 -590 -35220
rect -270 -35255 -130 -35220
rect -790 -36755 -590 -36720
rect -270 -36755 -130 -36720
rect -790 -38255 -590 -38220
rect -270 -38255 -130 -38220
rect -790 -39755 -590 -39720
rect -270 -39755 -130 -39720
rect -790 -41255 -590 -41220
rect -270 -41255 -130 -41220
rect -790 -42755 -590 -42720
rect -270 -42755 -130 -42720
rect -790 -44255 -590 -44220
rect -270 -44255 -130 -44220
rect -790 -45755 -590 -45720
rect -270 -45755 -130 -45720
rect -790 -47255 -590 -47220
rect -270 -47255 -130 -47220
rect -790 -48755 -590 -48720
rect -270 -48755 -130 -48720
rect -790 -50255 -590 -50220
rect -270 -50255 -130 -50220
rect -790 -51755 -590 -51720
rect -270 -51755 -130 -51720
rect -790 -53255 -590 -53220
rect -270 -53255 -130 -53220
rect -790 -54755 -590 -54720
rect -270 -54755 -130 -54720
rect -790 -56255 -590 -56220
rect -270 -56255 -130 -56220
rect -790 -57755 -590 -57720
rect -270 -57755 -130 -57720
rect -790 -59255 -590 -59220
rect -270 -59255 -130 -59220
rect -790 -60755 -590 -60720
rect -270 -60755 -130 -60720
rect -790 -62255 -590 -62220
rect -270 -62255 -130 -62220
rect -790 -63755 -590 -63720
rect -270 -63755 -130 -63720
rect -790 -65255 -590 -65220
rect -270 -65255 -130 -65220
rect -790 -66755 -590 -66720
rect -270 -66755 -130 -66720
rect -790 -68255 -590 -68220
rect -270 -68255 -130 -68220
rect -790 -69755 -590 -69720
rect -270 -69755 -130 -69720
rect -790 -71255 -590 -71220
rect -270 -71255 -130 -71220
rect -790 -72755 -590 -72720
rect -270 -72755 -130 -72720
rect -790 -74255 -590 -74220
rect -270 -74255 -130 -74220
rect -790 -75755 -590 -75720
rect -270 -75755 -130 -75720
rect -790 -77255 -590 -77220
rect -270 -77255 -130 -77220
rect -790 -78755 -590 -78720
rect -270 -78755 -130 -78720
rect -790 -80255 -590 -80220
rect -270 -80255 -130 -80220
rect -790 -81755 -590 -81720
rect -270 -81755 -130 -81720
rect -790 -83255 -590 -83220
rect -270 -83255 -130 -83220
rect -790 -84755 -590 -84720
rect -270 -84755 -130 -84720
rect -790 -86255 -590 -86220
rect -270 -86255 -130 -86220
rect -790 -87755 -590 -87720
rect -270 -87755 -130 -87720
rect -790 -89255 -590 -89220
rect -270 -89255 -130 -89220
rect -790 -90755 -590 -90720
rect -270 -90755 -130 -90720
rect -790 -92255 -590 -92220
rect -270 -92255 -130 -92220
rect -790 -93755 -590 -93720
rect -270 -93755 -130 -93720
rect -790 -95255 -590 -95220
rect -270 -95255 -130 -95220
rect -790 -96755 -590 -96720
rect -270 -96755 -130 -96720
rect -790 -98255 -590 -98220
rect -270 -98255 -130 -98220
rect -790 -99755 -590 -99720
rect -270 -99755 -130 -99720
rect -790 -101255 -590 -101220
rect -270 -101255 -130 -101220
rect -790 -102755 -590 -102720
rect -270 -102755 -130 -102720
rect -790 -104255 -590 -104220
rect -270 -104255 -130 -104220
rect -790 -105755 -590 -105720
rect -270 -105755 -130 -105720
rect -790 -107255 -590 -107220
rect -270 -107255 -130 -107220
rect -790 -108755 -590 -108720
rect -270 -108755 -130 -108720
rect -790 -110255 -590 -110220
rect -270 -110255 -130 -110220
rect -790 -111755 -590 -111720
rect -270 -111755 -130 -111720
rect -790 -113255 -590 -113220
rect -270 -113255 -130 -113220
rect -790 -114755 -590 -114720
rect -270 -114755 -130 -114720
rect -790 -116255 -590 -116220
rect -270 -116255 -130 -116220
rect -790 -117755 -590 -117720
rect -270 -117755 -130 -117720
rect 280 -118600 1060 -118565
rect 1780 -118600 2560 -118565
rect 3280 -118600 4060 -118565
rect 4780 -118600 5560 -118565
rect 6280 -118600 7060 -118565
rect 7780 -118600 8560 -118565
rect 9280 -118600 10060 -118565
rect 10780 -118600 11560 -118565
rect 12280 -118600 13060 -118565
rect 13780 -118600 14560 -118565
rect 15280 -118600 16060 -118565
rect 16780 -118600 17560 -118565
rect 18280 -118600 19060 -118565
rect 19780 -118600 20560 -118565
rect 21280 -118600 22060 -118565
rect 22780 -118600 23560 -118565
rect 24280 -118600 25060 -118565
rect 25780 -118600 26560 -118565
rect 27280 -118600 28060 -118565
rect 28780 -118600 29560 -118565
rect 30280 -118600 31060 -118565
rect 31780 -118600 32560 -118565
rect 33280 -118600 34060 -118565
rect 34780 -118600 35560 -118565
rect 36280 -118600 37060 -118565
rect 37780 -118600 38560 -118565
rect 39280 -118600 40060 -118565
rect 40780 -118600 41560 -118565
rect 42280 -118600 43060 -118565
rect 43780 -118600 44560 -118565
rect 45280 -118600 46060 -118565
rect 46780 -118600 47560 -118565
rect 48280 -118600 49060 -118565
rect 49780 -118600 50560 -118565
rect 51280 -118600 52060 -118565
rect 52780 -118600 53560 -118565
rect 54280 -118600 55060 -118565
rect 55780 -118600 56560 -118565
rect 57280 -118600 58060 -118565
rect 58780 -118600 59560 -118565
rect 60280 -118600 61060 -118565
rect 61780 -118600 62560 -118565
rect 63280 -118600 64060 -118565
rect 64780 -118600 65560 -118565
rect 66280 -118600 67060 -118565
rect 67780 -118600 68560 -118565
rect 69280 -118600 70060 -118565
rect 70780 -118600 71560 -118565
rect 72280 -118600 73060 -118565
rect 73780 -118600 74560 -118565
rect 75280 -118600 76060 -118565
rect 76780 -118600 77560 -118565
rect 78280 -118600 79060 -118565
rect 79780 -118600 80560 -118565
rect 81280 -118600 82060 -118565
rect 82780 -118600 83560 -118565
rect 84280 -118600 85060 -118565
rect 85780 -118600 86560 -118565
rect 87280 -118600 88060 -118565
rect 88780 -118600 89560 -118565
rect 90280 -118600 91060 -118565
rect 91780 -118600 92560 -118565
rect 93280 -118600 94060 -118565
rect 94780 -118600 95560 -118565
rect 96280 -118600 97060 -118565
rect 97780 -118600 98560 -118565
rect 99280 -118600 100060 -118565
rect 100780 -118600 101560 -118565
rect 102280 -118600 103060 -118565
rect 103780 -118600 104560 -118565
rect 105280 -118600 106060 -118565
rect 106780 -118600 107560 -118565
rect 108280 -118600 109060 -118565
rect 109780 -118600 110560 -118565
rect 111280 -118600 112060 -118565
rect 112780 -118600 113560 -118565
rect 114280 -118600 115060 -118565
rect 115780 -118600 116560 -118565
rect 117280 -118600 118060 -118565
rect 118780 -118600 119560 -118565
rect 120 -118850 210 -118750
rect 1620 -118850 1710 -118750
rect 3120 -118850 3210 -118750
rect 4620 -118850 4710 -118750
rect 6120 -118850 6210 -118750
rect 7620 -118850 7710 -118750
rect 9120 -118850 9210 -118750
rect 10620 -118850 10710 -118750
rect 12120 -118850 12210 -118750
rect 13620 -118850 13710 -118750
rect 15120 -118850 15210 -118750
rect 16620 -118850 16710 -118750
rect 18120 -118850 18210 -118750
rect 19620 -118850 19710 -118750
rect 21120 -118850 21210 -118750
rect 22620 -118850 22710 -118750
rect 24120 -118850 24210 -118750
rect 25620 -118850 25710 -118750
rect 27120 -118850 27210 -118750
rect 28620 -118850 28710 -118750
rect 30120 -118850 30210 -118750
rect 31620 -118850 31710 -118750
rect 33120 -118850 33210 -118750
rect 34620 -118850 34710 -118750
rect 36120 -118850 36210 -118750
rect 37620 -118850 37710 -118750
rect 39120 -118850 39210 -118750
rect 40620 -118850 40710 -118750
rect 42120 -118850 42210 -118750
rect 43620 -118850 43710 -118750
rect 45120 -118850 45210 -118750
rect 46620 -118850 46710 -118750
rect 48120 -118850 48210 -118750
rect 49620 -118850 49710 -118750
rect 51120 -118850 51210 -118750
rect 52620 -118850 52710 -118750
rect 54120 -118850 54210 -118750
rect 55620 -118850 55710 -118750
rect 57120 -118850 57210 -118750
rect 58620 -118850 58710 -118750
rect 60120 -118850 60210 -118750
rect 61620 -118850 61710 -118750
rect 63120 -118850 63210 -118750
rect 64620 -118850 64710 -118750
rect 66120 -118850 66210 -118750
rect 67620 -118850 67710 -118750
rect 69120 -118850 69210 -118750
rect 70620 -118850 70710 -118750
rect 72120 -118850 72210 -118750
rect 73620 -118850 73710 -118750
rect 75120 -118850 75210 -118750
rect 76620 -118850 76710 -118750
rect 78120 -118850 78210 -118750
rect 79620 -118850 79710 -118750
rect 81120 -118850 81210 -118750
rect 82620 -118850 82710 -118750
rect 84120 -118850 84210 -118750
rect 85620 -118850 85710 -118750
rect 87120 -118850 87210 -118750
rect 88620 -118850 88710 -118750
rect 90120 -118850 90210 -118750
rect 91620 -118850 91710 -118750
rect 93120 -118850 93210 -118750
rect 94620 -118850 94710 -118750
rect 96120 -118850 96210 -118750
rect 97620 -118850 97710 -118750
rect 99120 -118850 99210 -118750
rect 100620 -118850 100710 -118750
rect 102120 -118850 102210 -118750
rect 103620 -118850 103710 -118750
rect 105120 -118850 105210 -118750
rect 106620 -118850 106710 -118750
rect 108120 -118850 108210 -118750
rect 109620 -118850 109710 -118750
rect 111120 -118850 111210 -118750
rect 112620 -118850 112710 -118750
rect 114120 -118850 114210 -118750
rect 115620 -118850 115710 -118750
rect 117120 -118850 117210 -118750
rect 118620 -118850 118710 -118750
rect 280 -118990 1060 -118960
rect 1060 -118990 1780 -118960
rect 1780 -118990 2560 -118960
rect 2560 -118990 3280 -118960
rect 3280 -118990 4060 -118960
rect 4060 -118990 4780 -118960
rect 4780 -118990 5560 -118960
rect 5560 -118990 6280 -118960
rect 6280 -118990 7060 -118960
rect 7060 -118990 7780 -118960
rect 7780 -118990 8560 -118960
rect 8560 -118990 9280 -118960
rect 9280 -118990 10060 -118960
rect 10060 -118990 10780 -118960
rect 10780 -118990 11560 -118960
rect 11560 -118990 12280 -118960
rect 12280 -118990 13060 -118960
rect 13060 -118990 13780 -118960
rect 13780 -118990 14560 -118960
rect 14560 -118990 15280 -118960
rect 15280 -118990 16060 -118960
rect 16060 -118990 16780 -118960
rect 16780 -118990 17560 -118960
rect 17560 -118990 18280 -118960
rect 18280 -118990 19060 -118960
rect 19060 -118990 19780 -118960
rect 19780 -118990 20560 -118960
rect 20560 -118990 21280 -118960
rect 21280 -118990 22060 -118960
rect 22060 -118990 22780 -118960
rect 22780 -118990 23560 -118960
rect 23560 -118990 24280 -118960
rect 24280 -118990 25060 -118960
rect 25060 -118990 25780 -118960
rect 25780 -118990 26560 -118960
rect 26560 -118990 27280 -118960
rect 27280 -118990 28060 -118960
rect 28060 -118990 28780 -118960
rect 28780 -118990 29560 -118960
rect 29560 -118990 30280 -118960
rect 30280 -118990 31060 -118960
rect 31060 -118990 31780 -118960
rect 31780 -118990 32560 -118960
rect 32560 -118990 33280 -118960
rect 33280 -118990 34060 -118960
rect 34060 -118990 34780 -118960
rect 34780 -118990 35560 -118960
rect 35560 -118990 36280 -118960
rect 36280 -118990 37060 -118960
rect 37060 -118990 37780 -118960
rect 37780 -118990 38560 -118960
rect 38560 -118990 39280 -118960
rect 39280 -118990 40060 -118960
rect 40060 -118990 40780 -118960
rect 40780 -118990 41560 -118960
rect 41560 -118990 42280 -118960
rect 42280 -118990 43060 -118960
rect 43060 -118990 43780 -118960
rect 43780 -118990 44560 -118960
rect 44560 -118990 45280 -118960
rect 45280 -118990 46060 -118960
rect 46060 -118990 46780 -118960
rect 46780 -118990 47560 -118960
rect 47560 -118990 48280 -118960
rect 48280 -118990 49060 -118960
rect 49060 -118990 49780 -118960
rect 49780 -118990 50560 -118960
rect 50560 -118990 51280 -118960
rect 51280 -118990 52060 -118960
rect 52060 -118990 52780 -118960
rect 52780 -118990 53560 -118960
rect 53560 -118990 54280 -118960
rect 54280 -118990 55060 -118960
rect 55060 -118990 55780 -118960
rect 55780 -118990 56560 -118960
rect 56560 -118990 57280 -118960
rect 57280 -118990 58060 -118960
rect 58060 -118990 58780 -118960
rect 58780 -118990 59560 -118960
rect 59560 -118990 60280 -118960
rect 60280 -118990 61060 -118960
rect 61060 -118990 61780 -118960
rect 61780 -118990 62560 -118960
rect 62560 -118990 63280 -118960
rect 63280 -118990 64060 -118960
rect 64060 -118990 64780 -118960
rect 64780 -118990 65560 -118960
rect 65560 -118990 66280 -118960
rect 66280 -118990 67060 -118960
rect 67060 -118990 67780 -118960
rect 67780 -118990 68560 -118960
rect 68560 -118990 69280 -118960
rect 69280 -118990 70060 -118960
rect 70060 -118990 70780 -118960
rect 70780 -118990 71560 -118960
rect 71560 -118990 72280 -118960
rect 72280 -118990 73060 -118960
rect 73060 -118990 73780 -118960
rect 73780 -118990 74560 -118960
rect 74560 -118990 75280 -118960
rect 75280 -118990 76060 -118960
rect 76060 -118990 76780 -118960
rect 76780 -118990 77560 -118960
rect 77560 -118990 78280 -118960
rect 78280 -118990 79060 -118960
rect 79060 -118990 79780 -118960
rect 79780 -118990 80560 -118960
rect 80560 -118990 81280 -118960
rect 81280 -118990 82060 -118960
rect 82060 -118990 82780 -118960
rect 82780 -118990 83560 -118960
rect 83560 -118990 84280 -118960
rect 84280 -118990 85060 -118960
rect 85060 -118990 85780 -118960
rect 85780 -118990 86560 -118960
rect 86560 -118990 87280 -118960
rect 87280 -118990 88060 -118960
rect 88060 -118990 88780 -118960
rect 88780 -118990 89560 -118960
rect 89560 -118990 90280 -118960
rect 90280 -118990 91060 -118960
rect 91060 -118990 91780 -118960
rect 91780 -118990 92560 -118960
rect 92560 -118990 93280 -118960
rect 93280 -118990 94060 -118960
rect 94060 -118990 94780 -118960
rect 94780 -118990 95560 -118960
rect 95560 -118990 96280 -118960
rect 96280 -118990 97060 -118960
rect 97060 -118990 97780 -118960
rect 97780 -118990 98560 -118960
rect 98560 -118990 99280 -118960
rect 99280 -118990 100060 -118960
rect 100060 -118990 100780 -118960
rect 100780 -118990 101560 -118960
rect 101560 -118990 102280 -118960
rect 102280 -118990 103060 -118960
rect 103060 -118990 103780 -118960
rect 103780 -118990 104560 -118960
rect 104560 -118990 105280 -118960
rect 105280 -118990 106060 -118960
rect 106060 -118990 106780 -118960
rect 106780 -118990 107560 -118960
rect 107560 -118990 108280 -118960
rect 108280 -118990 109060 -118960
rect 109060 -118990 109780 -118960
rect 109780 -118990 110560 -118960
rect 110560 -118990 111280 -118960
rect 111280 -118990 112060 -118960
rect 112060 -118990 112780 -118960
rect 112780 -118990 113560 -118960
rect 113560 -118990 114280 -118960
rect 114280 -118990 115060 -118960
rect 115060 -118990 115780 -118960
rect 115780 -118990 116560 -118960
rect 116560 -118990 117280 -118960
rect 117280 -118990 118060 -118960
rect 118060 -118990 118780 -118960
rect 118780 -118990 119560 -118960
rect 119560 -118990 120370 -118960
rect 280 -119040 120370 -118990
<< metal2 >>
rect 0 2020 120000 2075
rect -1500 1725 -445 1730
rect -1500 1680 -960 1725
rect -450 1680 -445 1725
rect -1500 1675 -445 1680
rect -1500 780 -500 785
rect -1500 745 -790 780
rect -590 745 -500 780
rect -1500 740 -500 745
rect -375 115 -320 2000
rect 240 1825 295 1830
rect 240 1780 245 1825
rect 290 1780 295 1825
rect 240 1775 295 1780
rect 20 1725 75 1730
rect 20 1680 25 1725
rect 70 1680 75 1725
rect 20 1675 75 1680
rect 30 1500 65 1675
rect 250 1500 285 1775
rect 510 1500 545 2020
rect 1740 1825 1795 1830
rect 1740 1780 1745 1825
rect 1790 1780 1795 1825
rect 1740 1775 1795 1780
rect 1520 1725 1575 1730
rect 1520 1680 1525 1725
rect 1570 1680 1575 1725
rect 1520 1675 1575 1680
rect 1530 1500 1565 1675
rect 1750 1500 1785 1775
rect 2010 1500 2045 2020
rect 3240 1825 3295 1830
rect 3240 1780 3245 1825
rect 3290 1780 3295 1825
rect 3240 1775 3295 1780
rect 3020 1725 3075 1730
rect 3020 1680 3025 1725
rect 3070 1680 3075 1725
rect 3020 1675 3075 1680
rect 3030 1500 3065 1675
rect 3250 1500 3285 1775
rect 3510 1500 3545 2020
rect 4740 1825 4795 1830
rect 4740 1780 4745 1825
rect 4790 1780 4795 1825
rect 4740 1775 4795 1780
rect 4520 1725 4575 1730
rect 4520 1680 4525 1725
rect 4570 1680 4575 1725
rect 4520 1675 4575 1680
rect 4530 1500 4565 1675
rect 4750 1500 4785 1775
rect 5010 1500 5045 2020
rect 6240 1825 6295 1830
rect 6240 1780 6245 1825
rect 6290 1780 6295 1825
rect 6240 1775 6295 1780
rect 6020 1725 6075 1730
rect 6020 1680 6025 1725
rect 6070 1680 6075 1725
rect 6020 1675 6075 1680
rect 6030 1500 6065 1675
rect 6250 1500 6285 1775
rect 6510 1500 6545 2020
rect 7740 1825 7795 1830
rect 7740 1780 7745 1825
rect 7790 1780 7795 1825
rect 7740 1775 7795 1780
rect 7520 1725 7575 1730
rect 7520 1680 7525 1725
rect 7570 1680 7575 1725
rect 7520 1675 7575 1680
rect 7530 1500 7565 1675
rect 7750 1500 7785 1775
rect 8010 1500 8045 2020
rect 9240 1825 9295 1830
rect 9240 1780 9245 1825
rect 9290 1780 9295 1825
rect 9240 1775 9295 1780
rect 9020 1725 9075 1730
rect 9020 1680 9025 1725
rect 9070 1680 9075 1725
rect 9020 1675 9075 1680
rect 9030 1500 9065 1675
rect 9250 1500 9285 1775
rect 9510 1500 9545 2020
rect 10740 1825 10795 1830
rect 10740 1780 10745 1825
rect 10790 1780 10795 1825
rect 10740 1775 10795 1780
rect 10520 1725 10575 1730
rect 10520 1680 10525 1725
rect 10570 1680 10575 1725
rect 10520 1675 10575 1680
rect 10530 1500 10565 1675
rect 10750 1500 10785 1775
rect 11010 1500 11045 2020
rect 12240 1825 12295 1830
rect 12240 1780 12245 1825
rect 12290 1780 12295 1825
rect 12240 1775 12295 1780
rect 12020 1725 12075 1730
rect 12020 1680 12025 1725
rect 12070 1680 12075 1725
rect 12020 1675 12075 1680
rect 12030 1500 12065 1675
rect 12250 1500 12285 1775
rect 12510 1500 12545 2020
rect 13740 1825 13795 1830
rect 13740 1780 13745 1825
rect 13790 1780 13795 1825
rect 13740 1775 13795 1780
rect 13520 1725 13575 1730
rect 13520 1680 13525 1725
rect 13570 1680 13575 1725
rect 13520 1675 13575 1680
rect 13530 1500 13565 1675
rect 13750 1500 13785 1775
rect 14010 1500 14045 2020
rect 15240 1825 15295 1830
rect 15240 1780 15245 1825
rect 15290 1780 15295 1825
rect 15240 1775 15295 1780
rect 15020 1725 15075 1730
rect 15020 1680 15025 1725
rect 15070 1680 15075 1725
rect 15020 1675 15075 1680
rect 15030 1500 15065 1675
rect 15250 1500 15285 1775
rect 15510 1500 15545 2020
rect 16740 1825 16795 1830
rect 16740 1780 16745 1825
rect 16790 1780 16795 1825
rect 16740 1775 16795 1780
rect 16520 1725 16575 1730
rect 16520 1680 16525 1725
rect 16570 1680 16575 1725
rect 16520 1675 16575 1680
rect 16530 1500 16565 1675
rect 16750 1500 16785 1775
rect 17010 1500 17045 2020
rect 18240 1825 18295 1830
rect 18240 1780 18245 1825
rect 18290 1780 18295 1825
rect 18240 1775 18295 1780
rect 18020 1725 18075 1730
rect 18020 1680 18025 1725
rect 18070 1680 18075 1725
rect 18020 1675 18075 1680
rect 18030 1500 18065 1675
rect 18250 1500 18285 1775
rect 18510 1500 18545 2020
rect 19740 1825 19795 1830
rect 19740 1780 19745 1825
rect 19790 1780 19795 1825
rect 19740 1775 19795 1780
rect 19520 1725 19575 1730
rect 19520 1680 19525 1725
rect 19570 1680 19575 1725
rect 19520 1675 19575 1680
rect 19530 1500 19565 1675
rect 19750 1500 19785 1775
rect 20010 1500 20045 2020
rect 21240 1825 21295 1830
rect 21240 1780 21245 1825
rect 21290 1780 21295 1825
rect 21240 1775 21295 1780
rect 21020 1725 21075 1730
rect 21020 1680 21025 1725
rect 21070 1680 21075 1725
rect 21020 1675 21075 1680
rect 21030 1500 21065 1675
rect 21250 1500 21285 1775
rect 21510 1500 21545 2020
rect 22740 1825 22795 1830
rect 22740 1780 22745 1825
rect 22790 1780 22795 1825
rect 22740 1775 22795 1780
rect 22520 1725 22575 1730
rect 22520 1680 22525 1725
rect 22570 1680 22575 1725
rect 22520 1675 22575 1680
rect 22530 1500 22565 1675
rect 22750 1500 22785 1775
rect 23010 1500 23045 2020
rect 24240 1825 24295 1830
rect 24240 1780 24245 1825
rect 24290 1780 24295 1825
rect 24240 1775 24295 1780
rect 24020 1725 24075 1730
rect 24020 1680 24025 1725
rect 24070 1680 24075 1725
rect 24020 1675 24075 1680
rect 24030 1500 24065 1675
rect 24250 1500 24285 1775
rect 24510 1500 24545 2020
rect 25740 1825 25795 1830
rect 25740 1780 25745 1825
rect 25790 1780 25795 1825
rect 25740 1775 25795 1780
rect 25520 1725 25575 1730
rect 25520 1680 25525 1725
rect 25570 1680 25575 1725
rect 25520 1675 25575 1680
rect 25530 1500 25565 1675
rect 25750 1500 25785 1775
rect 26010 1500 26045 2020
rect 27240 1825 27295 1830
rect 27240 1780 27245 1825
rect 27290 1780 27295 1825
rect 27240 1775 27295 1780
rect 27020 1725 27075 1730
rect 27020 1680 27025 1725
rect 27070 1680 27075 1725
rect 27020 1675 27075 1680
rect 27030 1500 27065 1675
rect 27250 1500 27285 1775
rect 27510 1500 27545 2020
rect 28740 1825 28795 1830
rect 28740 1780 28745 1825
rect 28790 1780 28795 1825
rect 28740 1775 28795 1780
rect 28520 1725 28575 1730
rect 28520 1680 28525 1725
rect 28570 1680 28575 1725
rect 28520 1675 28575 1680
rect 28530 1500 28565 1675
rect 28750 1500 28785 1775
rect 29010 1500 29045 2020
rect 30240 1825 30295 1830
rect 30240 1780 30245 1825
rect 30290 1780 30295 1825
rect 30240 1775 30295 1780
rect 30020 1725 30075 1730
rect 30020 1680 30025 1725
rect 30070 1680 30075 1725
rect 30020 1675 30075 1680
rect 30030 1500 30065 1675
rect 30250 1500 30285 1775
rect 30510 1500 30545 2020
rect 31740 1825 31795 1830
rect 31740 1780 31745 1825
rect 31790 1780 31795 1825
rect 31740 1775 31795 1780
rect 31520 1725 31575 1730
rect 31520 1680 31525 1725
rect 31570 1680 31575 1725
rect 31520 1675 31575 1680
rect 31530 1500 31565 1675
rect 31750 1500 31785 1775
rect 32010 1500 32045 2020
rect 33240 1825 33295 1830
rect 33240 1780 33245 1825
rect 33290 1780 33295 1825
rect 33240 1775 33295 1780
rect 33020 1725 33075 1730
rect 33020 1680 33025 1725
rect 33070 1680 33075 1725
rect 33020 1675 33075 1680
rect 33030 1500 33065 1675
rect 33250 1500 33285 1775
rect 33510 1500 33545 2020
rect 34740 1825 34795 1830
rect 34740 1780 34745 1825
rect 34790 1780 34795 1825
rect 34740 1775 34795 1780
rect 34520 1725 34575 1730
rect 34520 1680 34525 1725
rect 34570 1680 34575 1725
rect 34520 1675 34575 1680
rect 34530 1500 34565 1675
rect 34750 1500 34785 1775
rect 35010 1500 35045 2020
rect 36240 1825 36295 1830
rect 36240 1780 36245 1825
rect 36290 1780 36295 1825
rect 36240 1775 36295 1780
rect 36020 1725 36075 1730
rect 36020 1680 36025 1725
rect 36070 1680 36075 1725
rect 36020 1675 36075 1680
rect 36030 1500 36065 1675
rect 36250 1500 36285 1775
rect 36510 1500 36545 2020
rect 37740 1825 37795 1830
rect 37740 1780 37745 1825
rect 37790 1780 37795 1825
rect 37740 1775 37795 1780
rect 37520 1725 37575 1730
rect 37520 1680 37525 1725
rect 37570 1680 37575 1725
rect 37520 1675 37575 1680
rect 37530 1500 37565 1675
rect 37750 1500 37785 1775
rect 38010 1500 38045 2020
rect 39240 1825 39295 1830
rect 39240 1780 39245 1825
rect 39290 1780 39295 1825
rect 39240 1775 39295 1780
rect 39020 1725 39075 1730
rect 39020 1680 39025 1725
rect 39070 1680 39075 1725
rect 39020 1675 39075 1680
rect 39030 1500 39065 1675
rect 39250 1500 39285 1775
rect 39510 1500 39545 2020
rect 40740 1825 40795 1830
rect 40740 1780 40745 1825
rect 40790 1780 40795 1825
rect 40740 1775 40795 1780
rect 40520 1725 40575 1730
rect 40520 1680 40525 1725
rect 40570 1680 40575 1725
rect 40520 1675 40575 1680
rect 40530 1500 40565 1675
rect 40750 1500 40785 1775
rect 41010 1500 41045 2020
rect 42240 1825 42295 1830
rect 42240 1780 42245 1825
rect 42290 1780 42295 1825
rect 42240 1775 42295 1780
rect 42020 1725 42075 1730
rect 42020 1680 42025 1725
rect 42070 1680 42075 1725
rect 42020 1675 42075 1680
rect 42030 1500 42065 1675
rect 42250 1500 42285 1775
rect 42510 1500 42545 2020
rect 43740 1825 43795 1830
rect 43740 1780 43745 1825
rect 43790 1780 43795 1825
rect 43740 1775 43795 1780
rect 43520 1725 43575 1730
rect 43520 1680 43525 1725
rect 43570 1680 43575 1725
rect 43520 1675 43575 1680
rect 43530 1500 43565 1675
rect 43750 1500 43785 1775
rect 44010 1500 44045 2020
rect 45240 1825 45295 1830
rect 45240 1780 45245 1825
rect 45290 1780 45295 1825
rect 45240 1775 45295 1780
rect 45020 1725 45075 1730
rect 45020 1680 45025 1725
rect 45070 1680 45075 1725
rect 45020 1675 45075 1680
rect 45030 1500 45065 1675
rect 45250 1500 45285 1775
rect 45510 1500 45545 2020
rect 46740 1825 46795 1830
rect 46740 1780 46745 1825
rect 46790 1780 46795 1825
rect 46740 1775 46795 1780
rect 46520 1725 46575 1730
rect 46520 1680 46525 1725
rect 46570 1680 46575 1725
rect 46520 1675 46575 1680
rect 46530 1500 46565 1675
rect 46750 1500 46785 1775
rect 47010 1500 47045 2020
rect 48240 1825 48295 1830
rect 48240 1780 48245 1825
rect 48290 1780 48295 1825
rect 48240 1775 48295 1780
rect 48020 1725 48075 1730
rect 48020 1680 48025 1725
rect 48070 1680 48075 1725
rect 48020 1675 48075 1680
rect 48030 1500 48065 1675
rect 48250 1500 48285 1775
rect 48510 1500 48545 2020
rect 49740 1825 49795 1830
rect 49740 1780 49745 1825
rect 49790 1780 49795 1825
rect 49740 1775 49795 1780
rect 49520 1725 49575 1730
rect 49520 1680 49525 1725
rect 49570 1680 49575 1725
rect 49520 1675 49575 1680
rect 49530 1500 49565 1675
rect 49750 1500 49785 1775
rect 50010 1500 50045 2020
rect 51240 1825 51295 1830
rect 51240 1780 51245 1825
rect 51290 1780 51295 1825
rect 51240 1775 51295 1780
rect 51020 1725 51075 1730
rect 51020 1680 51025 1725
rect 51070 1680 51075 1725
rect 51020 1675 51075 1680
rect 51030 1500 51065 1675
rect 51250 1500 51285 1775
rect 51510 1500 51545 2020
rect 52740 1825 52795 1830
rect 52740 1780 52745 1825
rect 52790 1780 52795 1825
rect 52740 1775 52795 1780
rect 52520 1725 52575 1730
rect 52520 1680 52525 1725
rect 52570 1680 52575 1725
rect 52520 1675 52575 1680
rect 52530 1500 52565 1675
rect 52750 1500 52785 1775
rect 53010 1500 53045 2020
rect 54240 1825 54295 1830
rect 54240 1780 54245 1825
rect 54290 1780 54295 1825
rect 54240 1775 54295 1780
rect 54020 1725 54075 1730
rect 54020 1680 54025 1725
rect 54070 1680 54075 1725
rect 54020 1675 54075 1680
rect 54030 1500 54065 1675
rect 54250 1500 54285 1775
rect 54510 1500 54545 2020
rect 55740 1825 55795 1830
rect 55740 1780 55745 1825
rect 55790 1780 55795 1825
rect 55740 1775 55795 1780
rect 55520 1725 55575 1730
rect 55520 1680 55525 1725
rect 55570 1680 55575 1725
rect 55520 1675 55575 1680
rect 55530 1500 55565 1675
rect 55750 1500 55785 1775
rect 56010 1500 56045 2020
rect 57240 1825 57295 1830
rect 57240 1780 57245 1825
rect 57290 1780 57295 1825
rect 57240 1775 57295 1780
rect 57020 1725 57075 1730
rect 57020 1680 57025 1725
rect 57070 1680 57075 1725
rect 57020 1675 57075 1680
rect 57030 1500 57065 1675
rect 57250 1500 57285 1775
rect 57510 1500 57545 2020
rect 58740 1825 58795 1830
rect 58740 1780 58745 1825
rect 58790 1780 58795 1825
rect 58740 1775 58795 1780
rect 58520 1725 58575 1730
rect 58520 1680 58525 1725
rect 58570 1680 58575 1725
rect 58520 1675 58575 1680
rect 58530 1500 58565 1675
rect 58750 1500 58785 1775
rect 59010 1500 59045 2020
rect 60240 1825 60295 1830
rect 60240 1780 60245 1825
rect 60290 1780 60295 1825
rect 60240 1775 60295 1780
rect 60020 1725 60075 1730
rect 60020 1680 60025 1725
rect 60070 1680 60075 1725
rect 60020 1675 60075 1680
rect 60030 1500 60065 1675
rect 60250 1500 60285 1775
rect 60510 1500 60545 2020
rect 61740 1825 61795 1830
rect 61740 1780 61745 1825
rect 61790 1780 61795 1825
rect 61740 1775 61795 1780
rect 61520 1725 61575 1730
rect 61520 1680 61525 1725
rect 61570 1680 61575 1725
rect 61520 1675 61575 1680
rect 61530 1500 61565 1675
rect 61750 1500 61785 1775
rect 62010 1500 62045 2020
rect 63240 1825 63295 1830
rect 63240 1780 63245 1825
rect 63290 1780 63295 1825
rect 63240 1775 63295 1780
rect 63020 1725 63075 1730
rect 63020 1680 63025 1725
rect 63070 1680 63075 1725
rect 63020 1675 63075 1680
rect 63030 1500 63065 1675
rect 63250 1500 63285 1775
rect 63510 1500 63545 2020
rect 64740 1825 64795 1830
rect 64740 1780 64745 1825
rect 64790 1780 64795 1825
rect 64740 1775 64795 1780
rect 64520 1725 64575 1730
rect 64520 1680 64525 1725
rect 64570 1680 64575 1725
rect 64520 1675 64575 1680
rect 64530 1500 64565 1675
rect 64750 1500 64785 1775
rect 65010 1500 65045 2020
rect 66240 1825 66295 1830
rect 66240 1780 66245 1825
rect 66290 1780 66295 1825
rect 66240 1775 66295 1780
rect 66020 1725 66075 1730
rect 66020 1680 66025 1725
rect 66070 1680 66075 1725
rect 66020 1675 66075 1680
rect 66030 1500 66065 1675
rect 66250 1500 66285 1775
rect 66510 1500 66545 2020
rect 67740 1825 67795 1830
rect 67740 1780 67745 1825
rect 67790 1780 67795 1825
rect 67740 1775 67795 1780
rect 67520 1725 67575 1730
rect 67520 1680 67525 1725
rect 67570 1680 67575 1725
rect 67520 1675 67575 1680
rect 67530 1500 67565 1675
rect 67750 1500 67785 1775
rect 68010 1500 68045 2020
rect 69240 1825 69295 1830
rect 69240 1780 69245 1825
rect 69290 1780 69295 1825
rect 69240 1775 69295 1780
rect 69020 1725 69075 1730
rect 69020 1680 69025 1725
rect 69070 1680 69075 1725
rect 69020 1675 69075 1680
rect 69030 1500 69065 1675
rect 69250 1500 69285 1775
rect 69510 1500 69545 2020
rect 70740 1825 70795 1830
rect 70740 1780 70745 1825
rect 70790 1780 70795 1825
rect 70740 1775 70795 1780
rect 70520 1725 70575 1730
rect 70520 1680 70525 1725
rect 70570 1680 70575 1725
rect 70520 1675 70575 1680
rect 70530 1500 70565 1675
rect 70750 1500 70785 1775
rect 71010 1500 71045 2020
rect 72240 1825 72295 1830
rect 72240 1780 72245 1825
rect 72290 1780 72295 1825
rect 72240 1775 72295 1780
rect 72020 1725 72075 1730
rect 72020 1680 72025 1725
rect 72070 1680 72075 1725
rect 72020 1675 72075 1680
rect 72030 1500 72065 1675
rect 72250 1500 72285 1775
rect 72510 1500 72545 2020
rect 73740 1825 73795 1830
rect 73740 1780 73745 1825
rect 73790 1780 73795 1825
rect 73740 1775 73795 1780
rect 73520 1725 73575 1730
rect 73520 1680 73525 1725
rect 73570 1680 73575 1725
rect 73520 1675 73575 1680
rect 73530 1500 73565 1675
rect 73750 1500 73785 1775
rect 74010 1500 74045 2020
rect 75240 1825 75295 1830
rect 75240 1780 75245 1825
rect 75290 1780 75295 1825
rect 75240 1775 75295 1780
rect 75020 1725 75075 1730
rect 75020 1680 75025 1725
rect 75070 1680 75075 1725
rect 75020 1675 75075 1680
rect 75030 1500 75065 1675
rect 75250 1500 75285 1775
rect 75510 1500 75545 2020
rect 76740 1825 76795 1830
rect 76740 1780 76745 1825
rect 76790 1780 76795 1825
rect 76740 1775 76795 1780
rect 76520 1725 76575 1730
rect 76520 1680 76525 1725
rect 76570 1680 76575 1725
rect 76520 1675 76575 1680
rect 76530 1500 76565 1675
rect 76750 1500 76785 1775
rect 77010 1500 77045 2020
rect 78240 1825 78295 1830
rect 78240 1780 78245 1825
rect 78290 1780 78295 1825
rect 78240 1775 78295 1780
rect 78020 1725 78075 1730
rect 78020 1680 78025 1725
rect 78070 1680 78075 1725
rect 78020 1675 78075 1680
rect 78030 1500 78065 1675
rect 78250 1500 78285 1775
rect 78510 1500 78545 2020
rect 79740 1825 79795 1830
rect 79740 1780 79745 1825
rect 79790 1780 79795 1825
rect 79740 1775 79795 1780
rect 79520 1725 79575 1730
rect 79520 1680 79525 1725
rect 79570 1680 79575 1725
rect 79520 1675 79575 1680
rect 79530 1500 79565 1675
rect 79750 1500 79785 1775
rect 80010 1500 80045 2020
rect 81240 1825 81295 1830
rect 81240 1780 81245 1825
rect 81290 1780 81295 1825
rect 81240 1775 81295 1780
rect 81020 1725 81075 1730
rect 81020 1680 81025 1725
rect 81070 1680 81075 1725
rect 81020 1675 81075 1680
rect 81030 1500 81065 1675
rect 81250 1500 81285 1775
rect 81510 1500 81545 2020
rect 82740 1825 82795 1830
rect 82740 1780 82745 1825
rect 82790 1780 82795 1825
rect 82740 1775 82795 1780
rect 82520 1725 82575 1730
rect 82520 1680 82525 1725
rect 82570 1680 82575 1725
rect 82520 1675 82575 1680
rect 82530 1500 82565 1675
rect 82750 1500 82785 1775
rect 83010 1500 83045 2020
rect 84240 1825 84295 1830
rect 84240 1780 84245 1825
rect 84290 1780 84295 1825
rect 84240 1775 84295 1780
rect 84020 1725 84075 1730
rect 84020 1680 84025 1725
rect 84070 1680 84075 1725
rect 84020 1675 84075 1680
rect 84030 1500 84065 1675
rect 84250 1500 84285 1775
rect 84510 1500 84545 2020
rect 85740 1825 85795 1830
rect 85740 1780 85745 1825
rect 85790 1780 85795 1825
rect 85740 1775 85795 1780
rect 85520 1725 85575 1730
rect 85520 1680 85525 1725
rect 85570 1680 85575 1725
rect 85520 1675 85575 1680
rect 85530 1500 85565 1675
rect 85750 1500 85785 1775
rect 86010 1500 86045 2020
rect 87240 1825 87295 1830
rect 87240 1780 87245 1825
rect 87290 1780 87295 1825
rect 87240 1775 87295 1780
rect 87020 1725 87075 1730
rect 87020 1680 87025 1725
rect 87070 1680 87075 1725
rect 87020 1675 87075 1680
rect 87030 1500 87065 1675
rect 87250 1500 87285 1775
rect 87510 1500 87545 2020
rect 88740 1825 88795 1830
rect 88740 1780 88745 1825
rect 88790 1780 88795 1825
rect 88740 1775 88795 1780
rect 88520 1725 88575 1730
rect 88520 1680 88525 1725
rect 88570 1680 88575 1725
rect 88520 1675 88575 1680
rect 88530 1500 88565 1675
rect 88750 1500 88785 1775
rect 89010 1500 89045 2020
rect 90240 1825 90295 1830
rect 90240 1780 90245 1825
rect 90290 1780 90295 1825
rect 90240 1775 90295 1780
rect 90020 1725 90075 1730
rect 90020 1680 90025 1725
rect 90070 1680 90075 1725
rect 90020 1675 90075 1680
rect 90030 1500 90065 1675
rect 90250 1500 90285 1775
rect 90510 1500 90545 2020
rect 91740 1825 91795 1830
rect 91740 1780 91745 1825
rect 91790 1780 91795 1825
rect 91740 1775 91795 1780
rect 91520 1725 91575 1730
rect 91520 1680 91525 1725
rect 91570 1680 91575 1725
rect 91520 1675 91575 1680
rect 91530 1500 91565 1675
rect 91750 1500 91785 1775
rect 92010 1500 92045 2020
rect 93240 1825 93295 1830
rect 93240 1780 93245 1825
rect 93290 1780 93295 1825
rect 93240 1775 93295 1780
rect 93020 1725 93075 1730
rect 93020 1680 93025 1725
rect 93070 1680 93075 1725
rect 93020 1675 93075 1680
rect 93030 1500 93065 1675
rect 93250 1500 93285 1775
rect 93510 1500 93545 2020
rect 94740 1825 94795 1830
rect 94740 1780 94745 1825
rect 94790 1780 94795 1825
rect 94740 1775 94795 1780
rect 94520 1725 94575 1730
rect 94520 1680 94525 1725
rect 94570 1680 94575 1725
rect 94520 1675 94575 1680
rect 94530 1500 94565 1675
rect 94750 1500 94785 1775
rect 95010 1500 95045 2020
rect 96240 1825 96295 1830
rect 96240 1780 96245 1825
rect 96290 1780 96295 1825
rect 96240 1775 96295 1780
rect 96020 1725 96075 1730
rect 96020 1680 96025 1725
rect 96070 1680 96075 1725
rect 96020 1675 96075 1680
rect 96030 1500 96065 1675
rect 96250 1500 96285 1775
rect 96510 1500 96545 2020
rect 97740 1825 97795 1830
rect 97740 1780 97745 1825
rect 97790 1780 97795 1825
rect 97740 1775 97795 1780
rect 97520 1725 97575 1730
rect 97520 1680 97525 1725
rect 97570 1680 97575 1725
rect 97520 1675 97575 1680
rect 97530 1500 97565 1675
rect 97750 1500 97785 1775
rect 98010 1500 98045 2020
rect 99240 1825 99295 1830
rect 99240 1780 99245 1825
rect 99290 1780 99295 1825
rect 99240 1775 99295 1780
rect 99020 1725 99075 1730
rect 99020 1680 99025 1725
rect 99070 1680 99075 1725
rect 99020 1675 99075 1680
rect 99030 1500 99065 1675
rect 99250 1500 99285 1775
rect 99510 1500 99545 2020
rect 100740 1825 100795 1830
rect 100740 1780 100745 1825
rect 100790 1780 100795 1825
rect 100740 1775 100795 1780
rect 100520 1725 100575 1730
rect 100520 1680 100525 1725
rect 100570 1680 100575 1725
rect 100520 1675 100575 1680
rect 100530 1500 100565 1675
rect 100750 1500 100785 1775
rect 101010 1500 101045 2020
rect 102240 1825 102295 1830
rect 102240 1780 102245 1825
rect 102290 1780 102295 1825
rect 102240 1775 102295 1780
rect 102020 1725 102075 1730
rect 102020 1680 102025 1725
rect 102070 1680 102075 1725
rect 102020 1675 102075 1680
rect 102030 1500 102065 1675
rect 102250 1500 102285 1775
rect 102510 1500 102545 2020
rect 103740 1825 103795 1830
rect 103740 1780 103745 1825
rect 103790 1780 103795 1825
rect 103740 1775 103795 1780
rect 103520 1725 103575 1730
rect 103520 1680 103525 1725
rect 103570 1680 103575 1725
rect 103520 1675 103575 1680
rect 103530 1500 103565 1675
rect 103750 1500 103785 1775
rect 104010 1500 104045 2020
rect 105240 1825 105295 1830
rect 105240 1780 105245 1825
rect 105290 1780 105295 1825
rect 105240 1775 105295 1780
rect 105020 1725 105075 1730
rect 105020 1680 105025 1725
rect 105070 1680 105075 1725
rect 105020 1675 105075 1680
rect 105030 1500 105065 1675
rect 105250 1500 105285 1775
rect 105510 1500 105545 2020
rect 106740 1825 106795 1830
rect 106740 1780 106745 1825
rect 106790 1780 106795 1825
rect 106740 1775 106795 1780
rect 106520 1725 106575 1730
rect 106520 1680 106525 1725
rect 106570 1680 106575 1725
rect 106520 1675 106575 1680
rect 106530 1500 106565 1675
rect 106750 1500 106785 1775
rect 107010 1500 107045 2020
rect 108240 1825 108295 1830
rect 108240 1780 108245 1825
rect 108290 1780 108295 1825
rect 108240 1775 108295 1780
rect 108020 1725 108075 1730
rect 108020 1680 108025 1725
rect 108070 1680 108075 1725
rect 108020 1675 108075 1680
rect 108030 1500 108065 1675
rect 108250 1500 108285 1775
rect 108510 1500 108545 2020
rect 109740 1825 109795 1830
rect 109740 1780 109745 1825
rect 109790 1780 109795 1825
rect 109740 1775 109795 1780
rect 109520 1725 109575 1730
rect 109520 1680 109525 1725
rect 109570 1680 109575 1725
rect 109520 1675 109575 1680
rect 109530 1500 109565 1675
rect 109750 1500 109785 1775
rect 110010 1500 110045 2020
rect 111240 1825 111295 1830
rect 111240 1780 111245 1825
rect 111290 1780 111295 1825
rect 111240 1775 111295 1780
rect 111020 1725 111075 1730
rect 111020 1680 111025 1725
rect 111070 1680 111075 1725
rect 111020 1675 111075 1680
rect 111030 1500 111065 1675
rect 111250 1500 111285 1775
rect 111510 1500 111545 2020
rect 112740 1825 112795 1830
rect 112740 1780 112745 1825
rect 112790 1780 112795 1825
rect 112740 1775 112795 1780
rect 112520 1725 112575 1730
rect 112520 1680 112525 1725
rect 112570 1680 112575 1725
rect 112520 1675 112575 1680
rect 112530 1500 112565 1675
rect 112750 1500 112785 1775
rect 113010 1500 113045 2020
rect 114240 1825 114295 1830
rect 114240 1780 114245 1825
rect 114290 1780 114295 1825
rect 114240 1775 114295 1780
rect 114020 1725 114075 1730
rect 114020 1680 114025 1725
rect 114070 1680 114075 1725
rect 114020 1675 114075 1680
rect 114030 1500 114065 1675
rect 114250 1500 114285 1775
rect 114510 1500 114545 2020
rect 115740 1825 115795 1830
rect 115740 1780 115745 1825
rect 115790 1780 115795 1825
rect 115740 1775 115795 1780
rect 115520 1725 115575 1730
rect 115520 1680 115525 1725
rect 115570 1680 115575 1725
rect 115520 1675 115575 1680
rect 115530 1500 115565 1675
rect 115750 1500 115785 1775
rect 116010 1500 116045 2020
rect 117240 1825 117295 1830
rect 117240 1780 117245 1825
rect 117290 1780 117295 1825
rect 117240 1775 117295 1780
rect 117020 1725 117075 1730
rect 117020 1680 117025 1725
rect 117070 1680 117075 1725
rect 117020 1675 117075 1680
rect 117030 1500 117065 1675
rect 117250 1500 117285 1775
rect 117510 1500 117545 2020
rect 118740 1825 118795 1830
rect 118740 1780 118745 1825
rect 118790 1780 118795 1825
rect 118740 1775 118795 1780
rect 118520 1725 118575 1730
rect 118520 1680 118525 1725
rect 118570 1680 118575 1725
rect 118520 1675 118575 1680
rect 118530 1500 118565 1675
rect 118750 1500 118785 1775
rect 119010 1500 119045 2020
rect -280 780 -130 785
rect -280 745 -270 780
rect -280 740 -130 745
rect -375 80 -370 115
rect -325 80 -320 115
rect -1500 -720 -500 -715
rect -1500 -755 -790 -720
rect -590 -755 -500 -720
rect -1500 -760 -500 -755
rect -375 -1385 -320 80
rect -280 -720 -130 -715
rect -280 -755 -270 -720
rect -280 -760 -130 -755
rect -375 -1420 -370 -1385
rect -325 -1420 -320 -1385
rect -1500 -2220 -500 -2215
rect -1500 -2255 -790 -2220
rect -590 -2255 -500 -2220
rect -1500 -2260 -500 -2255
rect -375 -2885 -320 -1420
rect -280 -2220 -130 -2215
rect -280 -2255 -270 -2220
rect -280 -2260 -130 -2255
rect -375 -2920 -370 -2885
rect -325 -2920 -320 -2885
rect -1500 -3720 -500 -3715
rect -1500 -3755 -790 -3720
rect -590 -3755 -500 -3720
rect -1500 -3760 -500 -3755
rect -375 -4385 -320 -2920
rect -280 -3720 -130 -3715
rect -280 -3755 -270 -3720
rect -280 -3760 -130 -3755
rect -375 -4420 -370 -4385
rect -325 -4420 -320 -4385
rect -1500 -5220 -500 -5215
rect -1500 -5255 -790 -5220
rect -590 -5255 -500 -5220
rect -1500 -5260 -500 -5255
rect -375 -5885 -320 -4420
rect -280 -5220 -130 -5215
rect -280 -5255 -270 -5220
rect -280 -5260 -130 -5255
rect -375 -5920 -370 -5885
rect -325 -5920 -320 -5885
rect -1500 -6720 -500 -6715
rect -1500 -6755 -790 -6720
rect -590 -6755 -500 -6720
rect -1500 -6760 -500 -6755
rect -375 -7385 -320 -5920
rect -280 -6720 -130 -6715
rect -280 -6755 -270 -6720
rect -280 -6760 -130 -6755
rect -375 -7420 -370 -7385
rect -325 -7420 -320 -7385
rect -1500 -8220 -500 -8215
rect -1500 -8255 -790 -8220
rect -590 -8255 -500 -8220
rect -1500 -8260 -500 -8255
rect -375 -8885 -320 -7420
rect -280 -8220 -130 -8215
rect -280 -8255 -270 -8220
rect -280 -8260 -130 -8255
rect -375 -8920 -370 -8885
rect -325 -8920 -320 -8885
rect -1500 -9720 -500 -9715
rect -1500 -9755 -790 -9720
rect -590 -9755 -500 -9720
rect -1500 -9760 -500 -9755
rect -375 -10385 -320 -8920
rect -280 -9720 -130 -9715
rect -280 -9755 -270 -9720
rect -280 -9760 -130 -9755
rect -375 -10420 -370 -10385
rect -325 -10420 -320 -10385
rect -1500 -11220 -500 -11215
rect -1500 -11255 -790 -11220
rect -590 -11255 -500 -11220
rect -1500 -11260 -500 -11255
rect -375 -11885 -320 -10420
rect -280 -11220 -130 -11215
rect -280 -11255 -270 -11220
rect -280 -11260 -130 -11255
rect -375 -11920 -370 -11885
rect -325 -11920 -320 -11885
rect -1500 -12720 -500 -12715
rect -1500 -12755 -790 -12720
rect -590 -12755 -500 -12720
rect -1500 -12760 -500 -12755
rect -375 -13385 -320 -11920
rect -280 -12720 -130 -12715
rect -280 -12755 -270 -12720
rect -280 -12760 -130 -12755
rect -375 -13420 -370 -13385
rect -325 -13420 -320 -13385
rect -1500 -14220 -500 -14215
rect -1500 -14255 -790 -14220
rect -590 -14255 -500 -14220
rect -1500 -14260 -500 -14255
rect -375 -14885 -320 -13420
rect -280 -14220 -130 -14215
rect -280 -14255 -270 -14220
rect -280 -14260 -130 -14255
rect -375 -14920 -370 -14885
rect -325 -14920 -320 -14885
rect -1500 -15720 -500 -15715
rect -1500 -15755 -790 -15720
rect -590 -15755 -500 -15720
rect -1500 -15760 -500 -15755
rect -375 -16385 -320 -14920
rect -280 -15720 -130 -15715
rect -280 -15755 -270 -15720
rect -280 -15760 -130 -15755
rect -375 -16420 -370 -16385
rect -325 -16420 -320 -16385
rect -1500 -17220 -500 -17215
rect -1500 -17255 -790 -17220
rect -590 -17255 -500 -17220
rect -1500 -17260 -500 -17255
rect -375 -17885 -320 -16420
rect -280 -17220 -130 -17215
rect -280 -17255 -270 -17220
rect -280 -17260 -130 -17255
rect -375 -17920 -370 -17885
rect -325 -17920 -320 -17885
rect -1500 -18720 -500 -18715
rect -1500 -18755 -790 -18720
rect -590 -18755 -500 -18720
rect -1500 -18760 -500 -18755
rect -375 -19385 -320 -17920
rect -280 -18720 -130 -18715
rect -280 -18755 -270 -18720
rect -280 -18760 -130 -18755
rect -375 -19420 -370 -19385
rect -325 -19420 -320 -19385
rect -1500 -20220 -500 -20215
rect -1500 -20255 -790 -20220
rect -590 -20255 -500 -20220
rect -1500 -20260 -500 -20255
rect -375 -20885 -320 -19420
rect -280 -20220 -130 -20215
rect -280 -20255 -270 -20220
rect -280 -20260 -130 -20255
rect -375 -20920 -370 -20885
rect -325 -20920 -320 -20885
rect -1500 -21720 -500 -21715
rect -1500 -21755 -790 -21720
rect -590 -21755 -500 -21720
rect -1500 -21760 -500 -21755
rect -375 -22385 -320 -20920
rect -280 -21720 -130 -21715
rect -280 -21755 -270 -21720
rect -280 -21760 -130 -21755
rect -375 -22420 -370 -22385
rect -325 -22420 -320 -22385
rect -1500 -23220 -500 -23215
rect -1500 -23255 -790 -23220
rect -590 -23255 -500 -23220
rect -1500 -23260 -500 -23255
rect -375 -23885 -320 -22420
rect -280 -23220 -130 -23215
rect -280 -23255 -270 -23220
rect -280 -23260 -130 -23255
rect -375 -23920 -370 -23885
rect -325 -23920 -320 -23885
rect -1500 -24720 -500 -24715
rect -1500 -24755 -790 -24720
rect -590 -24755 -500 -24720
rect -1500 -24760 -500 -24755
rect -375 -25385 -320 -23920
rect -280 -24720 -130 -24715
rect -280 -24755 -270 -24720
rect -280 -24760 -130 -24755
rect -375 -25420 -370 -25385
rect -325 -25420 -320 -25385
rect -1500 -26220 -500 -26215
rect -1500 -26255 -790 -26220
rect -590 -26255 -500 -26220
rect -1500 -26260 -500 -26255
rect -375 -26885 -320 -25420
rect -280 -26220 -130 -26215
rect -280 -26255 -270 -26220
rect -280 -26260 -130 -26255
rect -375 -26920 -370 -26885
rect -325 -26920 -320 -26885
rect -1500 -27720 -500 -27715
rect -1500 -27755 -790 -27720
rect -590 -27755 -500 -27720
rect -1500 -27760 -500 -27755
rect -375 -28385 -320 -26920
rect -280 -27720 -130 -27715
rect -280 -27755 -270 -27720
rect -280 -27760 -130 -27755
rect -375 -28420 -370 -28385
rect -325 -28420 -320 -28385
rect -1500 -29220 -500 -29215
rect -1500 -29255 -790 -29220
rect -590 -29255 -500 -29220
rect -1500 -29260 -500 -29255
rect -375 -29885 -320 -28420
rect -280 -29220 -130 -29215
rect -280 -29255 -270 -29220
rect -280 -29260 -130 -29255
rect -375 -29920 -370 -29885
rect -325 -29920 -320 -29885
rect -1500 -30720 -500 -30715
rect -1500 -30755 -790 -30720
rect -590 -30755 -500 -30720
rect -1500 -30760 -500 -30755
rect -375 -31385 -320 -29920
rect -280 -30720 -130 -30715
rect -280 -30755 -270 -30720
rect -280 -30760 -130 -30755
rect -375 -31420 -370 -31385
rect -325 -31420 -320 -31385
rect -1500 -32220 -500 -32215
rect -1500 -32255 -790 -32220
rect -590 -32255 -500 -32220
rect -1500 -32260 -500 -32255
rect -375 -32885 -320 -31420
rect -280 -32220 -130 -32215
rect -280 -32255 -270 -32220
rect -280 -32260 -130 -32255
rect -375 -32920 -370 -32885
rect -325 -32920 -320 -32885
rect -1500 -33720 -500 -33715
rect -1500 -33755 -790 -33720
rect -590 -33755 -500 -33720
rect -1500 -33760 -500 -33755
rect -375 -34385 -320 -32920
rect -280 -33720 -130 -33715
rect -280 -33755 -270 -33720
rect -280 -33760 -130 -33755
rect -375 -34420 -370 -34385
rect -325 -34420 -320 -34385
rect -1500 -35220 -500 -35215
rect -1500 -35255 -790 -35220
rect -590 -35255 -500 -35220
rect -1500 -35260 -500 -35255
rect -375 -35885 -320 -34420
rect -280 -35220 -130 -35215
rect -280 -35255 -270 -35220
rect -280 -35260 -130 -35255
rect -375 -35920 -370 -35885
rect -325 -35920 -320 -35885
rect -1500 -36720 -500 -36715
rect -1500 -36755 -790 -36720
rect -590 -36755 -500 -36720
rect -1500 -36760 -500 -36755
rect -375 -37385 -320 -35920
rect -280 -36720 -130 -36715
rect -280 -36755 -270 -36720
rect -280 -36760 -130 -36755
rect -375 -37420 -370 -37385
rect -325 -37420 -320 -37385
rect -1500 -38220 -500 -38215
rect -1500 -38255 -790 -38220
rect -590 -38255 -500 -38220
rect -1500 -38260 -500 -38255
rect -375 -38885 -320 -37420
rect -280 -38220 -130 -38215
rect -280 -38255 -270 -38220
rect -280 -38260 -130 -38255
rect -375 -38920 -370 -38885
rect -325 -38920 -320 -38885
rect -1500 -39720 -500 -39715
rect -1500 -39755 -790 -39720
rect -590 -39755 -500 -39720
rect -1500 -39760 -500 -39755
rect -375 -40385 -320 -38920
rect -280 -39720 -130 -39715
rect -280 -39755 -270 -39720
rect -280 -39760 -130 -39755
rect -375 -40420 -370 -40385
rect -325 -40420 -320 -40385
rect -1500 -41220 -500 -41215
rect -1500 -41255 -790 -41220
rect -590 -41255 -500 -41220
rect -1500 -41260 -500 -41255
rect -375 -41885 -320 -40420
rect -280 -41220 -130 -41215
rect -280 -41255 -270 -41220
rect -280 -41260 -130 -41255
rect -375 -41920 -370 -41885
rect -325 -41920 -320 -41885
rect -1500 -42720 -500 -42715
rect -1500 -42755 -790 -42720
rect -590 -42755 -500 -42720
rect -1500 -42760 -500 -42755
rect -375 -43385 -320 -41920
rect -280 -42720 -130 -42715
rect -280 -42755 -270 -42720
rect -280 -42760 -130 -42755
rect -375 -43420 -370 -43385
rect -325 -43420 -320 -43385
rect -1500 -44220 -500 -44215
rect -1500 -44255 -790 -44220
rect -590 -44255 -500 -44220
rect -1500 -44260 -500 -44255
rect -375 -44885 -320 -43420
rect -280 -44220 -130 -44215
rect -280 -44255 -270 -44220
rect -280 -44260 -130 -44255
rect -375 -44920 -370 -44885
rect -325 -44920 -320 -44885
rect -1500 -45720 -500 -45715
rect -1500 -45755 -790 -45720
rect -590 -45755 -500 -45720
rect -1500 -45760 -500 -45755
rect -375 -46385 -320 -44920
rect -280 -45720 -130 -45715
rect -280 -45755 -270 -45720
rect -280 -45760 -130 -45755
rect -375 -46420 -370 -46385
rect -325 -46420 -320 -46385
rect -1500 -47220 -500 -47215
rect -1500 -47255 -790 -47220
rect -590 -47255 -500 -47220
rect -1500 -47260 -500 -47255
rect -375 -47885 -320 -46420
rect -280 -47220 -130 -47215
rect -280 -47255 -270 -47220
rect -280 -47260 -130 -47255
rect -375 -47920 -370 -47885
rect -325 -47920 -320 -47885
rect -1500 -48720 -500 -48715
rect -1500 -48755 -790 -48720
rect -590 -48755 -500 -48720
rect -1500 -48760 -500 -48755
rect -375 -49385 -320 -47920
rect -280 -48720 -130 -48715
rect -280 -48755 -270 -48720
rect -280 -48760 -130 -48755
rect -375 -49420 -370 -49385
rect -325 -49420 -320 -49385
rect -1500 -50220 -500 -50215
rect -1500 -50255 -790 -50220
rect -590 -50255 -500 -50220
rect -1500 -50260 -500 -50255
rect -375 -50885 -320 -49420
rect -280 -50220 -130 -50215
rect -280 -50255 -270 -50220
rect -280 -50260 -130 -50255
rect -375 -50920 -370 -50885
rect -325 -50920 -320 -50885
rect -1500 -51720 -500 -51715
rect -1500 -51755 -790 -51720
rect -590 -51755 -500 -51720
rect -1500 -51760 -500 -51755
rect -375 -52385 -320 -50920
rect -280 -51720 -130 -51715
rect -280 -51755 -270 -51720
rect -280 -51760 -130 -51755
rect -375 -52420 -370 -52385
rect -325 -52420 -320 -52385
rect -1500 -53220 -500 -53215
rect -1500 -53255 -790 -53220
rect -590 -53255 -500 -53220
rect -1500 -53260 -500 -53255
rect -375 -53885 -320 -52420
rect -280 -53220 -130 -53215
rect -280 -53255 -270 -53220
rect -280 -53260 -130 -53255
rect -375 -53920 -370 -53885
rect -325 -53920 -320 -53885
rect -1500 -54720 -500 -54715
rect -1500 -54755 -790 -54720
rect -590 -54755 -500 -54720
rect -1500 -54760 -500 -54755
rect -375 -55385 -320 -53920
rect -280 -54720 -130 -54715
rect -280 -54755 -270 -54720
rect -280 -54760 -130 -54755
rect -375 -55420 -370 -55385
rect -325 -55420 -320 -55385
rect -1500 -56220 -500 -56215
rect -1500 -56255 -790 -56220
rect -590 -56255 -500 -56220
rect -1500 -56260 -500 -56255
rect -375 -56885 -320 -55420
rect -280 -56220 -130 -56215
rect -280 -56255 -270 -56220
rect -280 -56260 -130 -56255
rect -375 -56920 -370 -56885
rect -325 -56920 -320 -56885
rect -1500 -57720 -500 -57715
rect -1500 -57755 -790 -57720
rect -590 -57755 -500 -57720
rect -1500 -57760 -500 -57755
rect -375 -58385 -320 -56920
rect -280 -57720 -130 -57715
rect -280 -57755 -270 -57720
rect -280 -57760 -130 -57755
rect -375 -58420 -370 -58385
rect -325 -58420 -320 -58385
rect -1500 -59220 -500 -59215
rect -1500 -59255 -790 -59220
rect -590 -59255 -500 -59220
rect -1500 -59260 -500 -59255
rect -375 -59885 -320 -58420
rect -280 -59220 -130 -59215
rect -280 -59255 -270 -59220
rect -280 -59260 -130 -59255
rect -375 -59920 -370 -59885
rect -325 -59920 -320 -59885
rect -1500 -60720 -500 -60715
rect -1500 -60755 -790 -60720
rect -590 -60755 -500 -60720
rect -1500 -60760 -500 -60755
rect -375 -61385 -320 -59920
rect -280 -60720 -130 -60715
rect -280 -60755 -270 -60720
rect -280 -60760 -130 -60755
rect -375 -61420 -370 -61385
rect -325 -61420 -320 -61385
rect -1500 -62220 -500 -62215
rect -1500 -62255 -790 -62220
rect -590 -62255 -500 -62220
rect -1500 -62260 -500 -62255
rect -375 -62885 -320 -61420
rect -280 -62220 -130 -62215
rect -280 -62255 -270 -62220
rect -280 -62260 -130 -62255
rect -375 -62920 -370 -62885
rect -325 -62920 -320 -62885
rect -1500 -63720 -500 -63715
rect -1500 -63755 -790 -63720
rect -590 -63755 -500 -63720
rect -1500 -63760 -500 -63755
rect -375 -64385 -320 -62920
rect -280 -63720 -130 -63715
rect -280 -63755 -270 -63720
rect -280 -63760 -130 -63755
rect -375 -64420 -370 -64385
rect -325 -64420 -320 -64385
rect -1500 -65220 -500 -65215
rect -1500 -65255 -790 -65220
rect -590 -65255 -500 -65220
rect -1500 -65260 -500 -65255
rect -375 -65885 -320 -64420
rect -280 -65220 -130 -65215
rect -280 -65255 -270 -65220
rect -280 -65260 -130 -65255
rect -375 -65920 -370 -65885
rect -325 -65920 -320 -65885
rect -1500 -66720 -500 -66715
rect -1500 -66755 -790 -66720
rect -590 -66755 -500 -66720
rect -1500 -66760 -500 -66755
rect -375 -67385 -320 -65920
rect -280 -66720 -130 -66715
rect -280 -66755 -270 -66720
rect -280 -66760 -130 -66755
rect -375 -67420 -370 -67385
rect -325 -67420 -320 -67385
rect -1500 -68220 -500 -68215
rect -1500 -68255 -790 -68220
rect -590 -68255 -500 -68220
rect -1500 -68260 -500 -68255
rect -375 -68885 -320 -67420
rect -280 -68220 -130 -68215
rect -280 -68255 -270 -68220
rect -280 -68260 -130 -68255
rect -375 -68920 -370 -68885
rect -325 -68920 -320 -68885
rect -1500 -69720 -500 -69715
rect -1500 -69755 -790 -69720
rect -590 -69755 -500 -69720
rect -1500 -69760 -500 -69755
rect -375 -70385 -320 -68920
rect -280 -69720 -130 -69715
rect -280 -69755 -270 -69720
rect -280 -69760 -130 -69755
rect -375 -70420 -370 -70385
rect -325 -70420 -320 -70385
rect -1500 -71220 -500 -71215
rect -1500 -71255 -790 -71220
rect -590 -71255 -500 -71220
rect -1500 -71260 -500 -71255
rect -375 -71885 -320 -70420
rect -280 -71220 -130 -71215
rect -280 -71255 -270 -71220
rect -280 -71260 -130 -71255
rect -375 -71920 -370 -71885
rect -325 -71920 -320 -71885
rect -1500 -72720 -500 -72715
rect -1500 -72755 -790 -72720
rect -590 -72755 -500 -72720
rect -1500 -72760 -500 -72755
rect -375 -73385 -320 -71920
rect -280 -72720 -130 -72715
rect -280 -72755 -270 -72720
rect -280 -72760 -130 -72755
rect -375 -73420 -370 -73385
rect -325 -73420 -320 -73385
rect -1500 -74220 -500 -74215
rect -1500 -74255 -790 -74220
rect -590 -74255 -500 -74220
rect -1500 -74260 -500 -74255
rect -375 -74885 -320 -73420
rect -280 -74220 -130 -74215
rect -280 -74255 -270 -74220
rect -280 -74260 -130 -74255
rect -375 -74920 -370 -74885
rect -325 -74920 -320 -74885
rect -1500 -75720 -500 -75715
rect -1500 -75755 -790 -75720
rect -590 -75755 -500 -75720
rect -1500 -75760 -500 -75755
rect -375 -76385 -320 -74920
rect -280 -75720 -130 -75715
rect -280 -75755 -270 -75720
rect -280 -75760 -130 -75755
rect -375 -76420 -370 -76385
rect -325 -76420 -320 -76385
rect -1500 -77220 -500 -77215
rect -1500 -77255 -790 -77220
rect -590 -77255 -500 -77220
rect -1500 -77260 -500 -77255
rect -375 -77885 -320 -76420
rect -280 -77220 -130 -77215
rect -280 -77255 -270 -77220
rect -280 -77260 -130 -77255
rect -375 -77920 -370 -77885
rect -325 -77920 -320 -77885
rect -1500 -78720 -500 -78715
rect -1500 -78755 -790 -78720
rect -590 -78755 -500 -78720
rect -1500 -78760 -500 -78755
rect -375 -79385 -320 -77920
rect -280 -78720 -130 -78715
rect -280 -78755 -270 -78720
rect -280 -78760 -130 -78755
rect -375 -79420 -370 -79385
rect -325 -79420 -320 -79385
rect -1500 -80220 -500 -80215
rect -1500 -80255 -790 -80220
rect -590 -80255 -500 -80220
rect -1500 -80260 -500 -80255
rect -375 -80885 -320 -79420
rect -280 -80220 -130 -80215
rect -280 -80255 -270 -80220
rect -280 -80260 -130 -80255
rect -375 -80920 -370 -80885
rect -325 -80920 -320 -80885
rect -1500 -81720 -500 -81715
rect -1500 -81755 -790 -81720
rect -590 -81755 -500 -81720
rect -1500 -81760 -500 -81755
rect -375 -82385 -320 -80920
rect -280 -81720 -130 -81715
rect -280 -81755 -270 -81720
rect -280 -81760 -130 -81755
rect -375 -82420 -370 -82385
rect -325 -82420 -320 -82385
rect -1500 -83220 -500 -83215
rect -1500 -83255 -790 -83220
rect -590 -83255 -500 -83220
rect -1500 -83260 -500 -83255
rect -375 -83885 -320 -82420
rect -280 -83220 -130 -83215
rect -280 -83255 -270 -83220
rect -280 -83260 -130 -83255
rect -375 -83920 -370 -83885
rect -325 -83920 -320 -83885
rect -1500 -84720 -500 -84715
rect -1500 -84755 -790 -84720
rect -590 -84755 -500 -84720
rect -1500 -84760 -500 -84755
rect -375 -85385 -320 -83920
rect -280 -84720 -130 -84715
rect -280 -84755 -270 -84720
rect -280 -84760 -130 -84755
rect -375 -85420 -370 -85385
rect -325 -85420 -320 -85385
rect -1500 -86220 -500 -86215
rect -1500 -86255 -790 -86220
rect -590 -86255 -500 -86220
rect -1500 -86260 -500 -86255
rect -375 -86885 -320 -85420
rect -280 -86220 -130 -86215
rect -280 -86255 -270 -86220
rect -280 -86260 -130 -86255
rect -375 -86920 -370 -86885
rect -325 -86920 -320 -86885
rect -1500 -87720 -500 -87715
rect -1500 -87755 -790 -87720
rect -590 -87755 -500 -87720
rect -1500 -87760 -500 -87755
rect -375 -88385 -320 -86920
rect -280 -87720 -130 -87715
rect -280 -87755 -270 -87720
rect -280 -87760 -130 -87755
rect -375 -88420 -370 -88385
rect -325 -88420 -320 -88385
rect -1500 -89220 -500 -89215
rect -1500 -89255 -790 -89220
rect -590 -89255 -500 -89220
rect -1500 -89260 -500 -89255
rect -375 -89885 -320 -88420
rect -280 -89220 -130 -89215
rect -280 -89255 -270 -89220
rect -280 -89260 -130 -89255
rect -375 -89920 -370 -89885
rect -325 -89920 -320 -89885
rect -1500 -90720 -500 -90715
rect -1500 -90755 -790 -90720
rect -590 -90755 -500 -90720
rect -1500 -90760 -500 -90755
rect -375 -91385 -320 -89920
rect -280 -90720 -130 -90715
rect -280 -90755 -270 -90720
rect -280 -90760 -130 -90755
rect -375 -91420 -370 -91385
rect -325 -91420 -320 -91385
rect -1500 -92220 -500 -92215
rect -1500 -92255 -790 -92220
rect -590 -92255 -500 -92220
rect -1500 -92260 -500 -92255
rect -375 -92885 -320 -91420
rect -280 -92220 -130 -92215
rect -280 -92255 -270 -92220
rect -280 -92260 -130 -92255
rect -375 -92920 -370 -92885
rect -325 -92920 -320 -92885
rect -1500 -93720 -500 -93715
rect -1500 -93755 -790 -93720
rect -590 -93755 -500 -93720
rect -1500 -93760 -500 -93755
rect -375 -94385 -320 -92920
rect -280 -93720 -130 -93715
rect -280 -93755 -270 -93720
rect -280 -93760 -130 -93755
rect -375 -94420 -370 -94385
rect -325 -94420 -320 -94385
rect -1500 -95220 -500 -95215
rect -1500 -95255 -790 -95220
rect -590 -95255 -500 -95220
rect -1500 -95260 -500 -95255
rect -375 -95885 -320 -94420
rect -280 -95220 -130 -95215
rect -280 -95255 -270 -95220
rect -280 -95260 -130 -95255
rect -375 -95920 -370 -95885
rect -325 -95920 -320 -95885
rect -1500 -96720 -500 -96715
rect -1500 -96755 -790 -96720
rect -590 -96755 -500 -96720
rect -1500 -96760 -500 -96755
rect -375 -97385 -320 -95920
rect -280 -96720 -130 -96715
rect -280 -96755 -270 -96720
rect -280 -96760 -130 -96755
rect -375 -97420 -370 -97385
rect -325 -97420 -320 -97385
rect -1500 -98220 -500 -98215
rect -1500 -98255 -790 -98220
rect -590 -98255 -500 -98220
rect -1500 -98260 -500 -98255
rect -375 -98885 -320 -97420
rect -280 -98220 -130 -98215
rect -280 -98255 -270 -98220
rect -280 -98260 -130 -98255
rect -375 -98920 -370 -98885
rect -325 -98920 -320 -98885
rect -1500 -99720 -500 -99715
rect -1500 -99755 -790 -99720
rect -590 -99755 -500 -99720
rect -1500 -99760 -500 -99755
rect -375 -100385 -320 -98920
rect -280 -99720 -130 -99715
rect -280 -99755 -270 -99720
rect -280 -99760 -130 -99755
rect -375 -100420 -370 -100385
rect -325 -100420 -320 -100385
rect -1500 -101220 -500 -101215
rect -1500 -101255 -790 -101220
rect -590 -101255 -500 -101220
rect -1500 -101260 -500 -101255
rect -375 -101885 -320 -100420
rect -280 -101220 -130 -101215
rect -280 -101255 -270 -101220
rect -280 -101260 -130 -101255
rect -375 -101920 -370 -101885
rect -325 -101920 -320 -101885
rect -1500 -102720 -500 -102715
rect -1500 -102755 -790 -102720
rect -590 -102755 -500 -102720
rect -1500 -102760 -500 -102755
rect -375 -103385 -320 -101920
rect -280 -102720 -130 -102715
rect -280 -102755 -270 -102720
rect -280 -102760 -130 -102755
rect -375 -103420 -370 -103385
rect -325 -103420 -320 -103385
rect -1500 -104220 -500 -104215
rect -1500 -104255 -790 -104220
rect -590 -104255 -500 -104220
rect -1500 -104260 -500 -104255
rect -375 -104885 -320 -103420
rect -280 -104220 -130 -104215
rect -280 -104255 -270 -104220
rect -280 -104260 -130 -104255
rect -375 -104920 -370 -104885
rect -325 -104920 -320 -104885
rect -1500 -105720 -500 -105715
rect -1500 -105755 -790 -105720
rect -590 -105755 -500 -105720
rect -1500 -105760 -500 -105755
rect -375 -106385 -320 -104920
rect -280 -105720 -130 -105715
rect -280 -105755 -270 -105720
rect -280 -105760 -130 -105755
rect -375 -106420 -370 -106385
rect -325 -106420 -320 -106385
rect -1500 -107220 -500 -107215
rect -1500 -107255 -790 -107220
rect -590 -107255 -500 -107220
rect -1500 -107260 -500 -107255
rect -375 -107885 -320 -106420
rect -280 -107220 -130 -107215
rect -280 -107255 -270 -107220
rect -280 -107260 -130 -107255
rect -375 -107920 -370 -107885
rect -325 -107920 -320 -107885
rect -1500 -108720 -500 -108715
rect -1500 -108755 -790 -108720
rect -590 -108755 -500 -108720
rect -1500 -108760 -500 -108755
rect -375 -109385 -320 -107920
rect -280 -108720 -130 -108715
rect -280 -108755 -270 -108720
rect -280 -108760 -130 -108755
rect -375 -109420 -370 -109385
rect -325 -109420 -320 -109385
rect -1500 -110220 -500 -110215
rect -1500 -110255 -790 -110220
rect -590 -110255 -500 -110220
rect -1500 -110260 -500 -110255
rect -375 -110885 -320 -109420
rect -280 -110220 -130 -110215
rect -280 -110255 -270 -110220
rect -280 -110260 -130 -110255
rect -375 -110920 -370 -110885
rect -325 -110920 -320 -110885
rect -1500 -111720 -500 -111715
rect -1500 -111755 -790 -111720
rect -590 -111755 -500 -111720
rect -1500 -111760 -500 -111755
rect -375 -112385 -320 -110920
rect -280 -111720 -130 -111715
rect -280 -111755 -270 -111720
rect -280 -111760 -130 -111755
rect -375 -112420 -370 -112385
rect -325 -112420 -320 -112385
rect -1500 -113220 -500 -113215
rect -1500 -113255 -790 -113220
rect -590 -113255 -500 -113220
rect -1500 -113260 -500 -113255
rect -375 -113885 -320 -112420
rect -280 -113220 -130 -113215
rect -280 -113255 -270 -113220
rect -280 -113260 -130 -113255
rect -375 -113920 -370 -113885
rect -325 -113920 -320 -113885
rect -1500 -114720 -500 -114715
rect -1500 -114755 -790 -114720
rect -590 -114755 -500 -114720
rect -1500 -114760 -500 -114755
rect -375 -115385 -320 -113920
rect -280 -114720 -130 -114715
rect -280 -114755 -270 -114720
rect -280 -114760 -130 -114755
rect -375 -115420 -370 -115385
rect -325 -115420 -320 -115385
rect -1500 -116220 -500 -116215
rect -1500 -116255 -790 -116220
rect -590 -116255 -500 -116220
rect -1500 -116260 -500 -116255
rect -375 -116885 -320 -115420
rect -280 -116220 -130 -116215
rect -280 -116255 -270 -116220
rect -280 -116260 -130 -116255
rect -375 -116920 -370 -116885
rect -325 -116920 -320 -116885
rect -1500 -117720 -500 -117715
rect -1500 -117755 -790 -117720
rect -590 -117755 -500 -117720
rect -1500 -117760 -500 -117755
rect -375 -118385 -320 -116920
rect -280 -117720 -130 -117715
rect -280 -117755 -270 -117720
rect -280 -117760 -130 -117755
rect -375 -118420 -370 -118385
rect -325 -118420 -320 -118385
rect -375 -118500 -320 -118420
rect 270 -118540 1390 -118530
rect 270 -118600 280 -118540
rect 1380 -118590 1390 -118540
rect 1060 -118600 1390 -118590
rect 1770 -118540 2890 -118530
rect 1770 -118600 1780 -118540
rect 2880 -118590 2890 -118540
rect 2560 -118600 2890 -118590
rect 3270 -118540 4390 -118530
rect 3270 -118600 3280 -118540
rect 4380 -118590 4390 -118540
rect 4060 -118600 4390 -118590
rect 4770 -118540 5890 -118530
rect 4770 -118600 4780 -118540
rect 5880 -118590 5890 -118540
rect 5560 -118600 5890 -118590
rect 6270 -118540 7390 -118530
rect 6270 -118600 6280 -118540
rect 7380 -118590 7390 -118540
rect 7060 -118600 7390 -118590
rect 7770 -118540 8890 -118530
rect 7770 -118600 7780 -118540
rect 8880 -118590 8890 -118540
rect 8560 -118600 8890 -118590
rect 9270 -118540 10390 -118530
rect 9270 -118600 9280 -118540
rect 10380 -118590 10390 -118540
rect 10060 -118600 10390 -118590
rect 10770 -118540 11890 -118530
rect 10770 -118600 10780 -118540
rect 11880 -118590 11890 -118540
rect 11560 -118600 11890 -118590
rect 12270 -118540 13390 -118530
rect 12270 -118600 12280 -118540
rect 13380 -118590 13390 -118540
rect 13060 -118600 13390 -118590
rect 13770 -118540 14890 -118530
rect 13770 -118600 13780 -118540
rect 14880 -118590 14890 -118540
rect 14560 -118600 14890 -118590
rect 15270 -118540 16390 -118530
rect 15270 -118600 15280 -118540
rect 16380 -118590 16390 -118540
rect 16060 -118600 16390 -118590
rect 16770 -118540 17890 -118530
rect 16770 -118600 16780 -118540
rect 17880 -118590 17890 -118540
rect 17560 -118600 17890 -118590
rect 18270 -118540 19390 -118530
rect 18270 -118600 18280 -118540
rect 19380 -118590 19390 -118540
rect 19060 -118600 19390 -118590
rect 19770 -118540 20890 -118530
rect 19770 -118600 19780 -118540
rect 20880 -118590 20890 -118540
rect 20560 -118600 20890 -118590
rect 21270 -118540 22390 -118530
rect 21270 -118600 21280 -118540
rect 22380 -118590 22390 -118540
rect 22060 -118600 22390 -118590
rect 22770 -118540 23890 -118530
rect 22770 -118600 22780 -118540
rect 23880 -118590 23890 -118540
rect 23560 -118600 23890 -118590
rect 24270 -118540 25390 -118530
rect 24270 -118600 24280 -118540
rect 25380 -118590 25390 -118540
rect 25060 -118600 25390 -118590
rect 25770 -118540 26890 -118530
rect 25770 -118600 25780 -118540
rect 26880 -118590 26890 -118540
rect 26560 -118600 26890 -118590
rect 27270 -118540 28390 -118530
rect 27270 -118600 27280 -118540
rect 28380 -118590 28390 -118540
rect 28060 -118600 28390 -118590
rect 28770 -118540 29890 -118530
rect 28770 -118600 28780 -118540
rect 29880 -118590 29890 -118540
rect 29560 -118600 29890 -118590
rect 30270 -118540 31390 -118530
rect 30270 -118600 30280 -118540
rect 31380 -118590 31390 -118540
rect 31060 -118600 31390 -118590
rect 31770 -118540 32890 -118530
rect 31770 -118600 31780 -118540
rect 32880 -118590 32890 -118540
rect 32560 -118600 32890 -118590
rect 33270 -118540 34390 -118530
rect 33270 -118600 33280 -118540
rect 34380 -118590 34390 -118540
rect 34060 -118600 34390 -118590
rect 34770 -118540 35890 -118530
rect 34770 -118600 34780 -118540
rect 35880 -118590 35890 -118540
rect 35560 -118600 35890 -118590
rect 36270 -118540 37390 -118530
rect 36270 -118600 36280 -118540
rect 37380 -118590 37390 -118540
rect 37060 -118600 37390 -118590
rect 37770 -118540 38890 -118530
rect 37770 -118600 37780 -118540
rect 38880 -118590 38890 -118540
rect 38560 -118600 38890 -118590
rect 39270 -118540 40390 -118530
rect 39270 -118600 39280 -118540
rect 40380 -118590 40390 -118540
rect 40060 -118600 40390 -118590
rect 40770 -118540 41890 -118530
rect 40770 -118600 40780 -118540
rect 41880 -118590 41890 -118540
rect 41560 -118600 41890 -118590
rect 42270 -118540 43390 -118530
rect 42270 -118600 42280 -118540
rect 43380 -118590 43390 -118540
rect 43060 -118600 43390 -118590
rect 43770 -118540 44890 -118530
rect 43770 -118600 43780 -118540
rect 44880 -118590 44890 -118540
rect 44560 -118600 44890 -118590
rect 45270 -118540 46390 -118530
rect 45270 -118600 45280 -118540
rect 46380 -118590 46390 -118540
rect 46060 -118600 46390 -118590
rect 46770 -118540 47890 -118530
rect 46770 -118600 46780 -118540
rect 47880 -118590 47890 -118540
rect 47560 -118600 47890 -118590
rect 48270 -118540 49390 -118530
rect 48270 -118600 48280 -118540
rect 49380 -118590 49390 -118540
rect 49060 -118600 49390 -118590
rect 49770 -118540 50890 -118530
rect 49770 -118600 49780 -118540
rect 50880 -118590 50890 -118540
rect 50560 -118600 50890 -118590
rect 51270 -118540 52390 -118530
rect 51270 -118600 51280 -118540
rect 52380 -118590 52390 -118540
rect 52060 -118600 52390 -118590
rect 52770 -118540 53890 -118530
rect 52770 -118600 52780 -118540
rect 53880 -118590 53890 -118540
rect 53560 -118600 53890 -118590
rect 54270 -118540 55390 -118530
rect 54270 -118600 54280 -118540
rect 55380 -118590 55390 -118540
rect 55060 -118600 55390 -118590
rect 55770 -118540 56890 -118530
rect 55770 -118600 55780 -118540
rect 56880 -118590 56890 -118540
rect 56560 -118600 56890 -118590
rect 57270 -118540 58390 -118530
rect 57270 -118600 57280 -118540
rect 58380 -118590 58390 -118540
rect 58060 -118600 58390 -118590
rect 58770 -118540 59890 -118530
rect 58770 -118600 58780 -118540
rect 59880 -118590 59890 -118540
rect 59560 -118600 59890 -118590
rect 60270 -118540 61390 -118530
rect 60270 -118600 60280 -118540
rect 61380 -118590 61390 -118540
rect 61060 -118600 61390 -118590
rect 61770 -118540 62890 -118530
rect 61770 -118600 61780 -118540
rect 62880 -118590 62890 -118540
rect 62560 -118600 62890 -118590
rect 63270 -118540 64390 -118530
rect 63270 -118600 63280 -118540
rect 64380 -118590 64390 -118540
rect 64060 -118600 64390 -118590
rect 64770 -118540 65890 -118530
rect 64770 -118600 64780 -118540
rect 65880 -118590 65890 -118540
rect 65560 -118600 65890 -118590
rect 66270 -118540 67390 -118530
rect 66270 -118600 66280 -118540
rect 67380 -118590 67390 -118540
rect 67060 -118600 67390 -118590
rect 67770 -118540 68890 -118530
rect 67770 -118600 67780 -118540
rect 68880 -118590 68890 -118540
rect 68560 -118600 68890 -118590
rect 69270 -118540 70390 -118530
rect 69270 -118600 69280 -118540
rect 70380 -118590 70390 -118540
rect 70060 -118600 70390 -118590
rect 70770 -118540 71890 -118530
rect 70770 -118600 70780 -118540
rect 71880 -118590 71890 -118540
rect 71560 -118600 71890 -118590
rect 72270 -118540 73390 -118530
rect 72270 -118600 72280 -118540
rect 73380 -118590 73390 -118540
rect 73060 -118600 73390 -118590
rect 73770 -118540 74890 -118530
rect 73770 -118600 73780 -118540
rect 74880 -118590 74890 -118540
rect 74560 -118600 74890 -118590
rect 75270 -118540 76390 -118530
rect 75270 -118600 75280 -118540
rect 76380 -118590 76390 -118540
rect 76060 -118600 76390 -118590
rect 76770 -118540 77890 -118530
rect 76770 -118600 76780 -118540
rect 77880 -118590 77890 -118540
rect 77560 -118600 77890 -118590
rect 78270 -118540 79390 -118530
rect 78270 -118600 78280 -118540
rect 79380 -118590 79390 -118540
rect 79060 -118600 79390 -118590
rect 79770 -118540 80890 -118530
rect 79770 -118600 79780 -118540
rect 80880 -118590 80890 -118540
rect 80560 -118600 80890 -118590
rect 81270 -118540 82390 -118530
rect 81270 -118600 81280 -118540
rect 82380 -118590 82390 -118540
rect 82060 -118600 82390 -118590
rect 82770 -118540 83890 -118530
rect 82770 -118600 82780 -118540
rect 83880 -118590 83890 -118540
rect 83560 -118600 83890 -118590
rect 84270 -118540 85390 -118530
rect 84270 -118600 84280 -118540
rect 85380 -118590 85390 -118540
rect 85060 -118600 85390 -118590
rect 85770 -118540 86890 -118530
rect 85770 -118600 85780 -118540
rect 86880 -118590 86890 -118540
rect 86560 -118600 86890 -118590
rect 87270 -118540 88390 -118530
rect 87270 -118600 87280 -118540
rect 88380 -118590 88390 -118540
rect 88060 -118600 88390 -118590
rect 88770 -118540 89890 -118530
rect 88770 -118600 88780 -118540
rect 89880 -118590 89890 -118540
rect 89560 -118600 89890 -118590
rect 90270 -118540 91390 -118530
rect 90270 -118600 90280 -118540
rect 91380 -118590 91390 -118540
rect 91060 -118600 91390 -118590
rect 91770 -118540 92890 -118530
rect 91770 -118600 91780 -118540
rect 92880 -118590 92890 -118540
rect 92560 -118600 92890 -118590
rect 93270 -118540 94390 -118530
rect 93270 -118600 93280 -118540
rect 94380 -118590 94390 -118540
rect 94060 -118600 94390 -118590
rect 94770 -118540 95890 -118530
rect 94770 -118600 94780 -118540
rect 95880 -118590 95890 -118540
rect 95560 -118600 95890 -118590
rect 96270 -118540 97390 -118530
rect 96270 -118600 96280 -118540
rect 97380 -118590 97390 -118540
rect 97060 -118600 97390 -118590
rect 97770 -118540 98890 -118530
rect 97770 -118600 97780 -118540
rect 98880 -118590 98890 -118540
rect 98560 -118600 98890 -118590
rect 99270 -118540 100390 -118530
rect 99270 -118600 99280 -118540
rect 100380 -118590 100390 -118540
rect 100060 -118600 100390 -118590
rect 100770 -118540 101890 -118530
rect 100770 -118600 100780 -118540
rect 101880 -118590 101890 -118540
rect 101560 -118600 101890 -118590
rect 102270 -118540 103390 -118530
rect 102270 -118600 102280 -118540
rect 103380 -118590 103390 -118540
rect 103060 -118600 103390 -118590
rect 103770 -118540 104890 -118530
rect 103770 -118600 103780 -118540
rect 104880 -118590 104890 -118540
rect 104560 -118600 104890 -118590
rect 105270 -118540 106390 -118530
rect 105270 -118600 105280 -118540
rect 106380 -118590 106390 -118540
rect 106060 -118600 106390 -118590
rect 106770 -118540 107890 -118530
rect 106770 -118600 106780 -118540
rect 107880 -118590 107890 -118540
rect 107560 -118600 107890 -118590
rect 108270 -118540 109390 -118530
rect 108270 -118600 108280 -118540
rect 109380 -118590 109390 -118540
rect 109060 -118600 109390 -118590
rect 109770 -118540 110890 -118530
rect 109770 -118600 109780 -118540
rect 110880 -118590 110890 -118540
rect 110560 -118600 110890 -118590
rect 111270 -118540 112390 -118530
rect 111270 -118600 111280 -118540
rect 112380 -118590 112390 -118540
rect 112060 -118600 112390 -118590
rect 112770 -118540 113890 -118530
rect 112770 -118600 112780 -118540
rect 113880 -118590 113890 -118540
rect 113560 -118600 113890 -118590
rect 114270 -118540 115390 -118530
rect 114270 -118600 114280 -118540
rect 115380 -118590 115390 -118540
rect 115060 -118600 115390 -118590
rect 115770 -118540 116890 -118530
rect 115770 -118600 115780 -118540
rect 116880 -118590 116890 -118540
rect 116560 -118600 116890 -118590
rect 117270 -118540 118390 -118530
rect 117270 -118600 117280 -118540
rect 118380 -118590 118390 -118540
rect 118060 -118600 118390 -118590
rect 118770 -118540 119890 -118530
rect 118770 -118600 118780 -118540
rect 119880 -118590 119890 -118540
rect 119560 -118600 119890 -118590
rect 110 -118750 220 -118745
rect 110 -118850 120 -118750
rect 210 -118850 220 -118750
rect 110 -118855 220 -118850
rect 1610 -118750 1720 -118745
rect 1610 -118850 1620 -118750
rect 1710 -118850 1720 -118750
rect 1610 -118855 1720 -118850
rect 3110 -118750 3220 -118745
rect 3110 -118850 3120 -118750
rect 3210 -118850 3220 -118750
rect 3110 -118855 3220 -118850
rect 4610 -118750 4720 -118745
rect 4610 -118850 4620 -118750
rect 4710 -118850 4720 -118750
rect 4610 -118855 4720 -118850
rect 6110 -118750 6220 -118745
rect 6110 -118850 6120 -118750
rect 6210 -118850 6220 -118750
rect 6110 -118855 6220 -118850
rect 7610 -118750 7720 -118745
rect 7610 -118850 7620 -118750
rect 7710 -118850 7720 -118750
rect 7610 -118855 7720 -118850
rect 9110 -118750 9220 -118745
rect 9110 -118850 9120 -118750
rect 9210 -118850 9220 -118750
rect 9110 -118855 9220 -118850
rect 10610 -118750 10720 -118745
rect 10610 -118850 10620 -118750
rect 10710 -118850 10720 -118750
rect 10610 -118855 10720 -118850
rect 12110 -118750 12220 -118745
rect 12110 -118850 12120 -118750
rect 12210 -118850 12220 -118750
rect 12110 -118855 12220 -118850
rect 13610 -118750 13720 -118745
rect 13610 -118850 13620 -118750
rect 13710 -118850 13720 -118750
rect 13610 -118855 13720 -118850
rect 15110 -118750 15220 -118745
rect 15110 -118850 15120 -118750
rect 15210 -118850 15220 -118750
rect 15110 -118855 15220 -118850
rect 16610 -118750 16720 -118745
rect 16610 -118850 16620 -118750
rect 16710 -118850 16720 -118750
rect 16610 -118855 16720 -118850
rect 18110 -118750 18220 -118745
rect 18110 -118850 18120 -118750
rect 18210 -118850 18220 -118750
rect 18110 -118855 18220 -118850
rect 19610 -118750 19720 -118745
rect 19610 -118850 19620 -118750
rect 19710 -118850 19720 -118750
rect 19610 -118855 19720 -118850
rect 21110 -118750 21220 -118745
rect 21110 -118850 21120 -118750
rect 21210 -118850 21220 -118750
rect 21110 -118855 21220 -118850
rect 22610 -118750 22720 -118745
rect 22610 -118850 22620 -118750
rect 22710 -118850 22720 -118750
rect 22610 -118855 22720 -118850
rect 24110 -118750 24220 -118745
rect 24110 -118850 24120 -118750
rect 24210 -118850 24220 -118750
rect 24110 -118855 24220 -118850
rect 25610 -118750 25720 -118745
rect 25610 -118850 25620 -118750
rect 25710 -118850 25720 -118750
rect 25610 -118855 25720 -118850
rect 27110 -118750 27220 -118745
rect 27110 -118850 27120 -118750
rect 27210 -118850 27220 -118750
rect 27110 -118855 27220 -118850
rect 28610 -118750 28720 -118745
rect 28610 -118850 28620 -118750
rect 28710 -118850 28720 -118750
rect 28610 -118855 28720 -118850
rect 30110 -118750 30220 -118745
rect 30110 -118850 30120 -118750
rect 30210 -118850 30220 -118750
rect 30110 -118855 30220 -118850
rect 31610 -118750 31720 -118745
rect 31610 -118850 31620 -118750
rect 31710 -118850 31720 -118750
rect 31610 -118855 31720 -118850
rect 33110 -118750 33220 -118745
rect 33110 -118850 33120 -118750
rect 33210 -118850 33220 -118750
rect 33110 -118855 33220 -118850
rect 34610 -118750 34720 -118745
rect 34610 -118850 34620 -118750
rect 34710 -118850 34720 -118750
rect 34610 -118855 34720 -118850
rect 36110 -118750 36220 -118745
rect 36110 -118850 36120 -118750
rect 36210 -118850 36220 -118750
rect 36110 -118855 36220 -118850
rect 37610 -118750 37720 -118745
rect 37610 -118850 37620 -118750
rect 37710 -118850 37720 -118750
rect 37610 -118855 37720 -118850
rect 39110 -118750 39220 -118745
rect 39110 -118850 39120 -118750
rect 39210 -118850 39220 -118750
rect 39110 -118855 39220 -118850
rect 40610 -118750 40720 -118745
rect 40610 -118850 40620 -118750
rect 40710 -118850 40720 -118750
rect 40610 -118855 40720 -118850
rect 42110 -118750 42220 -118745
rect 42110 -118850 42120 -118750
rect 42210 -118850 42220 -118750
rect 42110 -118855 42220 -118850
rect 43610 -118750 43720 -118745
rect 43610 -118850 43620 -118750
rect 43710 -118850 43720 -118750
rect 43610 -118855 43720 -118850
rect 45110 -118750 45220 -118745
rect 45110 -118850 45120 -118750
rect 45210 -118850 45220 -118750
rect 45110 -118855 45220 -118850
rect 46610 -118750 46720 -118745
rect 46610 -118850 46620 -118750
rect 46710 -118850 46720 -118750
rect 46610 -118855 46720 -118850
rect 48110 -118750 48220 -118745
rect 48110 -118850 48120 -118750
rect 48210 -118850 48220 -118750
rect 48110 -118855 48220 -118850
rect 49610 -118750 49720 -118745
rect 49610 -118850 49620 -118750
rect 49710 -118850 49720 -118750
rect 49610 -118855 49720 -118850
rect 51110 -118750 51220 -118745
rect 51110 -118850 51120 -118750
rect 51210 -118850 51220 -118750
rect 51110 -118855 51220 -118850
rect 52610 -118750 52720 -118745
rect 52610 -118850 52620 -118750
rect 52710 -118850 52720 -118750
rect 52610 -118855 52720 -118850
rect 54110 -118750 54220 -118745
rect 54110 -118850 54120 -118750
rect 54210 -118850 54220 -118750
rect 54110 -118855 54220 -118850
rect 55610 -118750 55720 -118745
rect 55610 -118850 55620 -118750
rect 55710 -118850 55720 -118750
rect 55610 -118855 55720 -118850
rect 57110 -118750 57220 -118745
rect 57110 -118850 57120 -118750
rect 57210 -118850 57220 -118750
rect 57110 -118855 57220 -118850
rect 58610 -118750 58720 -118745
rect 58610 -118850 58620 -118750
rect 58710 -118850 58720 -118750
rect 58610 -118855 58720 -118850
rect 60110 -118750 60220 -118745
rect 60110 -118850 60120 -118750
rect 60210 -118850 60220 -118750
rect 60110 -118855 60220 -118850
rect 61610 -118750 61720 -118745
rect 61610 -118850 61620 -118750
rect 61710 -118850 61720 -118750
rect 61610 -118855 61720 -118850
rect 63110 -118750 63220 -118745
rect 63110 -118850 63120 -118750
rect 63210 -118850 63220 -118750
rect 63110 -118855 63220 -118850
rect 64610 -118750 64720 -118745
rect 64610 -118850 64620 -118750
rect 64710 -118850 64720 -118750
rect 64610 -118855 64720 -118850
rect 66110 -118750 66220 -118745
rect 66110 -118850 66120 -118750
rect 66210 -118850 66220 -118750
rect 66110 -118855 66220 -118850
rect 67610 -118750 67720 -118745
rect 67610 -118850 67620 -118750
rect 67710 -118850 67720 -118750
rect 67610 -118855 67720 -118850
rect 69110 -118750 69220 -118745
rect 69110 -118850 69120 -118750
rect 69210 -118850 69220 -118750
rect 69110 -118855 69220 -118850
rect 70610 -118750 70720 -118745
rect 70610 -118850 70620 -118750
rect 70710 -118850 70720 -118750
rect 70610 -118855 70720 -118850
rect 72110 -118750 72220 -118745
rect 72110 -118850 72120 -118750
rect 72210 -118850 72220 -118750
rect 72110 -118855 72220 -118850
rect 73610 -118750 73720 -118745
rect 73610 -118850 73620 -118750
rect 73710 -118850 73720 -118750
rect 73610 -118855 73720 -118850
rect 75110 -118750 75220 -118745
rect 75110 -118850 75120 -118750
rect 75210 -118850 75220 -118750
rect 75110 -118855 75220 -118850
rect 76610 -118750 76720 -118745
rect 76610 -118850 76620 -118750
rect 76710 -118850 76720 -118750
rect 76610 -118855 76720 -118850
rect 78110 -118750 78220 -118745
rect 78110 -118850 78120 -118750
rect 78210 -118850 78220 -118750
rect 78110 -118855 78220 -118850
rect 79610 -118750 79720 -118745
rect 79610 -118850 79620 -118750
rect 79710 -118850 79720 -118750
rect 79610 -118855 79720 -118850
rect 81110 -118750 81220 -118745
rect 81110 -118850 81120 -118750
rect 81210 -118850 81220 -118750
rect 81110 -118855 81220 -118850
rect 82610 -118750 82720 -118745
rect 82610 -118850 82620 -118750
rect 82710 -118850 82720 -118750
rect 82610 -118855 82720 -118850
rect 84110 -118750 84220 -118745
rect 84110 -118850 84120 -118750
rect 84210 -118850 84220 -118750
rect 84110 -118855 84220 -118850
rect 85610 -118750 85720 -118745
rect 85610 -118850 85620 -118750
rect 85710 -118850 85720 -118750
rect 85610 -118855 85720 -118850
rect 87110 -118750 87220 -118745
rect 87110 -118850 87120 -118750
rect 87210 -118850 87220 -118750
rect 87110 -118855 87220 -118850
rect 88610 -118750 88720 -118745
rect 88610 -118850 88620 -118750
rect 88710 -118850 88720 -118750
rect 88610 -118855 88720 -118850
rect 90110 -118750 90220 -118745
rect 90110 -118850 90120 -118750
rect 90210 -118850 90220 -118750
rect 90110 -118855 90220 -118850
rect 91610 -118750 91720 -118745
rect 91610 -118850 91620 -118750
rect 91710 -118850 91720 -118750
rect 91610 -118855 91720 -118850
rect 93110 -118750 93220 -118745
rect 93110 -118850 93120 -118750
rect 93210 -118850 93220 -118750
rect 93110 -118855 93220 -118850
rect 94610 -118750 94720 -118745
rect 94610 -118850 94620 -118750
rect 94710 -118850 94720 -118750
rect 94610 -118855 94720 -118850
rect 96110 -118750 96220 -118745
rect 96110 -118850 96120 -118750
rect 96210 -118850 96220 -118750
rect 96110 -118855 96220 -118850
rect 97610 -118750 97720 -118745
rect 97610 -118850 97620 -118750
rect 97710 -118850 97720 -118750
rect 97610 -118855 97720 -118850
rect 99110 -118750 99220 -118745
rect 99110 -118850 99120 -118750
rect 99210 -118850 99220 -118750
rect 99110 -118855 99220 -118850
rect 100610 -118750 100720 -118745
rect 100610 -118850 100620 -118750
rect 100710 -118850 100720 -118750
rect 100610 -118855 100720 -118850
rect 102110 -118750 102220 -118745
rect 102110 -118850 102120 -118750
rect 102210 -118850 102220 -118750
rect 102110 -118855 102220 -118850
rect 103610 -118750 103720 -118745
rect 103610 -118850 103620 -118750
rect 103710 -118850 103720 -118750
rect 103610 -118855 103720 -118850
rect 105110 -118750 105220 -118745
rect 105110 -118850 105120 -118750
rect 105210 -118850 105220 -118750
rect 105110 -118855 105220 -118850
rect 106610 -118750 106720 -118745
rect 106610 -118850 106620 -118750
rect 106710 -118850 106720 -118750
rect 106610 -118855 106720 -118850
rect 108110 -118750 108220 -118745
rect 108110 -118850 108120 -118750
rect 108210 -118850 108220 -118750
rect 108110 -118855 108220 -118850
rect 109610 -118750 109720 -118745
rect 109610 -118850 109620 -118750
rect 109710 -118850 109720 -118750
rect 109610 -118855 109720 -118850
rect 111110 -118750 111220 -118745
rect 111110 -118850 111120 -118750
rect 111210 -118850 111220 -118750
rect 111110 -118855 111220 -118850
rect 112610 -118750 112720 -118745
rect 112610 -118850 112620 -118750
rect 112710 -118850 112720 -118750
rect 112610 -118855 112720 -118850
rect 114110 -118750 114220 -118745
rect 114110 -118850 114120 -118750
rect 114210 -118850 114220 -118750
rect 114110 -118855 114220 -118850
rect 115610 -118750 115720 -118745
rect 115610 -118850 115620 -118750
rect 115710 -118850 115720 -118750
rect 115610 -118855 115720 -118850
rect 117110 -118750 117220 -118745
rect 117110 -118850 117120 -118750
rect 117210 -118850 117220 -118750
rect 117110 -118855 117220 -118850
rect 118610 -118750 118720 -118745
rect 118610 -118850 118620 -118750
rect 118710 -118850 118720 -118750
rect 118610 -118855 118720 -118850
rect 270 -118960 120370 -118950
rect 270 -119040 280 -118960
rect 270 -119050 120370 -119040
<< via2 >>
rect 245 1780 290 1825
rect 1745 1780 1790 1825
rect 3245 1780 3290 1825
rect 4745 1780 4790 1825
rect 6245 1780 6290 1825
rect 7745 1780 7790 1825
rect 9245 1780 9290 1825
rect 10745 1780 10790 1825
rect 12245 1780 12290 1825
rect 13745 1780 13790 1825
rect 15245 1780 15290 1825
rect 16745 1780 16790 1825
rect 18245 1780 18290 1825
rect 19745 1780 19790 1825
rect 21245 1780 21290 1825
rect 22745 1780 22790 1825
rect 24245 1780 24290 1825
rect 25745 1780 25790 1825
rect 27245 1780 27290 1825
rect 28745 1780 28790 1825
rect 30245 1780 30290 1825
rect 31745 1780 31790 1825
rect 33245 1780 33290 1825
rect 34745 1780 34790 1825
rect 36245 1780 36290 1825
rect 37745 1780 37790 1825
rect 39245 1780 39290 1825
rect 40745 1780 40790 1825
rect 42245 1780 42290 1825
rect 43745 1780 43790 1825
rect 45245 1780 45290 1825
rect 46745 1780 46790 1825
rect 48245 1780 48290 1825
rect 49745 1780 49790 1825
rect 51245 1780 51290 1825
rect 52745 1780 52790 1825
rect 54245 1780 54290 1825
rect 55745 1780 55790 1825
rect 57245 1780 57290 1825
rect 58745 1780 58790 1825
rect 60245 1780 60290 1825
rect 61745 1780 61790 1825
rect 63245 1780 63290 1825
rect 64745 1780 64790 1825
rect 66245 1780 66290 1825
rect 67745 1780 67790 1825
rect 69245 1780 69290 1825
rect 70745 1780 70790 1825
rect 72245 1780 72290 1825
rect 73745 1780 73790 1825
rect 75245 1780 75290 1825
rect 76745 1780 76790 1825
rect 78245 1780 78290 1825
rect 79745 1780 79790 1825
rect 81245 1780 81290 1825
rect 82745 1780 82790 1825
rect 84245 1780 84290 1825
rect 85745 1780 85790 1825
rect 87245 1780 87290 1825
rect 88745 1780 88790 1825
rect 90245 1780 90290 1825
rect 91745 1780 91790 1825
rect 93245 1780 93290 1825
rect 94745 1780 94790 1825
rect 96245 1780 96290 1825
rect 97745 1780 97790 1825
rect 99245 1780 99290 1825
rect 100745 1780 100790 1825
rect 102245 1780 102290 1825
rect 103745 1780 103790 1825
rect 105245 1780 105290 1825
rect 106745 1780 106790 1825
rect 108245 1780 108290 1825
rect 109745 1780 109790 1825
rect 111245 1780 111290 1825
rect 112745 1780 112790 1825
rect 114245 1780 114290 1825
rect 115745 1780 115790 1825
rect 117245 1780 117290 1825
rect 118745 1780 118790 1825
rect -270 745 -130 780
rect -370 80 -325 115
rect -270 -755 -130 -720
rect -370 -1420 -325 -1385
rect -270 -2255 -130 -2220
rect -370 -2920 -325 -2885
rect -270 -3755 -130 -3720
rect -370 -4420 -325 -4385
rect -270 -5255 -130 -5220
rect -370 -5920 -325 -5885
rect -270 -6755 -130 -6720
rect -370 -7420 -325 -7385
rect -270 -8255 -130 -8220
rect -370 -8920 -325 -8885
rect -270 -9755 -130 -9720
rect -370 -10420 -325 -10385
rect -270 -11255 -130 -11220
rect -370 -11920 -325 -11885
rect -270 -12755 -130 -12720
rect -370 -13420 -325 -13385
rect -270 -14255 -130 -14220
rect -370 -14920 -325 -14885
rect -270 -15755 -130 -15720
rect -370 -16420 -325 -16385
rect -270 -17255 -130 -17220
rect -370 -17920 -325 -17885
rect -270 -18755 -130 -18720
rect -370 -19420 -325 -19385
rect -270 -20255 -130 -20220
rect -370 -20920 -325 -20885
rect -270 -21755 -130 -21720
rect -370 -22420 -325 -22385
rect -270 -23255 -130 -23220
rect -370 -23920 -325 -23885
rect -270 -24755 -130 -24720
rect -370 -25420 -325 -25385
rect -270 -26255 -130 -26220
rect -370 -26920 -325 -26885
rect -270 -27755 -130 -27720
rect -370 -28420 -325 -28385
rect -270 -29255 -130 -29220
rect -370 -29920 -325 -29885
rect -270 -30755 -130 -30720
rect -370 -31420 -325 -31385
rect -270 -32255 -130 -32220
rect -370 -32920 -325 -32885
rect -270 -33755 -130 -33720
rect -370 -34420 -325 -34385
rect -270 -35255 -130 -35220
rect -370 -35920 -325 -35885
rect -270 -36755 -130 -36720
rect -370 -37420 -325 -37385
rect -270 -38255 -130 -38220
rect -370 -38920 -325 -38885
rect -270 -39755 -130 -39720
rect -370 -40420 -325 -40385
rect -270 -41255 -130 -41220
rect -370 -41920 -325 -41885
rect -270 -42755 -130 -42720
rect -370 -43420 -325 -43385
rect -270 -44255 -130 -44220
rect -370 -44920 -325 -44885
rect -270 -45755 -130 -45720
rect -370 -46420 -325 -46385
rect -270 -47255 -130 -47220
rect -370 -47920 -325 -47885
rect -270 -48755 -130 -48720
rect -370 -49420 -325 -49385
rect -270 -50255 -130 -50220
rect -370 -50920 -325 -50885
rect -270 -51755 -130 -51720
rect -370 -52420 -325 -52385
rect -270 -53255 -130 -53220
rect -370 -53920 -325 -53885
rect -270 -54755 -130 -54720
rect -370 -55420 -325 -55385
rect -270 -56255 -130 -56220
rect -370 -56920 -325 -56885
rect -270 -57755 -130 -57720
rect -370 -58420 -325 -58385
rect -270 -59255 -130 -59220
rect -370 -59920 -325 -59885
rect -270 -60755 -130 -60720
rect -370 -61420 -325 -61385
rect -270 -62255 -130 -62220
rect -370 -62920 -325 -62885
rect -270 -63755 -130 -63720
rect -370 -64420 -325 -64385
rect -270 -65255 -130 -65220
rect -370 -65920 -325 -65885
rect -270 -66755 -130 -66720
rect -370 -67420 -325 -67385
rect -270 -68255 -130 -68220
rect -370 -68920 -325 -68885
rect -270 -69755 -130 -69720
rect -370 -70420 -325 -70385
rect -270 -71255 -130 -71220
rect -370 -71920 -325 -71885
rect -270 -72755 -130 -72720
rect -370 -73420 -325 -73385
rect -270 -74255 -130 -74220
rect -370 -74920 -325 -74885
rect -270 -75755 -130 -75720
rect -370 -76420 -325 -76385
rect -270 -77255 -130 -77220
rect -370 -77920 -325 -77885
rect -270 -78755 -130 -78720
rect -370 -79420 -325 -79385
rect -270 -80255 -130 -80220
rect -370 -80920 -325 -80885
rect -270 -81755 -130 -81720
rect -370 -82420 -325 -82385
rect -270 -83255 -130 -83220
rect -370 -83920 -325 -83885
rect -270 -84755 -130 -84720
rect -370 -85420 -325 -85385
rect -270 -86255 -130 -86220
rect -370 -86920 -325 -86885
rect -270 -87755 -130 -87720
rect -370 -88420 -325 -88385
rect -270 -89255 -130 -89220
rect -370 -89920 -325 -89885
rect -270 -90755 -130 -90720
rect -370 -91420 -325 -91385
rect -270 -92255 -130 -92220
rect -370 -92920 -325 -92885
rect -270 -93755 -130 -93720
rect -370 -94420 -325 -94385
rect -270 -95255 -130 -95220
rect -370 -95920 -325 -95885
rect -270 -96755 -130 -96720
rect -370 -97420 -325 -97385
rect -270 -98255 -130 -98220
rect -370 -98920 -325 -98885
rect -270 -99755 -130 -99720
rect -370 -100420 -325 -100385
rect -270 -101255 -130 -101220
rect -370 -101920 -325 -101885
rect -270 -102755 -130 -102720
rect -370 -103420 -325 -103385
rect -270 -104255 -130 -104220
rect -370 -104920 -325 -104885
rect -270 -105755 -130 -105720
rect -370 -106420 -325 -106385
rect -270 -107255 -130 -107220
rect -370 -107920 -325 -107885
rect -270 -108755 -130 -108720
rect -370 -109420 -325 -109385
rect -270 -110255 -130 -110220
rect -370 -110920 -325 -110885
rect -270 -111755 -130 -111720
rect -370 -112420 -325 -112385
rect -270 -113255 -130 -113220
rect -370 -113920 -325 -113885
rect -270 -114755 -130 -114720
rect -370 -115420 -325 -115385
rect -270 -116255 -130 -116220
rect -370 -116920 -325 -116885
rect -270 -117755 -130 -117720
rect -370 -118420 -325 -118385
rect 280 -118565 1380 -118540
rect 280 -118590 1060 -118565
rect 1060 -118590 1380 -118565
rect 1780 -118565 2880 -118540
rect 1780 -118590 2560 -118565
rect 2560 -118590 2880 -118565
rect 3280 -118565 4380 -118540
rect 3280 -118590 4060 -118565
rect 4060 -118590 4380 -118565
rect 4780 -118565 5880 -118540
rect 4780 -118590 5560 -118565
rect 5560 -118590 5880 -118565
rect 6280 -118565 7380 -118540
rect 6280 -118590 7060 -118565
rect 7060 -118590 7380 -118565
rect 7780 -118565 8880 -118540
rect 7780 -118590 8560 -118565
rect 8560 -118590 8880 -118565
rect 9280 -118565 10380 -118540
rect 9280 -118590 10060 -118565
rect 10060 -118590 10380 -118565
rect 10780 -118565 11880 -118540
rect 10780 -118590 11560 -118565
rect 11560 -118590 11880 -118565
rect 12280 -118565 13380 -118540
rect 12280 -118590 13060 -118565
rect 13060 -118590 13380 -118565
rect 13780 -118565 14880 -118540
rect 13780 -118590 14560 -118565
rect 14560 -118590 14880 -118565
rect 15280 -118565 16380 -118540
rect 15280 -118590 16060 -118565
rect 16060 -118590 16380 -118565
rect 16780 -118565 17880 -118540
rect 16780 -118590 17560 -118565
rect 17560 -118590 17880 -118565
rect 18280 -118565 19380 -118540
rect 18280 -118590 19060 -118565
rect 19060 -118590 19380 -118565
rect 19780 -118565 20880 -118540
rect 19780 -118590 20560 -118565
rect 20560 -118590 20880 -118565
rect 21280 -118565 22380 -118540
rect 21280 -118590 22060 -118565
rect 22060 -118590 22380 -118565
rect 22780 -118565 23880 -118540
rect 22780 -118590 23560 -118565
rect 23560 -118590 23880 -118565
rect 24280 -118565 25380 -118540
rect 24280 -118590 25060 -118565
rect 25060 -118590 25380 -118565
rect 25780 -118565 26880 -118540
rect 25780 -118590 26560 -118565
rect 26560 -118590 26880 -118565
rect 27280 -118565 28380 -118540
rect 27280 -118590 28060 -118565
rect 28060 -118590 28380 -118565
rect 28780 -118565 29880 -118540
rect 28780 -118590 29560 -118565
rect 29560 -118590 29880 -118565
rect 30280 -118565 31380 -118540
rect 30280 -118590 31060 -118565
rect 31060 -118590 31380 -118565
rect 31780 -118565 32880 -118540
rect 31780 -118590 32560 -118565
rect 32560 -118590 32880 -118565
rect 33280 -118565 34380 -118540
rect 33280 -118590 34060 -118565
rect 34060 -118590 34380 -118565
rect 34780 -118565 35880 -118540
rect 34780 -118590 35560 -118565
rect 35560 -118590 35880 -118565
rect 36280 -118565 37380 -118540
rect 36280 -118590 37060 -118565
rect 37060 -118590 37380 -118565
rect 37780 -118565 38880 -118540
rect 37780 -118590 38560 -118565
rect 38560 -118590 38880 -118565
rect 39280 -118565 40380 -118540
rect 39280 -118590 40060 -118565
rect 40060 -118590 40380 -118565
rect 40780 -118565 41880 -118540
rect 40780 -118590 41560 -118565
rect 41560 -118590 41880 -118565
rect 42280 -118565 43380 -118540
rect 42280 -118590 43060 -118565
rect 43060 -118590 43380 -118565
rect 43780 -118565 44880 -118540
rect 43780 -118590 44560 -118565
rect 44560 -118590 44880 -118565
rect 45280 -118565 46380 -118540
rect 45280 -118590 46060 -118565
rect 46060 -118590 46380 -118565
rect 46780 -118565 47880 -118540
rect 46780 -118590 47560 -118565
rect 47560 -118590 47880 -118565
rect 48280 -118565 49380 -118540
rect 48280 -118590 49060 -118565
rect 49060 -118590 49380 -118565
rect 49780 -118565 50880 -118540
rect 49780 -118590 50560 -118565
rect 50560 -118590 50880 -118565
rect 51280 -118565 52380 -118540
rect 51280 -118590 52060 -118565
rect 52060 -118590 52380 -118565
rect 52780 -118565 53880 -118540
rect 52780 -118590 53560 -118565
rect 53560 -118590 53880 -118565
rect 54280 -118565 55380 -118540
rect 54280 -118590 55060 -118565
rect 55060 -118590 55380 -118565
rect 55780 -118565 56880 -118540
rect 55780 -118590 56560 -118565
rect 56560 -118590 56880 -118565
rect 57280 -118565 58380 -118540
rect 57280 -118590 58060 -118565
rect 58060 -118590 58380 -118565
rect 58780 -118565 59880 -118540
rect 58780 -118590 59560 -118565
rect 59560 -118590 59880 -118565
rect 60280 -118565 61380 -118540
rect 60280 -118590 61060 -118565
rect 61060 -118590 61380 -118565
rect 61780 -118565 62880 -118540
rect 61780 -118590 62560 -118565
rect 62560 -118590 62880 -118565
rect 63280 -118565 64380 -118540
rect 63280 -118590 64060 -118565
rect 64060 -118590 64380 -118565
rect 64780 -118565 65880 -118540
rect 64780 -118590 65560 -118565
rect 65560 -118590 65880 -118565
rect 66280 -118565 67380 -118540
rect 66280 -118590 67060 -118565
rect 67060 -118590 67380 -118565
rect 67780 -118565 68880 -118540
rect 67780 -118590 68560 -118565
rect 68560 -118590 68880 -118565
rect 69280 -118565 70380 -118540
rect 69280 -118590 70060 -118565
rect 70060 -118590 70380 -118565
rect 70780 -118565 71880 -118540
rect 70780 -118590 71560 -118565
rect 71560 -118590 71880 -118565
rect 72280 -118565 73380 -118540
rect 72280 -118590 73060 -118565
rect 73060 -118590 73380 -118565
rect 73780 -118565 74880 -118540
rect 73780 -118590 74560 -118565
rect 74560 -118590 74880 -118565
rect 75280 -118565 76380 -118540
rect 75280 -118590 76060 -118565
rect 76060 -118590 76380 -118565
rect 76780 -118565 77880 -118540
rect 76780 -118590 77560 -118565
rect 77560 -118590 77880 -118565
rect 78280 -118565 79380 -118540
rect 78280 -118590 79060 -118565
rect 79060 -118590 79380 -118565
rect 79780 -118565 80880 -118540
rect 79780 -118590 80560 -118565
rect 80560 -118590 80880 -118565
rect 81280 -118565 82380 -118540
rect 81280 -118590 82060 -118565
rect 82060 -118590 82380 -118565
rect 82780 -118565 83880 -118540
rect 82780 -118590 83560 -118565
rect 83560 -118590 83880 -118565
rect 84280 -118565 85380 -118540
rect 84280 -118590 85060 -118565
rect 85060 -118590 85380 -118565
rect 85780 -118565 86880 -118540
rect 85780 -118590 86560 -118565
rect 86560 -118590 86880 -118565
rect 87280 -118565 88380 -118540
rect 87280 -118590 88060 -118565
rect 88060 -118590 88380 -118565
rect 88780 -118565 89880 -118540
rect 88780 -118590 89560 -118565
rect 89560 -118590 89880 -118565
rect 90280 -118565 91380 -118540
rect 90280 -118590 91060 -118565
rect 91060 -118590 91380 -118565
rect 91780 -118565 92880 -118540
rect 91780 -118590 92560 -118565
rect 92560 -118590 92880 -118565
rect 93280 -118565 94380 -118540
rect 93280 -118590 94060 -118565
rect 94060 -118590 94380 -118565
rect 94780 -118565 95880 -118540
rect 94780 -118590 95560 -118565
rect 95560 -118590 95880 -118565
rect 96280 -118565 97380 -118540
rect 96280 -118590 97060 -118565
rect 97060 -118590 97380 -118565
rect 97780 -118565 98880 -118540
rect 97780 -118590 98560 -118565
rect 98560 -118590 98880 -118565
rect 99280 -118565 100380 -118540
rect 99280 -118590 100060 -118565
rect 100060 -118590 100380 -118565
rect 100780 -118565 101880 -118540
rect 100780 -118590 101560 -118565
rect 101560 -118590 101880 -118565
rect 102280 -118565 103380 -118540
rect 102280 -118590 103060 -118565
rect 103060 -118590 103380 -118565
rect 103780 -118565 104880 -118540
rect 103780 -118590 104560 -118565
rect 104560 -118590 104880 -118565
rect 105280 -118565 106380 -118540
rect 105280 -118590 106060 -118565
rect 106060 -118590 106380 -118565
rect 106780 -118565 107880 -118540
rect 106780 -118590 107560 -118565
rect 107560 -118590 107880 -118565
rect 108280 -118565 109380 -118540
rect 108280 -118590 109060 -118565
rect 109060 -118590 109380 -118565
rect 109780 -118565 110880 -118540
rect 109780 -118590 110560 -118565
rect 110560 -118590 110880 -118565
rect 111280 -118565 112380 -118540
rect 111280 -118590 112060 -118565
rect 112060 -118590 112380 -118565
rect 112780 -118565 113880 -118540
rect 112780 -118590 113560 -118565
rect 113560 -118590 113880 -118565
rect 114280 -118565 115380 -118540
rect 114280 -118590 115060 -118565
rect 115060 -118590 115380 -118565
rect 115780 -118565 116880 -118540
rect 115780 -118590 116560 -118565
rect 116560 -118590 116880 -118565
rect 117280 -118565 118380 -118540
rect 117280 -118590 118060 -118565
rect 118060 -118590 118380 -118565
rect 118780 -118565 119880 -118540
rect 118780 -118590 119560 -118565
rect 119560 -118590 119880 -118565
rect 120 -118850 210 -118750
rect 1620 -118850 1710 -118750
rect 3120 -118850 3210 -118750
rect 4620 -118850 4710 -118750
rect 6120 -118850 6210 -118750
rect 7620 -118850 7710 -118750
rect 9120 -118850 9210 -118750
rect 10620 -118850 10710 -118750
rect 12120 -118850 12210 -118750
rect 13620 -118850 13710 -118750
rect 15120 -118850 15210 -118750
rect 16620 -118850 16710 -118750
rect 18120 -118850 18210 -118750
rect 19620 -118850 19710 -118750
rect 21120 -118850 21210 -118750
rect 22620 -118850 22710 -118750
rect 24120 -118850 24210 -118750
rect 25620 -118850 25710 -118750
rect 27120 -118850 27210 -118750
rect 28620 -118850 28710 -118750
rect 30120 -118850 30210 -118750
rect 31620 -118850 31710 -118750
rect 33120 -118850 33210 -118750
rect 34620 -118850 34710 -118750
rect 36120 -118850 36210 -118750
rect 37620 -118850 37710 -118750
rect 39120 -118850 39210 -118750
rect 40620 -118850 40710 -118750
rect 42120 -118850 42210 -118750
rect 43620 -118850 43710 -118750
rect 45120 -118850 45210 -118750
rect 46620 -118850 46710 -118750
rect 48120 -118850 48210 -118750
rect 49620 -118850 49710 -118750
rect 51120 -118850 51210 -118750
rect 52620 -118850 52710 -118750
rect 54120 -118850 54210 -118750
rect 55620 -118850 55710 -118750
rect 57120 -118850 57210 -118750
rect 58620 -118850 58710 -118750
rect 60120 -118850 60210 -118750
rect 61620 -118850 61710 -118750
rect 63120 -118850 63210 -118750
rect 64620 -118850 64710 -118750
rect 66120 -118850 66210 -118750
rect 67620 -118850 67710 -118750
rect 69120 -118850 69210 -118750
rect 70620 -118850 70710 -118750
rect 72120 -118850 72210 -118750
rect 73620 -118850 73710 -118750
rect 75120 -118850 75210 -118750
rect 76620 -118850 76710 -118750
rect 78120 -118850 78210 -118750
rect 79620 -118850 79710 -118750
rect 81120 -118850 81210 -118750
rect 82620 -118850 82710 -118750
rect 84120 -118850 84210 -118750
rect 85620 -118850 85710 -118750
rect 87120 -118850 87210 -118750
rect 88620 -118850 88710 -118750
rect 90120 -118850 90210 -118750
rect 91620 -118850 91710 -118750
rect 93120 -118850 93210 -118750
rect 94620 -118850 94710 -118750
rect 96120 -118850 96210 -118750
rect 97620 -118850 97710 -118750
rect 99120 -118850 99210 -118750
rect 100620 -118850 100710 -118750
rect 102120 -118850 102210 -118750
rect 103620 -118850 103710 -118750
rect 105120 -118850 105210 -118750
rect 106620 -118850 106710 -118750
rect 108120 -118850 108210 -118750
rect 109620 -118850 109710 -118750
rect 111120 -118850 111210 -118750
rect 112620 -118850 112710 -118750
rect 114120 -118850 114210 -118750
rect 115620 -118850 115710 -118750
rect 117120 -118850 117210 -118750
rect 118620 -118850 118710 -118750
<< metal3 >>
rect -600 1420 -555 2500
rect 240 1825 295 1830
rect 240 1780 245 1825
rect 290 1780 295 1825
rect 240 1775 295 1780
rect 1740 1825 1795 1830
rect 1740 1780 1745 1825
rect 1790 1780 1795 1825
rect 1740 1775 1795 1780
rect 3240 1825 3295 1830
rect 3240 1780 3245 1825
rect 3290 1780 3295 1825
rect 3240 1775 3295 1780
rect 4740 1825 4795 1830
rect 4740 1780 4745 1825
rect 4790 1780 4795 1825
rect 4740 1775 4795 1780
rect 6240 1825 6295 1830
rect 6240 1780 6245 1825
rect 6290 1780 6295 1825
rect 6240 1775 6295 1780
rect 7740 1825 7795 1830
rect 7740 1780 7745 1825
rect 7790 1780 7795 1825
rect 7740 1775 7795 1780
rect 9240 1825 9295 1830
rect 9240 1780 9245 1825
rect 9290 1780 9295 1825
rect 9240 1775 9295 1780
rect 10740 1825 10795 1830
rect 10740 1780 10745 1825
rect 10790 1780 10795 1825
rect 10740 1775 10795 1780
rect 12240 1825 12295 1830
rect 12240 1780 12245 1825
rect 12290 1780 12295 1825
rect 12240 1775 12295 1780
rect 13740 1825 13795 1830
rect 13740 1780 13745 1825
rect 13790 1780 13795 1825
rect 13740 1775 13795 1780
rect 15240 1825 15295 1830
rect 15240 1780 15245 1825
rect 15290 1780 15295 1825
rect 15240 1775 15295 1780
rect 16740 1825 16795 1830
rect 16740 1780 16745 1825
rect 16790 1780 16795 1825
rect 16740 1775 16795 1780
rect 18240 1825 18295 1830
rect 18240 1780 18245 1825
rect 18290 1780 18295 1825
rect 18240 1775 18295 1780
rect 19740 1825 19795 1830
rect 19740 1780 19745 1825
rect 19790 1780 19795 1825
rect 19740 1775 19795 1780
rect 21240 1825 21295 1830
rect 21240 1780 21245 1825
rect 21290 1780 21295 1825
rect 21240 1775 21295 1780
rect 22740 1825 22795 1830
rect 22740 1780 22745 1825
rect 22790 1780 22795 1825
rect 22740 1775 22795 1780
rect 24240 1825 24295 1830
rect 24240 1780 24245 1825
rect 24290 1780 24295 1825
rect 24240 1775 24295 1780
rect 25740 1825 25795 1830
rect 25740 1780 25745 1825
rect 25790 1780 25795 1825
rect 25740 1775 25795 1780
rect 27240 1825 27295 1830
rect 27240 1780 27245 1825
rect 27290 1780 27295 1825
rect 27240 1775 27295 1780
rect 28740 1825 28795 1830
rect 28740 1780 28745 1825
rect 28790 1780 28795 1825
rect 28740 1775 28795 1780
rect 30240 1825 30295 1830
rect 30240 1780 30245 1825
rect 30290 1780 30295 1825
rect 30240 1775 30295 1780
rect 31740 1825 31795 1830
rect 31740 1780 31745 1825
rect 31790 1780 31795 1825
rect 31740 1775 31795 1780
rect 33240 1825 33295 1830
rect 33240 1780 33245 1825
rect 33290 1780 33295 1825
rect 33240 1775 33295 1780
rect 34740 1825 34795 1830
rect 34740 1780 34745 1825
rect 34790 1780 34795 1825
rect 34740 1775 34795 1780
rect 36240 1825 36295 1830
rect 36240 1780 36245 1825
rect 36290 1780 36295 1825
rect 36240 1775 36295 1780
rect 37740 1825 37795 1830
rect 37740 1780 37745 1825
rect 37790 1780 37795 1825
rect 37740 1775 37795 1780
rect 39240 1825 39295 1830
rect 39240 1780 39245 1825
rect 39290 1780 39295 1825
rect 39240 1775 39295 1780
rect 40740 1825 40795 1830
rect 40740 1780 40745 1825
rect 40790 1780 40795 1825
rect 40740 1775 40795 1780
rect 42240 1825 42295 1830
rect 42240 1780 42245 1825
rect 42290 1780 42295 1825
rect 42240 1775 42295 1780
rect 43740 1825 43795 1830
rect 43740 1780 43745 1825
rect 43790 1780 43795 1825
rect 43740 1775 43795 1780
rect 45240 1825 45295 1830
rect 45240 1780 45245 1825
rect 45290 1780 45295 1825
rect 45240 1775 45295 1780
rect 46740 1825 46795 1830
rect 46740 1780 46745 1825
rect 46790 1780 46795 1825
rect 46740 1775 46795 1780
rect 48240 1825 48295 1830
rect 48240 1780 48245 1825
rect 48290 1780 48295 1825
rect 48240 1775 48295 1780
rect 49740 1825 49795 1830
rect 49740 1780 49745 1825
rect 49790 1780 49795 1825
rect 49740 1775 49795 1780
rect 51240 1825 51295 1830
rect 51240 1780 51245 1825
rect 51290 1780 51295 1825
rect 51240 1775 51295 1780
rect 52740 1825 52795 1830
rect 52740 1780 52745 1825
rect 52790 1780 52795 1825
rect 52740 1775 52795 1780
rect 54240 1825 54295 1830
rect 54240 1780 54245 1825
rect 54290 1780 54295 1825
rect 54240 1775 54295 1780
rect 55740 1825 55795 1830
rect 55740 1780 55745 1825
rect 55790 1780 55795 1825
rect 55740 1775 55795 1780
rect 57240 1825 57295 1830
rect 57240 1780 57245 1825
rect 57290 1780 57295 1825
rect 57240 1775 57295 1780
rect 58740 1825 58795 1830
rect 58740 1780 58745 1825
rect 58790 1780 58795 1825
rect 58740 1775 58795 1780
rect 60240 1825 60295 1830
rect 60240 1780 60245 1825
rect 60290 1780 60295 1825
rect 60240 1775 60295 1780
rect 61740 1825 61795 1830
rect 61740 1780 61745 1825
rect 61790 1780 61795 1825
rect 61740 1775 61795 1780
rect 63240 1825 63295 1830
rect 63240 1780 63245 1825
rect 63290 1780 63295 1825
rect 63240 1775 63295 1780
rect 64740 1825 64795 1830
rect 64740 1780 64745 1825
rect 64790 1780 64795 1825
rect 64740 1775 64795 1780
rect 66240 1825 66295 1830
rect 66240 1780 66245 1825
rect 66290 1780 66295 1825
rect 66240 1775 66295 1780
rect 67740 1825 67795 1830
rect 67740 1780 67745 1825
rect 67790 1780 67795 1825
rect 67740 1775 67795 1780
rect 69240 1825 69295 1830
rect 69240 1780 69245 1825
rect 69290 1780 69295 1825
rect 69240 1775 69295 1780
rect 70740 1825 70795 1830
rect 70740 1780 70745 1825
rect 70790 1780 70795 1825
rect 70740 1775 70795 1780
rect 72240 1825 72295 1830
rect 72240 1780 72245 1825
rect 72290 1780 72295 1825
rect 72240 1775 72295 1780
rect 73740 1825 73795 1830
rect 73740 1780 73745 1825
rect 73790 1780 73795 1825
rect 73740 1775 73795 1780
rect 75240 1825 75295 1830
rect 75240 1780 75245 1825
rect 75290 1780 75295 1825
rect 75240 1775 75295 1780
rect 76740 1825 76795 1830
rect 76740 1780 76745 1825
rect 76790 1780 76795 1825
rect 76740 1775 76795 1780
rect 78240 1825 78295 1830
rect 78240 1780 78245 1825
rect 78290 1780 78295 1825
rect 78240 1775 78295 1780
rect 79740 1825 79795 1830
rect 79740 1780 79745 1825
rect 79790 1780 79795 1825
rect 79740 1775 79795 1780
rect 81240 1825 81295 1830
rect 81240 1780 81245 1825
rect 81290 1780 81295 1825
rect 81240 1775 81295 1780
rect 82740 1825 82795 1830
rect 82740 1780 82745 1825
rect 82790 1780 82795 1825
rect 82740 1775 82795 1780
rect 84240 1825 84295 1830
rect 84240 1780 84245 1825
rect 84290 1780 84295 1825
rect 84240 1775 84295 1780
rect 85740 1825 85795 1830
rect 85740 1780 85745 1825
rect 85790 1780 85795 1825
rect 85740 1775 85795 1780
rect 87240 1825 87295 1830
rect 87240 1780 87245 1825
rect 87290 1780 87295 1825
rect 87240 1775 87295 1780
rect 88740 1825 88795 1830
rect 88740 1780 88745 1825
rect 88790 1780 88795 1825
rect 88740 1775 88795 1780
rect 90240 1825 90295 1830
rect 90240 1780 90245 1825
rect 90290 1780 90295 1825
rect 90240 1775 90295 1780
rect 91740 1825 91795 1830
rect 91740 1780 91745 1825
rect 91790 1780 91795 1825
rect 91740 1775 91795 1780
rect 93240 1825 93295 1830
rect 93240 1780 93245 1825
rect 93290 1780 93295 1825
rect 93240 1775 93295 1780
rect 94740 1825 94795 1830
rect 94740 1780 94745 1825
rect 94790 1780 94795 1825
rect 94740 1775 94795 1780
rect 96240 1825 96295 1830
rect 96240 1780 96245 1825
rect 96290 1780 96295 1825
rect 96240 1775 96295 1780
rect 97740 1825 97795 1830
rect 97740 1780 97745 1825
rect 97790 1780 97795 1825
rect 97740 1775 97795 1780
rect 99240 1825 99295 1830
rect 99240 1780 99245 1825
rect 99290 1780 99295 1825
rect 99240 1775 99295 1780
rect 100740 1825 100795 1830
rect 100740 1780 100745 1825
rect 100790 1780 100795 1825
rect 100740 1775 100795 1780
rect 102240 1825 102295 1830
rect 102240 1780 102245 1825
rect 102290 1780 102295 1825
rect 102240 1775 102295 1780
rect 103740 1825 103795 1830
rect 103740 1780 103745 1825
rect 103790 1780 103795 1825
rect 103740 1775 103795 1780
rect 105240 1825 105295 1830
rect 105240 1780 105245 1825
rect 105290 1780 105295 1825
rect 105240 1775 105295 1780
rect 106740 1825 106795 1830
rect 106740 1780 106745 1825
rect 106790 1780 106795 1825
rect 106740 1775 106795 1780
rect 108240 1825 108295 1830
rect 108240 1780 108245 1825
rect 108290 1780 108295 1825
rect 108240 1775 108295 1780
rect 109740 1825 109795 1830
rect 109740 1780 109745 1825
rect 109790 1780 109795 1825
rect 109740 1775 109795 1780
rect 111240 1825 111295 1830
rect 111240 1780 111245 1825
rect 111290 1780 111295 1825
rect 111240 1775 111295 1780
rect 112740 1825 112795 1830
rect 112740 1780 112745 1825
rect 112790 1780 112795 1825
rect 112740 1775 112795 1780
rect 114240 1825 114295 1830
rect 114240 1780 114245 1825
rect 114290 1780 114295 1825
rect 114240 1775 114295 1780
rect 115740 1825 115795 1830
rect 115740 1780 115745 1825
rect 115790 1780 115795 1825
rect 115740 1775 115795 1780
rect 117240 1825 117295 1830
rect 117240 1780 117245 1825
rect 117290 1780 117295 1825
rect 117240 1775 117295 1780
rect 118740 1825 118795 1830
rect 118740 1780 118745 1825
rect 118790 1780 118795 1825
rect 118740 1775 118795 1780
rect -600 1375 100 1420
rect -600 -80 -555 1375
rect -240 1275 -185 1280
rect -240 1270 260 1275
rect -240 1235 -235 1270
rect -190 1235 260 1270
rect -240 1230 260 1235
rect -240 1225 -185 1230
rect -280 780 220 785
rect -280 745 -270 780
rect -130 745 220 780
rect -280 740 220 745
rect -380 115 20 125
rect -380 80 -370 115
rect -325 80 20 115
rect -375 70 -320 80
rect -600 -125 100 -80
rect -600 -1580 -555 -125
rect -240 -225 -185 -220
rect -240 -230 260 -225
rect -240 -265 -235 -230
rect -190 -265 260 -230
rect -240 -270 260 -265
rect -240 -275 -185 -270
rect -280 -720 220 -715
rect -280 -755 -270 -720
rect -130 -755 220 -720
rect -280 -760 220 -755
rect -380 -1385 20 -1375
rect -380 -1420 -370 -1385
rect -325 -1420 20 -1385
rect -375 -1430 -320 -1420
rect -600 -1625 100 -1580
rect -600 -3080 -555 -1625
rect -240 -1725 -185 -1720
rect -240 -1730 260 -1725
rect -240 -1765 -235 -1730
rect -190 -1765 260 -1730
rect -240 -1770 260 -1765
rect -240 -1775 -185 -1770
rect -280 -2220 220 -2215
rect -280 -2255 -270 -2220
rect -130 -2255 220 -2220
rect -280 -2260 220 -2255
rect -380 -2885 20 -2875
rect -380 -2920 -370 -2885
rect -325 -2920 20 -2885
rect -375 -2930 -320 -2920
rect -600 -3125 100 -3080
rect -600 -4580 -555 -3125
rect -240 -3225 -185 -3220
rect -240 -3230 260 -3225
rect -240 -3265 -235 -3230
rect -190 -3265 260 -3230
rect -240 -3270 260 -3265
rect -240 -3275 -185 -3270
rect -280 -3720 220 -3715
rect -280 -3755 -270 -3720
rect -130 -3755 220 -3720
rect -280 -3760 220 -3755
rect -380 -4385 20 -4375
rect -380 -4420 -370 -4385
rect -325 -4420 20 -4385
rect -375 -4430 -320 -4420
rect -600 -4625 100 -4580
rect -600 -6080 -555 -4625
rect -240 -4725 -185 -4720
rect -240 -4730 260 -4725
rect -240 -4765 -235 -4730
rect -190 -4765 260 -4730
rect -240 -4770 260 -4765
rect -240 -4775 -185 -4770
rect -280 -5220 220 -5215
rect -280 -5255 -270 -5220
rect -130 -5255 220 -5220
rect -280 -5260 220 -5255
rect -380 -5885 20 -5875
rect -380 -5920 -370 -5885
rect -325 -5920 20 -5885
rect -375 -5930 -320 -5920
rect -600 -6125 100 -6080
rect -600 -7580 -555 -6125
rect -240 -6225 -185 -6220
rect -240 -6230 260 -6225
rect -240 -6265 -235 -6230
rect -190 -6265 260 -6230
rect -240 -6270 260 -6265
rect -240 -6275 -185 -6270
rect -280 -6720 220 -6715
rect -280 -6755 -270 -6720
rect -130 -6755 220 -6720
rect -280 -6760 220 -6755
rect -380 -7385 20 -7375
rect -380 -7420 -370 -7385
rect -325 -7420 20 -7385
rect -375 -7430 -320 -7420
rect -600 -7625 100 -7580
rect -600 -9080 -555 -7625
rect -240 -7725 -185 -7720
rect -240 -7730 260 -7725
rect -240 -7765 -235 -7730
rect -190 -7765 260 -7730
rect -240 -7770 260 -7765
rect -240 -7775 -185 -7770
rect -280 -8220 220 -8215
rect -280 -8255 -270 -8220
rect -130 -8255 220 -8220
rect -280 -8260 220 -8255
rect -380 -8885 20 -8875
rect -380 -8920 -370 -8885
rect -325 -8920 20 -8885
rect -375 -8930 -320 -8920
rect -600 -9125 100 -9080
rect -600 -10580 -555 -9125
rect -240 -9225 -185 -9220
rect -240 -9230 260 -9225
rect -240 -9265 -235 -9230
rect -190 -9265 260 -9230
rect -240 -9270 260 -9265
rect -240 -9275 -185 -9270
rect -280 -9720 220 -9715
rect -280 -9755 -270 -9720
rect -130 -9755 220 -9720
rect -280 -9760 220 -9755
rect -380 -10385 20 -10375
rect -380 -10420 -370 -10385
rect -325 -10420 20 -10385
rect -375 -10430 -320 -10420
rect -600 -10625 100 -10580
rect -600 -12080 -555 -10625
rect -240 -10725 -185 -10720
rect -240 -10730 260 -10725
rect -240 -10765 -235 -10730
rect -190 -10765 260 -10730
rect -240 -10770 260 -10765
rect -240 -10775 -185 -10770
rect -280 -11220 220 -11215
rect -280 -11255 -270 -11220
rect -130 -11255 220 -11220
rect -280 -11260 220 -11255
rect -380 -11885 20 -11875
rect -380 -11920 -370 -11885
rect -325 -11920 20 -11885
rect -375 -11930 -320 -11920
rect -600 -12125 100 -12080
rect -600 -13580 -555 -12125
rect -240 -12225 -185 -12220
rect -240 -12230 260 -12225
rect -240 -12265 -235 -12230
rect -190 -12265 260 -12230
rect -240 -12270 260 -12265
rect -240 -12275 -185 -12270
rect -280 -12720 220 -12715
rect -280 -12755 -270 -12720
rect -130 -12755 220 -12720
rect -280 -12760 220 -12755
rect -380 -13385 20 -13375
rect -380 -13420 -370 -13385
rect -325 -13420 20 -13385
rect -375 -13430 -320 -13420
rect -600 -13625 100 -13580
rect -600 -15080 -555 -13625
rect -240 -13725 -185 -13720
rect -240 -13730 260 -13725
rect -240 -13765 -235 -13730
rect -190 -13765 260 -13730
rect -240 -13770 260 -13765
rect -240 -13775 -185 -13770
rect -280 -14220 220 -14215
rect -280 -14255 -270 -14220
rect -130 -14255 220 -14220
rect -280 -14260 220 -14255
rect -380 -14885 20 -14875
rect -380 -14920 -370 -14885
rect -325 -14920 20 -14885
rect -375 -14930 -320 -14920
rect -600 -15125 100 -15080
rect -600 -16580 -555 -15125
rect -240 -15225 -185 -15220
rect -240 -15230 260 -15225
rect -240 -15265 -235 -15230
rect -190 -15265 260 -15230
rect -240 -15270 260 -15265
rect -240 -15275 -185 -15270
rect -280 -15720 220 -15715
rect -280 -15755 -270 -15720
rect -130 -15755 220 -15720
rect -280 -15760 220 -15755
rect -380 -16385 20 -16375
rect -380 -16420 -370 -16385
rect -325 -16420 20 -16385
rect -375 -16430 -320 -16420
rect -600 -16625 100 -16580
rect -600 -18080 -555 -16625
rect -240 -16725 -185 -16720
rect -240 -16730 260 -16725
rect -240 -16765 -235 -16730
rect -190 -16765 260 -16730
rect -240 -16770 260 -16765
rect -240 -16775 -185 -16770
rect -280 -17220 220 -17215
rect -280 -17255 -270 -17220
rect -130 -17255 220 -17220
rect -280 -17260 220 -17255
rect -380 -17885 20 -17875
rect -380 -17920 -370 -17885
rect -325 -17920 20 -17885
rect -375 -17930 -320 -17920
rect -600 -18125 100 -18080
rect -600 -19580 -555 -18125
rect -240 -18225 -185 -18220
rect -240 -18230 260 -18225
rect -240 -18265 -235 -18230
rect -190 -18265 260 -18230
rect -240 -18270 260 -18265
rect -240 -18275 -185 -18270
rect -280 -18720 220 -18715
rect -280 -18755 -270 -18720
rect -130 -18755 220 -18720
rect -280 -18760 220 -18755
rect -380 -19385 20 -19375
rect -380 -19420 -370 -19385
rect -325 -19420 20 -19385
rect -375 -19430 -320 -19420
rect -600 -19625 100 -19580
rect -600 -21080 -555 -19625
rect -240 -19725 -185 -19720
rect -240 -19730 260 -19725
rect -240 -19765 -235 -19730
rect -190 -19765 260 -19730
rect -240 -19770 260 -19765
rect -240 -19775 -185 -19770
rect -280 -20220 220 -20215
rect -280 -20255 -270 -20220
rect -130 -20255 220 -20220
rect -280 -20260 220 -20255
rect -380 -20885 20 -20875
rect -380 -20920 -370 -20885
rect -325 -20920 20 -20885
rect -375 -20930 -320 -20920
rect -600 -21125 100 -21080
rect -600 -22580 -555 -21125
rect -240 -21225 -185 -21220
rect -240 -21230 260 -21225
rect -240 -21265 -235 -21230
rect -190 -21265 260 -21230
rect -240 -21270 260 -21265
rect -240 -21275 -185 -21270
rect -280 -21720 220 -21715
rect -280 -21755 -270 -21720
rect -130 -21755 220 -21720
rect -280 -21760 220 -21755
rect -380 -22385 20 -22375
rect -380 -22420 -370 -22385
rect -325 -22420 20 -22385
rect -375 -22430 -320 -22420
rect -600 -22625 100 -22580
rect -600 -24080 -555 -22625
rect -240 -22725 -185 -22720
rect -240 -22730 260 -22725
rect -240 -22765 -235 -22730
rect -190 -22765 260 -22730
rect -240 -22770 260 -22765
rect -240 -22775 -185 -22770
rect -280 -23220 220 -23215
rect -280 -23255 -270 -23220
rect -130 -23255 220 -23220
rect -280 -23260 220 -23255
rect -380 -23885 20 -23875
rect -380 -23920 -370 -23885
rect -325 -23920 20 -23885
rect -375 -23930 -320 -23920
rect -600 -24125 100 -24080
rect -600 -25580 -555 -24125
rect -240 -24225 -185 -24220
rect -240 -24230 260 -24225
rect -240 -24265 -235 -24230
rect -190 -24265 260 -24230
rect -240 -24270 260 -24265
rect -240 -24275 -185 -24270
rect -280 -24720 220 -24715
rect -280 -24755 -270 -24720
rect -130 -24755 220 -24720
rect -280 -24760 220 -24755
rect -380 -25385 20 -25375
rect -380 -25420 -370 -25385
rect -325 -25420 20 -25385
rect -375 -25430 -320 -25420
rect -600 -25625 100 -25580
rect -600 -27080 -555 -25625
rect -240 -25725 -185 -25720
rect -240 -25730 260 -25725
rect -240 -25765 -235 -25730
rect -190 -25765 260 -25730
rect -240 -25770 260 -25765
rect -240 -25775 -185 -25770
rect -280 -26220 220 -26215
rect -280 -26255 -270 -26220
rect -130 -26255 220 -26220
rect -280 -26260 220 -26255
rect -380 -26885 20 -26875
rect -380 -26920 -370 -26885
rect -325 -26920 20 -26885
rect -375 -26930 -320 -26920
rect -600 -27125 100 -27080
rect -600 -28580 -555 -27125
rect -240 -27225 -185 -27220
rect -240 -27230 260 -27225
rect -240 -27265 -235 -27230
rect -190 -27265 260 -27230
rect -240 -27270 260 -27265
rect -240 -27275 -185 -27270
rect -280 -27720 220 -27715
rect -280 -27755 -270 -27720
rect -130 -27755 220 -27720
rect -280 -27760 220 -27755
rect -380 -28385 20 -28375
rect -380 -28420 -370 -28385
rect -325 -28420 20 -28385
rect -375 -28430 -320 -28420
rect -600 -28625 100 -28580
rect -600 -30080 -555 -28625
rect -240 -28725 -185 -28720
rect -240 -28730 260 -28725
rect -240 -28765 -235 -28730
rect -190 -28765 260 -28730
rect -240 -28770 260 -28765
rect -240 -28775 -185 -28770
rect -280 -29220 220 -29215
rect -280 -29255 -270 -29220
rect -130 -29255 220 -29220
rect -280 -29260 220 -29255
rect -380 -29885 20 -29875
rect -380 -29920 -370 -29885
rect -325 -29920 20 -29885
rect -375 -29930 -320 -29920
rect -600 -30125 100 -30080
rect -600 -31580 -555 -30125
rect -240 -30225 -185 -30220
rect -240 -30230 260 -30225
rect -240 -30265 -235 -30230
rect -190 -30265 260 -30230
rect -240 -30270 260 -30265
rect -240 -30275 -185 -30270
rect -280 -30720 220 -30715
rect -280 -30755 -270 -30720
rect -130 -30755 220 -30720
rect -280 -30760 220 -30755
rect -380 -31385 20 -31375
rect -380 -31420 -370 -31385
rect -325 -31420 20 -31385
rect -375 -31430 -320 -31420
rect -600 -31625 100 -31580
rect -600 -33080 -555 -31625
rect -240 -31725 -185 -31720
rect -240 -31730 260 -31725
rect -240 -31765 -235 -31730
rect -190 -31765 260 -31730
rect -240 -31770 260 -31765
rect -240 -31775 -185 -31770
rect -280 -32220 220 -32215
rect -280 -32255 -270 -32220
rect -130 -32255 220 -32220
rect -280 -32260 220 -32255
rect -380 -32885 20 -32875
rect -380 -32920 -370 -32885
rect -325 -32920 20 -32885
rect -375 -32930 -320 -32920
rect -600 -33125 100 -33080
rect -600 -34580 -555 -33125
rect -240 -33225 -185 -33220
rect -240 -33230 260 -33225
rect -240 -33265 -235 -33230
rect -190 -33265 260 -33230
rect -240 -33270 260 -33265
rect -240 -33275 -185 -33270
rect -280 -33720 220 -33715
rect -280 -33755 -270 -33720
rect -130 -33755 220 -33720
rect -280 -33760 220 -33755
rect -380 -34385 20 -34375
rect -380 -34420 -370 -34385
rect -325 -34420 20 -34385
rect -375 -34430 -320 -34420
rect -600 -34625 100 -34580
rect -600 -36080 -555 -34625
rect -240 -34725 -185 -34720
rect -240 -34730 260 -34725
rect -240 -34765 -235 -34730
rect -190 -34765 260 -34730
rect -240 -34770 260 -34765
rect -240 -34775 -185 -34770
rect -280 -35220 220 -35215
rect -280 -35255 -270 -35220
rect -130 -35255 220 -35220
rect -280 -35260 220 -35255
rect -380 -35885 20 -35875
rect -380 -35920 -370 -35885
rect -325 -35920 20 -35885
rect -375 -35930 -320 -35920
rect -600 -36125 100 -36080
rect -600 -37580 -555 -36125
rect -240 -36225 -185 -36220
rect -240 -36230 260 -36225
rect -240 -36265 -235 -36230
rect -190 -36265 260 -36230
rect -240 -36270 260 -36265
rect -240 -36275 -185 -36270
rect -280 -36720 220 -36715
rect -280 -36755 -270 -36720
rect -130 -36755 220 -36720
rect -280 -36760 220 -36755
rect -380 -37385 20 -37375
rect -380 -37420 -370 -37385
rect -325 -37420 20 -37385
rect -375 -37430 -320 -37420
rect -600 -37625 100 -37580
rect -600 -39080 -555 -37625
rect -240 -37725 -185 -37720
rect -240 -37730 260 -37725
rect -240 -37765 -235 -37730
rect -190 -37765 260 -37730
rect -240 -37770 260 -37765
rect -240 -37775 -185 -37770
rect -280 -38220 220 -38215
rect -280 -38255 -270 -38220
rect -130 -38255 220 -38220
rect -280 -38260 220 -38255
rect -380 -38885 20 -38875
rect -380 -38920 -370 -38885
rect -325 -38920 20 -38885
rect -375 -38930 -320 -38920
rect -600 -39125 100 -39080
rect -600 -40580 -555 -39125
rect -240 -39225 -185 -39220
rect -240 -39230 260 -39225
rect -240 -39265 -235 -39230
rect -190 -39265 260 -39230
rect -240 -39270 260 -39265
rect -240 -39275 -185 -39270
rect -280 -39720 220 -39715
rect -280 -39755 -270 -39720
rect -130 -39755 220 -39720
rect -280 -39760 220 -39755
rect -380 -40385 20 -40375
rect -380 -40420 -370 -40385
rect -325 -40420 20 -40385
rect -375 -40430 -320 -40420
rect -600 -40625 100 -40580
rect -600 -42080 -555 -40625
rect -240 -40725 -185 -40720
rect -240 -40730 260 -40725
rect -240 -40765 -235 -40730
rect -190 -40765 260 -40730
rect -240 -40770 260 -40765
rect -240 -40775 -185 -40770
rect -280 -41220 220 -41215
rect -280 -41255 -270 -41220
rect -130 -41255 220 -41220
rect -280 -41260 220 -41255
rect -380 -41885 20 -41875
rect -380 -41920 -370 -41885
rect -325 -41920 20 -41885
rect -375 -41930 -320 -41920
rect -600 -42125 100 -42080
rect -600 -43580 -555 -42125
rect -240 -42225 -185 -42220
rect -240 -42230 260 -42225
rect -240 -42265 -235 -42230
rect -190 -42265 260 -42230
rect -240 -42270 260 -42265
rect -240 -42275 -185 -42270
rect -280 -42720 220 -42715
rect -280 -42755 -270 -42720
rect -130 -42755 220 -42720
rect -280 -42760 220 -42755
rect -380 -43385 20 -43375
rect -380 -43420 -370 -43385
rect -325 -43420 20 -43385
rect -375 -43430 -320 -43420
rect -600 -43625 100 -43580
rect -600 -45080 -555 -43625
rect -240 -43725 -185 -43720
rect -240 -43730 260 -43725
rect -240 -43765 -235 -43730
rect -190 -43765 260 -43730
rect -240 -43770 260 -43765
rect -240 -43775 -185 -43770
rect -280 -44220 220 -44215
rect -280 -44255 -270 -44220
rect -130 -44255 220 -44220
rect -280 -44260 220 -44255
rect -380 -44885 20 -44875
rect -380 -44920 -370 -44885
rect -325 -44920 20 -44885
rect -375 -44930 -320 -44920
rect -600 -45125 100 -45080
rect -600 -46580 -555 -45125
rect -240 -45225 -185 -45220
rect -240 -45230 260 -45225
rect -240 -45265 -235 -45230
rect -190 -45265 260 -45230
rect -240 -45270 260 -45265
rect -240 -45275 -185 -45270
rect -280 -45720 220 -45715
rect -280 -45755 -270 -45720
rect -130 -45755 220 -45720
rect -280 -45760 220 -45755
rect -380 -46385 20 -46375
rect -380 -46420 -370 -46385
rect -325 -46420 20 -46385
rect -375 -46430 -320 -46420
rect -600 -46625 100 -46580
rect -600 -48080 -555 -46625
rect -240 -46725 -185 -46720
rect -240 -46730 260 -46725
rect -240 -46765 -235 -46730
rect -190 -46765 260 -46730
rect -240 -46770 260 -46765
rect -240 -46775 -185 -46770
rect -280 -47220 220 -47215
rect -280 -47255 -270 -47220
rect -130 -47255 220 -47220
rect -280 -47260 220 -47255
rect -380 -47885 20 -47875
rect -380 -47920 -370 -47885
rect -325 -47920 20 -47885
rect -375 -47930 -320 -47920
rect -600 -48125 100 -48080
rect -600 -49580 -555 -48125
rect -240 -48225 -185 -48220
rect -240 -48230 260 -48225
rect -240 -48265 -235 -48230
rect -190 -48265 260 -48230
rect -240 -48270 260 -48265
rect -240 -48275 -185 -48270
rect -280 -48720 220 -48715
rect -280 -48755 -270 -48720
rect -130 -48755 220 -48720
rect -280 -48760 220 -48755
rect -380 -49385 20 -49375
rect -380 -49420 -370 -49385
rect -325 -49420 20 -49385
rect -375 -49430 -320 -49420
rect -600 -49625 100 -49580
rect -600 -51080 -555 -49625
rect -240 -49725 -185 -49720
rect -240 -49730 260 -49725
rect -240 -49765 -235 -49730
rect -190 -49765 260 -49730
rect -240 -49770 260 -49765
rect -240 -49775 -185 -49770
rect -280 -50220 220 -50215
rect -280 -50255 -270 -50220
rect -130 -50255 220 -50220
rect -280 -50260 220 -50255
rect -380 -50885 20 -50875
rect -380 -50920 -370 -50885
rect -325 -50920 20 -50885
rect -375 -50930 -320 -50920
rect -600 -51125 100 -51080
rect -600 -52580 -555 -51125
rect -240 -51225 -185 -51220
rect -240 -51230 260 -51225
rect -240 -51265 -235 -51230
rect -190 -51265 260 -51230
rect -240 -51270 260 -51265
rect -240 -51275 -185 -51270
rect -280 -51720 220 -51715
rect -280 -51755 -270 -51720
rect -130 -51755 220 -51720
rect -280 -51760 220 -51755
rect -380 -52385 20 -52375
rect -380 -52420 -370 -52385
rect -325 -52420 20 -52385
rect -375 -52430 -320 -52420
rect -600 -52625 100 -52580
rect -600 -54080 -555 -52625
rect -240 -52725 -185 -52720
rect -240 -52730 260 -52725
rect -240 -52765 -235 -52730
rect -190 -52765 260 -52730
rect -240 -52770 260 -52765
rect -240 -52775 -185 -52770
rect -280 -53220 220 -53215
rect -280 -53255 -270 -53220
rect -130 -53255 220 -53220
rect -280 -53260 220 -53255
rect -380 -53885 20 -53875
rect -380 -53920 -370 -53885
rect -325 -53920 20 -53885
rect -375 -53930 -320 -53920
rect -600 -54125 100 -54080
rect -600 -55580 -555 -54125
rect -240 -54225 -185 -54220
rect -240 -54230 260 -54225
rect -240 -54265 -235 -54230
rect -190 -54265 260 -54230
rect -240 -54270 260 -54265
rect -240 -54275 -185 -54270
rect -280 -54720 220 -54715
rect -280 -54755 -270 -54720
rect -130 -54755 220 -54720
rect -280 -54760 220 -54755
rect -380 -55385 20 -55375
rect -380 -55420 -370 -55385
rect -325 -55420 20 -55385
rect -375 -55430 -320 -55420
rect -600 -55625 100 -55580
rect -600 -57080 -555 -55625
rect -240 -55725 -185 -55720
rect -240 -55730 260 -55725
rect -240 -55765 -235 -55730
rect -190 -55765 260 -55730
rect -240 -55770 260 -55765
rect -240 -55775 -185 -55770
rect -280 -56220 220 -56215
rect -280 -56255 -270 -56220
rect -130 -56255 220 -56220
rect -280 -56260 220 -56255
rect -380 -56885 20 -56875
rect -380 -56920 -370 -56885
rect -325 -56920 20 -56885
rect -375 -56930 -320 -56920
rect -600 -57125 100 -57080
rect -600 -58580 -555 -57125
rect -240 -57225 -185 -57220
rect -240 -57230 260 -57225
rect -240 -57265 -235 -57230
rect -190 -57265 260 -57230
rect -240 -57270 260 -57265
rect -240 -57275 -185 -57270
rect -280 -57720 220 -57715
rect -280 -57755 -270 -57720
rect -130 -57755 220 -57720
rect -280 -57760 220 -57755
rect -380 -58385 20 -58375
rect -380 -58420 -370 -58385
rect -325 -58420 20 -58385
rect -375 -58430 -320 -58420
rect -600 -58625 100 -58580
rect -600 -60080 -555 -58625
rect -240 -58725 -185 -58720
rect -240 -58730 260 -58725
rect -240 -58765 -235 -58730
rect -190 -58765 260 -58730
rect -240 -58770 260 -58765
rect -240 -58775 -185 -58770
rect -280 -59220 220 -59215
rect -280 -59255 -270 -59220
rect -130 -59255 220 -59220
rect -280 -59260 220 -59255
rect -380 -59885 20 -59875
rect -380 -59920 -370 -59885
rect -325 -59920 20 -59885
rect -375 -59930 -320 -59920
rect -600 -60125 100 -60080
rect -600 -61580 -555 -60125
rect -240 -60225 -185 -60220
rect -240 -60230 260 -60225
rect -240 -60265 -235 -60230
rect -190 -60265 260 -60230
rect -240 -60270 260 -60265
rect -240 -60275 -185 -60270
rect -280 -60720 220 -60715
rect -280 -60755 -270 -60720
rect -130 -60755 220 -60720
rect -280 -60760 220 -60755
rect -380 -61385 20 -61375
rect -380 -61420 -370 -61385
rect -325 -61420 20 -61385
rect -375 -61430 -320 -61420
rect -600 -61625 100 -61580
rect -600 -63080 -555 -61625
rect -240 -61725 -185 -61720
rect -240 -61730 260 -61725
rect -240 -61765 -235 -61730
rect -190 -61765 260 -61730
rect -240 -61770 260 -61765
rect -240 -61775 -185 -61770
rect -280 -62220 220 -62215
rect -280 -62255 -270 -62220
rect -130 -62255 220 -62220
rect -280 -62260 220 -62255
rect -380 -62885 20 -62875
rect -380 -62920 -370 -62885
rect -325 -62920 20 -62885
rect -375 -62930 -320 -62920
rect -600 -63125 100 -63080
rect -600 -64580 -555 -63125
rect -240 -63225 -185 -63220
rect -240 -63230 260 -63225
rect -240 -63265 -235 -63230
rect -190 -63265 260 -63230
rect -240 -63270 260 -63265
rect -240 -63275 -185 -63270
rect -280 -63720 220 -63715
rect -280 -63755 -270 -63720
rect -130 -63755 220 -63720
rect -280 -63760 220 -63755
rect -380 -64385 20 -64375
rect -380 -64420 -370 -64385
rect -325 -64420 20 -64385
rect -375 -64430 -320 -64420
rect -600 -64625 100 -64580
rect -600 -66080 -555 -64625
rect -240 -64725 -185 -64720
rect -240 -64730 260 -64725
rect -240 -64765 -235 -64730
rect -190 -64765 260 -64730
rect -240 -64770 260 -64765
rect -240 -64775 -185 -64770
rect -280 -65220 220 -65215
rect -280 -65255 -270 -65220
rect -130 -65255 220 -65220
rect -280 -65260 220 -65255
rect -380 -65885 20 -65875
rect -380 -65920 -370 -65885
rect -325 -65920 20 -65885
rect -375 -65930 -320 -65920
rect -600 -66125 100 -66080
rect -600 -67580 -555 -66125
rect -240 -66225 -185 -66220
rect -240 -66230 260 -66225
rect -240 -66265 -235 -66230
rect -190 -66265 260 -66230
rect -240 -66270 260 -66265
rect -240 -66275 -185 -66270
rect -280 -66720 220 -66715
rect -280 -66755 -270 -66720
rect -130 -66755 220 -66720
rect -280 -66760 220 -66755
rect -380 -67385 20 -67375
rect -380 -67420 -370 -67385
rect -325 -67420 20 -67385
rect -375 -67430 -320 -67420
rect -600 -67625 100 -67580
rect -600 -69080 -555 -67625
rect -240 -67725 -185 -67720
rect -240 -67730 260 -67725
rect -240 -67765 -235 -67730
rect -190 -67765 260 -67730
rect -240 -67770 260 -67765
rect -240 -67775 -185 -67770
rect -280 -68220 220 -68215
rect -280 -68255 -270 -68220
rect -130 -68255 220 -68220
rect -280 -68260 220 -68255
rect -380 -68885 20 -68875
rect -380 -68920 -370 -68885
rect -325 -68920 20 -68885
rect -375 -68930 -320 -68920
rect -600 -69125 100 -69080
rect -600 -70580 -555 -69125
rect -240 -69225 -185 -69220
rect -240 -69230 260 -69225
rect -240 -69265 -235 -69230
rect -190 -69265 260 -69230
rect -240 -69270 260 -69265
rect -240 -69275 -185 -69270
rect -280 -69720 220 -69715
rect -280 -69755 -270 -69720
rect -130 -69755 220 -69720
rect -280 -69760 220 -69755
rect -380 -70385 20 -70375
rect -380 -70420 -370 -70385
rect -325 -70420 20 -70385
rect -375 -70430 -320 -70420
rect -600 -70625 100 -70580
rect -600 -72080 -555 -70625
rect -240 -70725 -185 -70720
rect -240 -70730 260 -70725
rect -240 -70765 -235 -70730
rect -190 -70765 260 -70730
rect -240 -70770 260 -70765
rect -240 -70775 -185 -70770
rect -280 -71220 220 -71215
rect -280 -71255 -270 -71220
rect -130 -71255 220 -71220
rect -280 -71260 220 -71255
rect -380 -71885 20 -71875
rect -380 -71920 -370 -71885
rect -325 -71920 20 -71885
rect -375 -71930 -320 -71920
rect -600 -72125 100 -72080
rect -600 -73580 -555 -72125
rect -240 -72225 -185 -72220
rect -240 -72230 260 -72225
rect -240 -72265 -235 -72230
rect -190 -72265 260 -72230
rect -240 -72270 260 -72265
rect -240 -72275 -185 -72270
rect -280 -72720 220 -72715
rect -280 -72755 -270 -72720
rect -130 -72755 220 -72720
rect -280 -72760 220 -72755
rect -380 -73385 20 -73375
rect -380 -73420 -370 -73385
rect -325 -73420 20 -73385
rect -375 -73430 -320 -73420
rect -600 -73625 100 -73580
rect -600 -75080 -555 -73625
rect -240 -73725 -185 -73720
rect -240 -73730 260 -73725
rect -240 -73765 -235 -73730
rect -190 -73765 260 -73730
rect -240 -73770 260 -73765
rect -240 -73775 -185 -73770
rect -280 -74220 220 -74215
rect -280 -74255 -270 -74220
rect -130 -74255 220 -74220
rect -280 -74260 220 -74255
rect -380 -74885 20 -74875
rect -380 -74920 -370 -74885
rect -325 -74920 20 -74885
rect -375 -74930 -320 -74920
rect -600 -75125 100 -75080
rect -600 -76580 -555 -75125
rect -240 -75225 -185 -75220
rect -240 -75230 260 -75225
rect -240 -75265 -235 -75230
rect -190 -75265 260 -75230
rect -240 -75270 260 -75265
rect -240 -75275 -185 -75270
rect -280 -75720 220 -75715
rect -280 -75755 -270 -75720
rect -130 -75755 220 -75720
rect -280 -75760 220 -75755
rect -380 -76385 20 -76375
rect -380 -76420 -370 -76385
rect -325 -76420 20 -76385
rect -375 -76430 -320 -76420
rect -600 -76625 100 -76580
rect -600 -78080 -555 -76625
rect -240 -76725 -185 -76720
rect -240 -76730 260 -76725
rect -240 -76765 -235 -76730
rect -190 -76765 260 -76730
rect -240 -76770 260 -76765
rect -240 -76775 -185 -76770
rect -280 -77220 220 -77215
rect -280 -77255 -270 -77220
rect -130 -77255 220 -77220
rect -280 -77260 220 -77255
rect -380 -77885 20 -77875
rect -380 -77920 -370 -77885
rect -325 -77920 20 -77885
rect -375 -77930 -320 -77920
rect -600 -78125 100 -78080
rect -600 -79580 -555 -78125
rect -240 -78225 -185 -78220
rect -240 -78230 260 -78225
rect -240 -78265 -235 -78230
rect -190 -78265 260 -78230
rect -240 -78270 260 -78265
rect -240 -78275 -185 -78270
rect -280 -78720 220 -78715
rect -280 -78755 -270 -78720
rect -130 -78755 220 -78720
rect -280 -78760 220 -78755
rect -380 -79385 20 -79375
rect -380 -79420 -370 -79385
rect -325 -79420 20 -79385
rect -375 -79430 -320 -79420
rect -600 -79625 100 -79580
rect -600 -81080 -555 -79625
rect -240 -79725 -185 -79720
rect -240 -79730 260 -79725
rect -240 -79765 -235 -79730
rect -190 -79765 260 -79730
rect -240 -79770 260 -79765
rect -240 -79775 -185 -79770
rect -280 -80220 220 -80215
rect -280 -80255 -270 -80220
rect -130 -80255 220 -80220
rect -280 -80260 220 -80255
rect -380 -80885 20 -80875
rect -380 -80920 -370 -80885
rect -325 -80920 20 -80885
rect -375 -80930 -320 -80920
rect -600 -81125 100 -81080
rect -600 -82580 -555 -81125
rect -240 -81225 -185 -81220
rect -240 -81230 260 -81225
rect -240 -81265 -235 -81230
rect -190 -81265 260 -81230
rect -240 -81270 260 -81265
rect -240 -81275 -185 -81270
rect -280 -81720 220 -81715
rect -280 -81755 -270 -81720
rect -130 -81755 220 -81720
rect -280 -81760 220 -81755
rect -380 -82385 20 -82375
rect -380 -82420 -370 -82385
rect -325 -82420 20 -82385
rect -375 -82430 -320 -82420
rect -600 -82625 100 -82580
rect -600 -84080 -555 -82625
rect -240 -82725 -185 -82720
rect -240 -82730 260 -82725
rect -240 -82765 -235 -82730
rect -190 -82765 260 -82730
rect -240 -82770 260 -82765
rect -240 -82775 -185 -82770
rect -280 -83220 220 -83215
rect -280 -83255 -270 -83220
rect -130 -83255 220 -83220
rect -280 -83260 220 -83255
rect -380 -83885 20 -83875
rect -380 -83920 -370 -83885
rect -325 -83920 20 -83885
rect -375 -83930 -320 -83920
rect -600 -84125 100 -84080
rect -600 -85580 -555 -84125
rect -240 -84225 -185 -84220
rect -240 -84230 260 -84225
rect -240 -84265 -235 -84230
rect -190 -84265 260 -84230
rect -240 -84270 260 -84265
rect -240 -84275 -185 -84270
rect -280 -84720 220 -84715
rect -280 -84755 -270 -84720
rect -130 -84755 220 -84720
rect -280 -84760 220 -84755
rect -380 -85385 20 -85375
rect -380 -85420 -370 -85385
rect -325 -85420 20 -85385
rect -375 -85430 -320 -85420
rect -600 -85625 100 -85580
rect -600 -87080 -555 -85625
rect -240 -85725 -185 -85720
rect -240 -85730 260 -85725
rect -240 -85765 -235 -85730
rect -190 -85765 260 -85730
rect -240 -85770 260 -85765
rect -240 -85775 -185 -85770
rect -280 -86220 220 -86215
rect -280 -86255 -270 -86220
rect -130 -86255 220 -86220
rect -280 -86260 220 -86255
rect -380 -86885 20 -86875
rect -380 -86920 -370 -86885
rect -325 -86920 20 -86885
rect -375 -86930 -320 -86920
rect -600 -87125 100 -87080
rect -600 -88580 -555 -87125
rect -240 -87225 -185 -87220
rect -240 -87230 260 -87225
rect -240 -87265 -235 -87230
rect -190 -87265 260 -87230
rect -240 -87270 260 -87265
rect -240 -87275 -185 -87270
rect -280 -87720 220 -87715
rect -280 -87755 -270 -87720
rect -130 -87755 220 -87720
rect -280 -87760 220 -87755
rect -380 -88385 20 -88375
rect -380 -88420 -370 -88385
rect -325 -88420 20 -88385
rect -375 -88430 -320 -88420
rect -600 -88625 100 -88580
rect -600 -90080 -555 -88625
rect -240 -88725 -185 -88720
rect -240 -88730 260 -88725
rect -240 -88765 -235 -88730
rect -190 -88765 260 -88730
rect -240 -88770 260 -88765
rect -240 -88775 -185 -88770
rect -280 -89220 220 -89215
rect -280 -89255 -270 -89220
rect -130 -89255 220 -89220
rect -280 -89260 220 -89255
rect -380 -89885 20 -89875
rect -380 -89920 -370 -89885
rect -325 -89920 20 -89885
rect -375 -89930 -320 -89920
rect -600 -90125 100 -90080
rect -600 -91580 -555 -90125
rect -240 -90225 -185 -90220
rect -240 -90230 260 -90225
rect -240 -90265 -235 -90230
rect -190 -90265 260 -90230
rect -240 -90270 260 -90265
rect -240 -90275 -185 -90270
rect -280 -90720 220 -90715
rect -280 -90755 -270 -90720
rect -130 -90755 220 -90720
rect -280 -90760 220 -90755
rect -380 -91385 20 -91375
rect -380 -91420 -370 -91385
rect -325 -91420 20 -91385
rect -375 -91430 -320 -91420
rect -600 -91625 100 -91580
rect -600 -93080 -555 -91625
rect -240 -91725 -185 -91720
rect -240 -91730 260 -91725
rect -240 -91765 -235 -91730
rect -190 -91765 260 -91730
rect -240 -91770 260 -91765
rect -240 -91775 -185 -91770
rect -280 -92220 220 -92215
rect -280 -92255 -270 -92220
rect -130 -92255 220 -92220
rect -280 -92260 220 -92255
rect -380 -92885 20 -92875
rect -380 -92920 -370 -92885
rect -325 -92920 20 -92885
rect -375 -92930 -320 -92920
rect -600 -93125 100 -93080
rect -600 -94580 -555 -93125
rect -240 -93225 -185 -93220
rect -240 -93230 260 -93225
rect -240 -93265 -235 -93230
rect -190 -93265 260 -93230
rect -240 -93270 260 -93265
rect -240 -93275 -185 -93270
rect -280 -93720 220 -93715
rect -280 -93755 -270 -93720
rect -130 -93755 220 -93720
rect -280 -93760 220 -93755
rect -380 -94385 20 -94375
rect -380 -94420 -370 -94385
rect -325 -94420 20 -94385
rect -375 -94430 -320 -94420
rect -600 -94625 100 -94580
rect -600 -96080 -555 -94625
rect -240 -94725 -185 -94720
rect -240 -94730 260 -94725
rect -240 -94765 -235 -94730
rect -190 -94765 260 -94730
rect -240 -94770 260 -94765
rect -240 -94775 -185 -94770
rect -280 -95220 220 -95215
rect -280 -95255 -270 -95220
rect -130 -95255 220 -95220
rect -280 -95260 220 -95255
rect -380 -95885 20 -95875
rect -380 -95920 -370 -95885
rect -325 -95920 20 -95885
rect -375 -95930 -320 -95920
rect -600 -96125 100 -96080
rect -600 -97580 -555 -96125
rect -240 -96225 -185 -96220
rect -240 -96230 260 -96225
rect -240 -96265 -235 -96230
rect -190 -96265 260 -96230
rect -240 -96270 260 -96265
rect -240 -96275 -185 -96270
rect -280 -96720 220 -96715
rect -280 -96755 -270 -96720
rect -130 -96755 220 -96720
rect -280 -96760 220 -96755
rect -380 -97385 20 -97375
rect -380 -97420 -370 -97385
rect -325 -97420 20 -97385
rect -375 -97430 -320 -97420
rect -600 -97625 100 -97580
rect -600 -99080 -555 -97625
rect -240 -97725 -185 -97720
rect -240 -97730 260 -97725
rect -240 -97765 -235 -97730
rect -190 -97765 260 -97730
rect -240 -97770 260 -97765
rect -240 -97775 -185 -97770
rect -280 -98220 220 -98215
rect -280 -98255 -270 -98220
rect -130 -98255 220 -98220
rect -280 -98260 220 -98255
rect -380 -98885 20 -98875
rect -380 -98920 -370 -98885
rect -325 -98920 20 -98885
rect -375 -98930 -320 -98920
rect -600 -99125 100 -99080
rect -600 -100580 -555 -99125
rect -240 -99225 -185 -99220
rect -240 -99230 260 -99225
rect -240 -99265 -235 -99230
rect -190 -99265 260 -99230
rect -240 -99270 260 -99265
rect -240 -99275 -185 -99270
rect -280 -99720 220 -99715
rect -280 -99755 -270 -99720
rect -130 -99755 220 -99720
rect -280 -99760 220 -99755
rect -380 -100385 20 -100375
rect -380 -100420 -370 -100385
rect -325 -100420 20 -100385
rect -375 -100430 -320 -100420
rect -600 -100625 100 -100580
rect -600 -102080 -555 -100625
rect -240 -100725 -185 -100720
rect -240 -100730 260 -100725
rect -240 -100765 -235 -100730
rect -190 -100765 260 -100730
rect -240 -100770 260 -100765
rect -240 -100775 -185 -100770
rect -280 -101220 220 -101215
rect -280 -101255 -270 -101220
rect -130 -101255 220 -101220
rect -280 -101260 220 -101255
rect -380 -101885 20 -101875
rect -380 -101920 -370 -101885
rect -325 -101920 20 -101885
rect -375 -101930 -320 -101920
rect -600 -102125 100 -102080
rect -600 -103580 -555 -102125
rect -240 -102225 -185 -102220
rect -240 -102230 260 -102225
rect -240 -102265 -235 -102230
rect -190 -102265 260 -102230
rect -240 -102270 260 -102265
rect -240 -102275 -185 -102270
rect -280 -102720 220 -102715
rect -280 -102755 -270 -102720
rect -130 -102755 220 -102720
rect -280 -102760 220 -102755
rect -380 -103385 20 -103375
rect -380 -103420 -370 -103385
rect -325 -103420 20 -103385
rect -375 -103430 -320 -103420
rect -600 -103625 100 -103580
rect -600 -105080 -555 -103625
rect -240 -103725 -185 -103720
rect -240 -103730 260 -103725
rect -240 -103765 -235 -103730
rect -190 -103765 260 -103730
rect -240 -103770 260 -103765
rect -240 -103775 -185 -103770
rect -280 -104220 220 -104215
rect -280 -104255 -270 -104220
rect -130 -104255 220 -104220
rect -280 -104260 220 -104255
rect -380 -104885 20 -104875
rect -380 -104920 -370 -104885
rect -325 -104920 20 -104885
rect -375 -104930 -320 -104920
rect -600 -105125 100 -105080
rect -600 -106580 -555 -105125
rect -240 -105225 -185 -105220
rect -240 -105230 260 -105225
rect -240 -105265 -235 -105230
rect -190 -105265 260 -105230
rect -240 -105270 260 -105265
rect -240 -105275 -185 -105270
rect -280 -105720 220 -105715
rect -280 -105755 -270 -105720
rect -130 -105755 220 -105720
rect -280 -105760 220 -105755
rect -380 -106385 20 -106375
rect -380 -106420 -370 -106385
rect -325 -106420 20 -106385
rect -375 -106430 -320 -106420
rect -600 -106625 100 -106580
rect -600 -108080 -555 -106625
rect -240 -106725 -185 -106720
rect -240 -106730 260 -106725
rect -240 -106765 -235 -106730
rect -190 -106765 260 -106730
rect -240 -106770 260 -106765
rect -240 -106775 -185 -106770
rect -280 -107220 220 -107215
rect -280 -107255 -270 -107220
rect -130 -107255 220 -107220
rect -280 -107260 220 -107255
rect -380 -107885 20 -107875
rect -380 -107920 -370 -107885
rect -325 -107920 20 -107885
rect -375 -107930 -320 -107920
rect -600 -108125 100 -108080
rect -600 -109580 -555 -108125
rect -240 -108225 -185 -108220
rect -240 -108230 260 -108225
rect -240 -108265 -235 -108230
rect -190 -108265 260 -108230
rect -240 -108270 260 -108265
rect -240 -108275 -185 -108270
rect -280 -108720 220 -108715
rect -280 -108755 -270 -108720
rect -130 -108755 220 -108720
rect -280 -108760 220 -108755
rect -380 -109385 20 -109375
rect -380 -109420 -370 -109385
rect -325 -109420 20 -109385
rect -375 -109430 -320 -109420
rect -600 -109625 100 -109580
rect -600 -111080 -555 -109625
rect -240 -109725 -185 -109720
rect -240 -109730 260 -109725
rect -240 -109765 -235 -109730
rect -190 -109765 260 -109730
rect -240 -109770 260 -109765
rect -240 -109775 -185 -109770
rect -280 -110220 220 -110215
rect -280 -110255 -270 -110220
rect -130 -110255 220 -110220
rect -280 -110260 220 -110255
rect -380 -110885 20 -110875
rect -380 -110920 -370 -110885
rect -325 -110920 20 -110885
rect -375 -110930 -320 -110920
rect -600 -111125 100 -111080
rect -600 -112580 -555 -111125
rect -240 -111225 -185 -111220
rect -240 -111230 260 -111225
rect -240 -111265 -235 -111230
rect -190 -111265 260 -111230
rect -240 -111270 260 -111265
rect -240 -111275 -185 -111270
rect -280 -111720 220 -111715
rect -280 -111755 -270 -111720
rect -130 -111755 220 -111720
rect -280 -111760 220 -111755
rect -380 -112385 20 -112375
rect -380 -112420 -370 -112385
rect -325 -112420 20 -112385
rect -375 -112430 -320 -112420
rect -600 -112625 100 -112580
rect -600 -114080 -555 -112625
rect -240 -112725 -185 -112720
rect -240 -112730 260 -112725
rect -240 -112765 -235 -112730
rect -190 -112765 260 -112730
rect -240 -112770 260 -112765
rect -240 -112775 -185 -112770
rect -280 -113220 220 -113215
rect -280 -113255 -270 -113220
rect -130 -113255 220 -113220
rect -280 -113260 220 -113255
rect -380 -113885 20 -113875
rect -380 -113920 -370 -113885
rect -325 -113920 20 -113885
rect -375 -113930 -320 -113920
rect -600 -114125 100 -114080
rect -600 -115580 -555 -114125
rect -240 -114225 -185 -114220
rect -240 -114230 260 -114225
rect -240 -114265 -235 -114230
rect -190 -114265 260 -114230
rect -240 -114270 260 -114265
rect -240 -114275 -185 -114270
rect -280 -114720 220 -114715
rect -280 -114755 -270 -114720
rect -130 -114755 220 -114720
rect -280 -114760 220 -114755
rect -380 -115385 20 -115375
rect -380 -115420 -370 -115385
rect -325 -115420 20 -115385
rect -375 -115430 -320 -115420
rect -600 -115625 100 -115580
rect -600 -117080 -555 -115625
rect -240 -115725 -185 -115720
rect -240 -115730 260 -115725
rect -240 -115765 -235 -115730
rect -190 -115765 260 -115730
rect -240 -115770 260 -115765
rect -240 -115775 -185 -115770
rect -280 -116220 220 -116215
rect -280 -116255 -270 -116220
rect -130 -116255 220 -116220
rect -280 -116260 220 -116255
rect -380 -116885 20 -116875
rect -380 -116920 -370 -116885
rect -325 -116920 20 -116885
rect -375 -116930 -320 -116920
rect -600 -117125 100 -117080
rect -600 -117500 -555 -117125
rect -240 -117225 -185 -117220
rect -240 -117230 260 -117225
rect -240 -117265 -235 -117230
rect -190 -117265 260 -117230
rect -240 -117270 260 -117265
rect -240 -117275 -185 -117270
rect -280 -117720 220 -117715
rect -280 -117755 -270 -117720
rect -130 -117755 220 -117720
rect -280 -117760 220 -117755
rect -380 -118385 20 -118375
rect -380 -118420 -370 -118385
rect -325 -118420 20 -118385
rect -375 -118430 -320 -118420
rect 270 -118540 1390 -118530
rect 270 -118590 280 -118540
rect 1380 -118590 1390 -118540
rect 270 -118600 1390 -118590
rect 1770 -118540 2890 -118530
rect 1770 -118590 1780 -118540
rect 2880 -118590 2890 -118540
rect 1770 -118600 2890 -118590
rect 3270 -118540 4390 -118530
rect 3270 -118590 3280 -118540
rect 4380 -118590 4390 -118540
rect 3270 -118600 4390 -118590
rect 4770 -118540 5890 -118530
rect 4770 -118590 4780 -118540
rect 5880 -118590 5890 -118540
rect 4770 -118600 5890 -118590
rect 6270 -118540 7390 -118530
rect 6270 -118590 6280 -118540
rect 7380 -118590 7390 -118540
rect 6270 -118600 7390 -118590
rect 7770 -118540 8890 -118530
rect 7770 -118590 7780 -118540
rect 8880 -118590 8890 -118540
rect 7770 -118600 8890 -118590
rect 9270 -118540 10390 -118530
rect 9270 -118590 9280 -118540
rect 10380 -118590 10390 -118540
rect 9270 -118600 10390 -118590
rect 10770 -118540 11890 -118530
rect 10770 -118590 10780 -118540
rect 11880 -118590 11890 -118540
rect 10770 -118600 11890 -118590
rect 12270 -118540 13390 -118530
rect 12270 -118590 12280 -118540
rect 13380 -118590 13390 -118540
rect 12270 -118600 13390 -118590
rect 13770 -118540 14890 -118530
rect 13770 -118590 13780 -118540
rect 14880 -118590 14890 -118540
rect 13770 -118600 14890 -118590
rect 15270 -118540 16390 -118530
rect 15270 -118590 15280 -118540
rect 16380 -118590 16390 -118540
rect 15270 -118600 16390 -118590
rect 16770 -118540 17890 -118530
rect 16770 -118590 16780 -118540
rect 17880 -118590 17890 -118540
rect 16770 -118600 17890 -118590
rect 18270 -118540 19390 -118530
rect 18270 -118590 18280 -118540
rect 19380 -118590 19390 -118540
rect 18270 -118600 19390 -118590
rect 19770 -118540 20890 -118530
rect 19770 -118590 19780 -118540
rect 20880 -118590 20890 -118540
rect 19770 -118600 20890 -118590
rect 21270 -118540 22390 -118530
rect 21270 -118590 21280 -118540
rect 22380 -118590 22390 -118540
rect 21270 -118600 22390 -118590
rect 22770 -118540 23890 -118530
rect 22770 -118590 22780 -118540
rect 23880 -118590 23890 -118540
rect 22770 -118600 23890 -118590
rect 24270 -118540 25390 -118530
rect 24270 -118590 24280 -118540
rect 25380 -118590 25390 -118540
rect 24270 -118600 25390 -118590
rect 25770 -118540 26890 -118530
rect 25770 -118590 25780 -118540
rect 26880 -118590 26890 -118540
rect 25770 -118600 26890 -118590
rect 27270 -118540 28390 -118530
rect 27270 -118590 27280 -118540
rect 28380 -118590 28390 -118540
rect 27270 -118600 28390 -118590
rect 28770 -118540 29890 -118530
rect 28770 -118590 28780 -118540
rect 29880 -118590 29890 -118540
rect 28770 -118600 29890 -118590
rect 30270 -118540 31390 -118530
rect 30270 -118590 30280 -118540
rect 31380 -118590 31390 -118540
rect 30270 -118600 31390 -118590
rect 31770 -118540 32890 -118530
rect 31770 -118590 31780 -118540
rect 32880 -118590 32890 -118540
rect 31770 -118600 32890 -118590
rect 33270 -118540 34390 -118530
rect 33270 -118590 33280 -118540
rect 34380 -118590 34390 -118540
rect 33270 -118600 34390 -118590
rect 34770 -118540 35890 -118530
rect 34770 -118590 34780 -118540
rect 35880 -118590 35890 -118540
rect 34770 -118600 35890 -118590
rect 36270 -118540 37390 -118530
rect 36270 -118590 36280 -118540
rect 37380 -118590 37390 -118540
rect 36270 -118600 37390 -118590
rect 37770 -118540 38890 -118530
rect 37770 -118590 37780 -118540
rect 38880 -118590 38890 -118540
rect 37770 -118600 38890 -118590
rect 39270 -118540 40390 -118530
rect 39270 -118590 39280 -118540
rect 40380 -118590 40390 -118540
rect 39270 -118600 40390 -118590
rect 40770 -118540 41890 -118530
rect 40770 -118590 40780 -118540
rect 41880 -118590 41890 -118540
rect 40770 -118600 41890 -118590
rect 42270 -118540 43390 -118530
rect 42270 -118590 42280 -118540
rect 43380 -118590 43390 -118540
rect 42270 -118600 43390 -118590
rect 43770 -118540 44890 -118530
rect 43770 -118590 43780 -118540
rect 44880 -118590 44890 -118540
rect 43770 -118600 44890 -118590
rect 45270 -118540 46390 -118530
rect 45270 -118590 45280 -118540
rect 46380 -118590 46390 -118540
rect 45270 -118600 46390 -118590
rect 46770 -118540 47890 -118530
rect 46770 -118590 46780 -118540
rect 47880 -118590 47890 -118540
rect 46770 -118600 47890 -118590
rect 48270 -118540 49390 -118530
rect 48270 -118590 48280 -118540
rect 49380 -118590 49390 -118540
rect 48270 -118600 49390 -118590
rect 49770 -118540 50890 -118530
rect 49770 -118590 49780 -118540
rect 50880 -118590 50890 -118540
rect 49770 -118600 50890 -118590
rect 51270 -118540 52390 -118530
rect 51270 -118590 51280 -118540
rect 52380 -118590 52390 -118540
rect 51270 -118600 52390 -118590
rect 52770 -118540 53890 -118530
rect 52770 -118590 52780 -118540
rect 53880 -118590 53890 -118540
rect 52770 -118600 53890 -118590
rect 54270 -118540 55390 -118530
rect 54270 -118590 54280 -118540
rect 55380 -118590 55390 -118540
rect 54270 -118600 55390 -118590
rect 55770 -118540 56890 -118530
rect 55770 -118590 55780 -118540
rect 56880 -118590 56890 -118540
rect 55770 -118600 56890 -118590
rect 57270 -118540 58390 -118530
rect 57270 -118590 57280 -118540
rect 58380 -118590 58390 -118540
rect 57270 -118600 58390 -118590
rect 58770 -118540 59890 -118530
rect 58770 -118590 58780 -118540
rect 59880 -118590 59890 -118540
rect 58770 -118600 59890 -118590
rect 60270 -118540 61390 -118530
rect 60270 -118590 60280 -118540
rect 61380 -118590 61390 -118540
rect 60270 -118600 61390 -118590
rect 61770 -118540 62890 -118530
rect 61770 -118590 61780 -118540
rect 62880 -118590 62890 -118540
rect 61770 -118600 62890 -118590
rect 63270 -118540 64390 -118530
rect 63270 -118590 63280 -118540
rect 64380 -118590 64390 -118540
rect 63270 -118600 64390 -118590
rect 64770 -118540 65890 -118530
rect 64770 -118590 64780 -118540
rect 65880 -118590 65890 -118540
rect 64770 -118600 65890 -118590
rect 66270 -118540 67390 -118530
rect 66270 -118590 66280 -118540
rect 67380 -118590 67390 -118540
rect 66270 -118600 67390 -118590
rect 67770 -118540 68890 -118530
rect 67770 -118590 67780 -118540
rect 68880 -118590 68890 -118540
rect 67770 -118600 68890 -118590
rect 69270 -118540 70390 -118530
rect 69270 -118590 69280 -118540
rect 70380 -118590 70390 -118540
rect 69270 -118600 70390 -118590
rect 70770 -118540 71890 -118530
rect 70770 -118590 70780 -118540
rect 71880 -118590 71890 -118540
rect 70770 -118600 71890 -118590
rect 72270 -118540 73390 -118530
rect 72270 -118590 72280 -118540
rect 73380 -118590 73390 -118540
rect 72270 -118600 73390 -118590
rect 73770 -118540 74890 -118530
rect 73770 -118590 73780 -118540
rect 74880 -118590 74890 -118540
rect 73770 -118600 74890 -118590
rect 75270 -118540 76390 -118530
rect 75270 -118590 75280 -118540
rect 76380 -118590 76390 -118540
rect 75270 -118600 76390 -118590
rect 76770 -118540 77890 -118530
rect 76770 -118590 76780 -118540
rect 77880 -118590 77890 -118540
rect 76770 -118600 77890 -118590
rect 78270 -118540 79390 -118530
rect 78270 -118590 78280 -118540
rect 79380 -118590 79390 -118540
rect 78270 -118600 79390 -118590
rect 79770 -118540 80890 -118530
rect 79770 -118590 79780 -118540
rect 80880 -118590 80890 -118540
rect 79770 -118600 80890 -118590
rect 81270 -118540 82390 -118530
rect 81270 -118590 81280 -118540
rect 82380 -118590 82390 -118540
rect 81270 -118600 82390 -118590
rect 82770 -118540 83890 -118530
rect 82770 -118590 82780 -118540
rect 83880 -118590 83890 -118540
rect 82770 -118600 83890 -118590
rect 84270 -118540 85390 -118530
rect 84270 -118590 84280 -118540
rect 85380 -118590 85390 -118540
rect 84270 -118600 85390 -118590
rect 85770 -118540 86890 -118530
rect 85770 -118590 85780 -118540
rect 86880 -118590 86890 -118540
rect 85770 -118600 86890 -118590
rect 87270 -118540 88390 -118530
rect 87270 -118590 87280 -118540
rect 88380 -118590 88390 -118540
rect 87270 -118600 88390 -118590
rect 88770 -118540 89890 -118530
rect 88770 -118590 88780 -118540
rect 89880 -118590 89890 -118540
rect 88770 -118600 89890 -118590
rect 90270 -118540 91390 -118530
rect 90270 -118590 90280 -118540
rect 91380 -118590 91390 -118540
rect 90270 -118600 91390 -118590
rect 91770 -118540 92890 -118530
rect 91770 -118590 91780 -118540
rect 92880 -118590 92890 -118540
rect 91770 -118600 92890 -118590
rect 93270 -118540 94390 -118530
rect 93270 -118590 93280 -118540
rect 94380 -118590 94390 -118540
rect 93270 -118600 94390 -118590
rect 94770 -118540 95890 -118530
rect 94770 -118590 94780 -118540
rect 95880 -118590 95890 -118540
rect 94770 -118600 95890 -118590
rect 96270 -118540 97390 -118530
rect 96270 -118590 96280 -118540
rect 97380 -118590 97390 -118540
rect 96270 -118600 97390 -118590
rect 97770 -118540 98890 -118530
rect 97770 -118590 97780 -118540
rect 98880 -118590 98890 -118540
rect 97770 -118600 98890 -118590
rect 99270 -118540 100390 -118530
rect 99270 -118590 99280 -118540
rect 100380 -118590 100390 -118540
rect 99270 -118600 100390 -118590
rect 100770 -118540 101890 -118530
rect 100770 -118590 100780 -118540
rect 101880 -118590 101890 -118540
rect 100770 -118600 101890 -118590
rect 102270 -118540 103390 -118530
rect 102270 -118590 102280 -118540
rect 103380 -118590 103390 -118540
rect 102270 -118600 103390 -118590
rect 103770 -118540 104890 -118530
rect 103770 -118590 103780 -118540
rect 104880 -118590 104890 -118540
rect 103770 -118600 104890 -118590
rect 105270 -118540 106390 -118530
rect 105270 -118590 105280 -118540
rect 106380 -118590 106390 -118540
rect 105270 -118600 106390 -118590
rect 106770 -118540 107890 -118530
rect 106770 -118590 106780 -118540
rect 107880 -118590 107890 -118540
rect 106770 -118600 107890 -118590
rect 108270 -118540 109390 -118530
rect 108270 -118590 108280 -118540
rect 109380 -118590 109390 -118540
rect 108270 -118600 109390 -118590
rect 109770 -118540 110890 -118530
rect 109770 -118590 109780 -118540
rect 110880 -118590 110890 -118540
rect 109770 -118600 110890 -118590
rect 111270 -118540 112390 -118530
rect 111270 -118590 111280 -118540
rect 112380 -118590 112390 -118540
rect 111270 -118600 112390 -118590
rect 112770 -118540 113890 -118530
rect 112770 -118590 112780 -118540
rect 113880 -118590 113890 -118540
rect 112770 -118600 113890 -118590
rect 114270 -118540 115390 -118530
rect 114270 -118590 114280 -118540
rect 115380 -118590 115390 -118540
rect 114270 -118600 115390 -118590
rect 115770 -118540 116890 -118530
rect 115770 -118590 115780 -118540
rect 116880 -118590 116890 -118540
rect 115770 -118600 116890 -118590
rect 117270 -118540 118390 -118530
rect 117270 -118590 117280 -118540
rect 118380 -118590 118390 -118540
rect 117270 -118600 118390 -118590
rect 118770 -118540 119890 -118530
rect 118770 -118590 118780 -118540
rect 119880 -118590 119890 -118540
rect 118770 -118600 119890 -118590
rect 110 -118750 220 -118745
rect 110 -118850 120 -118750
rect 210 -118850 220 -118750
rect 110 -118855 220 -118850
rect 1610 -118750 1720 -118745
rect 1610 -118850 1620 -118750
rect 1710 -118850 1720 -118750
rect 1610 -118855 1720 -118850
rect 3110 -118750 3220 -118745
rect 3110 -118850 3120 -118750
rect 3210 -118850 3220 -118750
rect 3110 -118855 3220 -118850
rect 4610 -118750 4720 -118745
rect 4610 -118850 4620 -118750
rect 4710 -118850 4720 -118750
rect 4610 -118855 4720 -118850
rect 6110 -118750 6220 -118745
rect 6110 -118850 6120 -118750
rect 6210 -118850 6220 -118750
rect 6110 -118855 6220 -118850
rect 7610 -118750 7720 -118745
rect 7610 -118850 7620 -118750
rect 7710 -118850 7720 -118750
rect 7610 -118855 7720 -118850
rect 9110 -118750 9220 -118745
rect 9110 -118850 9120 -118750
rect 9210 -118850 9220 -118750
rect 9110 -118855 9220 -118850
rect 10610 -118750 10720 -118745
rect 10610 -118850 10620 -118750
rect 10710 -118850 10720 -118750
rect 10610 -118855 10720 -118850
rect 12110 -118750 12220 -118745
rect 12110 -118850 12120 -118750
rect 12210 -118850 12220 -118750
rect 12110 -118855 12220 -118850
rect 13610 -118750 13720 -118745
rect 13610 -118850 13620 -118750
rect 13710 -118850 13720 -118750
rect 13610 -118855 13720 -118850
rect 15110 -118750 15220 -118745
rect 15110 -118850 15120 -118750
rect 15210 -118850 15220 -118750
rect 15110 -118855 15220 -118850
rect 16610 -118750 16720 -118745
rect 16610 -118850 16620 -118750
rect 16710 -118850 16720 -118750
rect 16610 -118855 16720 -118850
rect 18110 -118750 18220 -118745
rect 18110 -118850 18120 -118750
rect 18210 -118850 18220 -118750
rect 18110 -118855 18220 -118850
rect 19610 -118750 19720 -118745
rect 19610 -118850 19620 -118750
rect 19710 -118850 19720 -118750
rect 19610 -118855 19720 -118850
rect 21110 -118750 21220 -118745
rect 21110 -118850 21120 -118750
rect 21210 -118850 21220 -118750
rect 21110 -118855 21220 -118850
rect 22610 -118750 22720 -118745
rect 22610 -118850 22620 -118750
rect 22710 -118850 22720 -118750
rect 22610 -118855 22720 -118850
rect 24110 -118750 24220 -118745
rect 24110 -118850 24120 -118750
rect 24210 -118850 24220 -118750
rect 24110 -118855 24220 -118850
rect 25610 -118750 25720 -118745
rect 25610 -118850 25620 -118750
rect 25710 -118850 25720 -118750
rect 25610 -118855 25720 -118850
rect 27110 -118750 27220 -118745
rect 27110 -118850 27120 -118750
rect 27210 -118850 27220 -118750
rect 27110 -118855 27220 -118850
rect 28610 -118750 28720 -118745
rect 28610 -118850 28620 -118750
rect 28710 -118850 28720 -118750
rect 28610 -118855 28720 -118850
rect 30110 -118750 30220 -118745
rect 30110 -118850 30120 -118750
rect 30210 -118850 30220 -118750
rect 30110 -118855 30220 -118850
rect 31610 -118750 31720 -118745
rect 31610 -118850 31620 -118750
rect 31710 -118850 31720 -118750
rect 31610 -118855 31720 -118850
rect 33110 -118750 33220 -118745
rect 33110 -118850 33120 -118750
rect 33210 -118850 33220 -118750
rect 33110 -118855 33220 -118850
rect 34610 -118750 34720 -118745
rect 34610 -118850 34620 -118750
rect 34710 -118850 34720 -118750
rect 34610 -118855 34720 -118850
rect 36110 -118750 36220 -118745
rect 36110 -118850 36120 -118750
rect 36210 -118850 36220 -118750
rect 36110 -118855 36220 -118850
rect 37610 -118750 37720 -118745
rect 37610 -118850 37620 -118750
rect 37710 -118850 37720 -118750
rect 37610 -118855 37720 -118850
rect 39110 -118750 39220 -118745
rect 39110 -118850 39120 -118750
rect 39210 -118850 39220 -118750
rect 39110 -118855 39220 -118850
rect 40610 -118750 40720 -118745
rect 40610 -118850 40620 -118750
rect 40710 -118850 40720 -118750
rect 40610 -118855 40720 -118850
rect 42110 -118750 42220 -118745
rect 42110 -118850 42120 -118750
rect 42210 -118850 42220 -118750
rect 42110 -118855 42220 -118850
rect 43610 -118750 43720 -118745
rect 43610 -118850 43620 -118750
rect 43710 -118850 43720 -118750
rect 43610 -118855 43720 -118850
rect 45110 -118750 45220 -118745
rect 45110 -118850 45120 -118750
rect 45210 -118850 45220 -118750
rect 45110 -118855 45220 -118850
rect 46610 -118750 46720 -118745
rect 46610 -118850 46620 -118750
rect 46710 -118850 46720 -118750
rect 46610 -118855 46720 -118850
rect 48110 -118750 48220 -118745
rect 48110 -118850 48120 -118750
rect 48210 -118850 48220 -118750
rect 48110 -118855 48220 -118850
rect 49610 -118750 49720 -118745
rect 49610 -118850 49620 -118750
rect 49710 -118850 49720 -118750
rect 49610 -118855 49720 -118850
rect 51110 -118750 51220 -118745
rect 51110 -118850 51120 -118750
rect 51210 -118850 51220 -118750
rect 51110 -118855 51220 -118850
rect 52610 -118750 52720 -118745
rect 52610 -118850 52620 -118750
rect 52710 -118850 52720 -118750
rect 52610 -118855 52720 -118850
rect 54110 -118750 54220 -118745
rect 54110 -118850 54120 -118750
rect 54210 -118850 54220 -118750
rect 54110 -118855 54220 -118850
rect 55610 -118750 55720 -118745
rect 55610 -118850 55620 -118750
rect 55710 -118850 55720 -118750
rect 55610 -118855 55720 -118850
rect 57110 -118750 57220 -118745
rect 57110 -118850 57120 -118750
rect 57210 -118850 57220 -118750
rect 57110 -118855 57220 -118850
rect 58610 -118750 58720 -118745
rect 58610 -118850 58620 -118750
rect 58710 -118850 58720 -118750
rect 58610 -118855 58720 -118850
rect 60110 -118750 60220 -118745
rect 60110 -118850 60120 -118750
rect 60210 -118850 60220 -118750
rect 60110 -118855 60220 -118850
rect 61610 -118750 61720 -118745
rect 61610 -118850 61620 -118750
rect 61710 -118850 61720 -118750
rect 61610 -118855 61720 -118850
rect 63110 -118750 63220 -118745
rect 63110 -118850 63120 -118750
rect 63210 -118850 63220 -118750
rect 63110 -118855 63220 -118850
rect 64610 -118750 64720 -118745
rect 64610 -118850 64620 -118750
rect 64710 -118850 64720 -118750
rect 64610 -118855 64720 -118850
rect 66110 -118750 66220 -118745
rect 66110 -118850 66120 -118750
rect 66210 -118850 66220 -118750
rect 66110 -118855 66220 -118850
rect 67610 -118750 67720 -118745
rect 67610 -118850 67620 -118750
rect 67710 -118850 67720 -118750
rect 67610 -118855 67720 -118850
rect 69110 -118750 69220 -118745
rect 69110 -118850 69120 -118750
rect 69210 -118850 69220 -118750
rect 69110 -118855 69220 -118850
rect 70610 -118750 70720 -118745
rect 70610 -118850 70620 -118750
rect 70710 -118850 70720 -118750
rect 70610 -118855 70720 -118850
rect 72110 -118750 72220 -118745
rect 72110 -118850 72120 -118750
rect 72210 -118850 72220 -118750
rect 72110 -118855 72220 -118850
rect 73610 -118750 73720 -118745
rect 73610 -118850 73620 -118750
rect 73710 -118850 73720 -118750
rect 73610 -118855 73720 -118850
rect 75110 -118750 75220 -118745
rect 75110 -118850 75120 -118750
rect 75210 -118850 75220 -118750
rect 75110 -118855 75220 -118850
rect 76610 -118750 76720 -118745
rect 76610 -118850 76620 -118750
rect 76710 -118850 76720 -118750
rect 76610 -118855 76720 -118850
rect 78110 -118750 78220 -118745
rect 78110 -118850 78120 -118750
rect 78210 -118850 78220 -118750
rect 78110 -118855 78220 -118850
rect 79610 -118750 79720 -118745
rect 79610 -118850 79620 -118750
rect 79710 -118850 79720 -118750
rect 79610 -118855 79720 -118850
rect 81110 -118750 81220 -118745
rect 81110 -118850 81120 -118750
rect 81210 -118850 81220 -118750
rect 81110 -118855 81220 -118850
rect 82610 -118750 82720 -118745
rect 82610 -118850 82620 -118750
rect 82710 -118850 82720 -118750
rect 82610 -118855 82720 -118850
rect 84110 -118750 84220 -118745
rect 84110 -118850 84120 -118750
rect 84210 -118850 84220 -118750
rect 84110 -118855 84220 -118850
rect 85610 -118750 85720 -118745
rect 85610 -118850 85620 -118750
rect 85710 -118850 85720 -118750
rect 85610 -118855 85720 -118850
rect 87110 -118750 87220 -118745
rect 87110 -118850 87120 -118750
rect 87210 -118850 87220 -118750
rect 87110 -118855 87220 -118850
rect 88610 -118750 88720 -118745
rect 88610 -118850 88620 -118750
rect 88710 -118850 88720 -118750
rect 88610 -118855 88720 -118850
rect 90110 -118750 90220 -118745
rect 90110 -118850 90120 -118750
rect 90210 -118850 90220 -118750
rect 90110 -118855 90220 -118850
rect 91610 -118750 91720 -118745
rect 91610 -118850 91620 -118750
rect 91710 -118850 91720 -118750
rect 91610 -118855 91720 -118850
rect 93110 -118750 93220 -118745
rect 93110 -118850 93120 -118750
rect 93210 -118850 93220 -118750
rect 93110 -118855 93220 -118850
rect 94610 -118750 94720 -118745
rect 94610 -118850 94620 -118750
rect 94710 -118850 94720 -118750
rect 94610 -118855 94720 -118850
rect 96110 -118750 96220 -118745
rect 96110 -118850 96120 -118750
rect 96210 -118850 96220 -118750
rect 96110 -118855 96220 -118850
rect 97610 -118750 97720 -118745
rect 97610 -118850 97620 -118750
rect 97710 -118850 97720 -118750
rect 97610 -118855 97720 -118850
rect 99110 -118750 99220 -118745
rect 99110 -118850 99120 -118750
rect 99210 -118850 99220 -118750
rect 99110 -118855 99220 -118850
rect 100610 -118750 100720 -118745
rect 100610 -118850 100620 -118750
rect 100710 -118850 100720 -118750
rect 100610 -118855 100720 -118850
rect 102110 -118750 102220 -118745
rect 102110 -118850 102120 -118750
rect 102210 -118850 102220 -118750
rect 102110 -118855 102220 -118850
rect 103610 -118750 103720 -118745
rect 103610 -118850 103620 -118750
rect 103710 -118850 103720 -118750
rect 103610 -118855 103720 -118850
rect 105110 -118750 105220 -118745
rect 105110 -118850 105120 -118750
rect 105210 -118850 105220 -118750
rect 105110 -118855 105220 -118850
rect 106610 -118750 106720 -118745
rect 106610 -118850 106620 -118750
rect 106710 -118850 106720 -118750
rect 106610 -118855 106720 -118850
rect 108110 -118750 108220 -118745
rect 108110 -118850 108120 -118750
rect 108210 -118850 108220 -118750
rect 108110 -118855 108220 -118850
rect 109610 -118750 109720 -118745
rect 109610 -118850 109620 -118750
rect 109710 -118850 109720 -118750
rect 109610 -118855 109720 -118850
rect 111110 -118750 111220 -118745
rect 111110 -118850 111120 -118750
rect 111210 -118850 111220 -118750
rect 111110 -118855 111220 -118850
rect 112610 -118750 112720 -118745
rect 112610 -118850 112620 -118750
rect 112710 -118850 112720 -118750
rect 112610 -118855 112720 -118850
rect 114110 -118750 114220 -118745
rect 114110 -118850 114120 -118750
rect 114210 -118850 114220 -118750
rect 114110 -118855 114220 -118850
rect 115610 -118750 115720 -118745
rect 115610 -118850 115620 -118750
rect 115710 -118850 115720 -118750
rect 115610 -118855 115720 -118850
rect 117110 -118750 117220 -118745
rect 117110 -118850 117120 -118750
rect 117210 -118850 117220 -118750
rect 117110 -118855 117220 -118850
rect 118610 -118750 118720 -118745
rect 118610 -118850 118620 -118750
rect 118710 -118850 118720 -118750
rect 118610 -118855 118720 -118850
<< via3 >>
rect 245 1780 290 1825
rect 1745 1780 1790 1825
rect 3245 1780 3290 1825
rect 4745 1780 4790 1825
rect 6245 1780 6290 1825
rect 7745 1780 7790 1825
rect 9245 1780 9290 1825
rect 10745 1780 10790 1825
rect 12245 1780 12290 1825
rect 13745 1780 13790 1825
rect 15245 1780 15290 1825
rect 16745 1780 16790 1825
rect 18245 1780 18290 1825
rect 19745 1780 19790 1825
rect 21245 1780 21290 1825
rect 22745 1780 22790 1825
rect 24245 1780 24290 1825
rect 25745 1780 25790 1825
rect 27245 1780 27290 1825
rect 28745 1780 28790 1825
rect 30245 1780 30290 1825
rect 31745 1780 31790 1825
rect 33245 1780 33290 1825
rect 34745 1780 34790 1825
rect 36245 1780 36290 1825
rect 37745 1780 37790 1825
rect 39245 1780 39290 1825
rect 40745 1780 40790 1825
rect 42245 1780 42290 1825
rect 43745 1780 43790 1825
rect 45245 1780 45290 1825
rect 46745 1780 46790 1825
rect 48245 1780 48290 1825
rect 49745 1780 49790 1825
rect 51245 1780 51290 1825
rect 52745 1780 52790 1825
rect 54245 1780 54290 1825
rect 55745 1780 55790 1825
rect 57245 1780 57290 1825
rect 58745 1780 58790 1825
rect 60245 1780 60290 1825
rect 61745 1780 61790 1825
rect 63245 1780 63290 1825
rect 64745 1780 64790 1825
rect 66245 1780 66290 1825
rect 67745 1780 67790 1825
rect 69245 1780 69290 1825
rect 70745 1780 70790 1825
rect 72245 1780 72290 1825
rect 73745 1780 73790 1825
rect 75245 1780 75290 1825
rect 76745 1780 76790 1825
rect 78245 1780 78290 1825
rect 79745 1780 79790 1825
rect 81245 1780 81290 1825
rect 82745 1780 82790 1825
rect 84245 1780 84290 1825
rect 85745 1780 85790 1825
rect 87245 1780 87290 1825
rect 88745 1780 88790 1825
rect 90245 1780 90290 1825
rect 91745 1780 91790 1825
rect 93245 1780 93290 1825
rect 94745 1780 94790 1825
rect 96245 1780 96290 1825
rect 97745 1780 97790 1825
rect 99245 1780 99290 1825
rect 100745 1780 100790 1825
rect 102245 1780 102290 1825
rect 103745 1780 103790 1825
rect 105245 1780 105290 1825
rect 106745 1780 106790 1825
rect 108245 1780 108290 1825
rect 109745 1780 109790 1825
rect 111245 1780 111290 1825
rect 112745 1780 112790 1825
rect 114245 1780 114290 1825
rect 115745 1780 115790 1825
rect 117245 1780 117290 1825
rect 118745 1780 118790 1825
rect -235 1235 -190 1270
rect -235 -265 -190 -230
rect -235 -1765 -190 -1730
rect -235 -3265 -190 -3230
rect -235 -4765 -190 -4730
rect -235 -6265 -190 -6230
rect -235 -7765 -190 -7730
rect -235 -9265 -190 -9230
rect -235 -10765 -190 -10730
rect -235 -12265 -190 -12230
rect -235 -13765 -190 -13730
rect -235 -15265 -190 -15230
rect -235 -16765 -190 -16730
rect -235 -18265 -190 -18230
rect -235 -19765 -190 -19730
rect -235 -21265 -190 -21230
rect -235 -22765 -190 -22730
rect -235 -24265 -190 -24230
rect -235 -25765 -190 -25730
rect -235 -27265 -190 -27230
rect -235 -28765 -190 -28730
rect -235 -30265 -190 -30230
rect -235 -31765 -190 -31730
rect -235 -33265 -190 -33230
rect -235 -34765 -190 -34730
rect -235 -36265 -190 -36230
rect -235 -37765 -190 -37730
rect -235 -39265 -190 -39230
rect -235 -40765 -190 -40730
rect -235 -42265 -190 -42230
rect -235 -43765 -190 -43730
rect -235 -45265 -190 -45230
rect -235 -46765 -190 -46730
rect -235 -48265 -190 -48230
rect -235 -49765 -190 -49730
rect -235 -51265 -190 -51230
rect -235 -52765 -190 -52730
rect -235 -54265 -190 -54230
rect -235 -55765 -190 -55730
rect -235 -57265 -190 -57230
rect -235 -58765 -190 -58730
rect -235 -60265 -190 -60230
rect -235 -61765 -190 -61730
rect -235 -63265 -190 -63230
rect -235 -64765 -190 -64730
rect -235 -66265 -190 -66230
rect -235 -67765 -190 -67730
rect -235 -69265 -190 -69230
rect -235 -70765 -190 -70730
rect -235 -72265 -190 -72230
rect -235 -73765 -190 -73730
rect -235 -75265 -190 -75230
rect -235 -76765 -190 -76730
rect -235 -78265 -190 -78230
rect -235 -79765 -190 -79730
rect -235 -81265 -190 -81230
rect -235 -82765 -190 -82730
rect -235 -84265 -190 -84230
rect -235 -85765 -190 -85730
rect -235 -87265 -190 -87230
rect -235 -88765 -190 -88730
rect -235 -90265 -190 -90230
rect -235 -91765 -190 -91730
rect -235 -93265 -190 -93230
rect -235 -94765 -190 -94730
rect -235 -96265 -190 -96230
rect -235 -97765 -190 -97730
rect -235 -99265 -190 -99230
rect -235 -100765 -190 -100730
rect -235 -102265 -190 -102230
rect -235 -103765 -190 -103730
rect -235 -105265 -190 -105230
rect -235 -106765 -190 -106730
rect -235 -108265 -190 -108230
rect -235 -109765 -190 -109730
rect -235 -111265 -190 -111230
rect -235 -112765 -190 -112730
rect -235 -114265 -190 -114230
rect -235 -115765 -190 -115730
rect -235 -117265 -190 -117230
rect 280 -118590 1380 -118540
rect 1780 -118590 2880 -118540
rect 3280 -118590 4380 -118540
rect 4780 -118590 5880 -118540
rect 6280 -118590 7380 -118540
rect 7780 -118590 8880 -118540
rect 9280 -118590 10380 -118540
rect 10780 -118590 11880 -118540
rect 12280 -118590 13380 -118540
rect 13780 -118590 14880 -118540
rect 15280 -118590 16380 -118540
rect 16780 -118590 17880 -118540
rect 18280 -118590 19380 -118540
rect 19780 -118590 20880 -118540
rect 21280 -118590 22380 -118540
rect 22780 -118590 23880 -118540
rect 24280 -118590 25380 -118540
rect 25780 -118590 26880 -118540
rect 27280 -118590 28380 -118540
rect 28780 -118590 29880 -118540
rect 30280 -118590 31380 -118540
rect 31780 -118590 32880 -118540
rect 33280 -118590 34380 -118540
rect 34780 -118590 35880 -118540
rect 36280 -118590 37380 -118540
rect 37780 -118590 38880 -118540
rect 39280 -118590 40380 -118540
rect 40780 -118590 41880 -118540
rect 42280 -118590 43380 -118540
rect 43780 -118590 44880 -118540
rect 45280 -118590 46380 -118540
rect 46780 -118590 47880 -118540
rect 48280 -118590 49380 -118540
rect 49780 -118590 50880 -118540
rect 51280 -118590 52380 -118540
rect 52780 -118590 53880 -118540
rect 54280 -118590 55380 -118540
rect 55780 -118590 56880 -118540
rect 57280 -118590 58380 -118540
rect 58780 -118590 59880 -118540
rect 60280 -118590 61380 -118540
rect 61780 -118590 62880 -118540
rect 63280 -118590 64380 -118540
rect 64780 -118590 65880 -118540
rect 66280 -118590 67380 -118540
rect 67780 -118590 68880 -118540
rect 69280 -118590 70380 -118540
rect 70780 -118590 71880 -118540
rect 72280 -118590 73380 -118540
rect 73780 -118590 74880 -118540
rect 75280 -118590 76380 -118540
rect 76780 -118590 77880 -118540
rect 78280 -118590 79380 -118540
rect 79780 -118590 80880 -118540
rect 81280 -118590 82380 -118540
rect 82780 -118590 83880 -118540
rect 84280 -118590 85380 -118540
rect 85780 -118590 86880 -118540
rect 87280 -118590 88380 -118540
rect 88780 -118590 89880 -118540
rect 90280 -118590 91380 -118540
rect 91780 -118590 92880 -118540
rect 93280 -118590 94380 -118540
rect 94780 -118590 95880 -118540
rect 96280 -118590 97380 -118540
rect 97780 -118590 98880 -118540
rect 99280 -118590 100380 -118540
rect 100780 -118590 101880 -118540
rect 102280 -118590 103380 -118540
rect 103780 -118590 104880 -118540
rect 105280 -118590 106380 -118540
rect 106780 -118590 107880 -118540
rect 108280 -118590 109380 -118540
rect 109780 -118590 110880 -118540
rect 111280 -118590 112380 -118540
rect 112780 -118590 113880 -118540
rect 114280 -118590 115380 -118540
rect 115780 -118590 116880 -118540
rect 117280 -118590 118380 -118540
rect 118780 -118590 119880 -118540
rect 120 -118850 210 -118750
rect 1620 -118850 1710 -118750
rect 3120 -118850 3210 -118750
rect 4620 -118850 4710 -118750
rect 6120 -118850 6210 -118750
rect 7620 -118850 7710 -118750
rect 9120 -118850 9210 -118750
rect 10620 -118850 10710 -118750
rect 12120 -118850 12210 -118750
rect 13620 -118850 13710 -118750
rect 15120 -118850 15210 -118750
rect 16620 -118850 16710 -118750
rect 18120 -118850 18210 -118750
rect 19620 -118850 19710 -118750
rect 21120 -118850 21210 -118750
rect 22620 -118850 22710 -118750
rect 24120 -118850 24210 -118750
rect 25620 -118850 25710 -118750
rect 27120 -118850 27210 -118750
rect 28620 -118850 28710 -118750
rect 30120 -118850 30210 -118750
rect 31620 -118850 31710 -118750
rect 33120 -118850 33210 -118750
rect 34620 -118850 34710 -118750
rect 36120 -118850 36210 -118750
rect 37620 -118850 37710 -118750
rect 39120 -118850 39210 -118750
rect 40620 -118850 40710 -118750
rect 42120 -118850 42210 -118750
rect 43620 -118850 43710 -118750
rect 45120 -118850 45210 -118750
rect 46620 -118850 46710 -118750
rect 48120 -118850 48210 -118750
rect 49620 -118850 49710 -118750
rect 51120 -118850 51210 -118750
rect 52620 -118850 52710 -118750
rect 54120 -118850 54210 -118750
rect 55620 -118850 55710 -118750
rect 57120 -118850 57210 -118750
rect 58620 -118850 58710 -118750
rect 60120 -118850 60210 -118750
rect 61620 -118850 61710 -118750
rect 63120 -118850 63210 -118750
rect 64620 -118850 64710 -118750
rect 66120 -118850 66210 -118750
rect 67620 -118850 67710 -118750
rect 69120 -118850 69210 -118750
rect 70620 -118850 70710 -118750
rect 72120 -118850 72210 -118750
rect 73620 -118850 73710 -118750
rect 75120 -118850 75210 -118750
rect 76620 -118850 76710 -118750
rect 78120 -118850 78210 -118750
rect 79620 -118850 79710 -118750
rect 81120 -118850 81210 -118750
rect 82620 -118850 82710 -118750
rect 84120 -118850 84210 -118750
rect 85620 -118850 85710 -118750
rect 87120 -118850 87210 -118750
rect 88620 -118850 88710 -118750
rect 90120 -118850 90210 -118750
rect 91620 -118850 91710 -118750
rect 93120 -118850 93210 -118750
rect 94620 -118850 94710 -118750
rect 96120 -118850 96210 -118750
rect 97620 -118850 97710 -118750
rect 99120 -118850 99210 -118750
rect 100620 -118850 100710 -118750
rect 102120 -118850 102210 -118750
rect 103620 -118850 103710 -118750
rect 105120 -118850 105210 -118750
rect 106620 -118850 106710 -118750
rect 108120 -118850 108210 -118750
rect 109620 -118850 109710 -118750
rect 111120 -118850 111210 -118750
rect 112620 -118850 112710 -118750
rect 114120 -118850 114210 -118750
rect 115620 -118850 115710 -118750
rect 117120 -118850 117210 -118750
rect 118620 -118850 118710 -118750
<< metal4 >>
rect -1500 1825 119600 1830
rect -1500 1780 245 1825
rect 290 1780 1745 1825
rect 1790 1780 3245 1825
rect 3290 1780 4745 1825
rect 4790 1780 6245 1825
rect 6290 1780 7745 1825
rect 7790 1780 9245 1825
rect 9290 1780 10745 1825
rect 10790 1780 12245 1825
rect 12290 1780 13745 1825
rect 13790 1780 15245 1825
rect 15290 1780 16745 1825
rect 16790 1780 18245 1825
rect 18290 1780 19745 1825
rect 19790 1780 21245 1825
rect 21290 1780 22745 1825
rect 22790 1780 24245 1825
rect 24290 1780 25745 1825
rect 25790 1780 27245 1825
rect 27290 1780 28745 1825
rect 28790 1780 30245 1825
rect 30290 1780 31745 1825
rect 31790 1780 33245 1825
rect 33290 1780 34745 1825
rect 34790 1780 36245 1825
rect 36290 1780 37745 1825
rect 37790 1780 39245 1825
rect 39290 1780 40745 1825
rect 40790 1780 42245 1825
rect 42290 1780 43745 1825
rect 43790 1780 45245 1825
rect 45290 1780 46745 1825
rect 46790 1780 48245 1825
rect 48290 1780 49745 1825
rect 49790 1780 51245 1825
rect 51290 1780 52745 1825
rect 52790 1780 54245 1825
rect 54290 1780 55745 1825
rect 55790 1780 57245 1825
rect 57290 1780 58745 1825
rect 58790 1780 60245 1825
rect 60290 1780 61745 1825
rect 61790 1780 63245 1825
rect 63290 1780 64745 1825
rect 64790 1780 66245 1825
rect 66290 1780 67745 1825
rect 67790 1780 69245 1825
rect 69290 1780 70745 1825
rect 70790 1780 72245 1825
rect 72290 1780 73745 1825
rect 73790 1780 75245 1825
rect 75290 1780 76745 1825
rect 76790 1780 78245 1825
rect 78290 1780 79745 1825
rect 79790 1780 81245 1825
rect 81290 1780 82745 1825
rect 82790 1780 84245 1825
rect 84290 1780 85745 1825
rect 85790 1780 87245 1825
rect 87290 1780 88745 1825
rect 88790 1780 90245 1825
rect 90290 1780 91745 1825
rect 91790 1780 93245 1825
rect 93290 1780 94745 1825
rect 94790 1780 96245 1825
rect 96290 1780 97745 1825
rect 97790 1780 99245 1825
rect 99290 1780 100745 1825
rect 100790 1780 102245 1825
rect 102290 1780 103745 1825
rect 103790 1780 105245 1825
rect 105290 1780 106745 1825
rect 106790 1780 108245 1825
rect 108290 1780 109745 1825
rect 109790 1780 111245 1825
rect 111290 1780 112745 1825
rect 112790 1780 114245 1825
rect 114290 1780 115745 1825
rect 115790 1780 117245 1825
rect 117290 1780 118745 1825
rect 118790 1780 119600 1825
rect -1500 1775 119600 1780
rect -240 1270 -185 1300
rect -240 1235 -235 1270
rect -190 1235 -185 1270
rect -240 -230 -185 1235
rect -240 -265 -235 -230
rect -190 -265 -185 -230
rect -240 -1730 -185 -265
rect -240 -1765 -235 -1730
rect -190 -1765 -185 -1730
rect -240 -3230 -185 -1765
rect -240 -3265 -235 -3230
rect -190 -3265 -185 -3230
rect -240 -4730 -185 -3265
rect -240 -4765 -235 -4730
rect -190 -4765 -185 -4730
rect -240 -6230 -185 -4765
rect -240 -6265 -235 -6230
rect -190 -6265 -185 -6230
rect -240 -7730 -185 -6265
rect -240 -7765 -235 -7730
rect -190 -7765 -185 -7730
rect -240 -9230 -185 -7765
rect -240 -9265 -235 -9230
rect -190 -9265 -185 -9230
rect -240 -10730 -185 -9265
rect -240 -10765 -235 -10730
rect -190 -10765 -185 -10730
rect -240 -12230 -185 -10765
rect -240 -12265 -235 -12230
rect -190 -12265 -185 -12230
rect -240 -13730 -185 -12265
rect -240 -13765 -235 -13730
rect -190 -13765 -185 -13730
rect -240 -15230 -185 -13765
rect -240 -15265 -235 -15230
rect -190 -15265 -185 -15230
rect -240 -16730 -185 -15265
rect -240 -16765 -235 -16730
rect -190 -16765 -185 -16730
rect -240 -18230 -185 -16765
rect -240 -18265 -235 -18230
rect -190 -18265 -185 -18230
rect -240 -19730 -185 -18265
rect -240 -19765 -235 -19730
rect -190 -19765 -185 -19730
rect -240 -21230 -185 -19765
rect -240 -21265 -235 -21230
rect -190 -21265 -185 -21230
rect -240 -22730 -185 -21265
rect -240 -22765 -235 -22730
rect -190 -22765 -185 -22730
rect -240 -24230 -185 -22765
rect -240 -24265 -235 -24230
rect -190 -24265 -185 -24230
rect -240 -25730 -185 -24265
rect -240 -25765 -235 -25730
rect -190 -25765 -185 -25730
rect -240 -27230 -185 -25765
rect -240 -27265 -235 -27230
rect -190 -27265 -185 -27230
rect -240 -28730 -185 -27265
rect -240 -28765 -235 -28730
rect -190 -28765 -185 -28730
rect -240 -30230 -185 -28765
rect -240 -30265 -235 -30230
rect -190 -30265 -185 -30230
rect -240 -31730 -185 -30265
rect -240 -31765 -235 -31730
rect -190 -31765 -185 -31730
rect -240 -33230 -185 -31765
rect -240 -33265 -235 -33230
rect -190 -33265 -185 -33230
rect -240 -34730 -185 -33265
rect -240 -34765 -235 -34730
rect -190 -34765 -185 -34730
rect -240 -36230 -185 -34765
rect -240 -36265 -235 -36230
rect -190 -36265 -185 -36230
rect -240 -37730 -185 -36265
rect -240 -37765 -235 -37730
rect -190 -37765 -185 -37730
rect -240 -39230 -185 -37765
rect -240 -39265 -235 -39230
rect -190 -39265 -185 -39230
rect -240 -40730 -185 -39265
rect -240 -40765 -235 -40730
rect -190 -40765 -185 -40730
rect -240 -42230 -185 -40765
rect -240 -42265 -235 -42230
rect -190 -42265 -185 -42230
rect -240 -43730 -185 -42265
rect -240 -43765 -235 -43730
rect -190 -43765 -185 -43730
rect -240 -45230 -185 -43765
rect -240 -45265 -235 -45230
rect -190 -45265 -185 -45230
rect -240 -46730 -185 -45265
rect -240 -46765 -235 -46730
rect -190 -46765 -185 -46730
rect -240 -48230 -185 -46765
rect -240 -48265 -235 -48230
rect -190 -48265 -185 -48230
rect -240 -49730 -185 -48265
rect -240 -49765 -235 -49730
rect -190 -49765 -185 -49730
rect -240 -51230 -185 -49765
rect -240 -51265 -235 -51230
rect -190 -51265 -185 -51230
rect -240 -52730 -185 -51265
rect -240 -52765 -235 -52730
rect -190 -52765 -185 -52730
rect -240 -54230 -185 -52765
rect -240 -54265 -235 -54230
rect -190 -54265 -185 -54230
rect -240 -55730 -185 -54265
rect -240 -55765 -235 -55730
rect -190 -55765 -185 -55730
rect -240 -57230 -185 -55765
rect -240 -57265 -235 -57230
rect -190 -57265 -185 -57230
rect -240 -58730 -185 -57265
rect -240 -58765 -235 -58730
rect -190 -58765 -185 -58730
rect -240 -60230 -185 -58765
rect -240 -60265 -235 -60230
rect -190 -60265 -185 -60230
rect -240 -61730 -185 -60265
rect -240 -61765 -235 -61730
rect -190 -61765 -185 -61730
rect -240 -63230 -185 -61765
rect -240 -63265 -235 -63230
rect -190 -63265 -185 -63230
rect -240 -64730 -185 -63265
rect -240 -64765 -235 -64730
rect -190 -64765 -185 -64730
rect -240 -66230 -185 -64765
rect -240 -66265 -235 -66230
rect -190 -66265 -185 -66230
rect -240 -67730 -185 -66265
rect -240 -67765 -235 -67730
rect -190 -67765 -185 -67730
rect -240 -69230 -185 -67765
rect -240 -69265 -235 -69230
rect -190 -69265 -185 -69230
rect -240 -70730 -185 -69265
rect -240 -70765 -235 -70730
rect -190 -70765 -185 -70730
rect -240 -72230 -185 -70765
rect -240 -72265 -235 -72230
rect -190 -72265 -185 -72230
rect -240 -73730 -185 -72265
rect -240 -73765 -235 -73730
rect -190 -73765 -185 -73730
rect -240 -75230 -185 -73765
rect -240 -75265 -235 -75230
rect -190 -75265 -185 -75230
rect -240 -76730 -185 -75265
rect -240 -76765 -235 -76730
rect -190 -76765 -185 -76730
rect -240 -78230 -185 -76765
rect -240 -78265 -235 -78230
rect -190 -78265 -185 -78230
rect -240 -79730 -185 -78265
rect -240 -79765 -235 -79730
rect -190 -79765 -185 -79730
rect -240 -81230 -185 -79765
rect -240 -81265 -235 -81230
rect -190 -81265 -185 -81230
rect -240 -82730 -185 -81265
rect -240 -82765 -235 -82730
rect -190 -82765 -185 -82730
rect -240 -84230 -185 -82765
rect -240 -84265 -235 -84230
rect -190 -84265 -185 -84230
rect -240 -85730 -185 -84265
rect -240 -85765 -235 -85730
rect -190 -85765 -185 -85730
rect -240 -87230 -185 -85765
rect -240 -87265 -235 -87230
rect -190 -87265 -185 -87230
rect -240 -88730 -185 -87265
rect -240 -88765 -235 -88730
rect -190 -88765 -185 -88730
rect -240 -90230 -185 -88765
rect -240 -90265 -235 -90230
rect -190 -90265 -185 -90230
rect -240 -91730 -185 -90265
rect -240 -91765 -235 -91730
rect -190 -91765 -185 -91730
rect -240 -93230 -185 -91765
rect -240 -93265 -235 -93230
rect -190 -93265 -185 -93230
rect -240 -94730 -185 -93265
rect -240 -94765 -235 -94730
rect -190 -94765 -185 -94730
rect -240 -96230 -185 -94765
rect -240 -96265 -235 -96230
rect -190 -96265 -185 -96230
rect -240 -97730 -185 -96265
rect -240 -97765 -235 -97730
rect -190 -97765 -185 -97730
rect -240 -99230 -185 -97765
rect -240 -99265 -235 -99230
rect -190 -99265 -185 -99230
rect -240 -100730 -185 -99265
rect -240 -100765 -235 -100730
rect -190 -100765 -185 -100730
rect -240 -102230 -185 -100765
rect -240 -102265 -235 -102230
rect -190 -102265 -185 -102230
rect -240 -103730 -185 -102265
rect -240 -103765 -235 -103730
rect -190 -103765 -185 -103730
rect -240 -105230 -185 -103765
rect -240 -105265 -235 -105230
rect -190 -105265 -185 -105230
rect -240 -106730 -185 -105265
rect -240 -106765 -235 -106730
rect -190 -106765 -185 -106730
rect -240 -108230 -185 -106765
rect -240 -108265 -235 -108230
rect -190 -108265 -185 -108230
rect -240 -109730 -185 -108265
rect -240 -109765 -235 -109730
rect -190 -109765 -185 -109730
rect -240 -111230 -185 -109765
rect -240 -111265 -235 -111230
rect -190 -111265 -185 -111230
rect -240 -112730 -185 -111265
rect -240 -112765 -235 -112730
rect -190 -112765 -185 -112730
rect -240 -114230 -185 -112765
rect -240 -114265 -235 -114230
rect -190 -114265 -185 -114230
rect -240 -115730 -185 -114265
rect -240 -115765 -235 -115730
rect -190 -115765 -185 -115730
rect -240 -117230 -185 -115765
rect -240 -117265 -235 -117230
rect -190 -117265 -185 -117230
rect -240 -119300 -185 -117265
rect 1315 -118530 1390 -118500
rect 2815 -118530 2890 -118500
rect 4315 -118530 4390 -118500
rect 5815 -118530 5890 -118500
rect 7315 -118530 7390 -118500
rect 8815 -118530 8890 -118500
rect 10315 -118530 10390 -118500
rect 11815 -118530 11890 -118500
rect 13315 -118530 13390 -118500
rect 14815 -118530 14890 -118500
rect 16315 -118530 16390 -118500
rect 17815 -118530 17890 -118500
rect 19315 -118530 19390 -118500
rect 20815 -118530 20890 -118500
rect 22315 -118530 22390 -118500
rect 23815 -118530 23890 -118500
rect 25315 -118530 25390 -118500
rect 26815 -118530 26890 -118500
rect 28315 -118530 28390 -118500
rect 29815 -118530 29890 -118500
rect 31315 -118530 31390 -118500
rect 32815 -118530 32890 -118500
rect 34315 -118530 34390 -118500
rect 35815 -118530 35890 -118500
rect 37315 -118530 37390 -118500
rect 38815 -118530 38890 -118500
rect 40315 -118530 40390 -118500
rect 41815 -118530 41890 -118500
rect 43315 -118530 43390 -118500
rect 44815 -118530 44890 -118500
rect 46315 -118530 46390 -118500
rect 47815 -118530 47890 -118500
rect 49315 -118530 49390 -118500
rect 50815 -118530 50890 -118500
rect 52315 -118530 52390 -118500
rect 53815 -118530 53890 -118500
rect 55315 -118530 55390 -118500
rect 56815 -118530 56890 -118500
rect 58315 -118530 58390 -118500
rect 59815 -118530 59890 -118500
rect 61315 -118530 61390 -118500
rect 62815 -118530 62890 -118500
rect 64315 -118530 64390 -118500
rect 65815 -118530 65890 -118500
rect 67315 -118530 67390 -118500
rect 68815 -118530 68890 -118500
rect 70315 -118530 70390 -118500
rect 71815 -118530 71890 -118500
rect 73315 -118530 73390 -118500
rect 74815 -118530 74890 -118500
rect 76315 -118530 76390 -118500
rect 77815 -118530 77890 -118500
rect 79315 -118530 79390 -118500
rect 80815 -118530 80890 -118500
rect 82315 -118530 82390 -118500
rect 83815 -118530 83890 -118500
rect 85315 -118530 85390 -118500
rect 86815 -118530 86890 -118500
rect 88315 -118530 88390 -118500
rect 89815 -118530 89890 -118500
rect 91315 -118530 91390 -118500
rect 92815 -118530 92890 -118500
rect 94315 -118530 94390 -118500
rect 95815 -118530 95890 -118500
rect 97315 -118530 97390 -118500
rect 98815 -118530 98890 -118500
rect 100315 -118530 100390 -118500
rect 101815 -118530 101890 -118500
rect 103315 -118530 103390 -118500
rect 104815 -118530 104890 -118500
rect 106315 -118530 106390 -118500
rect 107815 -118530 107890 -118500
rect 109315 -118530 109390 -118500
rect 110815 -118530 110890 -118500
rect 112315 -118530 112390 -118500
rect 113815 -118530 113890 -118500
rect 115315 -118530 115390 -118500
rect 116815 -118530 116890 -118500
rect 118315 -118530 118390 -118500
rect 119815 -118530 119890 -118500
rect 270 -118540 1390 -118530
rect 270 -118590 280 -118540
rect 1380 -118590 1390 -118540
rect 270 -118600 1390 -118590
rect 1770 -118540 2890 -118530
rect 1770 -118590 1780 -118540
rect 2880 -118590 2890 -118540
rect 1770 -118600 2890 -118590
rect 3270 -118540 4390 -118530
rect 3270 -118590 3280 -118540
rect 4380 -118590 4390 -118540
rect 3270 -118600 4390 -118590
rect 4770 -118540 5890 -118530
rect 4770 -118590 4780 -118540
rect 5880 -118590 5890 -118540
rect 4770 -118600 5890 -118590
rect 6270 -118540 7390 -118530
rect 6270 -118590 6280 -118540
rect 7380 -118590 7390 -118540
rect 6270 -118600 7390 -118590
rect 7770 -118540 8890 -118530
rect 7770 -118590 7780 -118540
rect 8880 -118590 8890 -118540
rect 7770 -118600 8890 -118590
rect 9270 -118540 10390 -118530
rect 9270 -118590 9280 -118540
rect 10380 -118590 10390 -118540
rect 9270 -118600 10390 -118590
rect 10770 -118540 11890 -118530
rect 10770 -118590 10780 -118540
rect 11880 -118590 11890 -118540
rect 10770 -118600 11890 -118590
rect 12270 -118540 13390 -118530
rect 12270 -118590 12280 -118540
rect 13380 -118590 13390 -118540
rect 12270 -118600 13390 -118590
rect 13770 -118540 14890 -118530
rect 13770 -118590 13780 -118540
rect 14880 -118590 14890 -118540
rect 13770 -118600 14890 -118590
rect 15270 -118540 16390 -118530
rect 15270 -118590 15280 -118540
rect 16380 -118590 16390 -118540
rect 15270 -118600 16390 -118590
rect 16770 -118540 17890 -118530
rect 16770 -118590 16780 -118540
rect 17880 -118590 17890 -118540
rect 16770 -118600 17890 -118590
rect 18270 -118540 19390 -118530
rect 18270 -118590 18280 -118540
rect 19380 -118590 19390 -118540
rect 18270 -118600 19390 -118590
rect 19770 -118540 20890 -118530
rect 19770 -118590 19780 -118540
rect 20880 -118590 20890 -118540
rect 19770 -118600 20890 -118590
rect 21270 -118540 22390 -118530
rect 21270 -118590 21280 -118540
rect 22380 -118590 22390 -118540
rect 21270 -118600 22390 -118590
rect 22770 -118540 23890 -118530
rect 22770 -118590 22780 -118540
rect 23880 -118590 23890 -118540
rect 22770 -118600 23890 -118590
rect 24270 -118540 25390 -118530
rect 24270 -118590 24280 -118540
rect 25380 -118590 25390 -118540
rect 24270 -118600 25390 -118590
rect 25770 -118540 26890 -118530
rect 25770 -118590 25780 -118540
rect 26880 -118590 26890 -118540
rect 25770 -118600 26890 -118590
rect 27270 -118540 28390 -118530
rect 27270 -118590 27280 -118540
rect 28380 -118590 28390 -118540
rect 27270 -118600 28390 -118590
rect 28770 -118540 29890 -118530
rect 28770 -118590 28780 -118540
rect 29880 -118590 29890 -118540
rect 28770 -118600 29890 -118590
rect 30270 -118540 31390 -118530
rect 30270 -118590 30280 -118540
rect 31380 -118590 31390 -118540
rect 30270 -118600 31390 -118590
rect 31770 -118540 32890 -118530
rect 31770 -118590 31780 -118540
rect 32880 -118590 32890 -118540
rect 31770 -118600 32890 -118590
rect 33270 -118540 34390 -118530
rect 33270 -118590 33280 -118540
rect 34380 -118590 34390 -118540
rect 33270 -118600 34390 -118590
rect 34770 -118540 35890 -118530
rect 34770 -118590 34780 -118540
rect 35880 -118590 35890 -118540
rect 34770 -118600 35890 -118590
rect 36270 -118540 37390 -118530
rect 36270 -118590 36280 -118540
rect 37380 -118590 37390 -118540
rect 36270 -118600 37390 -118590
rect 37770 -118540 38890 -118530
rect 37770 -118590 37780 -118540
rect 38880 -118590 38890 -118540
rect 37770 -118600 38890 -118590
rect 39270 -118540 40390 -118530
rect 39270 -118590 39280 -118540
rect 40380 -118590 40390 -118540
rect 39270 -118600 40390 -118590
rect 40770 -118540 41890 -118530
rect 40770 -118590 40780 -118540
rect 41880 -118590 41890 -118540
rect 40770 -118600 41890 -118590
rect 42270 -118540 43390 -118530
rect 42270 -118590 42280 -118540
rect 43380 -118590 43390 -118540
rect 42270 -118600 43390 -118590
rect 43770 -118540 44890 -118530
rect 43770 -118590 43780 -118540
rect 44880 -118590 44890 -118540
rect 43770 -118600 44890 -118590
rect 45270 -118540 46390 -118530
rect 45270 -118590 45280 -118540
rect 46380 -118590 46390 -118540
rect 45270 -118600 46390 -118590
rect 46770 -118540 47890 -118530
rect 46770 -118590 46780 -118540
rect 47880 -118590 47890 -118540
rect 46770 -118600 47890 -118590
rect 48270 -118540 49390 -118530
rect 48270 -118590 48280 -118540
rect 49380 -118590 49390 -118540
rect 48270 -118600 49390 -118590
rect 49770 -118540 50890 -118530
rect 49770 -118590 49780 -118540
rect 50880 -118590 50890 -118540
rect 49770 -118600 50890 -118590
rect 51270 -118540 52390 -118530
rect 51270 -118590 51280 -118540
rect 52380 -118590 52390 -118540
rect 51270 -118600 52390 -118590
rect 52770 -118540 53890 -118530
rect 52770 -118590 52780 -118540
rect 53880 -118590 53890 -118540
rect 52770 -118600 53890 -118590
rect 54270 -118540 55390 -118530
rect 54270 -118590 54280 -118540
rect 55380 -118590 55390 -118540
rect 54270 -118600 55390 -118590
rect 55770 -118540 56890 -118530
rect 55770 -118590 55780 -118540
rect 56880 -118590 56890 -118540
rect 55770 -118600 56890 -118590
rect 57270 -118540 58390 -118530
rect 57270 -118590 57280 -118540
rect 58380 -118590 58390 -118540
rect 57270 -118600 58390 -118590
rect 58770 -118540 59890 -118530
rect 58770 -118590 58780 -118540
rect 59880 -118590 59890 -118540
rect 58770 -118600 59890 -118590
rect 60270 -118540 61390 -118530
rect 60270 -118590 60280 -118540
rect 61380 -118590 61390 -118540
rect 60270 -118600 61390 -118590
rect 61770 -118540 62890 -118530
rect 61770 -118590 61780 -118540
rect 62880 -118590 62890 -118540
rect 61770 -118600 62890 -118590
rect 63270 -118540 64390 -118530
rect 63270 -118590 63280 -118540
rect 64380 -118590 64390 -118540
rect 63270 -118600 64390 -118590
rect 64770 -118540 65890 -118530
rect 64770 -118590 64780 -118540
rect 65880 -118590 65890 -118540
rect 64770 -118600 65890 -118590
rect 66270 -118540 67390 -118530
rect 66270 -118590 66280 -118540
rect 67380 -118590 67390 -118540
rect 66270 -118600 67390 -118590
rect 67770 -118540 68890 -118530
rect 67770 -118590 67780 -118540
rect 68880 -118590 68890 -118540
rect 67770 -118600 68890 -118590
rect 69270 -118540 70390 -118530
rect 69270 -118590 69280 -118540
rect 70380 -118590 70390 -118540
rect 69270 -118600 70390 -118590
rect 70770 -118540 71890 -118530
rect 70770 -118590 70780 -118540
rect 71880 -118590 71890 -118540
rect 70770 -118600 71890 -118590
rect 72270 -118540 73390 -118530
rect 72270 -118590 72280 -118540
rect 73380 -118590 73390 -118540
rect 72270 -118600 73390 -118590
rect 73770 -118540 74890 -118530
rect 73770 -118590 73780 -118540
rect 74880 -118590 74890 -118540
rect 73770 -118600 74890 -118590
rect 75270 -118540 76390 -118530
rect 75270 -118590 75280 -118540
rect 76380 -118590 76390 -118540
rect 75270 -118600 76390 -118590
rect 76770 -118540 77890 -118530
rect 76770 -118590 76780 -118540
rect 77880 -118590 77890 -118540
rect 76770 -118600 77890 -118590
rect 78270 -118540 79390 -118530
rect 78270 -118590 78280 -118540
rect 79380 -118590 79390 -118540
rect 78270 -118600 79390 -118590
rect 79770 -118540 80890 -118530
rect 79770 -118590 79780 -118540
rect 80880 -118590 80890 -118540
rect 79770 -118600 80890 -118590
rect 81270 -118540 82390 -118530
rect 81270 -118590 81280 -118540
rect 82380 -118590 82390 -118540
rect 81270 -118600 82390 -118590
rect 82770 -118540 83890 -118530
rect 82770 -118590 82780 -118540
rect 83880 -118590 83890 -118540
rect 82770 -118600 83890 -118590
rect 84270 -118540 85390 -118530
rect 84270 -118590 84280 -118540
rect 85380 -118590 85390 -118540
rect 84270 -118600 85390 -118590
rect 85770 -118540 86890 -118530
rect 85770 -118590 85780 -118540
rect 86880 -118590 86890 -118540
rect 85770 -118600 86890 -118590
rect 87270 -118540 88390 -118530
rect 87270 -118590 87280 -118540
rect 88380 -118590 88390 -118540
rect 87270 -118600 88390 -118590
rect 88770 -118540 89890 -118530
rect 88770 -118590 88780 -118540
rect 89880 -118590 89890 -118540
rect 88770 -118600 89890 -118590
rect 90270 -118540 91390 -118530
rect 90270 -118590 90280 -118540
rect 91380 -118590 91390 -118540
rect 90270 -118600 91390 -118590
rect 91770 -118540 92890 -118530
rect 91770 -118590 91780 -118540
rect 92880 -118590 92890 -118540
rect 91770 -118600 92890 -118590
rect 93270 -118540 94390 -118530
rect 93270 -118590 93280 -118540
rect 94380 -118590 94390 -118540
rect 93270 -118600 94390 -118590
rect 94770 -118540 95890 -118530
rect 94770 -118590 94780 -118540
rect 95880 -118590 95890 -118540
rect 94770 -118600 95890 -118590
rect 96270 -118540 97390 -118530
rect 96270 -118590 96280 -118540
rect 97380 -118590 97390 -118540
rect 96270 -118600 97390 -118590
rect 97770 -118540 98890 -118530
rect 97770 -118590 97780 -118540
rect 98880 -118590 98890 -118540
rect 97770 -118600 98890 -118590
rect 99270 -118540 100390 -118530
rect 99270 -118590 99280 -118540
rect 100380 -118590 100390 -118540
rect 99270 -118600 100390 -118590
rect 100770 -118540 101890 -118530
rect 100770 -118590 100780 -118540
rect 101880 -118590 101890 -118540
rect 100770 -118600 101890 -118590
rect 102270 -118540 103390 -118530
rect 102270 -118590 102280 -118540
rect 103380 -118590 103390 -118540
rect 102270 -118600 103390 -118590
rect 103770 -118540 104890 -118530
rect 103770 -118590 103780 -118540
rect 104880 -118590 104890 -118540
rect 103770 -118600 104890 -118590
rect 105270 -118540 106390 -118530
rect 105270 -118590 105280 -118540
rect 106380 -118590 106390 -118540
rect 105270 -118600 106390 -118590
rect 106770 -118540 107890 -118530
rect 106770 -118590 106780 -118540
rect 107880 -118590 107890 -118540
rect 106770 -118600 107890 -118590
rect 108270 -118540 109390 -118530
rect 108270 -118590 108280 -118540
rect 109380 -118590 109390 -118540
rect 108270 -118600 109390 -118590
rect 109770 -118540 110890 -118530
rect 109770 -118590 109780 -118540
rect 110880 -118590 110890 -118540
rect 109770 -118600 110890 -118590
rect 111270 -118540 112390 -118530
rect 111270 -118590 111280 -118540
rect 112380 -118590 112390 -118540
rect 111270 -118600 112390 -118590
rect 112770 -118540 113890 -118530
rect 112770 -118590 112780 -118540
rect 113880 -118590 113890 -118540
rect 112770 -118600 113890 -118590
rect 114270 -118540 115390 -118530
rect 114270 -118590 114280 -118540
rect 115380 -118590 115390 -118540
rect 114270 -118600 115390 -118590
rect 115770 -118540 116890 -118530
rect 115770 -118590 115780 -118540
rect 116880 -118590 116890 -118540
rect 115770 -118600 116890 -118590
rect 117270 -118540 118390 -118530
rect 117270 -118590 117280 -118540
rect 118380 -118590 118390 -118540
rect 117270 -118600 118390 -118590
rect 118770 -118540 119890 -118530
rect 118770 -118590 118780 -118540
rect 119880 -118590 119890 -118540
rect 118770 -118600 119890 -118590
rect 110 -118750 220 -118745
rect 110 -118850 120 -118750
rect 210 -118850 220 -118750
rect 110 -119050 220 -118850
rect 1610 -118750 1720 -118745
rect 1610 -118850 1620 -118750
rect 1710 -118850 1720 -118750
rect 1610 -119050 1720 -118850
rect 3110 -118750 3220 -118745
rect 3110 -118850 3120 -118750
rect 3210 -118850 3220 -118750
rect 3110 -119050 3220 -118850
rect 4610 -118750 4720 -118745
rect 4610 -118850 4620 -118750
rect 4710 -118850 4720 -118750
rect 4610 -119050 4720 -118850
rect 6110 -118750 6220 -118745
rect 6110 -118850 6120 -118750
rect 6210 -118850 6220 -118750
rect 6110 -119050 6220 -118850
rect 7610 -118750 7720 -118745
rect 7610 -118850 7620 -118750
rect 7710 -118850 7720 -118750
rect 7610 -119050 7720 -118850
rect 9110 -118750 9220 -118745
rect 9110 -118850 9120 -118750
rect 9210 -118850 9220 -118750
rect 9110 -119050 9220 -118850
rect 10610 -118750 10720 -118745
rect 10610 -118850 10620 -118750
rect 10710 -118850 10720 -118750
rect 10610 -119050 10720 -118850
rect 12110 -118750 12220 -118745
rect 12110 -118850 12120 -118750
rect 12210 -118850 12220 -118750
rect 12110 -119050 12220 -118850
rect 13610 -118750 13720 -118745
rect 13610 -118850 13620 -118750
rect 13710 -118850 13720 -118750
rect 13610 -119050 13720 -118850
rect 15110 -118750 15220 -118745
rect 15110 -118850 15120 -118750
rect 15210 -118850 15220 -118750
rect 15110 -119050 15220 -118850
rect 16610 -118750 16720 -118745
rect 16610 -118850 16620 -118750
rect 16710 -118850 16720 -118750
rect 16610 -119050 16720 -118850
rect 18110 -118750 18220 -118745
rect 18110 -118850 18120 -118750
rect 18210 -118850 18220 -118750
rect 18110 -119050 18220 -118850
rect 19610 -118750 19720 -118745
rect 19610 -118850 19620 -118750
rect 19710 -118850 19720 -118750
rect 19610 -119050 19720 -118850
rect 21110 -118750 21220 -118745
rect 21110 -118850 21120 -118750
rect 21210 -118850 21220 -118750
rect 21110 -119050 21220 -118850
rect 22610 -118750 22720 -118745
rect 22610 -118850 22620 -118750
rect 22710 -118850 22720 -118750
rect 22610 -119050 22720 -118850
rect 24110 -118750 24220 -118745
rect 24110 -118850 24120 -118750
rect 24210 -118850 24220 -118750
rect 24110 -119050 24220 -118850
rect 25610 -118750 25720 -118745
rect 25610 -118850 25620 -118750
rect 25710 -118850 25720 -118750
rect 25610 -119050 25720 -118850
rect 27110 -118750 27220 -118745
rect 27110 -118850 27120 -118750
rect 27210 -118850 27220 -118750
rect 27110 -119050 27220 -118850
rect 28610 -118750 28720 -118745
rect 28610 -118850 28620 -118750
rect 28710 -118850 28720 -118750
rect 28610 -119050 28720 -118850
rect 30110 -118750 30220 -118745
rect 30110 -118850 30120 -118750
rect 30210 -118850 30220 -118750
rect 30110 -119050 30220 -118850
rect 31610 -118750 31720 -118745
rect 31610 -118850 31620 -118750
rect 31710 -118850 31720 -118750
rect 31610 -119050 31720 -118850
rect 33110 -118750 33220 -118745
rect 33110 -118850 33120 -118750
rect 33210 -118850 33220 -118750
rect 33110 -119050 33220 -118850
rect 34610 -118750 34720 -118745
rect 34610 -118850 34620 -118750
rect 34710 -118850 34720 -118750
rect 34610 -119050 34720 -118850
rect 36110 -118750 36220 -118745
rect 36110 -118850 36120 -118750
rect 36210 -118850 36220 -118750
rect 36110 -119050 36220 -118850
rect 37610 -118750 37720 -118745
rect 37610 -118850 37620 -118750
rect 37710 -118850 37720 -118750
rect 37610 -119050 37720 -118850
rect 39110 -118750 39220 -118745
rect 39110 -118850 39120 -118750
rect 39210 -118850 39220 -118750
rect 39110 -119050 39220 -118850
rect 40610 -118750 40720 -118745
rect 40610 -118850 40620 -118750
rect 40710 -118850 40720 -118750
rect 40610 -119050 40720 -118850
rect 42110 -118750 42220 -118745
rect 42110 -118850 42120 -118750
rect 42210 -118850 42220 -118750
rect 42110 -119050 42220 -118850
rect 43610 -118750 43720 -118745
rect 43610 -118850 43620 -118750
rect 43710 -118850 43720 -118750
rect 43610 -119050 43720 -118850
rect 45110 -118750 45220 -118745
rect 45110 -118850 45120 -118750
rect 45210 -118850 45220 -118750
rect 45110 -119050 45220 -118850
rect 46610 -118750 46720 -118745
rect 46610 -118850 46620 -118750
rect 46710 -118850 46720 -118750
rect 46610 -119050 46720 -118850
rect 48110 -118750 48220 -118745
rect 48110 -118850 48120 -118750
rect 48210 -118850 48220 -118750
rect 48110 -119050 48220 -118850
rect 49610 -118750 49720 -118745
rect 49610 -118850 49620 -118750
rect 49710 -118850 49720 -118750
rect 49610 -119050 49720 -118850
rect 51110 -118750 51220 -118745
rect 51110 -118850 51120 -118750
rect 51210 -118850 51220 -118750
rect 51110 -119050 51220 -118850
rect 52610 -118750 52720 -118745
rect 52610 -118850 52620 -118750
rect 52710 -118850 52720 -118750
rect 52610 -119050 52720 -118850
rect 54110 -118750 54220 -118745
rect 54110 -118850 54120 -118750
rect 54210 -118850 54220 -118750
rect 54110 -119050 54220 -118850
rect 55610 -118750 55720 -118745
rect 55610 -118850 55620 -118750
rect 55710 -118850 55720 -118750
rect 55610 -119050 55720 -118850
rect 57110 -118750 57220 -118745
rect 57110 -118850 57120 -118750
rect 57210 -118850 57220 -118750
rect 57110 -119050 57220 -118850
rect 58610 -118750 58720 -118745
rect 58610 -118850 58620 -118750
rect 58710 -118850 58720 -118750
rect 58610 -119050 58720 -118850
rect 60110 -118750 60220 -118745
rect 60110 -118850 60120 -118750
rect 60210 -118850 60220 -118750
rect 60110 -119050 60220 -118850
rect 61610 -118750 61720 -118745
rect 61610 -118850 61620 -118750
rect 61710 -118850 61720 -118750
rect 61610 -119050 61720 -118850
rect 63110 -118750 63220 -118745
rect 63110 -118850 63120 -118750
rect 63210 -118850 63220 -118750
rect 63110 -119050 63220 -118850
rect 64610 -118750 64720 -118745
rect 64610 -118850 64620 -118750
rect 64710 -118850 64720 -118750
rect 64610 -119050 64720 -118850
rect 66110 -118750 66220 -118745
rect 66110 -118850 66120 -118750
rect 66210 -118850 66220 -118750
rect 66110 -119050 66220 -118850
rect 67610 -118750 67720 -118745
rect 67610 -118850 67620 -118750
rect 67710 -118850 67720 -118750
rect 67610 -119050 67720 -118850
rect 69110 -118750 69220 -118745
rect 69110 -118850 69120 -118750
rect 69210 -118850 69220 -118750
rect 69110 -119050 69220 -118850
rect 70610 -118750 70720 -118745
rect 70610 -118850 70620 -118750
rect 70710 -118850 70720 -118750
rect 70610 -119050 70720 -118850
rect 72110 -118750 72220 -118745
rect 72110 -118850 72120 -118750
rect 72210 -118850 72220 -118750
rect 72110 -119050 72220 -118850
rect 73610 -118750 73720 -118745
rect 73610 -118850 73620 -118750
rect 73710 -118850 73720 -118750
rect 73610 -119050 73720 -118850
rect 75110 -118750 75220 -118745
rect 75110 -118850 75120 -118750
rect 75210 -118850 75220 -118750
rect 75110 -119050 75220 -118850
rect 76610 -118750 76720 -118745
rect 76610 -118850 76620 -118750
rect 76710 -118850 76720 -118750
rect 76610 -119050 76720 -118850
rect 78110 -118750 78220 -118745
rect 78110 -118850 78120 -118750
rect 78210 -118850 78220 -118750
rect 78110 -119050 78220 -118850
rect 79610 -118750 79720 -118745
rect 79610 -118850 79620 -118750
rect 79710 -118850 79720 -118750
rect 79610 -119050 79720 -118850
rect 81110 -118750 81220 -118745
rect 81110 -118850 81120 -118750
rect 81210 -118850 81220 -118750
rect 81110 -119050 81220 -118850
rect 82610 -118750 82720 -118745
rect 82610 -118850 82620 -118750
rect 82710 -118850 82720 -118750
rect 82610 -119050 82720 -118850
rect 84110 -118750 84220 -118745
rect 84110 -118850 84120 -118750
rect 84210 -118850 84220 -118750
rect 84110 -119050 84220 -118850
rect 85610 -118750 85720 -118745
rect 85610 -118850 85620 -118750
rect 85710 -118850 85720 -118750
rect 85610 -119050 85720 -118850
rect 87110 -118750 87220 -118745
rect 87110 -118850 87120 -118750
rect 87210 -118850 87220 -118750
rect 87110 -119050 87220 -118850
rect 88610 -118750 88720 -118745
rect 88610 -118850 88620 -118750
rect 88710 -118850 88720 -118750
rect 88610 -119050 88720 -118850
rect 90110 -118750 90220 -118745
rect 90110 -118850 90120 -118750
rect 90210 -118850 90220 -118750
rect 90110 -119050 90220 -118850
rect 91610 -118750 91720 -118745
rect 91610 -118850 91620 -118750
rect 91710 -118850 91720 -118750
rect 91610 -119050 91720 -118850
rect 93110 -118750 93220 -118745
rect 93110 -118850 93120 -118750
rect 93210 -118850 93220 -118750
rect 93110 -119050 93220 -118850
rect 94610 -118750 94720 -118745
rect 94610 -118850 94620 -118750
rect 94710 -118850 94720 -118750
rect 94610 -119050 94720 -118850
rect 96110 -118750 96220 -118745
rect 96110 -118850 96120 -118750
rect 96210 -118850 96220 -118750
rect 96110 -119050 96220 -118850
rect 97610 -118750 97720 -118745
rect 97610 -118850 97620 -118750
rect 97710 -118850 97720 -118750
rect 97610 -119050 97720 -118850
rect 99110 -118750 99220 -118745
rect 99110 -118850 99120 -118750
rect 99210 -118850 99220 -118750
rect 99110 -119050 99220 -118850
rect 100610 -118750 100720 -118745
rect 100610 -118850 100620 -118750
rect 100710 -118850 100720 -118750
rect 100610 -119050 100720 -118850
rect 102110 -118750 102220 -118745
rect 102110 -118850 102120 -118750
rect 102210 -118850 102220 -118750
rect 102110 -119050 102220 -118850
rect 103610 -118750 103720 -118745
rect 103610 -118850 103620 -118750
rect 103710 -118850 103720 -118750
rect 103610 -119050 103720 -118850
rect 105110 -118750 105220 -118745
rect 105110 -118850 105120 -118750
rect 105210 -118850 105220 -118750
rect 105110 -119050 105220 -118850
rect 106610 -118750 106720 -118745
rect 106610 -118850 106620 -118750
rect 106710 -118850 106720 -118750
rect 106610 -119050 106720 -118850
rect 108110 -118750 108220 -118745
rect 108110 -118850 108120 -118750
rect 108210 -118850 108220 -118750
rect 108110 -119050 108220 -118850
rect 109610 -118750 109720 -118745
rect 109610 -118850 109620 -118750
rect 109710 -118850 109720 -118750
rect 109610 -119050 109720 -118850
rect 111110 -118750 111220 -118745
rect 111110 -118850 111120 -118750
rect 111210 -118850 111220 -118750
rect 111110 -119050 111220 -118850
rect 112610 -118750 112720 -118745
rect 112610 -118850 112620 -118750
rect 112710 -118850 112720 -118750
rect 112610 -119050 112720 -118850
rect 114110 -118750 114220 -118745
rect 114110 -118850 114120 -118750
rect 114210 -118850 114220 -118750
rect 114110 -119050 114220 -118850
rect 115610 -118750 115720 -118745
rect 115610 -118850 115620 -118750
rect 115710 -118850 115720 -118750
rect 115610 -119050 115720 -118850
rect 117110 -118750 117220 -118745
rect 117110 -118850 117120 -118750
rect 117210 -118850 117220 -118750
rect 117110 -119050 117220 -118850
rect 118610 -118750 118720 -118745
rect 118610 -118850 118620 -118750
rect 118710 -118850 118720 -118750
rect 118610 -119050 118720 -118850
<< metal5 >>
rect -1000 1420 0 1580
rect 520 520 620 620
rect 2020 520 2120 620
rect 3520 520 3620 620
rect 5020 520 5120 620
rect 6520 520 6620 620
rect 8020 520 8120 620
rect 9520 520 9620 620
rect 11020 520 11120 620
rect 12520 520 12620 620
rect 14020 520 14120 620
rect 15520 520 15620 620
rect 17020 520 17120 620
rect 18520 520 18620 620
rect 20020 520 20120 620
rect 21520 520 21620 620
rect 23020 520 23120 620
rect 24520 520 24620 620
rect 26020 520 26120 620
rect 27520 520 27620 620
rect 29020 520 29120 620
rect 30520 520 30620 620
rect 32020 520 32120 620
rect 33520 520 33620 620
rect 35020 520 35120 620
rect 36520 520 36620 620
rect 38020 520 38120 620
rect 39520 520 39620 620
rect 41020 520 41120 620
rect 42520 520 42620 620
rect 44020 520 44120 620
rect 45520 520 45620 620
rect 47020 520 47120 620
rect 48520 520 48620 620
rect 50020 520 50120 620
rect 51520 520 51620 620
rect 53020 520 53120 620
rect 54520 520 54620 620
rect 56020 520 56120 620
rect 57520 520 57620 620
rect 59020 520 59120 620
rect 60520 520 60620 620
rect 62020 520 62120 620
rect 63520 520 63620 620
rect 65020 520 65120 620
rect 66520 520 66620 620
rect 68020 520 68120 620
rect 69520 520 69620 620
rect 71020 520 71120 620
rect 72520 520 72620 620
rect 74020 520 74120 620
rect 75520 520 75620 620
rect 77020 520 77120 620
rect 78520 520 78620 620
rect 80020 520 80120 620
rect 81520 520 81620 620
rect 83020 520 83120 620
rect 84520 520 84620 620
rect 86020 520 86120 620
rect 87520 520 87620 620
rect 89020 520 89120 620
rect 90520 520 90620 620
rect 92020 520 92120 620
rect 93520 520 93620 620
rect 95020 520 95120 620
rect 96520 520 96620 620
rect 98020 520 98120 620
rect 99520 520 99620 620
rect 101020 520 101120 620
rect 102520 520 102620 620
rect 104020 520 104120 620
rect 105520 520 105620 620
rect 107020 520 107120 620
rect 108520 520 108620 620
rect 110020 520 110120 620
rect 111520 520 111620 620
rect 113020 520 113120 620
rect 114520 520 114620 620
rect 116020 520 116120 620
rect 117520 520 117620 620
rect 119020 520 119120 620
rect 520 -980 620 -880
rect 2020 -980 2120 -880
rect 3520 -980 3620 -880
rect 5020 -980 5120 -880
rect 6520 -980 6620 -880
rect 8020 -980 8120 -880
rect 9520 -980 9620 -880
rect 11020 -980 11120 -880
rect 12520 -980 12620 -880
rect 14020 -980 14120 -880
rect 15520 -980 15620 -880
rect 17020 -980 17120 -880
rect 18520 -980 18620 -880
rect 20020 -980 20120 -880
rect 21520 -980 21620 -880
rect 23020 -980 23120 -880
rect 24520 -980 24620 -880
rect 26020 -980 26120 -880
rect 27520 -980 27620 -880
rect 29020 -980 29120 -880
rect 30520 -980 30620 -880
rect 32020 -980 32120 -880
rect 33520 -980 33620 -880
rect 35020 -980 35120 -880
rect 36520 -980 36620 -880
rect 38020 -980 38120 -880
rect 39520 -980 39620 -880
rect 41020 -980 41120 -880
rect 42520 -980 42620 -880
rect 44020 -980 44120 -880
rect 45520 -980 45620 -880
rect 47020 -980 47120 -880
rect 48520 -980 48620 -880
rect 50020 -980 50120 -880
rect 51520 -980 51620 -880
rect 53020 -980 53120 -880
rect 54520 -980 54620 -880
rect 56020 -980 56120 -880
rect 57520 -980 57620 -880
rect 59020 -980 59120 -880
rect 60520 -980 60620 -880
rect 62020 -980 62120 -880
rect 63520 -980 63620 -880
rect 65020 -980 65120 -880
rect 66520 -980 66620 -880
rect 68020 -980 68120 -880
rect 69520 -980 69620 -880
rect 71020 -980 71120 -880
rect 72520 -980 72620 -880
rect 74020 -980 74120 -880
rect 75520 -980 75620 -880
rect 77020 -980 77120 -880
rect 78520 -980 78620 -880
rect 80020 -980 80120 -880
rect 81520 -980 81620 -880
rect 83020 -980 83120 -880
rect 84520 -980 84620 -880
rect 86020 -980 86120 -880
rect 87520 -980 87620 -880
rect 89020 -980 89120 -880
rect 90520 -980 90620 -880
rect 92020 -980 92120 -880
rect 93520 -980 93620 -880
rect 95020 -980 95120 -880
rect 96520 -980 96620 -880
rect 98020 -980 98120 -880
rect 99520 -980 99620 -880
rect 101020 -980 101120 -880
rect 102520 -980 102620 -880
rect 104020 -980 104120 -880
rect 105520 -980 105620 -880
rect 107020 -980 107120 -880
rect 108520 -980 108620 -880
rect 110020 -980 110120 -880
rect 111520 -980 111620 -880
rect 113020 -980 113120 -880
rect 114520 -980 114620 -880
rect 116020 -980 116120 -880
rect 117520 -980 117620 -880
rect 119020 -980 119120 -880
rect 520 -2480 620 -2380
rect 2020 -2480 2120 -2380
rect 3520 -2480 3620 -2380
rect 5020 -2480 5120 -2380
rect 6520 -2480 6620 -2380
rect 8020 -2480 8120 -2380
rect 9520 -2480 9620 -2380
rect 11020 -2480 11120 -2380
rect 12520 -2480 12620 -2380
rect 14020 -2480 14120 -2380
rect 15520 -2480 15620 -2380
rect 17020 -2480 17120 -2380
rect 18520 -2480 18620 -2380
rect 20020 -2480 20120 -2380
rect 21520 -2480 21620 -2380
rect 23020 -2480 23120 -2380
rect 24520 -2480 24620 -2380
rect 26020 -2480 26120 -2380
rect 27520 -2480 27620 -2380
rect 29020 -2480 29120 -2380
rect 30520 -2480 30620 -2380
rect 32020 -2480 32120 -2380
rect 33520 -2480 33620 -2380
rect 35020 -2480 35120 -2380
rect 36520 -2480 36620 -2380
rect 38020 -2480 38120 -2380
rect 39520 -2480 39620 -2380
rect 41020 -2480 41120 -2380
rect 42520 -2480 42620 -2380
rect 44020 -2480 44120 -2380
rect 45520 -2480 45620 -2380
rect 47020 -2480 47120 -2380
rect 48520 -2480 48620 -2380
rect 50020 -2480 50120 -2380
rect 51520 -2480 51620 -2380
rect 53020 -2480 53120 -2380
rect 54520 -2480 54620 -2380
rect 56020 -2480 56120 -2380
rect 57520 -2480 57620 -2380
rect 59020 -2480 59120 -2380
rect 60520 -2480 60620 -2380
rect 62020 -2480 62120 -2380
rect 63520 -2480 63620 -2380
rect 65020 -2480 65120 -2380
rect 66520 -2480 66620 -2380
rect 68020 -2480 68120 -2380
rect 69520 -2480 69620 -2380
rect 71020 -2480 71120 -2380
rect 72520 -2480 72620 -2380
rect 74020 -2480 74120 -2380
rect 75520 -2480 75620 -2380
rect 77020 -2480 77120 -2380
rect 78520 -2480 78620 -2380
rect 80020 -2480 80120 -2380
rect 81520 -2480 81620 -2380
rect 83020 -2480 83120 -2380
rect 84520 -2480 84620 -2380
rect 86020 -2480 86120 -2380
rect 87520 -2480 87620 -2380
rect 89020 -2480 89120 -2380
rect 90520 -2480 90620 -2380
rect 92020 -2480 92120 -2380
rect 93520 -2480 93620 -2380
rect 95020 -2480 95120 -2380
rect 96520 -2480 96620 -2380
rect 98020 -2480 98120 -2380
rect 99520 -2480 99620 -2380
rect 101020 -2480 101120 -2380
rect 102520 -2480 102620 -2380
rect 104020 -2480 104120 -2380
rect 105520 -2480 105620 -2380
rect 107020 -2480 107120 -2380
rect 108520 -2480 108620 -2380
rect 110020 -2480 110120 -2380
rect 111520 -2480 111620 -2380
rect 113020 -2480 113120 -2380
rect 114520 -2480 114620 -2380
rect 116020 -2480 116120 -2380
rect 117520 -2480 117620 -2380
rect 119020 -2480 119120 -2380
rect 520 -3980 620 -3880
rect 2020 -3980 2120 -3880
rect 3520 -3980 3620 -3880
rect 5020 -3980 5120 -3880
rect 6520 -3980 6620 -3880
rect 8020 -3980 8120 -3880
rect 9520 -3980 9620 -3880
rect 11020 -3980 11120 -3880
rect 12520 -3980 12620 -3880
rect 14020 -3980 14120 -3880
rect 15520 -3980 15620 -3880
rect 17020 -3980 17120 -3880
rect 18520 -3980 18620 -3880
rect 20020 -3980 20120 -3880
rect 21520 -3980 21620 -3880
rect 23020 -3980 23120 -3880
rect 24520 -3980 24620 -3880
rect 26020 -3980 26120 -3880
rect 27520 -3980 27620 -3880
rect 29020 -3980 29120 -3880
rect 30520 -3980 30620 -3880
rect 32020 -3980 32120 -3880
rect 33520 -3980 33620 -3880
rect 35020 -3980 35120 -3880
rect 36520 -3980 36620 -3880
rect 38020 -3980 38120 -3880
rect 39520 -3980 39620 -3880
rect 41020 -3980 41120 -3880
rect 42520 -3980 42620 -3880
rect 44020 -3980 44120 -3880
rect 45520 -3980 45620 -3880
rect 47020 -3980 47120 -3880
rect 48520 -3980 48620 -3880
rect 50020 -3980 50120 -3880
rect 51520 -3980 51620 -3880
rect 53020 -3980 53120 -3880
rect 54520 -3980 54620 -3880
rect 56020 -3980 56120 -3880
rect 57520 -3980 57620 -3880
rect 59020 -3980 59120 -3880
rect 60520 -3980 60620 -3880
rect 62020 -3980 62120 -3880
rect 63520 -3980 63620 -3880
rect 65020 -3980 65120 -3880
rect 66520 -3980 66620 -3880
rect 68020 -3980 68120 -3880
rect 69520 -3980 69620 -3880
rect 71020 -3980 71120 -3880
rect 72520 -3980 72620 -3880
rect 74020 -3980 74120 -3880
rect 75520 -3980 75620 -3880
rect 77020 -3980 77120 -3880
rect 78520 -3980 78620 -3880
rect 80020 -3980 80120 -3880
rect 81520 -3980 81620 -3880
rect 83020 -3980 83120 -3880
rect 84520 -3980 84620 -3880
rect 86020 -3980 86120 -3880
rect 87520 -3980 87620 -3880
rect 89020 -3980 89120 -3880
rect 90520 -3980 90620 -3880
rect 92020 -3980 92120 -3880
rect 93520 -3980 93620 -3880
rect 95020 -3980 95120 -3880
rect 96520 -3980 96620 -3880
rect 98020 -3980 98120 -3880
rect 99520 -3980 99620 -3880
rect 101020 -3980 101120 -3880
rect 102520 -3980 102620 -3880
rect 104020 -3980 104120 -3880
rect 105520 -3980 105620 -3880
rect 107020 -3980 107120 -3880
rect 108520 -3980 108620 -3880
rect 110020 -3980 110120 -3880
rect 111520 -3980 111620 -3880
rect 113020 -3980 113120 -3880
rect 114520 -3980 114620 -3880
rect 116020 -3980 116120 -3880
rect 117520 -3980 117620 -3880
rect 119020 -3980 119120 -3880
rect 520 -5480 620 -5380
rect 2020 -5480 2120 -5380
rect 3520 -5480 3620 -5380
rect 5020 -5480 5120 -5380
rect 6520 -5480 6620 -5380
rect 8020 -5480 8120 -5380
rect 9520 -5480 9620 -5380
rect 11020 -5480 11120 -5380
rect 12520 -5480 12620 -5380
rect 14020 -5480 14120 -5380
rect 15520 -5480 15620 -5380
rect 17020 -5480 17120 -5380
rect 18520 -5480 18620 -5380
rect 20020 -5480 20120 -5380
rect 21520 -5480 21620 -5380
rect 23020 -5480 23120 -5380
rect 24520 -5480 24620 -5380
rect 26020 -5480 26120 -5380
rect 27520 -5480 27620 -5380
rect 29020 -5480 29120 -5380
rect 30520 -5480 30620 -5380
rect 32020 -5480 32120 -5380
rect 33520 -5480 33620 -5380
rect 35020 -5480 35120 -5380
rect 36520 -5480 36620 -5380
rect 38020 -5480 38120 -5380
rect 39520 -5480 39620 -5380
rect 41020 -5480 41120 -5380
rect 42520 -5480 42620 -5380
rect 44020 -5480 44120 -5380
rect 45520 -5480 45620 -5380
rect 47020 -5480 47120 -5380
rect 48520 -5480 48620 -5380
rect 50020 -5480 50120 -5380
rect 51520 -5480 51620 -5380
rect 53020 -5480 53120 -5380
rect 54520 -5480 54620 -5380
rect 56020 -5480 56120 -5380
rect 57520 -5480 57620 -5380
rect 59020 -5480 59120 -5380
rect 60520 -5480 60620 -5380
rect 62020 -5480 62120 -5380
rect 63520 -5480 63620 -5380
rect 65020 -5480 65120 -5380
rect 66520 -5480 66620 -5380
rect 68020 -5480 68120 -5380
rect 69520 -5480 69620 -5380
rect 71020 -5480 71120 -5380
rect 72520 -5480 72620 -5380
rect 74020 -5480 74120 -5380
rect 75520 -5480 75620 -5380
rect 77020 -5480 77120 -5380
rect 78520 -5480 78620 -5380
rect 80020 -5480 80120 -5380
rect 81520 -5480 81620 -5380
rect 83020 -5480 83120 -5380
rect 84520 -5480 84620 -5380
rect 86020 -5480 86120 -5380
rect 87520 -5480 87620 -5380
rect 89020 -5480 89120 -5380
rect 90520 -5480 90620 -5380
rect 92020 -5480 92120 -5380
rect 93520 -5480 93620 -5380
rect 95020 -5480 95120 -5380
rect 96520 -5480 96620 -5380
rect 98020 -5480 98120 -5380
rect 99520 -5480 99620 -5380
rect 101020 -5480 101120 -5380
rect 102520 -5480 102620 -5380
rect 104020 -5480 104120 -5380
rect 105520 -5480 105620 -5380
rect 107020 -5480 107120 -5380
rect 108520 -5480 108620 -5380
rect 110020 -5480 110120 -5380
rect 111520 -5480 111620 -5380
rect 113020 -5480 113120 -5380
rect 114520 -5480 114620 -5380
rect 116020 -5480 116120 -5380
rect 117520 -5480 117620 -5380
rect 119020 -5480 119120 -5380
rect 520 -6980 620 -6880
rect 2020 -6980 2120 -6880
rect 3520 -6980 3620 -6880
rect 5020 -6980 5120 -6880
rect 6520 -6980 6620 -6880
rect 8020 -6980 8120 -6880
rect 9520 -6980 9620 -6880
rect 11020 -6980 11120 -6880
rect 12520 -6980 12620 -6880
rect 14020 -6980 14120 -6880
rect 15520 -6980 15620 -6880
rect 17020 -6980 17120 -6880
rect 18520 -6980 18620 -6880
rect 20020 -6980 20120 -6880
rect 21520 -6980 21620 -6880
rect 23020 -6980 23120 -6880
rect 24520 -6980 24620 -6880
rect 26020 -6980 26120 -6880
rect 27520 -6980 27620 -6880
rect 29020 -6980 29120 -6880
rect 30520 -6980 30620 -6880
rect 32020 -6980 32120 -6880
rect 33520 -6980 33620 -6880
rect 35020 -6980 35120 -6880
rect 36520 -6980 36620 -6880
rect 38020 -6980 38120 -6880
rect 39520 -6980 39620 -6880
rect 41020 -6980 41120 -6880
rect 42520 -6980 42620 -6880
rect 44020 -6980 44120 -6880
rect 45520 -6980 45620 -6880
rect 47020 -6980 47120 -6880
rect 48520 -6980 48620 -6880
rect 50020 -6980 50120 -6880
rect 51520 -6980 51620 -6880
rect 53020 -6980 53120 -6880
rect 54520 -6980 54620 -6880
rect 56020 -6980 56120 -6880
rect 57520 -6980 57620 -6880
rect 59020 -6980 59120 -6880
rect 60520 -6980 60620 -6880
rect 62020 -6980 62120 -6880
rect 63520 -6980 63620 -6880
rect 65020 -6980 65120 -6880
rect 66520 -6980 66620 -6880
rect 68020 -6980 68120 -6880
rect 69520 -6980 69620 -6880
rect 71020 -6980 71120 -6880
rect 72520 -6980 72620 -6880
rect 74020 -6980 74120 -6880
rect 75520 -6980 75620 -6880
rect 77020 -6980 77120 -6880
rect 78520 -6980 78620 -6880
rect 80020 -6980 80120 -6880
rect 81520 -6980 81620 -6880
rect 83020 -6980 83120 -6880
rect 84520 -6980 84620 -6880
rect 86020 -6980 86120 -6880
rect 87520 -6980 87620 -6880
rect 89020 -6980 89120 -6880
rect 90520 -6980 90620 -6880
rect 92020 -6980 92120 -6880
rect 93520 -6980 93620 -6880
rect 95020 -6980 95120 -6880
rect 96520 -6980 96620 -6880
rect 98020 -6980 98120 -6880
rect 99520 -6980 99620 -6880
rect 101020 -6980 101120 -6880
rect 102520 -6980 102620 -6880
rect 104020 -6980 104120 -6880
rect 105520 -6980 105620 -6880
rect 107020 -6980 107120 -6880
rect 108520 -6980 108620 -6880
rect 110020 -6980 110120 -6880
rect 111520 -6980 111620 -6880
rect 113020 -6980 113120 -6880
rect 114520 -6980 114620 -6880
rect 116020 -6980 116120 -6880
rect 117520 -6980 117620 -6880
rect 119020 -6980 119120 -6880
rect 520 -8480 620 -8380
rect 2020 -8480 2120 -8380
rect 3520 -8480 3620 -8380
rect 5020 -8480 5120 -8380
rect 6520 -8480 6620 -8380
rect 8020 -8480 8120 -8380
rect 9520 -8480 9620 -8380
rect 11020 -8480 11120 -8380
rect 12520 -8480 12620 -8380
rect 14020 -8480 14120 -8380
rect 15520 -8480 15620 -8380
rect 17020 -8480 17120 -8380
rect 18520 -8480 18620 -8380
rect 20020 -8480 20120 -8380
rect 21520 -8480 21620 -8380
rect 23020 -8480 23120 -8380
rect 24520 -8480 24620 -8380
rect 26020 -8480 26120 -8380
rect 27520 -8480 27620 -8380
rect 29020 -8480 29120 -8380
rect 30520 -8480 30620 -8380
rect 32020 -8480 32120 -8380
rect 33520 -8480 33620 -8380
rect 35020 -8480 35120 -8380
rect 36520 -8480 36620 -8380
rect 38020 -8480 38120 -8380
rect 39520 -8480 39620 -8380
rect 41020 -8480 41120 -8380
rect 42520 -8480 42620 -8380
rect 44020 -8480 44120 -8380
rect 45520 -8480 45620 -8380
rect 47020 -8480 47120 -8380
rect 48520 -8480 48620 -8380
rect 50020 -8480 50120 -8380
rect 51520 -8480 51620 -8380
rect 53020 -8480 53120 -8380
rect 54520 -8480 54620 -8380
rect 56020 -8480 56120 -8380
rect 57520 -8480 57620 -8380
rect 59020 -8480 59120 -8380
rect 60520 -8480 60620 -8380
rect 62020 -8480 62120 -8380
rect 63520 -8480 63620 -8380
rect 65020 -8480 65120 -8380
rect 66520 -8480 66620 -8380
rect 68020 -8480 68120 -8380
rect 69520 -8480 69620 -8380
rect 71020 -8480 71120 -8380
rect 72520 -8480 72620 -8380
rect 74020 -8480 74120 -8380
rect 75520 -8480 75620 -8380
rect 77020 -8480 77120 -8380
rect 78520 -8480 78620 -8380
rect 80020 -8480 80120 -8380
rect 81520 -8480 81620 -8380
rect 83020 -8480 83120 -8380
rect 84520 -8480 84620 -8380
rect 86020 -8480 86120 -8380
rect 87520 -8480 87620 -8380
rect 89020 -8480 89120 -8380
rect 90520 -8480 90620 -8380
rect 92020 -8480 92120 -8380
rect 93520 -8480 93620 -8380
rect 95020 -8480 95120 -8380
rect 96520 -8480 96620 -8380
rect 98020 -8480 98120 -8380
rect 99520 -8480 99620 -8380
rect 101020 -8480 101120 -8380
rect 102520 -8480 102620 -8380
rect 104020 -8480 104120 -8380
rect 105520 -8480 105620 -8380
rect 107020 -8480 107120 -8380
rect 108520 -8480 108620 -8380
rect 110020 -8480 110120 -8380
rect 111520 -8480 111620 -8380
rect 113020 -8480 113120 -8380
rect 114520 -8480 114620 -8380
rect 116020 -8480 116120 -8380
rect 117520 -8480 117620 -8380
rect 119020 -8480 119120 -8380
rect 520 -9980 620 -9880
rect 2020 -9980 2120 -9880
rect 3520 -9980 3620 -9880
rect 5020 -9980 5120 -9880
rect 6520 -9980 6620 -9880
rect 8020 -9980 8120 -9880
rect 9520 -9980 9620 -9880
rect 11020 -9980 11120 -9880
rect 12520 -9980 12620 -9880
rect 14020 -9980 14120 -9880
rect 15520 -9980 15620 -9880
rect 17020 -9980 17120 -9880
rect 18520 -9980 18620 -9880
rect 20020 -9980 20120 -9880
rect 21520 -9980 21620 -9880
rect 23020 -9980 23120 -9880
rect 24520 -9980 24620 -9880
rect 26020 -9980 26120 -9880
rect 27520 -9980 27620 -9880
rect 29020 -9980 29120 -9880
rect 30520 -9980 30620 -9880
rect 32020 -9980 32120 -9880
rect 33520 -9980 33620 -9880
rect 35020 -9980 35120 -9880
rect 36520 -9980 36620 -9880
rect 38020 -9980 38120 -9880
rect 39520 -9980 39620 -9880
rect 41020 -9980 41120 -9880
rect 42520 -9980 42620 -9880
rect 44020 -9980 44120 -9880
rect 45520 -9980 45620 -9880
rect 47020 -9980 47120 -9880
rect 48520 -9980 48620 -9880
rect 50020 -9980 50120 -9880
rect 51520 -9980 51620 -9880
rect 53020 -9980 53120 -9880
rect 54520 -9980 54620 -9880
rect 56020 -9980 56120 -9880
rect 57520 -9980 57620 -9880
rect 59020 -9980 59120 -9880
rect 60520 -9980 60620 -9880
rect 62020 -9980 62120 -9880
rect 63520 -9980 63620 -9880
rect 65020 -9980 65120 -9880
rect 66520 -9980 66620 -9880
rect 68020 -9980 68120 -9880
rect 69520 -9980 69620 -9880
rect 71020 -9980 71120 -9880
rect 72520 -9980 72620 -9880
rect 74020 -9980 74120 -9880
rect 75520 -9980 75620 -9880
rect 77020 -9980 77120 -9880
rect 78520 -9980 78620 -9880
rect 80020 -9980 80120 -9880
rect 81520 -9980 81620 -9880
rect 83020 -9980 83120 -9880
rect 84520 -9980 84620 -9880
rect 86020 -9980 86120 -9880
rect 87520 -9980 87620 -9880
rect 89020 -9980 89120 -9880
rect 90520 -9980 90620 -9880
rect 92020 -9980 92120 -9880
rect 93520 -9980 93620 -9880
rect 95020 -9980 95120 -9880
rect 96520 -9980 96620 -9880
rect 98020 -9980 98120 -9880
rect 99520 -9980 99620 -9880
rect 101020 -9980 101120 -9880
rect 102520 -9980 102620 -9880
rect 104020 -9980 104120 -9880
rect 105520 -9980 105620 -9880
rect 107020 -9980 107120 -9880
rect 108520 -9980 108620 -9880
rect 110020 -9980 110120 -9880
rect 111520 -9980 111620 -9880
rect 113020 -9980 113120 -9880
rect 114520 -9980 114620 -9880
rect 116020 -9980 116120 -9880
rect 117520 -9980 117620 -9880
rect 119020 -9980 119120 -9880
rect 520 -11480 620 -11380
rect 2020 -11480 2120 -11380
rect 3520 -11480 3620 -11380
rect 5020 -11480 5120 -11380
rect 6520 -11480 6620 -11380
rect 8020 -11480 8120 -11380
rect 9520 -11480 9620 -11380
rect 11020 -11480 11120 -11380
rect 12520 -11480 12620 -11380
rect 14020 -11480 14120 -11380
rect 15520 -11480 15620 -11380
rect 17020 -11480 17120 -11380
rect 18520 -11480 18620 -11380
rect 20020 -11480 20120 -11380
rect 21520 -11480 21620 -11380
rect 23020 -11480 23120 -11380
rect 24520 -11480 24620 -11380
rect 26020 -11480 26120 -11380
rect 27520 -11480 27620 -11380
rect 29020 -11480 29120 -11380
rect 30520 -11480 30620 -11380
rect 32020 -11480 32120 -11380
rect 33520 -11480 33620 -11380
rect 35020 -11480 35120 -11380
rect 36520 -11480 36620 -11380
rect 38020 -11480 38120 -11380
rect 39520 -11480 39620 -11380
rect 41020 -11480 41120 -11380
rect 42520 -11480 42620 -11380
rect 44020 -11480 44120 -11380
rect 45520 -11480 45620 -11380
rect 47020 -11480 47120 -11380
rect 48520 -11480 48620 -11380
rect 50020 -11480 50120 -11380
rect 51520 -11480 51620 -11380
rect 53020 -11480 53120 -11380
rect 54520 -11480 54620 -11380
rect 56020 -11480 56120 -11380
rect 57520 -11480 57620 -11380
rect 59020 -11480 59120 -11380
rect 60520 -11480 60620 -11380
rect 62020 -11480 62120 -11380
rect 63520 -11480 63620 -11380
rect 65020 -11480 65120 -11380
rect 66520 -11480 66620 -11380
rect 68020 -11480 68120 -11380
rect 69520 -11480 69620 -11380
rect 71020 -11480 71120 -11380
rect 72520 -11480 72620 -11380
rect 74020 -11480 74120 -11380
rect 75520 -11480 75620 -11380
rect 77020 -11480 77120 -11380
rect 78520 -11480 78620 -11380
rect 80020 -11480 80120 -11380
rect 81520 -11480 81620 -11380
rect 83020 -11480 83120 -11380
rect 84520 -11480 84620 -11380
rect 86020 -11480 86120 -11380
rect 87520 -11480 87620 -11380
rect 89020 -11480 89120 -11380
rect 90520 -11480 90620 -11380
rect 92020 -11480 92120 -11380
rect 93520 -11480 93620 -11380
rect 95020 -11480 95120 -11380
rect 96520 -11480 96620 -11380
rect 98020 -11480 98120 -11380
rect 99520 -11480 99620 -11380
rect 101020 -11480 101120 -11380
rect 102520 -11480 102620 -11380
rect 104020 -11480 104120 -11380
rect 105520 -11480 105620 -11380
rect 107020 -11480 107120 -11380
rect 108520 -11480 108620 -11380
rect 110020 -11480 110120 -11380
rect 111520 -11480 111620 -11380
rect 113020 -11480 113120 -11380
rect 114520 -11480 114620 -11380
rect 116020 -11480 116120 -11380
rect 117520 -11480 117620 -11380
rect 119020 -11480 119120 -11380
rect 520 -12980 620 -12880
rect 2020 -12980 2120 -12880
rect 3520 -12980 3620 -12880
rect 5020 -12980 5120 -12880
rect 6520 -12980 6620 -12880
rect 8020 -12980 8120 -12880
rect 9520 -12980 9620 -12880
rect 11020 -12980 11120 -12880
rect 12520 -12980 12620 -12880
rect 14020 -12980 14120 -12880
rect 15520 -12980 15620 -12880
rect 17020 -12980 17120 -12880
rect 18520 -12980 18620 -12880
rect 20020 -12980 20120 -12880
rect 21520 -12980 21620 -12880
rect 23020 -12980 23120 -12880
rect 24520 -12980 24620 -12880
rect 26020 -12980 26120 -12880
rect 27520 -12980 27620 -12880
rect 29020 -12980 29120 -12880
rect 30520 -12980 30620 -12880
rect 32020 -12980 32120 -12880
rect 33520 -12980 33620 -12880
rect 35020 -12980 35120 -12880
rect 36520 -12980 36620 -12880
rect 38020 -12980 38120 -12880
rect 39520 -12980 39620 -12880
rect 41020 -12980 41120 -12880
rect 42520 -12980 42620 -12880
rect 44020 -12980 44120 -12880
rect 45520 -12980 45620 -12880
rect 47020 -12980 47120 -12880
rect 48520 -12980 48620 -12880
rect 50020 -12980 50120 -12880
rect 51520 -12980 51620 -12880
rect 53020 -12980 53120 -12880
rect 54520 -12980 54620 -12880
rect 56020 -12980 56120 -12880
rect 57520 -12980 57620 -12880
rect 59020 -12980 59120 -12880
rect 60520 -12980 60620 -12880
rect 62020 -12980 62120 -12880
rect 63520 -12980 63620 -12880
rect 65020 -12980 65120 -12880
rect 66520 -12980 66620 -12880
rect 68020 -12980 68120 -12880
rect 69520 -12980 69620 -12880
rect 71020 -12980 71120 -12880
rect 72520 -12980 72620 -12880
rect 74020 -12980 74120 -12880
rect 75520 -12980 75620 -12880
rect 77020 -12980 77120 -12880
rect 78520 -12980 78620 -12880
rect 80020 -12980 80120 -12880
rect 81520 -12980 81620 -12880
rect 83020 -12980 83120 -12880
rect 84520 -12980 84620 -12880
rect 86020 -12980 86120 -12880
rect 87520 -12980 87620 -12880
rect 89020 -12980 89120 -12880
rect 90520 -12980 90620 -12880
rect 92020 -12980 92120 -12880
rect 93520 -12980 93620 -12880
rect 95020 -12980 95120 -12880
rect 96520 -12980 96620 -12880
rect 98020 -12980 98120 -12880
rect 99520 -12980 99620 -12880
rect 101020 -12980 101120 -12880
rect 102520 -12980 102620 -12880
rect 104020 -12980 104120 -12880
rect 105520 -12980 105620 -12880
rect 107020 -12980 107120 -12880
rect 108520 -12980 108620 -12880
rect 110020 -12980 110120 -12880
rect 111520 -12980 111620 -12880
rect 113020 -12980 113120 -12880
rect 114520 -12980 114620 -12880
rect 116020 -12980 116120 -12880
rect 117520 -12980 117620 -12880
rect 119020 -12980 119120 -12880
rect 520 -14480 620 -14380
rect 2020 -14480 2120 -14380
rect 3520 -14480 3620 -14380
rect 5020 -14480 5120 -14380
rect 6520 -14480 6620 -14380
rect 8020 -14480 8120 -14380
rect 9520 -14480 9620 -14380
rect 11020 -14480 11120 -14380
rect 12520 -14480 12620 -14380
rect 14020 -14480 14120 -14380
rect 15520 -14480 15620 -14380
rect 17020 -14480 17120 -14380
rect 18520 -14480 18620 -14380
rect 20020 -14480 20120 -14380
rect 21520 -14480 21620 -14380
rect 23020 -14480 23120 -14380
rect 24520 -14480 24620 -14380
rect 26020 -14480 26120 -14380
rect 27520 -14480 27620 -14380
rect 29020 -14480 29120 -14380
rect 30520 -14480 30620 -14380
rect 32020 -14480 32120 -14380
rect 33520 -14480 33620 -14380
rect 35020 -14480 35120 -14380
rect 36520 -14480 36620 -14380
rect 38020 -14480 38120 -14380
rect 39520 -14480 39620 -14380
rect 41020 -14480 41120 -14380
rect 42520 -14480 42620 -14380
rect 44020 -14480 44120 -14380
rect 45520 -14480 45620 -14380
rect 47020 -14480 47120 -14380
rect 48520 -14480 48620 -14380
rect 50020 -14480 50120 -14380
rect 51520 -14480 51620 -14380
rect 53020 -14480 53120 -14380
rect 54520 -14480 54620 -14380
rect 56020 -14480 56120 -14380
rect 57520 -14480 57620 -14380
rect 59020 -14480 59120 -14380
rect 60520 -14480 60620 -14380
rect 62020 -14480 62120 -14380
rect 63520 -14480 63620 -14380
rect 65020 -14480 65120 -14380
rect 66520 -14480 66620 -14380
rect 68020 -14480 68120 -14380
rect 69520 -14480 69620 -14380
rect 71020 -14480 71120 -14380
rect 72520 -14480 72620 -14380
rect 74020 -14480 74120 -14380
rect 75520 -14480 75620 -14380
rect 77020 -14480 77120 -14380
rect 78520 -14480 78620 -14380
rect 80020 -14480 80120 -14380
rect 81520 -14480 81620 -14380
rect 83020 -14480 83120 -14380
rect 84520 -14480 84620 -14380
rect 86020 -14480 86120 -14380
rect 87520 -14480 87620 -14380
rect 89020 -14480 89120 -14380
rect 90520 -14480 90620 -14380
rect 92020 -14480 92120 -14380
rect 93520 -14480 93620 -14380
rect 95020 -14480 95120 -14380
rect 96520 -14480 96620 -14380
rect 98020 -14480 98120 -14380
rect 99520 -14480 99620 -14380
rect 101020 -14480 101120 -14380
rect 102520 -14480 102620 -14380
rect 104020 -14480 104120 -14380
rect 105520 -14480 105620 -14380
rect 107020 -14480 107120 -14380
rect 108520 -14480 108620 -14380
rect 110020 -14480 110120 -14380
rect 111520 -14480 111620 -14380
rect 113020 -14480 113120 -14380
rect 114520 -14480 114620 -14380
rect 116020 -14480 116120 -14380
rect 117520 -14480 117620 -14380
rect 119020 -14480 119120 -14380
rect 520 -15980 620 -15880
rect 2020 -15980 2120 -15880
rect 3520 -15980 3620 -15880
rect 5020 -15980 5120 -15880
rect 6520 -15980 6620 -15880
rect 8020 -15980 8120 -15880
rect 9520 -15980 9620 -15880
rect 11020 -15980 11120 -15880
rect 12520 -15980 12620 -15880
rect 14020 -15980 14120 -15880
rect 15520 -15980 15620 -15880
rect 17020 -15980 17120 -15880
rect 18520 -15980 18620 -15880
rect 20020 -15980 20120 -15880
rect 21520 -15980 21620 -15880
rect 23020 -15980 23120 -15880
rect 24520 -15980 24620 -15880
rect 26020 -15980 26120 -15880
rect 27520 -15980 27620 -15880
rect 29020 -15980 29120 -15880
rect 30520 -15980 30620 -15880
rect 32020 -15980 32120 -15880
rect 33520 -15980 33620 -15880
rect 35020 -15980 35120 -15880
rect 36520 -15980 36620 -15880
rect 38020 -15980 38120 -15880
rect 39520 -15980 39620 -15880
rect 41020 -15980 41120 -15880
rect 42520 -15980 42620 -15880
rect 44020 -15980 44120 -15880
rect 45520 -15980 45620 -15880
rect 47020 -15980 47120 -15880
rect 48520 -15980 48620 -15880
rect 50020 -15980 50120 -15880
rect 51520 -15980 51620 -15880
rect 53020 -15980 53120 -15880
rect 54520 -15980 54620 -15880
rect 56020 -15980 56120 -15880
rect 57520 -15980 57620 -15880
rect 59020 -15980 59120 -15880
rect 60520 -15980 60620 -15880
rect 62020 -15980 62120 -15880
rect 63520 -15980 63620 -15880
rect 65020 -15980 65120 -15880
rect 66520 -15980 66620 -15880
rect 68020 -15980 68120 -15880
rect 69520 -15980 69620 -15880
rect 71020 -15980 71120 -15880
rect 72520 -15980 72620 -15880
rect 74020 -15980 74120 -15880
rect 75520 -15980 75620 -15880
rect 77020 -15980 77120 -15880
rect 78520 -15980 78620 -15880
rect 80020 -15980 80120 -15880
rect 81520 -15980 81620 -15880
rect 83020 -15980 83120 -15880
rect 84520 -15980 84620 -15880
rect 86020 -15980 86120 -15880
rect 87520 -15980 87620 -15880
rect 89020 -15980 89120 -15880
rect 90520 -15980 90620 -15880
rect 92020 -15980 92120 -15880
rect 93520 -15980 93620 -15880
rect 95020 -15980 95120 -15880
rect 96520 -15980 96620 -15880
rect 98020 -15980 98120 -15880
rect 99520 -15980 99620 -15880
rect 101020 -15980 101120 -15880
rect 102520 -15980 102620 -15880
rect 104020 -15980 104120 -15880
rect 105520 -15980 105620 -15880
rect 107020 -15980 107120 -15880
rect 108520 -15980 108620 -15880
rect 110020 -15980 110120 -15880
rect 111520 -15980 111620 -15880
rect 113020 -15980 113120 -15880
rect 114520 -15980 114620 -15880
rect 116020 -15980 116120 -15880
rect 117520 -15980 117620 -15880
rect 119020 -15980 119120 -15880
rect 520 -17480 620 -17380
rect 2020 -17480 2120 -17380
rect 3520 -17480 3620 -17380
rect 5020 -17480 5120 -17380
rect 6520 -17480 6620 -17380
rect 8020 -17480 8120 -17380
rect 9520 -17480 9620 -17380
rect 11020 -17480 11120 -17380
rect 12520 -17480 12620 -17380
rect 14020 -17480 14120 -17380
rect 15520 -17480 15620 -17380
rect 17020 -17480 17120 -17380
rect 18520 -17480 18620 -17380
rect 20020 -17480 20120 -17380
rect 21520 -17480 21620 -17380
rect 23020 -17480 23120 -17380
rect 24520 -17480 24620 -17380
rect 26020 -17480 26120 -17380
rect 27520 -17480 27620 -17380
rect 29020 -17480 29120 -17380
rect 30520 -17480 30620 -17380
rect 32020 -17480 32120 -17380
rect 33520 -17480 33620 -17380
rect 35020 -17480 35120 -17380
rect 36520 -17480 36620 -17380
rect 38020 -17480 38120 -17380
rect 39520 -17480 39620 -17380
rect 41020 -17480 41120 -17380
rect 42520 -17480 42620 -17380
rect 44020 -17480 44120 -17380
rect 45520 -17480 45620 -17380
rect 47020 -17480 47120 -17380
rect 48520 -17480 48620 -17380
rect 50020 -17480 50120 -17380
rect 51520 -17480 51620 -17380
rect 53020 -17480 53120 -17380
rect 54520 -17480 54620 -17380
rect 56020 -17480 56120 -17380
rect 57520 -17480 57620 -17380
rect 59020 -17480 59120 -17380
rect 60520 -17480 60620 -17380
rect 62020 -17480 62120 -17380
rect 63520 -17480 63620 -17380
rect 65020 -17480 65120 -17380
rect 66520 -17480 66620 -17380
rect 68020 -17480 68120 -17380
rect 69520 -17480 69620 -17380
rect 71020 -17480 71120 -17380
rect 72520 -17480 72620 -17380
rect 74020 -17480 74120 -17380
rect 75520 -17480 75620 -17380
rect 77020 -17480 77120 -17380
rect 78520 -17480 78620 -17380
rect 80020 -17480 80120 -17380
rect 81520 -17480 81620 -17380
rect 83020 -17480 83120 -17380
rect 84520 -17480 84620 -17380
rect 86020 -17480 86120 -17380
rect 87520 -17480 87620 -17380
rect 89020 -17480 89120 -17380
rect 90520 -17480 90620 -17380
rect 92020 -17480 92120 -17380
rect 93520 -17480 93620 -17380
rect 95020 -17480 95120 -17380
rect 96520 -17480 96620 -17380
rect 98020 -17480 98120 -17380
rect 99520 -17480 99620 -17380
rect 101020 -17480 101120 -17380
rect 102520 -17480 102620 -17380
rect 104020 -17480 104120 -17380
rect 105520 -17480 105620 -17380
rect 107020 -17480 107120 -17380
rect 108520 -17480 108620 -17380
rect 110020 -17480 110120 -17380
rect 111520 -17480 111620 -17380
rect 113020 -17480 113120 -17380
rect 114520 -17480 114620 -17380
rect 116020 -17480 116120 -17380
rect 117520 -17480 117620 -17380
rect 119020 -17480 119120 -17380
rect 520 -18980 620 -18880
rect 2020 -18980 2120 -18880
rect 3520 -18980 3620 -18880
rect 5020 -18980 5120 -18880
rect 6520 -18980 6620 -18880
rect 8020 -18980 8120 -18880
rect 9520 -18980 9620 -18880
rect 11020 -18980 11120 -18880
rect 12520 -18980 12620 -18880
rect 14020 -18980 14120 -18880
rect 15520 -18980 15620 -18880
rect 17020 -18980 17120 -18880
rect 18520 -18980 18620 -18880
rect 20020 -18980 20120 -18880
rect 21520 -18980 21620 -18880
rect 23020 -18980 23120 -18880
rect 24520 -18980 24620 -18880
rect 26020 -18980 26120 -18880
rect 27520 -18980 27620 -18880
rect 29020 -18980 29120 -18880
rect 30520 -18980 30620 -18880
rect 32020 -18980 32120 -18880
rect 33520 -18980 33620 -18880
rect 35020 -18980 35120 -18880
rect 36520 -18980 36620 -18880
rect 38020 -18980 38120 -18880
rect 39520 -18980 39620 -18880
rect 41020 -18980 41120 -18880
rect 42520 -18980 42620 -18880
rect 44020 -18980 44120 -18880
rect 45520 -18980 45620 -18880
rect 47020 -18980 47120 -18880
rect 48520 -18980 48620 -18880
rect 50020 -18980 50120 -18880
rect 51520 -18980 51620 -18880
rect 53020 -18980 53120 -18880
rect 54520 -18980 54620 -18880
rect 56020 -18980 56120 -18880
rect 57520 -18980 57620 -18880
rect 59020 -18980 59120 -18880
rect 60520 -18980 60620 -18880
rect 62020 -18980 62120 -18880
rect 63520 -18980 63620 -18880
rect 65020 -18980 65120 -18880
rect 66520 -18980 66620 -18880
rect 68020 -18980 68120 -18880
rect 69520 -18980 69620 -18880
rect 71020 -18980 71120 -18880
rect 72520 -18980 72620 -18880
rect 74020 -18980 74120 -18880
rect 75520 -18980 75620 -18880
rect 77020 -18980 77120 -18880
rect 78520 -18980 78620 -18880
rect 80020 -18980 80120 -18880
rect 81520 -18980 81620 -18880
rect 83020 -18980 83120 -18880
rect 84520 -18980 84620 -18880
rect 86020 -18980 86120 -18880
rect 87520 -18980 87620 -18880
rect 89020 -18980 89120 -18880
rect 90520 -18980 90620 -18880
rect 92020 -18980 92120 -18880
rect 93520 -18980 93620 -18880
rect 95020 -18980 95120 -18880
rect 96520 -18980 96620 -18880
rect 98020 -18980 98120 -18880
rect 99520 -18980 99620 -18880
rect 101020 -18980 101120 -18880
rect 102520 -18980 102620 -18880
rect 104020 -18980 104120 -18880
rect 105520 -18980 105620 -18880
rect 107020 -18980 107120 -18880
rect 108520 -18980 108620 -18880
rect 110020 -18980 110120 -18880
rect 111520 -18980 111620 -18880
rect 113020 -18980 113120 -18880
rect 114520 -18980 114620 -18880
rect 116020 -18980 116120 -18880
rect 117520 -18980 117620 -18880
rect 119020 -18980 119120 -18880
rect 520 -20480 620 -20380
rect 2020 -20480 2120 -20380
rect 3520 -20480 3620 -20380
rect 5020 -20480 5120 -20380
rect 6520 -20480 6620 -20380
rect 8020 -20480 8120 -20380
rect 9520 -20480 9620 -20380
rect 11020 -20480 11120 -20380
rect 12520 -20480 12620 -20380
rect 14020 -20480 14120 -20380
rect 15520 -20480 15620 -20380
rect 17020 -20480 17120 -20380
rect 18520 -20480 18620 -20380
rect 20020 -20480 20120 -20380
rect 21520 -20480 21620 -20380
rect 23020 -20480 23120 -20380
rect 24520 -20480 24620 -20380
rect 26020 -20480 26120 -20380
rect 27520 -20480 27620 -20380
rect 29020 -20480 29120 -20380
rect 30520 -20480 30620 -20380
rect 32020 -20480 32120 -20380
rect 33520 -20480 33620 -20380
rect 35020 -20480 35120 -20380
rect 36520 -20480 36620 -20380
rect 38020 -20480 38120 -20380
rect 39520 -20480 39620 -20380
rect 41020 -20480 41120 -20380
rect 42520 -20480 42620 -20380
rect 44020 -20480 44120 -20380
rect 45520 -20480 45620 -20380
rect 47020 -20480 47120 -20380
rect 48520 -20480 48620 -20380
rect 50020 -20480 50120 -20380
rect 51520 -20480 51620 -20380
rect 53020 -20480 53120 -20380
rect 54520 -20480 54620 -20380
rect 56020 -20480 56120 -20380
rect 57520 -20480 57620 -20380
rect 59020 -20480 59120 -20380
rect 60520 -20480 60620 -20380
rect 62020 -20480 62120 -20380
rect 63520 -20480 63620 -20380
rect 65020 -20480 65120 -20380
rect 66520 -20480 66620 -20380
rect 68020 -20480 68120 -20380
rect 69520 -20480 69620 -20380
rect 71020 -20480 71120 -20380
rect 72520 -20480 72620 -20380
rect 74020 -20480 74120 -20380
rect 75520 -20480 75620 -20380
rect 77020 -20480 77120 -20380
rect 78520 -20480 78620 -20380
rect 80020 -20480 80120 -20380
rect 81520 -20480 81620 -20380
rect 83020 -20480 83120 -20380
rect 84520 -20480 84620 -20380
rect 86020 -20480 86120 -20380
rect 87520 -20480 87620 -20380
rect 89020 -20480 89120 -20380
rect 90520 -20480 90620 -20380
rect 92020 -20480 92120 -20380
rect 93520 -20480 93620 -20380
rect 95020 -20480 95120 -20380
rect 96520 -20480 96620 -20380
rect 98020 -20480 98120 -20380
rect 99520 -20480 99620 -20380
rect 101020 -20480 101120 -20380
rect 102520 -20480 102620 -20380
rect 104020 -20480 104120 -20380
rect 105520 -20480 105620 -20380
rect 107020 -20480 107120 -20380
rect 108520 -20480 108620 -20380
rect 110020 -20480 110120 -20380
rect 111520 -20480 111620 -20380
rect 113020 -20480 113120 -20380
rect 114520 -20480 114620 -20380
rect 116020 -20480 116120 -20380
rect 117520 -20480 117620 -20380
rect 119020 -20480 119120 -20380
rect 520 -21980 620 -21880
rect 2020 -21980 2120 -21880
rect 3520 -21980 3620 -21880
rect 5020 -21980 5120 -21880
rect 6520 -21980 6620 -21880
rect 8020 -21980 8120 -21880
rect 9520 -21980 9620 -21880
rect 11020 -21980 11120 -21880
rect 12520 -21980 12620 -21880
rect 14020 -21980 14120 -21880
rect 15520 -21980 15620 -21880
rect 17020 -21980 17120 -21880
rect 18520 -21980 18620 -21880
rect 20020 -21980 20120 -21880
rect 21520 -21980 21620 -21880
rect 23020 -21980 23120 -21880
rect 24520 -21980 24620 -21880
rect 26020 -21980 26120 -21880
rect 27520 -21980 27620 -21880
rect 29020 -21980 29120 -21880
rect 30520 -21980 30620 -21880
rect 32020 -21980 32120 -21880
rect 33520 -21980 33620 -21880
rect 35020 -21980 35120 -21880
rect 36520 -21980 36620 -21880
rect 38020 -21980 38120 -21880
rect 39520 -21980 39620 -21880
rect 41020 -21980 41120 -21880
rect 42520 -21980 42620 -21880
rect 44020 -21980 44120 -21880
rect 45520 -21980 45620 -21880
rect 47020 -21980 47120 -21880
rect 48520 -21980 48620 -21880
rect 50020 -21980 50120 -21880
rect 51520 -21980 51620 -21880
rect 53020 -21980 53120 -21880
rect 54520 -21980 54620 -21880
rect 56020 -21980 56120 -21880
rect 57520 -21980 57620 -21880
rect 59020 -21980 59120 -21880
rect 60520 -21980 60620 -21880
rect 62020 -21980 62120 -21880
rect 63520 -21980 63620 -21880
rect 65020 -21980 65120 -21880
rect 66520 -21980 66620 -21880
rect 68020 -21980 68120 -21880
rect 69520 -21980 69620 -21880
rect 71020 -21980 71120 -21880
rect 72520 -21980 72620 -21880
rect 74020 -21980 74120 -21880
rect 75520 -21980 75620 -21880
rect 77020 -21980 77120 -21880
rect 78520 -21980 78620 -21880
rect 80020 -21980 80120 -21880
rect 81520 -21980 81620 -21880
rect 83020 -21980 83120 -21880
rect 84520 -21980 84620 -21880
rect 86020 -21980 86120 -21880
rect 87520 -21980 87620 -21880
rect 89020 -21980 89120 -21880
rect 90520 -21980 90620 -21880
rect 92020 -21980 92120 -21880
rect 93520 -21980 93620 -21880
rect 95020 -21980 95120 -21880
rect 96520 -21980 96620 -21880
rect 98020 -21980 98120 -21880
rect 99520 -21980 99620 -21880
rect 101020 -21980 101120 -21880
rect 102520 -21980 102620 -21880
rect 104020 -21980 104120 -21880
rect 105520 -21980 105620 -21880
rect 107020 -21980 107120 -21880
rect 108520 -21980 108620 -21880
rect 110020 -21980 110120 -21880
rect 111520 -21980 111620 -21880
rect 113020 -21980 113120 -21880
rect 114520 -21980 114620 -21880
rect 116020 -21980 116120 -21880
rect 117520 -21980 117620 -21880
rect 119020 -21980 119120 -21880
rect 520 -23480 620 -23380
rect 2020 -23480 2120 -23380
rect 3520 -23480 3620 -23380
rect 5020 -23480 5120 -23380
rect 6520 -23480 6620 -23380
rect 8020 -23480 8120 -23380
rect 9520 -23480 9620 -23380
rect 11020 -23480 11120 -23380
rect 12520 -23480 12620 -23380
rect 14020 -23480 14120 -23380
rect 15520 -23480 15620 -23380
rect 17020 -23480 17120 -23380
rect 18520 -23480 18620 -23380
rect 20020 -23480 20120 -23380
rect 21520 -23480 21620 -23380
rect 23020 -23480 23120 -23380
rect 24520 -23480 24620 -23380
rect 26020 -23480 26120 -23380
rect 27520 -23480 27620 -23380
rect 29020 -23480 29120 -23380
rect 30520 -23480 30620 -23380
rect 32020 -23480 32120 -23380
rect 33520 -23480 33620 -23380
rect 35020 -23480 35120 -23380
rect 36520 -23480 36620 -23380
rect 38020 -23480 38120 -23380
rect 39520 -23480 39620 -23380
rect 41020 -23480 41120 -23380
rect 42520 -23480 42620 -23380
rect 44020 -23480 44120 -23380
rect 45520 -23480 45620 -23380
rect 47020 -23480 47120 -23380
rect 48520 -23480 48620 -23380
rect 50020 -23480 50120 -23380
rect 51520 -23480 51620 -23380
rect 53020 -23480 53120 -23380
rect 54520 -23480 54620 -23380
rect 56020 -23480 56120 -23380
rect 57520 -23480 57620 -23380
rect 59020 -23480 59120 -23380
rect 60520 -23480 60620 -23380
rect 62020 -23480 62120 -23380
rect 63520 -23480 63620 -23380
rect 65020 -23480 65120 -23380
rect 66520 -23480 66620 -23380
rect 68020 -23480 68120 -23380
rect 69520 -23480 69620 -23380
rect 71020 -23480 71120 -23380
rect 72520 -23480 72620 -23380
rect 74020 -23480 74120 -23380
rect 75520 -23480 75620 -23380
rect 77020 -23480 77120 -23380
rect 78520 -23480 78620 -23380
rect 80020 -23480 80120 -23380
rect 81520 -23480 81620 -23380
rect 83020 -23480 83120 -23380
rect 84520 -23480 84620 -23380
rect 86020 -23480 86120 -23380
rect 87520 -23480 87620 -23380
rect 89020 -23480 89120 -23380
rect 90520 -23480 90620 -23380
rect 92020 -23480 92120 -23380
rect 93520 -23480 93620 -23380
rect 95020 -23480 95120 -23380
rect 96520 -23480 96620 -23380
rect 98020 -23480 98120 -23380
rect 99520 -23480 99620 -23380
rect 101020 -23480 101120 -23380
rect 102520 -23480 102620 -23380
rect 104020 -23480 104120 -23380
rect 105520 -23480 105620 -23380
rect 107020 -23480 107120 -23380
rect 108520 -23480 108620 -23380
rect 110020 -23480 110120 -23380
rect 111520 -23480 111620 -23380
rect 113020 -23480 113120 -23380
rect 114520 -23480 114620 -23380
rect 116020 -23480 116120 -23380
rect 117520 -23480 117620 -23380
rect 119020 -23480 119120 -23380
rect 520 -24980 620 -24880
rect 2020 -24980 2120 -24880
rect 3520 -24980 3620 -24880
rect 5020 -24980 5120 -24880
rect 6520 -24980 6620 -24880
rect 8020 -24980 8120 -24880
rect 9520 -24980 9620 -24880
rect 11020 -24980 11120 -24880
rect 12520 -24980 12620 -24880
rect 14020 -24980 14120 -24880
rect 15520 -24980 15620 -24880
rect 17020 -24980 17120 -24880
rect 18520 -24980 18620 -24880
rect 20020 -24980 20120 -24880
rect 21520 -24980 21620 -24880
rect 23020 -24980 23120 -24880
rect 24520 -24980 24620 -24880
rect 26020 -24980 26120 -24880
rect 27520 -24980 27620 -24880
rect 29020 -24980 29120 -24880
rect 30520 -24980 30620 -24880
rect 32020 -24980 32120 -24880
rect 33520 -24980 33620 -24880
rect 35020 -24980 35120 -24880
rect 36520 -24980 36620 -24880
rect 38020 -24980 38120 -24880
rect 39520 -24980 39620 -24880
rect 41020 -24980 41120 -24880
rect 42520 -24980 42620 -24880
rect 44020 -24980 44120 -24880
rect 45520 -24980 45620 -24880
rect 47020 -24980 47120 -24880
rect 48520 -24980 48620 -24880
rect 50020 -24980 50120 -24880
rect 51520 -24980 51620 -24880
rect 53020 -24980 53120 -24880
rect 54520 -24980 54620 -24880
rect 56020 -24980 56120 -24880
rect 57520 -24980 57620 -24880
rect 59020 -24980 59120 -24880
rect 60520 -24980 60620 -24880
rect 62020 -24980 62120 -24880
rect 63520 -24980 63620 -24880
rect 65020 -24980 65120 -24880
rect 66520 -24980 66620 -24880
rect 68020 -24980 68120 -24880
rect 69520 -24980 69620 -24880
rect 71020 -24980 71120 -24880
rect 72520 -24980 72620 -24880
rect 74020 -24980 74120 -24880
rect 75520 -24980 75620 -24880
rect 77020 -24980 77120 -24880
rect 78520 -24980 78620 -24880
rect 80020 -24980 80120 -24880
rect 81520 -24980 81620 -24880
rect 83020 -24980 83120 -24880
rect 84520 -24980 84620 -24880
rect 86020 -24980 86120 -24880
rect 87520 -24980 87620 -24880
rect 89020 -24980 89120 -24880
rect 90520 -24980 90620 -24880
rect 92020 -24980 92120 -24880
rect 93520 -24980 93620 -24880
rect 95020 -24980 95120 -24880
rect 96520 -24980 96620 -24880
rect 98020 -24980 98120 -24880
rect 99520 -24980 99620 -24880
rect 101020 -24980 101120 -24880
rect 102520 -24980 102620 -24880
rect 104020 -24980 104120 -24880
rect 105520 -24980 105620 -24880
rect 107020 -24980 107120 -24880
rect 108520 -24980 108620 -24880
rect 110020 -24980 110120 -24880
rect 111520 -24980 111620 -24880
rect 113020 -24980 113120 -24880
rect 114520 -24980 114620 -24880
rect 116020 -24980 116120 -24880
rect 117520 -24980 117620 -24880
rect 119020 -24980 119120 -24880
rect 520 -26480 620 -26380
rect 2020 -26480 2120 -26380
rect 3520 -26480 3620 -26380
rect 5020 -26480 5120 -26380
rect 6520 -26480 6620 -26380
rect 8020 -26480 8120 -26380
rect 9520 -26480 9620 -26380
rect 11020 -26480 11120 -26380
rect 12520 -26480 12620 -26380
rect 14020 -26480 14120 -26380
rect 15520 -26480 15620 -26380
rect 17020 -26480 17120 -26380
rect 18520 -26480 18620 -26380
rect 20020 -26480 20120 -26380
rect 21520 -26480 21620 -26380
rect 23020 -26480 23120 -26380
rect 24520 -26480 24620 -26380
rect 26020 -26480 26120 -26380
rect 27520 -26480 27620 -26380
rect 29020 -26480 29120 -26380
rect 30520 -26480 30620 -26380
rect 32020 -26480 32120 -26380
rect 33520 -26480 33620 -26380
rect 35020 -26480 35120 -26380
rect 36520 -26480 36620 -26380
rect 38020 -26480 38120 -26380
rect 39520 -26480 39620 -26380
rect 41020 -26480 41120 -26380
rect 42520 -26480 42620 -26380
rect 44020 -26480 44120 -26380
rect 45520 -26480 45620 -26380
rect 47020 -26480 47120 -26380
rect 48520 -26480 48620 -26380
rect 50020 -26480 50120 -26380
rect 51520 -26480 51620 -26380
rect 53020 -26480 53120 -26380
rect 54520 -26480 54620 -26380
rect 56020 -26480 56120 -26380
rect 57520 -26480 57620 -26380
rect 59020 -26480 59120 -26380
rect 60520 -26480 60620 -26380
rect 62020 -26480 62120 -26380
rect 63520 -26480 63620 -26380
rect 65020 -26480 65120 -26380
rect 66520 -26480 66620 -26380
rect 68020 -26480 68120 -26380
rect 69520 -26480 69620 -26380
rect 71020 -26480 71120 -26380
rect 72520 -26480 72620 -26380
rect 74020 -26480 74120 -26380
rect 75520 -26480 75620 -26380
rect 77020 -26480 77120 -26380
rect 78520 -26480 78620 -26380
rect 80020 -26480 80120 -26380
rect 81520 -26480 81620 -26380
rect 83020 -26480 83120 -26380
rect 84520 -26480 84620 -26380
rect 86020 -26480 86120 -26380
rect 87520 -26480 87620 -26380
rect 89020 -26480 89120 -26380
rect 90520 -26480 90620 -26380
rect 92020 -26480 92120 -26380
rect 93520 -26480 93620 -26380
rect 95020 -26480 95120 -26380
rect 96520 -26480 96620 -26380
rect 98020 -26480 98120 -26380
rect 99520 -26480 99620 -26380
rect 101020 -26480 101120 -26380
rect 102520 -26480 102620 -26380
rect 104020 -26480 104120 -26380
rect 105520 -26480 105620 -26380
rect 107020 -26480 107120 -26380
rect 108520 -26480 108620 -26380
rect 110020 -26480 110120 -26380
rect 111520 -26480 111620 -26380
rect 113020 -26480 113120 -26380
rect 114520 -26480 114620 -26380
rect 116020 -26480 116120 -26380
rect 117520 -26480 117620 -26380
rect 119020 -26480 119120 -26380
rect 520 -27980 620 -27880
rect 2020 -27980 2120 -27880
rect 3520 -27980 3620 -27880
rect 5020 -27980 5120 -27880
rect 6520 -27980 6620 -27880
rect 8020 -27980 8120 -27880
rect 9520 -27980 9620 -27880
rect 11020 -27980 11120 -27880
rect 12520 -27980 12620 -27880
rect 14020 -27980 14120 -27880
rect 15520 -27980 15620 -27880
rect 17020 -27980 17120 -27880
rect 18520 -27980 18620 -27880
rect 20020 -27980 20120 -27880
rect 21520 -27980 21620 -27880
rect 23020 -27980 23120 -27880
rect 24520 -27980 24620 -27880
rect 26020 -27980 26120 -27880
rect 27520 -27980 27620 -27880
rect 29020 -27980 29120 -27880
rect 30520 -27980 30620 -27880
rect 32020 -27980 32120 -27880
rect 33520 -27980 33620 -27880
rect 35020 -27980 35120 -27880
rect 36520 -27980 36620 -27880
rect 38020 -27980 38120 -27880
rect 39520 -27980 39620 -27880
rect 41020 -27980 41120 -27880
rect 42520 -27980 42620 -27880
rect 44020 -27980 44120 -27880
rect 45520 -27980 45620 -27880
rect 47020 -27980 47120 -27880
rect 48520 -27980 48620 -27880
rect 50020 -27980 50120 -27880
rect 51520 -27980 51620 -27880
rect 53020 -27980 53120 -27880
rect 54520 -27980 54620 -27880
rect 56020 -27980 56120 -27880
rect 57520 -27980 57620 -27880
rect 59020 -27980 59120 -27880
rect 60520 -27980 60620 -27880
rect 62020 -27980 62120 -27880
rect 63520 -27980 63620 -27880
rect 65020 -27980 65120 -27880
rect 66520 -27980 66620 -27880
rect 68020 -27980 68120 -27880
rect 69520 -27980 69620 -27880
rect 71020 -27980 71120 -27880
rect 72520 -27980 72620 -27880
rect 74020 -27980 74120 -27880
rect 75520 -27980 75620 -27880
rect 77020 -27980 77120 -27880
rect 78520 -27980 78620 -27880
rect 80020 -27980 80120 -27880
rect 81520 -27980 81620 -27880
rect 83020 -27980 83120 -27880
rect 84520 -27980 84620 -27880
rect 86020 -27980 86120 -27880
rect 87520 -27980 87620 -27880
rect 89020 -27980 89120 -27880
rect 90520 -27980 90620 -27880
rect 92020 -27980 92120 -27880
rect 93520 -27980 93620 -27880
rect 95020 -27980 95120 -27880
rect 96520 -27980 96620 -27880
rect 98020 -27980 98120 -27880
rect 99520 -27980 99620 -27880
rect 101020 -27980 101120 -27880
rect 102520 -27980 102620 -27880
rect 104020 -27980 104120 -27880
rect 105520 -27980 105620 -27880
rect 107020 -27980 107120 -27880
rect 108520 -27980 108620 -27880
rect 110020 -27980 110120 -27880
rect 111520 -27980 111620 -27880
rect 113020 -27980 113120 -27880
rect 114520 -27980 114620 -27880
rect 116020 -27980 116120 -27880
rect 117520 -27980 117620 -27880
rect 119020 -27980 119120 -27880
rect 520 -29480 620 -29380
rect 2020 -29480 2120 -29380
rect 3520 -29480 3620 -29380
rect 5020 -29480 5120 -29380
rect 6520 -29480 6620 -29380
rect 8020 -29480 8120 -29380
rect 9520 -29480 9620 -29380
rect 11020 -29480 11120 -29380
rect 12520 -29480 12620 -29380
rect 14020 -29480 14120 -29380
rect 15520 -29480 15620 -29380
rect 17020 -29480 17120 -29380
rect 18520 -29480 18620 -29380
rect 20020 -29480 20120 -29380
rect 21520 -29480 21620 -29380
rect 23020 -29480 23120 -29380
rect 24520 -29480 24620 -29380
rect 26020 -29480 26120 -29380
rect 27520 -29480 27620 -29380
rect 29020 -29480 29120 -29380
rect 30520 -29480 30620 -29380
rect 32020 -29480 32120 -29380
rect 33520 -29480 33620 -29380
rect 35020 -29480 35120 -29380
rect 36520 -29480 36620 -29380
rect 38020 -29480 38120 -29380
rect 39520 -29480 39620 -29380
rect 41020 -29480 41120 -29380
rect 42520 -29480 42620 -29380
rect 44020 -29480 44120 -29380
rect 45520 -29480 45620 -29380
rect 47020 -29480 47120 -29380
rect 48520 -29480 48620 -29380
rect 50020 -29480 50120 -29380
rect 51520 -29480 51620 -29380
rect 53020 -29480 53120 -29380
rect 54520 -29480 54620 -29380
rect 56020 -29480 56120 -29380
rect 57520 -29480 57620 -29380
rect 59020 -29480 59120 -29380
rect 60520 -29480 60620 -29380
rect 62020 -29480 62120 -29380
rect 63520 -29480 63620 -29380
rect 65020 -29480 65120 -29380
rect 66520 -29480 66620 -29380
rect 68020 -29480 68120 -29380
rect 69520 -29480 69620 -29380
rect 71020 -29480 71120 -29380
rect 72520 -29480 72620 -29380
rect 74020 -29480 74120 -29380
rect 75520 -29480 75620 -29380
rect 77020 -29480 77120 -29380
rect 78520 -29480 78620 -29380
rect 80020 -29480 80120 -29380
rect 81520 -29480 81620 -29380
rect 83020 -29480 83120 -29380
rect 84520 -29480 84620 -29380
rect 86020 -29480 86120 -29380
rect 87520 -29480 87620 -29380
rect 89020 -29480 89120 -29380
rect 90520 -29480 90620 -29380
rect 92020 -29480 92120 -29380
rect 93520 -29480 93620 -29380
rect 95020 -29480 95120 -29380
rect 96520 -29480 96620 -29380
rect 98020 -29480 98120 -29380
rect 99520 -29480 99620 -29380
rect 101020 -29480 101120 -29380
rect 102520 -29480 102620 -29380
rect 104020 -29480 104120 -29380
rect 105520 -29480 105620 -29380
rect 107020 -29480 107120 -29380
rect 108520 -29480 108620 -29380
rect 110020 -29480 110120 -29380
rect 111520 -29480 111620 -29380
rect 113020 -29480 113120 -29380
rect 114520 -29480 114620 -29380
rect 116020 -29480 116120 -29380
rect 117520 -29480 117620 -29380
rect 119020 -29480 119120 -29380
rect 520 -30980 620 -30880
rect 2020 -30980 2120 -30880
rect 3520 -30980 3620 -30880
rect 5020 -30980 5120 -30880
rect 6520 -30980 6620 -30880
rect 8020 -30980 8120 -30880
rect 9520 -30980 9620 -30880
rect 11020 -30980 11120 -30880
rect 12520 -30980 12620 -30880
rect 14020 -30980 14120 -30880
rect 15520 -30980 15620 -30880
rect 17020 -30980 17120 -30880
rect 18520 -30980 18620 -30880
rect 20020 -30980 20120 -30880
rect 21520 -30980 21620 -30880
rect 23020 -30980 23120 -30880
rect 24520 -30980 24620 -30880
rect 26020 -30980 26120 -30880
rect 27520 -30980 27620 -30880
rect 29020 -30980 29120 -30880
rect 30520 -30980 30620 -30880
rect 32020 -30980 32120 -30880
rect 33520 -30980 33620 -30880
rect 35020 -30980 35120 -30880
rect 36520 -30980 36620 -30880
rect 38020 -30980 38120 -30880
rect 39520 -30980 39620 -30880
rect 41020 -30980 41120 -30880
rect 42520 -30980 42620 -30880
rect 44020 -30980 44120 -30880
rect 45520 -30980 45620 -30880
rect 47020 -30980 47120 -30880
rect 48520 -30980 48620 -30880
rect 50020 -30980 50120 -30880
rect 51520 -30980 51620 -30880
rect 53020 -30980 53120 -30880
rect 54520 -30980 54620 -30880
rect 56020 -30980 56120 -30880
rect 57520 -30980 57620 -30880
rect 59020 -30980 59120 -30880
rect 60520 -30980 60620 -30880
rect 62020 -30980 62120 -30880
rect 63520 -30980 63620 -30880
rect 65020 -30980 65120 -30880
rect 66520 -30980 66620 -30880
rect 68020 -30980 68120 -30880
rect 69520 -30980 69620 -30880
rect 71020 -30980 71120 -30880
rect 72520 -30980 72620 -30880
rect 74020 -30980 74120 -30880
rect 75520 -30980 75620 -30880
rect 77020 -30980 77120 -30880
rect 78520 -30980 78620 -30880
rect 80020 -30980 80120 -30880
rect 81520 -30980 81620 -30880
rect 83020 -30980 83120 -30880
rect 84520 -30980 84620 -30880
rect 86020 -30980 86120 -30880
rect 87520 -30980 87620 -30880
rect 89020 -30980 89120 -30880
rect 90520 -30980 90620 -30880
rect 92020 -30980 92120 -30880
rect 93520 -30980 93620 -30880
rect 95020 -30980 95120 -30880
rect 96520 -30980 96620 -30880
rect 98020 -30980 98120 -30880
rect 99520 -30980 99620 -30880
rect 101020 -30980 101120 -30880
rect 102520 -30980 102620 -30880
rect 104020 -30980 104120 -30880
rect 105520 -30980 105620 -30880
rect 107020 -30980 107120 -30880
rect 108520 -30980 108620 -30880
rect 110020 -30980 110120 -30880
rect 111520 -30980 111620 -30880
rect 113020 -30980 113120 -30880
rect 114520 -30980 114620 -30880
rect 116020 -30980 116120 -30880
rect 117520 -30980 117620 -30880
rect 119020 -30980 119120 -30880
rect 520 -32480 620 -32380
rect 2020 -32480 2120 -32380
rect 3520 -32480 3620 -32380
rect 5020 -32480 5120 -32380
rect 6520 -32480 6620 -32380
rect 8020 -32480 8120 -32380
rect 9520 -32480 9620 -32380
rect 11020 -32480 11120 -32380
rect 12520 -32480 12620 -32380
rect 14020 -32480 14120 -32380
rect 15520 -32480 15620 -32380
rect 17020 -32480 17120 -32380
rect 18520 -32480 18620 -32380
rect 20020 -32480 20120 -32380
rect 21520 -32480 21620 -32380
rect 23020 -32480 23120 -32380
rect 24520 -32480 24620 -32380
rect 26020 -32480 26120 -32380
rect 27520 -32480 27620 -32380
rect 29020 -32480 29120 -32380
rect 30520 -32480 30620 -32380
rect 32020 -32480 32120 -32380
rect 33520 -32480 33620 -32380
rect 35020 -32480 35120 -32380
rect 36520 -32480 36620 -32380
rect 38020 -32480 38120 -32380
rect 39520 -32480 39620 -32380
rect 41020 -32480 41120 -32380
rect 42520 -32480 42620 -32380
rect 44020 -32480 44120 -32380
rect 45520 -32480 45620 -32380
rect 47020 -32480 47120 -32380
rect 48520 -32480 48620 -32380
rect 50020 -32480 50120 -32380
rect 51520 -32480 51620 -32380
rect 53020 -32480 53120 -32380
rect 54520 -32480 54620 -32380
rect 56020 -32480 56120 -32380
rect 57520 -32480 57620 -32380
rect 59020 -32480 59120 -32380
rect 60520 -32480 60620 -32380
rect 62020 -32480 62120 -32380
rect 63520 -32480 63620 -32380
rect 65020 -32480 65120 -32380
rect 66520 -32480 66620 -32380
rect 68020 -32480 68120 -32380
rect 69520 -32480 69620 -32380
rect 71020 -32480 71120 -32380
rect 72520 -32480 72620 -32380
rect 74020 -32480 74120 -32380
rect 75520 -32480 75620 -32380
rect 77020 -32480 77120 -32380
rect 78520 -32480 78620 -32380
rect 80020 -32480 80120 -32380
rect 81520 -32480 81620 -32380
rect 83020 -32480 83120 -32380
rect 84520 -32480 84620 -32380
rect 86020 -32480 86120 -32380
rect 87520 -32480 87620 -32380
rect 89020 -32480 89120 -32380
rect 90520 -32480 90620 -32380
rect 92020 -32480 92120 -32380
rect 93520 -32480 93620 -32380
rect 95020 -32480 95120 -32380
rect 96520 -32480 96620 -32380
rect 98020 -32480 98120 -32380
rect 99520 -32480 99620 -32380
rect 101020 -32480 101120 -32380
rect 102520 -32480 102620 -32380
rect 104020 -32480 104120 -32380
rect 105520 -32480 105620 -32380
rect 107020 -32480 107120 -32380
rect 108520 -32480 108620 -32380
rect 110020 -32480 110120 -32380
rect 111520 -32480 111620 -32380
rect 113020 -32480 113120 -32380
rect 114520 -32480 114620 -32380
rect 116020 -32480 116120 -32380
rect 117520 -32480 117620 -32380
rect 119020 -32480 119120 -32380
rect 520 -33980 620 -33880
rect 2020 -33980 2120 -33880
rect 3520 -33980 3620 -33880
rect 5020 -33980 5120 -33880
rect 6520 -33980 6620 -33880
rect 8020 -33980 8120 -33880
rect 9520 -33980 9620 -33880
rect 11020 -33980 11120 -33880
rect 12520 -33980 12620 -33880
rect 14020 -33980 14120 -33880
rect 15520 -33980 15620 -33880
rect 17020 -33980 17120 -33880
rect 18520 -33980 18620 -33880
rect 20020 -33980 20120 -33880
rect 21520 -33980 21620 -33880
rect 23020 -33980 23120 -33880
rect 24520 -33980 24620 -33880
rect 26020 -33980 26120 -33880
rect 27520 -33980 27620 -33880
rect 29020 -33980 29120 -33880
rect 30520 -33980 30620 -33880
rect 32020 -33980 32120 -33880
rect 33520 -33980 33620 -33880
rect 35020 -33980 35120 -33880
rect 36520 -33980 36620 -33880
rect 38020 -33980 38120 -33880
rect 39520 -33980 39620 -33880
rect 41020 -33980 41120 -33880
rect 42520 -33980 42620 -33880
rect 44020 -33980 44120 -33880
rect 45520 -33980 45620 -33880
rect 47020 -33980 47120 -33880
rect 48520 -33980 48620 -33880
rect 50020 -33980 50120 -33880
rect 51520 -33980 51620 -33880
rect 53020 -33980 53120 -33880
rect 54520 -33980 54620 -33880
rect 56020 -33980 56120 -33880
rect 57520 -33980 57620 -33880
rect 59020 -33980 59120 -33880
rect 60520 -33980 60620 -33880
rect 62020 -33980 62120 -33880
rect 63520 -33980 63620 -33880
rect 65020 -33980 65120 -33880
rect 66520 -33980 66620 -33880
rect 68020 -33980 68120 -33880
rect 69520 -33980 69620 -33880
rect 71020 -33980 71120 -33880
rect 72520 -33980 72620 -33880
rect 74020 -33980 74120 -33880
rect 75520 -33980 75620 -33880
rect 77020 -33980 77120 -33880
rect 78520 -33980 78620 -33880
rect 80020 -33980 80120 -33880
rect 81520 -33980 81620 -33880
rect 83020 -33980 83120 -33880
rect 84520 -33980 84620 -33880
rect 86020 -33980 86120 -33880
rect 87520 -33980 87620 -33880
rect 89020 -33980 89120 -33880
rect 90520 -33980 90620 -33880
rect 92020 -33980 92120 -33880
rect 93520 -33980 93620 -33880
rect 95020 -33980 95120 -33880
rect 96520 -33980 96620 -33880
rect 98020 -33980 98120 -33880
rect 99520 -33980 99620 -33880
rect 101020 -33980 101120 -33880
rect 102520 -33980 102620 -33880
rect 104020 -33980 104120 -33880
rect 105520 -33980 105620 -33880
rect 107020 -33980 107120 -33880
rect 108520 -33980 108620 -33880
rect 110020 -33980 110120 -33880
rect 111520 -33980 111620 -33880
rect 113020 -33980 113120 -33880
rect 114520 -33980 114620 -33880
rect 116020 -33980 116120 -33880
rect 117520 -33980 117620 -33880
rect 119020 -33980 119120 -33880
rect 520 -35480 620 -35380
rect 2020 -35480 2120 -35380
rect 3520 -35480 3620 -35380
rect 5020 -35480 5120 -35380
rect 6520 -35480 6620 -35380
rect 8020 -35480 8120 -35380
rect 9520 -35480 9620 -35380
rect 11020 -35480 11120 -35380
rect 12520 -35480 12620 -35380
rect 14020 -35480 14120 -35380
rect 15520 -35480 15620 -35380
rect 17020 -35480 17120 -35380
rect 18520 -35480 18620 -35380
rect 20020 -35480 20120 -35380
rect 21520 -35480 21620 -35380
rect 23020 -35480 23120 -35380
rect 24520 -35480 24620 -35380
rect 26020 -35480 26120 -35380
rect 27520 -35480 27620 -35380
rect 29020 -35480 29120 -35380
rect 30520 -35480 30620 -35380
rect 32020 -35480 32120 -35380
rect 33520 -35480 33620 -35380
rect 35020 -35480 35120 -35380
rect 36520 -35480 36620 -35380
rect 38020 -35480 38120 -35380
rect 39520 -35480 39620 -35380
rect 41020 -35480 41120 -35380
rect 42520 -35480 42620 -35380
rect 44020 -35480 44120 -35380
rect 45520 -35480 45620 -35380
rect 47020 -35480 47120 -35380
rect 48520 -35480 48620 -35380
rect 50020 -35480 50120 -35380
rect 51520 -35480 51620 -35380
rect 53020 -35480 53120 -35380
rect 54520 -35480 54620 -35380
rect 56020 -35480 56120 -35380
rect 57520 -35480 57620 -35380
rect 59020 -35480 59120 -35380
rect 60520 -35480 60620 -35380
rect 62020 -35480 62120 -35380
rect 63520 -35480 63620 -35380
rect 65020 -35480 65120 -35380
rect 66520 -35480 66620 -35380
rect 68020 -35480 68120 -35380
rect 69520 -35480 69620 -35380
rect 71020 -35480 71120 -35380
rect 72520 -35480 72620 -35380
rect 74020 -35480 74120 -35380
rect 75520 -35480 75620 -35380
rect 77020 -35480 77120 -35380
rect 78520 -35480 78620 -35380
rect 80020 -35480 80120 -35380
rect 81520 -35480 81620 -35380
rect 83020 -35480 83120 -35380
rect 84520 -35480 84620 -35380
rect 86020 -35480 86120 -35380
rect 87520 -35480 87620 -35380
rect 89020 -35480 89120 -35380
rect 90520 -35480 90620 -35380
rect 92020 -35480 92120 -35380
rect 93520 -35480 93620 -35380
rect 95020 -35480 95120 -35380
rect 96520 -35480 96620 -35380
rect 98020 -35480 98120 -35380
rect 99520 -35480 99620 -35380
rect 101020 -35480 101120 -35380
rect 102520 -35480 102620 -35380
rect 104020 -35480 104120 -35380
rect 105520 -35480 105620 -35380
rect 107020 -35480 107120 -35380
rect 108520 -35480 108620 -35380
rect 110020 -35480 110120 -35380
rect 111520 -35480 111620 -35380
rect 113020 -35480 113120 -35380
rect 114520 -35480 114620 -35380
rect 116020 -35480 116120 -35380
rect 117520 -35480 117620 -35380
rect 119020 -35480 119120 -35380
rect 520 -36980 620 -36880
rect 2020 -36980 2120 -36880
rect 3520 -36980 3620 -36880
rect 5020 -36980 5120 -36880
rect 6520 -36980 6620 -36880
rect 8020 -36980 8120 -36880
rect 9520 -36980 9620 -36880
rect 11020 -36980 11120 -36880
rect 12520 -36980 12620 -36880
rect 14020 -36980 14120 -36880
rect 15520 -36980 15620 -36880
rect 17020 -36980 17120 -36880
rect 18520 -36980 18620 -36880
rect 20020 -36980 20120 -36880
rect 21520 -36980 21620 -36880
rect 23020 -36980 23120 -36880
rect 24520 -36980 24620 -36880
rect 26020 -36980 26120 -36880
rect 27520 -36980 27620 -36880
rect 29020 -36980 29120 -36880
rect 30520 -36980 30620 -36880
rect 32020 -36980 32120 -36880
rect 33520 -36980 33620 -36880
rect 35020 -36980 35120 -36880
rect 36520 -36980 36620 -36880
rect 38020 -36980 38120 -36880
rect 39520 -36980 39620 -36880
rect 41020 -36980 41120 -36880
rect 42520 -36980 42620 -36880
rect 44020 -36980 44120 -36880
rect 45520 -36980 45620 -36880
rect 47020 -36980 47120 -36880
rect 48520 -36980 48620 -36880
rect 50020 -36980 50120 -36880
rect 51520 -36980 51620 -36880
rect 53020 -36980 53120 -36880
rect 54520 -36980 54620 -36880
rect 56020 -36980 56120 -36880
rect 57520 -36980 57620 -36880
rect 59020 -36980 59120 -36880
rect 60520 -36980 60620 -36880
rect 62020 -36980 62120 -36880
rect 63520 -36980 63620 -36880
rect 65020 -36980 65120 -36880
rect 66520 -36980 66620 -36880
rect 68020 -36980 68120 -36880
rect 69520 -36980 69620 -36880
rect 71020 -36980 71120 -36880
rect 72520 -36980 72620 -36880
rect 74020 -36980 74120 -36880
rect 75520 -36980 75620 -36880
rect 77020 -36980 77120 -36880
rect 78520 -36980 78620 -36880
rect 80020 -36980 80120 -36880
rect 81520 -36980 81620 -36880
rect 83020 -36980 83120 -36880
rect 84520 -36980 84620 -36880
rect 86020 -36980 86120 -36880
rect 87520 -36980 87620 -36880
rect 89020 -36980 89120 -36880
rect 90520 -36980 90620 -36880
rect 92020 -36980 92120 -36880
rect 93520 -36980 93620 -36880
rect 95020 -36980 95120 -36880
rect 96520 -36980 96620 -36880
rect 98020 -36980 98120 -36880
rect 99520 -36980 99620 -36880
rect 101020 -36980 101120 -36880
rect 102520 -36980 102620 -36880
rect 104020 -36980 104120 -36880
rect 105520 -36980 105620 -36880
rect 107020 -36980 107120 -36880
rect 108520 -36980 108620 -36880
rect 110020 -36980 110120 -36880
rect 111520 -36980 111620 -36880
rect 113020 -36980 113120 -36880
rect 114520 -36980 114620 -36880
rect 116020 -36980 116120 -36880
rect 117520 -36980 117620 -36880
rect 119020 -36980 119120 -36880
rect 520 -38480 620 -38380
rect 2020 -38480 2120 -38380
rect 3520 -38480 3620 -38380
rect 5020 -38480 5120 -38380
rect 6520 -38480 6620 -38380
rect 8020 -38480 8120 -38380
rect 9520 -38480 9620 -38380
rect 11020 -38480 11120 -38380
rect 12520 -38480 12620 -38380
rect 14020 -38480 14120 -38380
rect 15520 -38480 15620 -38380
rect 17020 -38480 17120 -38380
rect 18520 -38480 18620 -38380
rect 20020 -38480 20120 -38380
rect 21520 -38480 21620 -38380
rect 23020 -38480 23120 -38380
rect 24520 -38480 24620 -38380
rect 26020 -38480 26120 -38380
rect 27520 -38480 27620 -38380
rect 29020 -38480 29120 -38380
rect 30520 -38480 30620 -38380
rect 32020 -38480 32120 -38380
rect 33520 -38480 33620 -38380
rect 35020 -38480 35120 -38380
rect 36520 -38480 36620 -38380
rect 38020 -38480 38120 -38380
rect 39520 -38480 39620 -38380
rect 41020 -38480 41120 -38380
rect 42520 -38480 42620 -38380
rect 44020 -38480 44120 -38380
rect 45520 -38480 45620 -38380
rect 47020 -38480 47120 -38380
rect 48520 -38480 48620 -38380
rect 50020 -38480 50120 -38380
rect 51520 -38480 51620 -38380
rect 53020 -38480 53120 -38380
rect 54520 -38480 54620 -38380
rect 56020 -38480 56120 -38380
rect 57520 -38480 57620 -38380
rect 59020 -38480 59120 -38380
rect 60520 -38480 60620 -38380
rect 62020 -38480 62120 -38380
rect 63520 -38480 63620 -38380
rect 65020 -38480 65120 -38380
rect 66520 -38480 66620 -38380
rect 68020 -38480 68120 -38380
rect 69520 -38480 69620 -38380
rect 71020 -38480 71120 -38380
rect 72520 -38480 72620 -38380
rect 74020 -38480 74120 -38380
rect 75520 -38480 75620 -38380
rect 77020 -38480 77120 -38380
rect 78520 -38480 78620 -38380
rect 80020 -38480 80120 -38380
rect 81520 -38480 81620 -38380
rect 83020 -38480 83120 -38380
rect 84520 -38480 84620 -38380
rect 86020 -38480 86120 -38380
rect 87520 -38480 87620 -38380
rect 89020 -38480 89120 -38380
rect 90520 -38480 90620 -38380
rect 92020 -38480 92120 -38380
rect 93520 -38480 93620 -38380
rect 95020 -38480 95120 -38380
rect 96520 -38480 96620 -38380
rect 98020 -38480 98120 -38380
rect 99520 -38480 99620 -38380
rect 101020 -38480 101120 -38380
rect 102520 -38480 102620 -38380
rect 104020 -38480 104120 -38380
rect 105520 -38480 105620 -38380
rect 107020 -38480 107120 -38380
rect 108520 -38480 108620 -38380
rect 110020 -38480 110120 -38380
rect 111520 -38480 111620 -38380
rect 113020 -38480 113120 -38380
rect 114520 -38480 114620 -38380
rect 116020 -38480 116120 -38380
rect 117520 -38480 117620 -38380
rect 119020 -38480 119120 -38380
rect 520 -39980 620 -39880
rect 2020 -39980 2120 -39880
rect 3520 -39980 3620 -39880
rect 5020 -39980 5120 -39880
rect 6520 -39980 6620 -39880
rect 8020 -39980 8120 -39880
rect 9520 -39980 9620 -39880
rect 11020 -39980 11120 -39880
rect 12520 -39980 12620 -39880
rect 14020 -39980 14120 -39880
rect 15520 -39980 15620 -39880
rect 17020 -39980 17120 -39880
rect 18520 -39980 18620 -39880
rect 20020 -39980 20120 -39880
rect 21520 -39980 21620 -39880
rect 23020 -39980 23120 -39880
rect 24520 -39980 24620 -39880
rect 26020 -39980 26120 -39880
rect 27520 -39980 27620 -39880
rect 29020 -39980 29120 -39880
rect 30520 -39980 30620 -39880
rect 32020 -39980 32120 -39880
rect 33520 -39980 33620 -39880
rect 35020 -39980 35120 -39880
rect 36520 -39980 36620 -39880
rect 38020 -39980 38120 -39880
rect 39520 -39980 39620 -39880
rect 41020 -39980 41120 -39880
rect 42520 -39980 42620 -39880
rect 44020 -39980 44120 -39880
rect 45520 -39980 45620 -39880
rect 47020 -39980 47120 -39880
rect 48520 -39980 48620 -39880
rect 50020 -39980 50120 -39880
rect 51520 -39980 51620 -39880
rect 53020 -39980 53120 -39880
rect 54520 -39980 54620 -39880
rect 56020 -39980 56120 -39880
rect 57520 -39980 57620 -39880
rect 59020 -39980 59120 -39880
rect 60520 -39980 60620 -39880
rect 62020 -39980 62120 -39880
rect 63520 -39980 63620 -39880
rect 65020 -39980 65120 -39880
rect 66520 -39980 66620 -39880
rect 68020 -39980 68120 -39880
rect 69520 -39980 69620 -39880
rect 71020 -39980 71120 -39880
rect 72520 -39980 72620 -39880
rect 74020 -39980 74120 -39880
rect 75520 -39980 75620 -39880
rect 77020 -39980 77120 -39880
rect 78520 -39980 78620 -39880
rect 80020 -39980 80120 -39880
rect 81520 -39980 81620 -39880
rect 83020 -39980 83120 -39880
rect 84520 -39980 84620 -39880
rect 86020 -39980 86120 -39880
rect 87520 -39980 87620 -39880
rect 89020 -39980 89120 -39880
rect 90520 -39980 90620 -39880
rect 92020 -39980 92120 -39880
rect 93520 -39980 93620 -39880
rect 95020 -39980 95120 -39880
rect 96520 -39980 96620 -39880
rect 98020 -39980 98120 -39880
rect 99520 -39980 99620 -39880
rect 101020 -39980 101120 -39880
rect 102520 -39980 102620 -39880
rect 104020 -39980 104120 -39880
rect 105520 -39980 105620 -39880
rect 107020 -39980 107120 -39880
rect 108520 -39980 108620 -39880
rect 110020 -39980 110120 -39880
rect 111520 -39980 111620 -39880
rect 113020 -39980 113120 -39880
rect 114520 -39980 114620 -39880
rect 116020 -39980 116120 -39880
rect 117520 -39980 117620 -39880
rect 119020 -39980 119120 -39880
rect 520 -41480 620 -41380
rect 2020 -41480 2120 -41380
rect 3520 -41480 3620 -41380
rect 5020 -41480 5120 -41380
rect 6520 -41480 6620 -41380
rect 8020 -41480 8120 -41380
rect 9520 -41480 9620 -41380
rect 11020 -41480 11120 -41380
rect 12520 -41480 12620 -41380
rect 14020 -41480 14120 -41380
rect 15520 -41480 15620 -41380
rect 17020 -41480 17120 -41380
rect 18520 -41480 18620 -41380
rect 20020 -41480 20120 -41380
rect 21520 -41480 21620 -41380
rect 23020 -41480 23120 -41380
rect 24520 -41480 24620 -41380
rect 26020 -41480 26120 -41380
rect 27520 -41480 27620 -41380
rect 29020 -41480 29120 -41380
rect 30520 -41480 30620 -41380
rect 32020 -41480 32120 -41380
rect 33520 -41480 33620 -41380
rect 35020 -41480 35120 -41380
rect 36520 -41480 36620 -41380
rect 38020 -41480 38120 -41380
rect 39520 -41480 39620 -41380
rect 41020 -41480 41120 -41380
rect 42520 -41480 42620 -41380
rect 44020 -41480 44120 -41380
rect 45520 -41480 45620 -41380
rect 47020 -41480 47120 -41380
rect 48520 -41480 48620 -41380
rect 50020 -41480 50120 -41380
rect 51520 -41480 51620 -41380
rect 53020 -41480 53120 -41380
rect 54520 -41480 54620 -41380
rect 56020 -41480 56120 -41380
rect 57520 -41480 57620 -41380
rect 59020 -41480 59120 -41380
rect 60520 -41480 60620 -41380
rect 62020 -41480 62120 -41380
rect 63520 -41480 63620 -41380
rect 65020 -41480 65120 -41380
rect 66520 -41480 66620 -41380
rect 68020 -41480 68120 -41380
rect 69520 -41480 69620 -41380
rect 71020 -41480 71120 -41380
rect 72520 -41480 72620 -41380
rect 74020 -41480 74120 -41380
rect 75520 -41480 75620 -41380
rect 77020 -41480 77120 -41380
rect 78520 -41480 78620 -41380
rect 80020 -41480 80120 -41380
rect 81520 -41480 81620 -41380
rect 83020 -41480 83120 -41380
rect 84520 -41480 84620 -41380
rect 86020 -41480 86120 -41380
rect 87520 -41480 87620 -41380
rect 89020 -41480 89120 -41380
rect 90520 -41480 90620 -41380
rect 92020 -41480 92120 -41380
rect 93520 -41480 93620 -41380
rect 95020 -41480 95120 -41380
rect 96520 -41480 96620 -41380
rect 98020 -41480 98120 -41380
rect 99520 -41480 99620 -41380
rect 101020 -41480 101120 -41380
rect 102520 -41480 102620 -41380
rect 104020 -41480 104120 -41380
rect 105520 -41480 105620 -41380
rect 107020 -41480 107120 -41380
rect 108520 -41480 108620 -41380
rect 110020 -41480 110120 -41380
rect 111520 -41480 111620 -41380
rect 113020 -41480 113120 -41380
rect 114520 -41480 114620 -41380
rect 116020 -41480 116120 -41380
rect 117520 -41480 117620 -41380
rect 119020 -41480 119120 -41380
rect 520 -42980 620 -42880
rect 2020 -42980 2120 -42880
rect 3520 -42980 3620 -42880
rect 5020 -42980 5120 -42880
rect 6520 -42980 6620 -42880
rect 8020 -42980 8120 -42880
rect 9520 -42980 9620 -42880
rect 11020 -42980 11120 -42880
rect 12520 -42980 12620 -42880
rect 14020 -42980 14120 -42880
rect 15520 -42980 15620 -42880
rect 17020 -42980 17120 -42880
rect 18520 -42980 18620 -42880
rect 20020 -42980 20120 -42880
rect 21520 -42980 21620 -42880
rect 23020 -42980 23120 -42880
rect 24520 -42980 24620 -42880
rect 26020 -42980 26120 -42880
rect 27520 -42980 27620 -42880
rect 29020 -42980 29120 -42880
rect 30520 -42980 30620 -42880
rect 32020 -42980 32120 -42880
rect 33520 -42980 33620 -42880
rect 35020 -42980 35120 -42880
rect 36520 -42980 36620 -42880
rect 38020 -42980 38120 -42880
rect 39520 -42980 39620 -42880
rect 41020 -42980 41120 -42880
rect 42520 -42980 42620 -42880
rect 44020 -42980 44120 -42880
rect 45520 -42980 45620 -42880
rect 47020 -42980 47120 -42880
rect 48520 -42980 48620 -42880
rect 50020 -42980 50120 -42880
rect 51520 -42980 51620 -42880
rect 53020 -42980 53120 -42880
rect 54520 -42980 54620 -42880
rect 56020 -42980 56120 -42880
rect 57520 -42980 57620 -42880
rect 59020 -42980 59120 -42880
rect 60520 -42980 60620 -42880
rect 62020 -42980 62120 -42880
rect 63520 -42980 63620 -42880
rect 65020 -42980 65120 -42880
rect 66520 -42980 66620 -42880
rect 68020 -42980 68120 -42880
rect 69520 -42980 69620 -42880
rect 71020 -42980 71120 -42880
rect 72520 -42980 72620 -42880
rect 74020 -42980 74120 -42880
rect 75520 -42980 75620 -42880
rect 77020 -42980 77120 -42880
rect 78520 -42980 78620 -42880
rect 80020 -42980 80120 -42880
rect 81520 -42980 81620 -42880
rect 83020 -42980 83120 -42880
rect 84520 -42980 84620 -42880
rect 86020 -42980 86120 -42880
rect 87520 -42980 87620 -42880
rect 89020 -42980 89120 -42880
rect 90520 -42980 90620 -42880
rect 92020 -42980 92120 -42880
rect 93520 -42980 93620 -42880
rect 95020 -42980 95120 -42880
rect 96520 -42980 96620 -42880
rect 98020 -42980 98120 -42880
rect 99520 -42980 99620 -42880
rect 101020 -42980 101120 -42880
rect 102520 -42980 102620 -42880
rect 104020 -42980 104120 -42880
rect 105520 -42980 105620 -42880
rect 107020 -42980 107120 -42880
rect 108520 -42980 108620 -42880
rect 110020 -42980 110120 -42880
rect 111520 -42980 111620 -42880
rect 113020 -42980 113120 -42880
rect 114520 -42980 114620 -42880
rect 116020 -42980 116120 -42880
rect 117520 -42980 117620 -42880
rect 119020 -42980 119120 -42880
rect 520 -44480 620 -44380
rect 2020 -44480 2120 -44380
rect 3520 -44480 3620 -44380
rect 5020 -44480 5120 -44380
rect 6520 -44480 6620 -44380
rect 8020 -44480 8120 -44380
rect 9520 -44480 9620 -44380
rect 11020 -44480 11120 -44380
rect 12520 -44480 12620 -44380
rect 14020 -44480 14120 -44380
rect 15520 -44480 15620 -44380
rect 17020 -44480 17120 -44380
rect 18520 -44480 18620 -44380
rect 20020 -44480 20120 -44380
rect 21520 -44480 21620 -44380
rect 23020 -44480 23120 -44380
rect 24520 -44480 24620 -44380
rect 26020 -44480 26120 -44380
rect 27520 -44480 27620 -44380
rect 29020 -44480 29120 -44380
rect 30520 -44480 30620 -44380
rect 32020 -44480 32120 -44380
rect 33520 -44480 33620 -44380
rect 35020 -44480 35120 -44380
rect 36520 -44480 36620 -44380
rect 38020 -44480 38120 -44380
rect 39520 -44480 39620 -44380
rect 41020 -44480 41120 -44380
rect 42520 -44480 42620 -44380
rect 44020 -44480 44120 -44380
rect 45520 -44480 45620 -44380
rect 47020 -44480 47120 -44380
rect 48520 -44480 48620 -44380
rect 50020 -44480 50120 -44380
rect 51520 -44480 51620 -44380
rect 53020 -44480 53120 -44380
rect 54520 -44480 54620 -44380
rect 56020 -44480 56120 -44380
rect 57520 -44480 57620 -44380
rect 59020 -44480 59120 -44380
rect 60520 -44480 60620 -44380
rect 62020 -44480 62120 -44380
rect 63520 -44480 63620 -44380
rect 65020 -44480 65120 -44380
rect 66520 -44480 66620 -44380
rect 68020 -44480 68120 -44380
rect 69520 -44480 69620 -44380
rect 71020 -44480 71120 -44380
rect 72520 -44480 72620 -44380
rect 74020 -44480 74120 -44380
rect 75520 -44480 75620 -44380
rect 77020 -44480 77120 -44380
rect 78520 -44480 78620 -44380
rect 80020 -44480 80120 -44380
rect 81520 -44480 81620 -44380
rect 83020 -44480 83120 -44380
rect 84520 -44480 84620 -44380
rect 86020 -44480 86120 -44380
rect 87520 -44480 87620 -44380
rect 89020 -44480 89120 -44380
rect 90520 -44480 90620 -44380
rect 92020 -44480 92120 -44380
rect 93520 -44480 93620 -44380
rect 95020 -44480 95120 -44380
rect 96520 -44480 96620 -44380
rect 98020 -44480 98120 -44380
rect 99520 -44480 99620 -44380
rect 101020 -44480 101120 -44380
rect 102520 -44480 102620 -44380
rect 104020 -44480 104120 -44380
rect 105520 -44480 105620 -44380
rect 107020 -44480 107120 -44380
rect 108520 -44480 108620 -44380
rect 110020 -44480 110120 -44380
rect 111520 -44480 111620 -44380
rect 113020 -44480 113120 -44380
rect 114520 -44480 114620 -44380
rect 116020 -44480 116120 -44380
rect 117520 -44480 117620 -44380
rect 119020 -44480 119120 -44380
rect 520 -45980 620 -45880
rect 2020 -45980 2120 -45880
rect 3520 -45980 3620 -45880
rect 5020 -45980 5120 -45880
rect 6520 -45980 6620 -45880
rect 8020 -45980 8120 -45880
rect 9520 -45980 9620 -45880
rect 11020 -45980 11120 -45880
rect 12520 -45980 12620 -45880
rect 14020 -45980 14120 -45880
rect 15520 -45980 15620 -45880
rect 17020 -45980 17120 -45880
rect 18520 -45980 18620 -45880
rect 20020 -45980 20120 -45880
rect 21520 -45980 21620 -45880
rect 23020 -45980 23120 -45880
rect 24520 -45980 24620 -45880
rect 26020 -45980 26120 -45880
rect 27520 -45980 27620 -45880
rect 29020 -45980 29120 -45880
rect 30520 -45980 30620 -45880
rect 32020 -45980 32120 -45880
rect 33520 -45980 33620 -45880
rect 35020 -45980 35120 -45880
rect 36520 -45980 36620 -45880
rect 38020 -45980 38120 -45880
rect 39520 -45980 39620 -45880
rect 41020 -45980 41120 -45880
rect 42520 -45980 42620 -45880
rect 44020 -45980 44120 -45880
rect 45520 -45980 45620 -45880
rect 47020 -45980 47120 -45880
rect 48520 -45980 48620 -45880
rect 50020 -45980 50120 -45880
rect 51520 -45980 51620 -45880
rect 53020 -45980 53120 -45880
rect 54520 -45980 54620 -45880
rect 56020 -45980 56120 -45880
rect 57520 -45980 57620 -45880
rect 59020 -45980 59120 -45880
rect 60520 -45980 60620 -45880
rect 62020 -45980 62120 -45880
rect 63520 -45980 63620 -45880
rect 65020 -45980 65120 -45880
rect 66520 -45980 66620 -45880
rect 68020 -45980 68120 -45880
rect 69520 -45980 69620 -45880
rect 71020 -45980 71120 -45880
rect 72520 -45980 72620 -45880
rect 74020 -45980 74120 -45880
rect 75520 -45980 75620 -45880
rect 77020 -45980 77120 -45880
rect 78520 -45980 78620 -45880
rect 80020 -45980 80120 -45880
rect 81520 -45980 81620 -45880
rect 83020 -45980 83120 -45880
rect 84520 -45980 84620 -45880
rect 86020 -45980 86120 -45880
rect 87520 -45980 87620 -45880
rect 89020 -45980 89120 -45880
rect 90520 -45980 90620 -45880
rect 92020 -45980 92120 -45880
rect 93520 -45980 93620 -45880
rect 95020 -45980 95120 -45880
rect 96520 -45980 96620 -45880
rect 98020 -45980 98120 -45880
rect 99520 -45980 99620 -45880
rect 101020 -45980 101120 -45880
rect 102520 -45980 102620 -45880
rect 104020 -45980 104120 -45880
rect 105520 -45980 105620 -45880
rect 107020 -45980 107120 -45880
rect 108520 -45980 108620 -45880
rect 110020 -45980 110120 -45880
rect 111520 -45980 111620 -45880
rect 113020 -45980 113120 -45880
rect 114520 -45980 114620 -45880
rect 116020 -45980 116120 -45880
rect 117520 -45980 117620 -45880
rect 119020 -45980 119120 -45880
rect 520 -47480 620 -47380
rect 2020 -47480 2120 -47380
rect 3520 -47480 3620 -47380
rect 5020 -47480 5120 -47380
rect 6520 -47480 6620 -47380
rect 8020 -47480 8120 -47380
rect 9520 -47480 9620 -47380
rect 11020 -47480 11120 -47380
rect 12520 -47480 12620 -47380
rect 14020 -47480 14120 -47380
rect 15520 -47480 15620 -47380
rect 17020 -47480 17120 -47380
rect 18520 -47480 18620 -47380
rect 20020 -47480 20120 -47380
rect 21520 -47480 21620 -47380
rect 23020 -47480 23120 -47380
rect 24520 -47480 24620 -47380
rect 26020 -47480 26120 -47380
rect 27520 -47480 27620 -47380
rect 29020 -47480 29120 -47380
rect 30520 -47480 30620 -47380
rect 32020 -47480 32120 -47380
rect 33520 -47480 33620 -47380
rect 35020 -47480 35120 -47380
rect 36520 -47480 36620 -47380
rect 38020 -47480 38120 -47380
rect 39520 -47480 39620 -47380
rect 41020 -47480 41120 -47380
rect 42520 -47480 42620 -47380
rect 44020 -47480 44120 -47380
rect 45520 -47480 45620 -47380
rect 47020 -47480 47120 -47380
rect 48520 -47480 48620 -47380
rect 50020 -47480 50120 -47380
rect 51520 -47480 51620 -47380
rect 53020 -47480 53120 -47380
rect 54520 -47480 54620 -47380
rect 56020 -47480 56120 -47380
rect 57520 -47480 57620 -47380
rect 59020 -47480 59120 -47380
rect 60520 -47480 60620 -47380
rect 62020 -47480 62120 -47380
rect 63520 -47480 63620 -47380
rect 65020 -47480 65120 -47380
rect 66520 -47480 66620 -47380
rect 68020 -47480 68120 -47380
rect 69520 -47480 69620 -47380
rect 71020 -47480 71120 -47380
rect 72520 -47480 72620 -47380
rect 74020 -47480 74120 -47380
rect 75520 -47480 75620 -47380
rect 77020 -47480 77120 -47380
rect 78520 -47480 78620 -47380
rect 80020 -47480 80120 -47380
rect 81520 -47480 81620 -47380
rect 83020 -47480 83120 -47380
rect 84520 -47480 84620 -47380
rect 86020 -47480 86120 -47380
rect 87520 -47480 87620 -47380
rect 89020 -47480 89120 -47380
rect 90520 -47480 90620 -47380
rect 92020 -47480 92120 -47380
rect 93520 -47480 93620 -47380
rect 95020 -47480 95120 -47380
rect 96520 -47480 96620 -47380
rect 98020 -47480 98120 -47380
rect 99520 -47480 99620 -47380
rect 101020 -47480 101120 -47380
rect 102520 -47480 102620 -47380
rect 104020 -47480 104120 -47380
rect 105520 -47480 105620 -47380
rect 107020 -47480 107120 -47380
rect 108520 -47480 108620 -47380
rect 110020 -47480 110120 -47380
rect 111520 -47480 111620 -47380
rect 113020 -47480 113120 -47380
rect 114520 -47480 114620 -47380
rect 116020 -47480 116120 -47380
rect 117520 -47480 117620 -47380
rect 119020 -47480 119120 -47380
rect 520 -48980 620 -48880
rect 2020 -48980 2120 -48880
rect 3520 -48980 3620 -48880
rect 5020 -48980 5120 -48880
rect 6520 -48980 6620 -48880
rect 8020 -48980 8120 -48880
rect 9520 -48980 9620 -48880
rect 11020 -48980 11120 -48880
rect 12520 -48980 12620 -48880
rect 14020 -48980 14120 -48880
rect 15520 -48980 15620 -48880
rect 17020 -48980 17120 -48880
rect 18520 -48980 18620 -48880
rect 20020 -48980 20120 -48880
rect 21520 -48980 21620 -48880
rect 23020 -48980 23120 -48880
rect 24520 -48980 24620 -48880
rect 26020 -48980 26120 -48880
rect 27520 -48980 27620 -48880
rect 29020 -48980 29120 -48880
rect 30520 -48980 30620 -48880
rect 32020 -48980 32120 -48880
rect 33520 -48980 33620 -48880
rect 35020 -48980 35120 -48880
rect 36520 -48980 36620 -48880
rect 38020 -48980 38120 -48880
rect 39520 -48980 39620 -48880
rect 41020 -48980 41120 -48880
rect 42520 -48980 42620 -48880
rect 44020 -48980 44120 -48880
rect 45520 -48980 45620 -48880
rect 47020 -48980 47120 -48880
rect 48520 -48980 48620 -48880
rect 50020 -48980 50120 -48880
rect 51520 -48980 51620 -48880
rect 53020 -48980 53120 -48880
rect 54520 -48980 54620 -48880
rect 56020 -48980 56120 -48880
rect 57520 -48980 57620 -48880
rect 59020 -48980 59120 -48880
rect 60520 -48980 60620 -48880
rect 62020 -48980 62120 -48880
rect 63520 -48980 63620 -48880
rect 65020 -48980 65120 -48880
rect 66520 -48980 66620 -48880
rect 68020 -48980 68120 -48880
rect 69520 -48980 69620 -48880
rect 71020 -48980 71120 -48880
rect 72520 -48980 72620 -48880
rect 74020 -48980 74120 -48880
rect 75520 -48980 75620 -48880
rect 77020 -48980 77120 -48880
rect 78520 -48980 78620 -48880
rect 80020 -48980 80120 -48880
rect 81520 -48980 81620 -48880
rect 83020 -48980 83120 -48880
rect 84520 -48980 84620 -48880
rect 86020 -48980 86120 -48880
rect 87520 -48980 87620 -48880
rect 89020 -48980 89120 -48880
rect 90520 -48980 90620 -48880
rect 92020 -48980 92120 -48880
rect 93520 -48980 93620 -48880
rect 95020 -48980 95120 -48880
rect 96520 -48980 96620 -48880
rect 98020 -48980 98120 -48880
rect 99520 -48980 99620 -48880
rect 101020 -48980 101120 -48880
rect 102520 -48980 102620 -48880
rect 104020 -48980 104120 -48880
rect 105520 -48980 105620 -48880
rect 107020 -48980 107120 -48880
rect 108520 -48980 108620 -48880
rect 110020 -48980 110120 -48880
rect 111520 -48980 111620 -48880
rect 113020 -48980 113120 -48880
rect 114520 -48980 114620 -48880
rect 116020 -48980 116120 -48880
rect 117520 -48980 117620 -48880
rect 119020 -48980 119120 -48880
rect 520 -50480 620 -50380
rect 2020 -50480 2120 -50380
rect 3520 -50480 3620 -50380
rect 5020 -50480 5120 -50380
rect 6520 -50480 6620 -50380
rect 8020 -50480 8120 -50380
rect 9520 -50480 9620 -50380
rect 11020 -50480 11120 -50380
rect 12520 -50480 12620 -50380
rect 14020 -50480 14120 -50380
rect 15520 -50480 15620 -50380
rect 17020 -50480 17120 -50380
rect 18520 -50480 18620 -50380
rect 20020 -50480 20120 -50380
rect 21520 -50480 21620 -50380
rect 23020 -50480 23120 -50380
rect 24520 -50480 24620 -50380
rect 26020 -50480 26120 -50380
rect 27520 -50480 27620 -50380
rect 29020 -50480 29120 -50380
rect 30520 -50480 30620 -50380
rect 32020 -50480 32120 -50380
rect 33520 -50480 33620 -50380
rect 35020 -50480 35120 -50380
rect 36520 -50480 36620 -50380
rect 38020 -50480 38120 -50380
rect 39520 -50480 39620 -50380
rect 41020 -50480 41120 -50380
rect 42520 -50480 42620 -50380
rect 44020 -50480 44120 -50380
rect 45520 -50480 45620 -50380
rect 47020 -50480 47120 -50380
rect 48520 -50480 48620 -50380
rect 50020 -50480 50120 -50380
rect 51520 -50480 51620 -50380
rect 53020 -50480 53120 -50380
rect 54520 -50480 54620 -50380
rect 56020 -50480 56120 -50380
rect 57520 -50480 57620 -50380
rect 59020 -50480 59120 -50380
rect 60520 -50480 60620 -50380
rect 62020 -50480 62120 -50380
rect 63520 -50480 63620 -50380
rect 65020 -50480 65120 -50380
rect 66520 -50480 66620 -50380
rect 68020 -50480 68120 -50380
rect 69520 -50480 69620 -50380
rect 71020 -50480 71120 -50380
rect 72520 -50480 72620 -50380
rect 74020 -50480 74120 -50380
rect 75520 -50480 75620 -50380
rect 77020 -50480 77120 -50380
rect 78520 -50480 78620 -50380
rect 80020 -50480 80120 -50380
rect 81520 -50480 81620 -50380
rect 83020 -50480 83120 -50380
rect 84520 -50480 84620 -50380
rect 86020 -50480 86120 -50380
rect 87520 -50480 87620 -50380
rect 89020 -50480 89120 -50380
rect 90520 -50480 90620 -50380
rect 92020 -50480 92120 -50380
rect 93520 -50480 93620 -50380
rect 95020 -50480 95120 -50380
rect 96520 -50480 96620 -50380
rect 98020 -50480 98120 -50380
rect 99520 -50480 99620 -50380
rect 101020 -50480 101120 -50380
rect 102520 -50480 102620 -50380
rect 104020 -50480 104120 -50380
rect 105520 -50480 105620 -50380
rect 107020 -50480 107120 -50380
rect 108520 -50480 108620 -50380
rect 110020 -50480 110120 -50380
rect 111520 -50480 111620 -50380
rect 113020 -50480 113120 -50380
rect 114520 -50480 114620 -50380
rect 116020 -50480 116120 -50380
rect 117520 -50480 117620 -50380
rect 119020 -50480 119120 -50380
rect 520 -51980 620 -51880
rect 2020 -51980 2120 -51880
rect 3520 -51980 3620 -51880
rect 5020 -51980 5120 -51880
rect 6520 -51980 6620 -51880
rect 8020 -51980 8120 -51880
rect 9520 -51980 9620 -51880
rect 11020 -51980 11120 -51880
rect 12520 -51980 12620 -51880
rect 14020 -51980 14120 -51880
rect 15520 -51980 15620 -51880
rect 17020 -51980 17120 -51880
rect 18520 -51980 18620 -51880
rect 20020 -51980 20120 -51880
rect 21520 -51980 21620 -51880
rect 23020 -51980 23120 -51880
rect 24520 -51980 24620 -51880
rect 26020 -51980 26120 -51880
rect 27520 -51980 27620 -51880
rect 29020 -51980 29120 -51880
rect 30520 -51980 30620 -51880
rect 32020 -51980 32120 -51880
rect 33520 -51980 33620 -51880
rect 35020 -51980 35120 -51880
rect 36520 -51980 36620 -51880
rect 38020 -51980 38120 -51880
rect 39520 -51980 39620 -51880
rect 41020 -51980 41120 -51880
rect 42520 -51980 42620 -51880
rect 44020 -51980 44120 -51880
rect 45520 -51980 45620 -51880
rect 47020 -51980 47120 -51880
rect 48520 -51980 48620 -51880
rect 50020 -51980 50120 -51880
rect 51520 -51980 51620 -51880
rect 53020 -51980 53120 -51880
rect 54520 -51980 54620 -51880
rect 56020 -51980 56120 -51880
rect 57520 -51980 57620 -51880
rect 59020 -51980 59120 -51880
rect 60520 -51980 60620 -51880
rect 62020 -51980 62120 -51880
rect 63520 -51980 63620 -51880
rect 65020 -51980 65120 -51880
rect 66520 -51980 66620 -51880
rect 68020 -51980 68120 -51880
rect 69520 -51980 69620 -51880
rect 71020 -51980 71120 -51880
rect 72520 -51980 72620 -51880
rect 74020 -51980 74120 -51880
rect 75520 -51980 75620 -51880
rect 77020 -51980 77120 -51880
rect 78520 -51980 78620 -51880
rect 80020 -51980 80120 -51880
rect 81520 -51980 81620 -51880
rect 83020 -51980 83120 -51880
rect 84520 -51980 84620 -51880
rect 86020 -51980 86120 -51880
rect 87520 -51980 87620 -51880
rect 89020 -51980 89120 -51880
rect 90520 -51980 90620 -51880
rect 92020 -51980 92120 -51880
rect 93520 -51980 93620 -51880
rect 95020 -51980 95120 -51880
rect 96520 -51980 96620 -51880
rect 98020 -51980 98120 -51880
rect 99520 -51980 99620 -51880
rect 101020 -51980 101120 -51880
rect 102520 -51980 102620 -51880
rect 104020 -51980 104120 -51880
rect 105520 -51980 105620 -51880
rect 107020 -51980 107120 -51880
rect 108520 -51980 108620 -51880
rect 110020 -51980 110120 -51880
rect 111520 -51980 111620 -51880
rect 113020 -51980 113120 -51880
rect 114520 -51980 114620 -51880
rect 116020 -51980 116120 -51880
rect 117520 -51980 117620 -51880
rect 119020 -51980 119120 -51880
rect 520 -53480 620 -53380
rect 2020 -53480 2120 -53380
rect 3520 -53480 3620 -53380
rect 5020 -53480 5120 -53380
rect 6520 -53480 6620 -53380
rect 8020 -53480 8120 -53380
rect 9520 -53480 9620 -53380
rect 11020 -53480 11120 -53380
rect 12520 -53480 12620 -53380
rect 14020 -53480 14120 -53380
rect 15520 -53480 15620 -53380
rect 17020 -53480 17120 -53380
rect 18520 -53480 18620 -53380
rect 20020 -53480 20120 -53380
rect 21520 -53480 21620 -53380
rect 23020 -53480 23120 -53380
rect 24520 -53480 24620 -53380
rect 26020 -53480 26120 -53380
rect 27520 -53480 27620 -53380
rect 29020 -53480 29120 -53380
rect 30520 -53480 30620 -53380
rect 32020 -53480 32120 -53380
rect 33520 -53480 33620 -53380
rect 35020 -53480 35120 -53380
rect 36520 -53480 36620 -53380
rect 38020 -53480 38120 -53380
rect 39520 -53480 39620 -53380
rect 41020 -53480 41120 -53380
rect 42520 -53480 42620 -53380
rect 44020 -53480 44120 -53380
rect 45520 -53480 45620 -53380
rect 47020 -53480 47120 -53380
rect 48520 -53480 48620 -53380
rect 50020 -53480 50120 -53380
rect 51520 -53480 51620 -53380
rect 53020 -53480 53120 -53380
rect 54520 -53480 54620 -53380
rect 56020 -53480 56120 -53380
rect 57520 -53480 57620 -53380
rect 59020 -53480 59120 -53380
rect 60520 -53480 60620 -53380
rect 62020 -53480 62120 -53380
rect 63520 -53480 63620 -53380
rect 65020 -53480 65120 -53380
rect 66520 -53480 66620 -53380
rect 68020 -53480 68120 -53380
rect 69520 -53480 69620 -53380
rect 71020 -53480 71120 -53380
rect 72520 -53480 72620 -53380
rect 74020 -53480 74120 -53380
rect 75520 -53480 75620 -53380
rect 77020 -53480 77120 -53380
rect 78520 -53480 78620 -53380
rect 80020 -53480 80120 -53380
rect 81520 -53480 81620 -53380
rect 83020 -53480 83120 -53380
rect 84520 -53480 84620 -53380
rect 86020 -53480 86120 -53380
rect 87520 -53480 87620 -53380
rect 89020 -53480 89120 -53380
rect 90520 -53480 90620 -53380
rect 92020 -53480 92120 -53380
rect 93520 -53480 93620 -53380
rect 95020 -53480 95120 -53380
rect 96520 -53480 96620 -53380
rect 98020 -53480 98120 -53380
rect 99520 -53480 99620 -53380
rect 101020 -53480 101120 -53380
rect 102520 -53480 102620 -53380
rect 104020 -53480 104120 -53380
rect 105520 -53480 105620 -53380
rect 107020 -53480 107120 -53380
rect 108520 -53480 108620 -53380
rect 110020 -53480 110120 -53380
rect 111520 -53480 111620 -53380
rect 113020 -53480 113120 -53380
rect 114520 -53480 114620 -53380
rect 116020 -53480 116120 -53380
rect 117520 -53480 117620 -53380
rect 119020 -53480 119120 -53380
rect 520 -54980 620 -54880
rect 2020 -54980 2120 -54880
rect 3520 -54980 3620 -54880
rect 5020 -54980 5120 -54880
rect 6520 -54980 6620 -54880
rect 8020 -54980 8120 -54880
rect 9520 -54980 9620 -54880
rect 11020 -54980 11120 -54880
rect 12520 -54980 12620 -54880
rect 14020 -54980 14120 -54880
rect 15520 -54980 15620 -54880
rect 17020 -54980 17120 -54880
rect 18520 -54980 18620 -54880
rect 20020 -54980 20120 -54880
rect 21520 -54980 21620 -54880
rect 23020 -54980 23120 -54880
rect 24520 -54980 24620 -54880
rect 26020 -54980 26120 -54880
rect 27520 -54980 27620 -54880
rect 29020 -54980 29120 -54880
rect 30520 -54980 30620 -54880
rect 32020 -54980 32120 -54880
rect 33520 -54980 33620 -54880
rect 35020 -54980 35120 -54880
rect 36520 -54980 36620 -54880
rect 38020 -54980 38120 -54880
rect 39520 -54980 39620 -54880
rect 41020 -54980 41120 -54880
rect 42520 -54980 42620 -54880
rect 44020 -54980 44120 -54880
rect 45520 -54980 45620 -54880
rect 47020 -54980 47120 -54880
rect 48520 -54980 48620 -54880
rect 50020 -54980 50120 -54880
rect 51520 -54980 51620 -54880
rect 53020 -54980 53120 -54880
rect 54520 -54980 54620 -54880
rect 56020 -54980 56120 -54880
rect 57520 -54980 57620 -54880
rect 59020 -54980 59120 -54880
rect 60520 -54980 60620 -54880
rect 62020 -54980 62120 -54880
rect 63520 -54980 63620 -54880
rect 65020 -54980 65120 -54880
rect 66520 -54980 66620 -54880
rect 68020 -54980 68120 -54880
rect 69520 -54980 69620 -54880
rect 71020 -54980 71120 -54880
rect 72520 -54980 72620 -54880
rect 74020 -54980 74120 -54880
rect 75520 -54980 75620 -54880
rect 77020 -54980 77120 -54880
rect 78520 -54980 78620 -54880
rect 80020 -54980 80120 -54880
rect 81520 -54980 81620 -54880
rect 83020 -54980 83120 -54880
rect 84520 -54980 84620 -54880
rect 86020 -54980 86120 -54880
rect 87520 -54980 87620 -54880
rect 89020 -54980 89120 -54880
rect 90520 -54980 90620 -54880
rect 92020 -54980 92120 -54880
rect 93520 -54980 93620 -54880
rect 95020 -54980 95120 -54880
rect 96520 -54980 96620 -54880
rect 98020 -54980 98120 -54880
rect 99520 -54980 99620 -54880
rect 101020 -54980 101120 -54880
rect 102520 -54980 102620 -54880
rect 104020 -54980 104120 -54880
rect 105520 -54980 105620 -54880
rect 107020 -54980 107120 -54880
rect 108520 -54980 108620 -54880
rect 110020 -54980 110120 -54880
rect 111520 -54980 111620 -54880
rect 113020 -54980 113120 -54880
rect 114520 -54980 114620 -54880
rect 116020 -54980 116120 -54880
rect 117520 -54980 117620 -54880
rect 119020 -54980 119120 -54880
rect 520 -56480 620 -56380
rect 2020 -56480 2120 -56380
rect 3520 -56480 3620 -56380
rect 5020 -56480 5120 -56380
rect 6520 -56480 6620 -56380
rect 8020 -56480 8120 -56380
rect 9520 -56480 9620 -56380
rect 11020 -56480 11120 -56380
rect 12520 -56480 12620 -56380
rect 14020 -56480 14120 -56380
rect 15520 -56480 15620 -56380
rect 17020 -56480 17120 -56380
rect 18520 -56480 18620 -56380
rect 20020 -56480 20120 -56380
rect 21520 -56480 21620 -56380
rect 23020 -56480 23120 -56380
rect 24520 -56480 24620 -56380
rect 26020 -56480 26120 -56380
rect 27520 -56480 27620 -56380
rect 29020 -56480 29120 -56380
rect 30520 -56480 30620 -56380
rect 32020 -56480 32120 -56380
rect 33520 -56480 33620 -56380
rect 35020 -56480 35120 -56380
rect 36520 -56480 36620 -56380
rect 38020 -56480 38120 -56380
rect 39520 -56480 39620 -56380
rect 41020 -56480 41120 -56380
rect 42520 -56480 42620 -56380
rect 44020 -56480 44120 -56380
rect 45520 -56480 45620 -56380
rect 47020 -56480 47120 -56380
rect 48520 -56480 48620 -56380
rect 50020 -56480 50120 -56380
rect 51520 -56480 51620 -56380
rect 53020 -56480 53120 -56380
rect 54520 -56480 54620 -56380
rect 56020 -56480 56120 -56380
rect 57520 -56480 57620 -56380
rect 59020 -56480 59120 -56380
rect 60520 -56480 60620 -56380
rect 62020 -56480 62120 -56380
rect 63520 -56480 63620 -56380
rect 65020 -56480 65120 -56380
rect 66520 -56480 66620 -56380
rect 68020 -56480 68120 -56380
rect 69520 -56480 69620 -56380
rect 71020 -56480 71120 -56380
rect 72520 -56480 72620 -56380
rect 74020 -56480 74120 -56380
rect 75520 -56480 75620 -56380
rect 77020 -56480 77120 -56380
rect 78520 -56480 78620 -56380
rect 80020 -56480 80120 -56380
rect 81520 -56480 81620 -56380
rect 83020 -56480 83120 -56380
rect 84520 -56480 84620 -56380
rect 86020 -56480 86120 -56380
rect 87520 -56480 87620 -56380
rect 89020 -56480 89120 -56380
rect 90520 -56480 90620 -56380
rect 92020 -56480 92120 -56380
rect 93520 -56480 93620 -56380
rect 95020 -56480 95120 -56380
rect 96520 -56480 96620 -56380
rect 98020 -56480 98120 -56380
rect 99520 -56480 99620 -56380
rect 101020 -56480 101120 -56380
rect 102520 -56480 102620 -56380
rect 104020 -56480 104120 -56380
rect 105520 -56480 105620 -56380
rect 107020 -56480 107120 -56380
rect 108520 -56480 108620 -56380
rect 110020 -56480 110120 -56380
rect 111520 -56480 111620 -56380
rect 113020 -56480 113120 -56380
rect 114520 -56480 114620 -56380
rect 116020 -56480 116120 -56380
rect 117520 -56480 117620 -56380
rect 119020 -56480 119120 -56380
rect 520 -57980 620 -57880
rect 2020 -57980 2120 -57880
rect 3520 -57980 3620 -57880
rect 5020 -57980 5120 -57880
rect 6520 -57980 6620 -57880
rect 8020 -57980 8120 -57880
rect 9520 -57980 9620 -57880
rect 11020 -57980 11120 -57880
rect 12520 -57980 12620 -57880
rect 14020 -57980 14120 -57880
rect 15520 -57980 15620 -57880
rect 17020 -57980 17120 -57880
rect 18520 -57980 18620 -57880
rect 20020 -57980 20120 -57880
rect 21520 -57980 21620 -57880
rect 23020 -57980 23120 -57880
rect 24520 -57980 24620 -57880
rect 26020 -57980 26120 -57880
rect 27520 -57980 27620 -57880
rect 29020 -57980 29120 -57880
rect 30520 -57980 30620 -57880
rect 32020 -57980 32120 -57880
rect 33520 -57980 33620 -57880
rect 35020 -57980 35120 -57880
rect 36520 -57980 36620 -57880
rect 38020 -57980 38120 -57880
rect 39520 -57980 39620 -57880
rect 41020 -57980 41120 -57880
rect 42520 -57980 42620 -57880
rect 44020 -57980 44120 -57880
rect 45520 -57980 45620 -57880
rect 47020 -57980 47120 -57880
rect 48520 -57980 48620 -57880
rect 50020 -57980 50120 -57880
rect 51520 -57980 51620 -57880
rect 53020 -57980 53120 -57880
rect 54520 -57980 54620 -57880
rect 56020 -57980 56120 -57880
rect 57520 -57980 57620 -57880
rect 59020 -57980 59120 -57880
rect 60520 -57980 60620 -57880
rect 62020 -57980 62120 -57880
rect 63520 -57980 63620 -57880
rect 65020 -57980 65120 -57880
rect 66520 -57980 66620 -57880
rect 68020 -57980 68120 -57880
rect 69520 -57980 69620 -57880
rect 71020 -57980 71120 -57880
rect 72520 -57980 72620 -57880
rect 74020 -57980 74120 -57880
rect 75520 -57980 75620 -57880
rect 77020 -57980 77120 -57880
rect 78520 -57980 78620 -57880
rect 80020 -57980 80120 -57880
rect 81520 -57980 81620 -57880
rect 83020 -57980 83120 -57880
rect 84520 -57980 84620 -57880
rect 86020 -57980 86120 -57880
rect 87520 -57980 87620 -57880
rect 89020 -57980 89120 -57880
rect 90520 -57980 90620 -57880
rect 92020 -57980 92120 -57880
rect 93520 -57980 93620 -57880
rect 95020 -57980 95120 -57880
rect 96520 -57980 96620 -57880
rect 98020 -57980 98120 -57880
rect 99520 -57980 99620 -57880
rect 101020 -57980 101120 -57880
rect 102520 -57980 102620 -57880
rect 104020 -57980 104120 -57880
rect 105520 -57980 105620 -57880
rect 107020 -57980 107120 -57880
rect 108520 -57980 108620 -57880
rect 110020 -57980 110120 -57880
rect 111520 -57980 111620 -57880
rect 113020 -57980 113120 -57880
rect 114520 -57980 114620 -57880
rect 116020 -57980 116120 -57880
rect 117520 -57980 117620 -57880
rect 119020 -57980 119120 -57880
rect 520 -59480 620 -59380
rect 2020 -59480 2120 -59380
rect 3520 -59480 3620 -59380
rect 5020 -59480 5120 -59380
rect 6520 -59480 6620 -59380
rect 8020 -59480 8120 -59380
rect 9520 -59480 9620 -59380
rect 11020 -59480 11120 -59380
rect 12520 -59480 12620 -59380
rect 14020 -59480 14120 -59380
rect 15520 -59480 15620 -59380
rect 17020 -59480 17120 -59380
rect 18520 -59480 18620 -59380
rect 20020 -59480 20120 -59380
rect 21520 -59480 21620 -59380
rect 23020 -59480 23120 -59380
rect 24520 -59480 24620 -59380
rect 26020 -59480 26120 -59380
rect 27520 -59480 27620 -59380
rect 29020 -59480 29120 -59380
rect 30520 -59480 30620 -59380
rect 32020 -59480 32120 -59380
rect 33520 -59480 33620 -59380
rect 35020 -59480 35120 -59380
rect 36520 -59480 36620 -59380
rect 38020 -59480 38120 -59380
rect 39520 -59480 39620 -59380
rect 41020 -59480 41120 -59380
rect 42520 -59480 42620 -59380
rect 44020 -59480 44120 -59380
rect 45520 -59480 45620 -59380
rect 47020 -59480 47120 -59380
rect 48520 -59480 48620 -59380
rect 50020 -59480 50120 -59380
rect 51520 -59480 51620 -59380
rect 53020 -59480 53120 -59380
rect 54520 -59480 54620 -59380
rect 56020 -59480 56120 -59380
rect 57520 -59480 57620 -59380
rect 59020 -59480 59120 -59380
rect 60520 -59480 60620 -59380
rect 62020 -59480 62120 -59380
rect 63520 -59480 63620 -59380
rect 65020 -59480 65120 -59380
rect 66520 -59480 66620 -59380
rect 68020 -59480 68120 -59380
rect 69520 -59480 69620 -59380
rect 71020 -59480 71120 -59380
rect 72520 -59480 72620 -59380
rect 74020 -59480 74120 -59380
rect 75520 -59480 75620 -59380
rect 77020 -59480 77120 -59380
rect 78520 -59480 78620 -59380
rect 80020 -59480 80120 -59380
rect 81520 -59480 81620 -59380
rect 83020 -59480 83120 -59380
rect 84520 -59480 84620 -59380
rect 86020 -59480 86120 -59380
rect 87520 -59480 87620 -59380
rect 89020 -59480 89120 -59380
rect 90520 -59480 90620 -59380
rect 92020 -59480 92120 -59380
rect 93520 -59480 93620 -59380
rect 95020 -59480 95120 -59380
rect 96520 -59480 96620 -59380
rect 98020 -59480 98120 -59380
rect 99520 -59480 99620 -59380
rect 101020 -59480 101120 -59380
rect 102520 -59480 102620 -59380
rect 104020 -59480 104120 -59380
rect 105520 -59480 105620 -59380
rect 107020 -59480 107120 -59380
rect 108520 -59480 108620 -59380
rect 110020 -59480 110120 -59380
rect 111520 -59480 111620 -59380
rect 113020 -59480 113120 -59380
rect 114520 -59480 114620 -59380
rect 116020 -59480 116120 -59380
rect 117520 -59480 117620 -59380
rect 119020 -59480 119120 -59380
rect 520 -60980 620 -60880
rect 2020 -60980 2120 -60880
rect 3520 -60980 3620 -60880
rect 5020 -60980 5120 -60880
rect 6520 -60980 6620 -60880
rect 8020 -60980 8120 -60880
rect 9520 -60980 9620 -60880
rect 11020 -60980 11120 -60880
rect 12520 -60980 12620 -60880
rect 14020 -60980 14120 -60880
rect 15520 -60980 15620 -60880
rect 17020 -60980 17120 -60880
rect 18520 -60980 18620 -60880
rect 20020 -60980 20120 -60880
rect 21520 -60980 21620 -60880
rect 23020 -60980 23120 -60880
rect 24520 -60980 24620 -60880
rect 26020 -60980 26120 -60880
rect 27520 -60980 27620 -60880
rect 29020 -60980 29120 -60880
rect 30520 -60980 30620 -60880
rect 32020 -60980 32120 -60880
rect 33520 -60980 33620 -60880
rect 35020 -60980 35120 -60880
rect 36520 -60980 36620 -60880
rect 38020 -60980 38120 -60880
rect 39520 -60980 39620 -60880
rect 41020 -60980 41120 -60880
rect 42520 -60980 42620 -60880
rect 44020 -60980 44120 -60880
rect 45520 -60980 45620 -60880
rect 47020 -60980 47120 -60880
rect 48520 -60980 48620 -60880
rect 50020 -60980 50120 -60880
rect 51520 -60980 51620 -60880
rect 53020 -60980 53120 -60880
rect 54520 -60980 54620 -60880
rect 56020 -60980 56120 -60880
rect 57520 -60980 57620 -60880
rect 59020 -60980 59120 -60880
rect 60520 -60980 60620 -60880
rect 62020 -60980 62120 -60880
rect 63520 -60980 63620 -60880
rect 65020 -60980 65120 -60880
rect 66520 -60980 66620 -60880
rect 68020 -60980 68120 -60880
rect 69520 -60980 69620 -60880
rect 71020 -60980 71120 -60880
rect 72520 -60980 72620 -60880
rect 74020 -60980 74120 -60880
rect 75520 -60980 75620 -60880
rect 77020 -60980 77120 -60880
rect 78520 -60980 78620 -60880
rect 80020 -60980 80120 -60880
rect 81520 -60980 81620 -60880
rect 83020 -60980 83120 -60880
rect 84520 -60980 84620 -60880
rect 86020 -60980 86120 -60880
rect 87520 -60980 87620 -60880
rect 89020 -60980 89120 -60880
rect 90520 -60980 90620 -60880
rect 92020 -60980 92120 -60880
rect 93520 -60980 93620 -60880
rect 95020 -60980 95120 -60880
rect 96520 -60980 96620 -60880
rect 98020 -60980 98120 -60880
rect 99520 -60980 99620 -60880
rect 101020 -60980 101120 -60880
rect 102520 -60980 102620 -60880
rect 104020 -60980 104120 -60880
rect 105520 -60980 105620 -60880
rect 107020 -60980 107120 -60880
rect 108520 -60980 108620 -60880
rect 110020 -60980 110120 -60880
rect 111520 -60980 111620 -60880
rect 113020 -60980 113120 -60880
rect 114520 -60980 114620 -60880
rect 116020 -60980 116120 -60880
rect 117520 -60980 117620 -60880
rect 119020 -60980 119120 -60880
rect 520 -62480 620 -62380
rect 2020 -62480 2120 -62380
rect 3520 -62480 3620 -62380
rect 5020 -62480 5120 -62380
rect 6520 -62480 6620 -62380
rect 8020 -62480 8120 -62380
rect 9520 -62480 9620 -62380
rect 11020 -62480 11120 -62380
rect 12520 -62480 12620 -62380
rect 14020 -62480 14120 -62380
rect 15520 -62480 15620 -62380
rect 17020 -62480 17120 -62380
rect 18520 -62480 18620 -62380
rect 20020 -62480 20120 -62380
rect 21520 -62480 21620 -62380
rect 23020 -62480 23120 -62380
rect 24520 -62480 24620 -62380
rect 26020 -62480 26120 -62380
rect 27520 -62480 27620 -62380
rect 29020 -62480 29120 -62380
rect 30520 -62480 30620 -62380
rect 32020 -62480 32120 -62380
rect 33520 -62480 33620 -62380
rect 35020 -62480 35120 -62380
rect 36520 -62480 36620 -62380
rect 38020 -62480 38120 -62380
rect 39520 -62480 39620 -62380
rect 41020 -62480 41120 -62380
rect 42520 -62480 42620 -62380
rect 44020 -62480 44120 -62380
rect 45520 -62480 45620 -62380
rect 47020 -62480 47120 -62380
rect 48520 -62480 48620 -62380
rect 50020 -62480 50120 -62380
rect 51520 -62480 51620 -62380
rect 53020 -62480 53120 -62380
rect 54520 -62480 54620 -62380
rect 56020 -62480 56120 -62380
rect 57520 -62480 57620 -62380
rect 59020 -62480 59120 -62380
rect 60520 -62480 60620 -62380
rect 62020 -62480 62120 -62380
rect 63520 -62480 63620 -62380
rect 65020 -62480 65120 -62380
rect 66520 -62480 66620 -62380
rect 68020 -62480 68120 -62380
rect 69520 -62480 69620 -62380
rect 71020 -62480 71120 -62380
rect 72520 -62480 72620 -62380
rect 74020 -62480 74120 -62380
rect 75520 -62480 75620 -62380
rect 77020 -62480 77120 -62380
rect 78520 -62480 78620 -62380
rect 80020 -62480 80120 -62380
rect 81520 -62480 81620 -62380
rect 83020 -62480 83120 -62380
rect 84520 -62480 84620 -62380
rect 86020 -62480 86120 -62380
rect 87520 -62480 87620 -62380
rect 89020 -62480 89120 -62380
rect 90520 -62480 90620 -62380
rect 92020 -62480 92120 -62380
rect 93520 -62480 93620 -62380
rect 95020 -62480 95120 -62380
rect 96520 -62480 96620 -62380
rect 98020 -62480 98120 -62380
rect 99520 -62480 99620 -62380
rect 101020 -62480 101120 -62380
rect 102520 -62480 102620 -62380
rect 104020 -62480 104120 -62380
rect 105520 -62480 105620 -62380
rect 107020 -62480 107120 -62380
rect 108520 -62480 108620 -62380
rect 110020 -62480 110120 -62380
rect 111520 -62480 111620 -62380
rect 113020 -62480 113120 -62380
rect 114520 -62480 114620 -62380
rect 116020 -62480 116120 -62380
rect 117520 -62480 117620 -62380
rect 119020 -62480 119120 -62380
rect 520 -63980 620 -63880
rect 2020 -63980 2120 -63880
rect 3520 -63980 3620 -63880
rect 5020 -63980 5120 -63880
rect 6520 -63980 6620 -63880
rect 8020 -63980 8120 -63880
rect 9520 -63980 9620 -63880
rect 11020 -63980 11120 -63880
rect 12520 -63980 12620 -63880
rect 14020 -63980 14120 -63880
rect 15520 -63980 15620 -63880
rect 17020 -63980 17120 -63880
rect 18520 -63980 18620 -63880
rect 20020 -63980 20120 -63880
rect 21520 -63980 21620 -63880
rect 23020 -63980 23120 -63880
rect 24520 -63980 24620 -63880
rect 26020 -63980 26120 -63880
rect 27520 -63980 27620 -63880
rect 29020 -63980 29120 -63880
rect 30520 -63980 30620 -63880
rect 32020 -63980 32120 -63880
rect 33520 -63980 33620 -63880
rect 35020 -63980 35120 -63880
rect 36520 -63980 36620 -63880
rect 38020 -63980 38120 -63880
rect 39520 -63980 39620 -63880
rect 41020 -63980 41120 -63880
rect 42520 -63980 42620 -63880
rect 44020 -63980 44120 -63880
rect 45520 -63980 45620 -63880
rect 47020 -63980 47120 -63880
rect 48520 -63980 48620 -63880
rect 50020 -63980 50120 -63880
rect 51520 -63980 51620 -63880
rect 53020 -63980 53120 -63880
rect 54520 -63980 54620 -63880
rect 56020 -63980 56120 -63880
rect 57520 -63980 57620 -63880
rect 59020 -63980 59120 -63880
rect 60520 -63980 60620 -63880
rect 62020 -63980 62120 -63880
rect 63520 -63980 63620 -63880
rect 65020 -63980 65120 -63880
rect 66520 -63980 66620 -63880
rect 68020 -63980 68120 -63880
rect 69520 -63980 69620 -63880
rect 71020 -63980 71120 -63880
rect 72520 -63980 72620 -63880
rect 74020 -63980 74120 -63880
rect 75520 -63980 75620 -63880
rect 77020 -63980 77120 -63880
rect 78520 -63980 78620 -63880
rect 80020 -63980 80120 -63880
rect 81520 -63980 81620 -63880
rect 83020 -63980 83120 -63880
rect 84520 -63980 84620 -63880
rect 86020 -63980 86120 -63880
rect 87520 -63980 87620 -63880
rect 89020 -63980 89120 -63880
rect 90520 -63980 90620 -63880
rect 92020 -63980 92120 -63880
rect 93520 -63980 93620 -63880
rect 95020 -63980 95120 -63880
rect 96520 -63980 96620 -63880
rect 98020 -63980 98120 -63880
rect 99520 -63980 99620 -63880
rect 101020 -63980 101120 -63880
rect 102520 -63980 102620 -63880
rect 104020 -63980 104120 -63880
rect 105520 -63980 105620 -63880
rect 107020 -63980 107120 -63880
rect 108520 -63980 108620 -63880
rect 110020 -63980 110120 -63880
rect 111520 -63980 111620 -63880
rect 113020 -63980 113120 -63880
rect 114520 -63980 114620 -63880
rect 116020 -63980 116120 -63880
rect 117520 -63980 117620 -63880
rect 119020 -63980 119120 -63880
rect 520 -65480 620 -65380
rect 2020 -65480 2120 -65380
rect 3520 -65480 3620 -65380
rect 5020 -65480 5120 -65380
rect 6520 -65480 6620 -65380
rect 8020 -65480 8120 -65380
rect 9520 -65480 9620 -65380
rect 11020 -65480 11120 -65380
rect 12520 -65480 12620 -65380
rect 14020 -65480 14120 -65380
rect 15520 -65480 15620 -65380
rect 17020 -65480 17120 -65380
rect 18520 -65480 18620 -65380
rect 20020 -65480 20120 -65380
rect 21520 -65480 21620 -65380
rect 23020 -65480 23120 -65380
rect 24520 -65480 24620 -65380
rect 26020 -65480 26120 -65380
rect 27520 -65480 27620 -65380
rect 29020 -65480 29120 -65380
rect 30520 -65480 30620 -65380
rect 32020 -65480 32120 -65380
rect 33520 -65480 33620 -65380
rect 35020 -65480 35120 -65380
rect 36520 -65480 36620 -65380
rect 38020 -65480 38120 -65380
rect 39520 -65480 39620 -65380
rect 41020 -65480 41120 -65380
rect 42520 -65480 42620 -65380
rect 44020 -65480 44120 -65380
rect 45520 -65480 45620 -65380
rect 47020 -65480 47120 -65380
rect 48520 -65480 48620 -65380
rect 50020 -65480 50120 -65380
rect 51520 -65480 51620 -65380
rect 53020 -65480 53120 -65380
rect 54520 -65480 54620 -65380
rect 56020 -65480 56120 -65380
rect 57520 -65480 57620 -65380
rect 59020 -65480 59120 -65380
rect 60520 -65480 60620 -65380
rect 62020 -65480 62120 -65380
rect 63520 -65480 63620 -65380
rect 65020 -65480 65120 -65380
rect 66520 -65480 66620 -65380
rect 68020 -65480 68120 -65380
rect 69520 -65480 69620 -65380
rect 71020 -65480 71120 -65380
rect 72520 -65480 72620 -65380
rect 74020 -65480 74120 -65380
rect 75520 -65480 75620 -65380
rect 77020 -65480 77120 -65380
rect 78520 -65480 78620 -65380
rect 80020 -65480 80120 -65380
rect 81520 -65480 81620 -65380
rect 83020 -65480 83120 -65380
rect 84520 -65480 84620 -65380
rect 86020 -65480 86120 -65380
rect 87520 -65480 87620 -65380
rect 89020 -65480 89120 -65380
rect 90520 -65480 90620 -65380
rect 92020 -65480 92120 -65380
rect 93520 -65480 93620 -65380
rect 95020 -65480 95120 -65380
rect 96520 -65480 96620 -65380
rect 98020 -65480 98120 -65380
rect 99520 -65480 99620 -65380
rect 101020 -65480 101120 -65380
rect 102520 -65480 102620 -65380
rect 104020 -65480 104120 -65380
rect 105520 -65480 105620 -65380
rect 107020 -65480 107120 -65380
rect 108520 -65480 108620 -65380
rect 110020 -65480 110120 -65380
rect 111520 -65480 111620 -65380
rect 113020 -65480 113120 -65380
rect 114520 -65480 114620 -65380
rect 116020 -65480 116120 -65380
rect 117520 -65480 117620 -65380
rect 119020 -65480 119120 -65380
rect 520 -66980 620 -66880
rect 2020 -66980 2120 -66880
rect 3520 -66980 3620 -66880
rect 5020 -66980 5120 -66880
rect 6520 -66980 6620 -66880
rect 8020 -66980 8120 -66880
rect 9520 -66980 9620 -66880
rect 11020 -66980 11120 -66880
rect 12520 -66980 12620 -66880
rect 14020 -66980 14120 -66880
rect 15520 -66980 15620 -66880
rect 17020 -66980 17120 -66880
rect 18520 -66980 18620 -66880
rect 20020 -66980 20120 -66880
rect 21520 -66980 21620 -66880
rect 23020 -66980 23120 -66880
rect 24520 -66980 24620 -66880
rect 26020 -66980 26120 -66880
rect 27520 -66980 27620 -66880
rect 29020 -66980 29120 -66880
rect 30520 -66980 30620 -66880
rect 32020 -66980 32120 -66880
rect 33520 -66980 33620 -66880
rect 35020 -66980 35120 -66880
rect 36520 -66980 36620 -66880
rect 38020 -66980 38120 -66880
rect 39520 -66980 39620 -66880
rect 41020 -66980 41120 -66880
rect 42520 -66980 42620 -66880
rect 44020 -66980 44120 -66880
rect 45520 -66980 45620 -66880
rect 47020 -66980 47120 -66880
rect 48520 -66980 48620 -66880
rect 50020 -66980 50120 -66880
rect 51520 -66980 51620 -66880
rect 53020 -66980 53120 -66880
rect 54520 -66980 54620 -66880
rect 56020 -66980 56120 -66880
rect 57520 -66980 57620 -66880
rect 59020 -66980 59120 -66880
rect 60520 -66980 60620 -66880
rect 62020 -66980 62120 -66880
rect 63520 -66980 63620 -66880
rect 65020 -66980 65120 -66880
rect 66520 -66980 66620 -66880
rect 68020 -66980 68120 -66880
rect 69520 -66980 69620 -66880
rect 71020 -66980 71120 -66880
rect 72520 -66980 72620 -66880
rect 74020 -66980 74120 -66880
rect 75520 -66980 75620 -66880
rect 77020 -66980 77120 -66880
rect 78520 -66980 78620 -66880
rect 80020 -66980 80120 -66880
rect 81520 -66980 81620 -66880
rect 83020 -66980 83120 -66880
rect 84520 -66980 84620 -66880
rect 86020 -66980 86120 -66880
rect 87520 -66980 87620 -66880
rect 89020 -66980 89120 -66880
rect 90520 -66980 90620 -66880
rect 92020 -66980 92120 -66880
rect 93520 -66980 93620 -66880
rect 95020 -66980 95120 -66880
rect 96520 -66980 96620 -66880
rect 98020 -66980 98120 -66880
rect 99520 -66980 99620 -66880
rect 101020 -66980 101120 -66880
rect 102520 -66980 102620 -66880
rect 104020 -66980 104120 -66880
rect 105520 -66980 105620 -66880
rect 107020 -66980 107120 -66880
rect 108520 -66980 108620 -66880
rect 110020 -66980 110120 -66880
rect 111520 -66980 111620 -66880
rect 113020 -66980 113120 -66880
rect 114520 -66980 114620 -66880
rect 116020 -66980 116120 -66880
rect 117520 -66980 117620 -66880
rect 119020 -66980 119120 -66880
rect 520 -68480 620 -68380
rect 2020 -68480 2120 -68380
rect 3520 -68480 3620 -68380
rect 5020 -68480 5120 -68380
rect 6520 -68480 6620 -68380
rect 8020 -68480 8120 -68380
rect 9520 -68480 9620 -68380
rect 11020 -68480 11120 -68380
rect 12520 -68480 12620 -68380
rect 14020 -68480 14120 -68380
rect 15520 -68480 15620 -68380
rect 17020 -68480 17120 -68380
rect 18520 -68480 18620 -68380
rect 20020 -68480 20120 -68380
rect 21520 -68480 21620 -68380
rect 23020 -68480 23120 -68380
rect 24520 -68480 24620 -68380
rect 26020 -68480 26120 -68380
rect 27520 -68480 27620 -68380
rect 29020 -68480 29120 -68380
rect 30520 -68480 30620 -68380
rect 32020 -68480 32120 -68380
rect 33520 -68480 33620 -68380
rect 35020 -68480 35120 -68380
rect 36520 -68480 36620 -68380
rect 38020 -68480 38120 -68380
rect 39520 -68480 39620 -68380
rect 41020 -68480 41120 -68380
rect 42520 -68480 42620 -68380
rect 44020 -68480 44120 -68380
rect 45520 -68480 45620 -68380
rect 47020 -68480 47120 -68380
rect 48520 -68480 48620 -68380
rect 50020 -68480 50120 -68380
rect 51520 -68480 51620 -68380
rect 53020 -68480 53120 -68380
rect 54520 -68480 54620 -68380
rect 56020 -68480 56120 -68380
rect 57520 -68480 57620 -68380
rect 59020 -68480 59120 -68380
rect 60520 -68480 60620 -68380
rect 62020 -68480 62120 -68380
rect 63520 -68480 63620 -68380
rect 65020 -68480 65120 -68380
rect 66520 -68480 66620 -68380
rect 68020 -68480 68120 -68380
rect 69520 -68480 69620 -68380
rect 71020 -68480 71120 -68380
rect 72520 -68480 72620 -68380
rect 74020 -68480 74120 -68380
rect 75520 -68480 75620 -68380
rect 77020 -68480 77120 -68380
rect 78520 -68480 78620 -68380
rect 80020 -68480 80120 -68380
rect 81520 -68480 81620 -68380
rect 83020 -68480 83120 -68380
rect 84520 -68480 84620 -68380
rect 86020 -68480 86120 -68380
rect 87520 -68480 87620 -68380
rect 89020 -68480 89120 -68380
rect 90520 -68480 90620 -68380
rect 92020 -68480 92120 -68380
rect 93520 -68480 93620 -68380
rect 95020 -68480 95120 -68380
rect 96520 -68480 96620 -68380
rect 98020 -68480 98120 -68380
rect 99520 -68480 99620 -68380
rect 101020 -68480 101120 -68380
rect 102520 -68480 102620 -68380
rect 104020 -68480 104120 -68380
rect 105520 -68480 105620 -68380
rect 107020 -68480 107120 -68380
rect 108520 -68480 108620 -68380
rect 110020 -68480 110120 -68380
rect 111520 -68480 111620 -68380
rect 113020 -68480 113120 -68380
rect 114520 -68480 114620 -68380
rect 116020 -68480 116120 -68380
rect 117520 -68480 117620 -68380
rect 119020 -68480 119120 -68380
rect 520 -69980 620 -69880
rect 2020 -69980 2120 -69880
rect 3520 -69980 3620 -69880
rect 5020 -69980 5120 -69880
rect 6520 -69980 6620 -69880
rect 8020 -69980 8120 -69880
rect 9520 -69980 9620 -69880
rect 11020 -69980 11120 -69880
rect 12520 -69980 12620 -69880
rect 14020 -69980 14120 -69880
rect 15520 -69980 15620 -69880
rect 17020 -69980 17120 -69880
rect 18520 -69980 18620 -69880
rect 20020 -69980 20120 -69880
rect 21520 -69980 21620 -69880
rect 23020 -69980 23120 -69880
rect 24520 -69980 24620 -69880
rect 26020 -69980 26120 -69880
rect 27520 -69980 27620 -69880
rect 29020 -69980 29120 -69880
rect 30520 -69980 30620 -69880
rect 32020 -69980 32120 -69880
rect 33520 -69980 33620 -69880
rect 35020 -69980 35120 -69880
rect 36520 -69980 36620 -69880
rect 38020 -69980 38120 -69880
rect 39520 -69980 39620 -69880
rect 41020 -69980 41120 -69880
rect 42520 -69980 42620 -69880
rect 44020 -69980 44120 -69880
rect 45520 -69980 45620 -69880
rect 47020 -69980 47120 -69880
rect 48520 -69980 48620 -69880
rect 50020 -69980 50120 -69880
rect 51520 -69980 51620 -69880
rect 53020 -69980 53120 -69880
rect 54520 -69980 54620 -69880
rect 56020 -69980 56120 -69880
rect 57520 -69980 57620 -69880
rect 59020 -69980 59120 -69880
rect 60520 -69980 60620 -69880
rect 62020 -69980 62120 -69880
rect 63520 -69980 63620 -69880
rect 65020 -69980 65120 -69880
rect 66520 -69980 66620 -69880
rect 68020 -69980 68120 -69880
rect 69520 -69980 69620 -69880
rect 71020 -69980 71120 -69880
rect 72520 -69980 72620 -69880
rect 74020 -69980 74120 -69880
rect 75520 -69980 75620 -69880
rect 77020 -69980 77120 -69880
rect 78520 -69980 78620 -69880
rect 80020 -69980 80120 -69880
rect 81520 -69980 81620 -69880
rect 83020 -69980 83120 -69880
rect 84520 -69980 84620 -69880
rect 86020 -69980 86120 -69880
rect 87520 -69980 87620 -69880
rect 89020 -69980 89120 -69880
rect 90520 -69980 90620 -69880
rect 92020 -69980 92120 -69880
rect 93520 -69980 93620 -69880
rect 95020 -69980 95120 -69880
rect 96520 -69980 96620 -69880
rect 98020 -69980 98120 -69880
rect 99520 -69980 99620 -69880
rect 101020 -69980 101120 -69880
rect 102520 -69980 102620 -69880
rect 104020 -69980 104120 -69880
rect 105520 -69980 105620 -69880
rect 107020 -69980 107120 -69880
rect 108520 -69980 108620 -69880
rect 110020 -69980 110120 -69880
rect 111520 -69980 111620 -69880
rect 113020 -69980 113120 -69880
rect 114520 -69980 114620 -69880
rect 116020 -69980 116120 -69880
rect 117520 -69980 117620 -69880
rect 119020 -69980 119120 -69880
rect 520 -71480 620 -71380
rect 2020 -71480 2120 -71380
rect 3520 -71480 3620 -71380
rect 5020 -71480 5120 -71380
rect 6520 -71480 6620 -71380
rect 8020 -71480 8120 -71380
rect 9520 -71480 9620 -71380
rect 11020 -71480 11120 -71380
rect 12520 -71480 12620 -71380
rect 14020 -71480 14120 -71380
rect 15520 -71480 15620 -71380
rect 17020 -71480 17120 -71380
rect 18520 -71480 18620 -71380
rect 20020 -71480 20120 -71380
rect 21520 -71480 21620 -71380
rect 23020 -71480 23120 -71380
rect 24520 -71480 24620 -71380
rect 26020 -71480 26120 -71380
rect 27520 -71480 27620 -71380
rect 29020 -71480 29120 -71380
rect 30520 -71480 30620 -71380
rect 32020 -71480 32120 -71380
rect 33520 -71480 33620 -71380
rect 35020 -71480 35120 -71380
rect 36520 -71480 36620 -71380
rect 38020 -71480 38120 -71380
rect 39520 -71480 39620 -71380
rect 41020 -71480 41120 -71380
rect 42520 -71480 42620 -71380
rect 44020 -71480 44120 -71380
rect 45520 -71480 45620 -71380
rect 47020 -71480 47120 -71380
rect 48520 -71480 48620 -71380
rect 50020 -71480 50120 -71380
rect 51520 -71480 51620 -71380
rect 53020 -71480 53120 -71380
rect 54520 -71480 54620 -71380
rect 56020 -71480 56120 -71380
rect 57520 -71480 57620 -71380
rect 59020 -71480 59120 -71380
rect 60520 -71480 60620 -71380
rect 62020 -71480 62120 -71380
rect 63520 -71480 63620 -71380
rect 65020 -71480 65120 -71380
rect 66520 -71480 66620 -71380
rect 68020 -71480 68120 -71380
rect 69520 -71480 69620 -71380
rect 71020 -71480 71120 -71380
rect 72520 -71480 72620 -71380
rect 74020 -71480 74120 -71380
rect 75520 -71480 75620 -71380
rect 77020 -71480 77120 -71380
rect 78520 -71480 78620 -71380
rect 80020 -71480 80120 -71380
rect 81520 -71480 81620 -71380
rect 83020 -71480 83120 -71380
rect 84520 -71480 84620 -71380
rect 86020 -71480 86120 -71380
rect 87520 -71480 87620 -71380
rect 89020 -71480 89120 -71380
rect 90520 -71480 90620 -71380
rect 92020 -71480 92120 -71380
rect 93520 -71480 93620 -71380
rect 95020 -71480 95120 -71380
rect 96520 -71480 96620 -71380
rect 98020 -71480 98120 -71380
rect 99520 -71480 99620 -71380
rect 101020 -71480 101120 -71380
rect 102520 -71480 102620 -71380
rect 104020 -71480 104120 -71380
rect 105520 -71480 105620 -71380
rect 107020 -71480 107120 -71380
rect 108520 -71480 108620 -71380
rect 110020 -71480 110120 -71380
rect 111520 -71480 111620 -71380
rect 113020 -71480 113120 -71380
rect 114520 -71480 114620 -71380
rect 116020 -71480 116120 -71380
rect 117520 -71480 117620 -71380
rect 119020 -71480 119120 -71380
rect 520 -72980 620 -72880
rect 2020 -72980 2120 -72880
rect 3520 -72980 3620 -72880
rect 5020 -72980 5120 -72880
rect 6520 -72980 6620 -72880
rect 8020 -72980 8120 -72880
rect 9520 -72980 9620 -72880
rect 11020 -72980 11120 -72880
rect 12520 -72980 12620 -72880
rect 14020 -72980 14120 -72880
rect 15520 -72980 15620 -72880
rect 17020 -72980 17120 -72880
rect 18520 -72980 18620 -72880
rect 20020 -72980 20120 -72880
rect 21520 -72980 21620 -72880
rect 23020 -72980 23120 -72880
rect 24520 -72980 24620 -72880
rect 26020 -72980 26120 -72880
rect 27520 -72980 27620 -72880
rect 29020 -72980 29120 -72880
rect 30520 -72980 30620 -72880
rect 32020 -72980 32120 -72880
rect 33520 -72980 33620 -72880
rect 35020 -72980 35120 -72880
rect 36520 -72980 36620 -72880
rect 38020 -72980 38120 -72880
rect 39520 -72980 39620 -72880
rect 41020 -72980 41120 -72880
rect 42520 -72980 42620 -72880
rect 44020 -72980 44120 -72880
rect 45520 -72980 45620 -72880
rect 47020 -72980 47120 -72880
rect 48520 -72980 48620 -72880
rect 50020 -72980 50120 -72880
rect 51520 -72980 51620 -72880
rect 53020 -72980 53120 -72880
rect 54520 -72980 54620 -72880
rect 56020 -72980 56120 -72880
rect 57520 -72980 57620 -72880
rect 59020 -72980 59120 -72880
rect 60520 -72980 60620 -72880
rect 62020 -72980 62120 -72880
rect 63520 -72980 63620 -72880
rect 65020 -72980 65120 -72880
rect 66520 -72980 66620 -72880
rect 68020 -72980 68120 -72880
rect 69520 -72980 69620 -72880
rect 71020 -72980 71120 -72880
rect 72520 -72980 72620 -72880
rect 74020 -72980 74120 -72880
rect 75520 -72980 75620 -72880
rect 77020 -72980 77120 -72880
rect 78520 -72980 78620 -72880
rect 80020 -72980 80120 -72880
rect 81520 -72980 81620 -72880
rect 83020 -72980 83120 -72880
rect 84520 -72980 84620 -72880
rect 86020 -72980 86120 -72880
rect 87520 -72980 87620 -72880
rect 89020 -72980 89120 -72880
rect 90520 -72980 90620 -72880
rect 92020 -72980 92120 -72880
rect 93520 -72980 93620 -72880
rect 95020 -72980 95120 -72880
rect 96520 -72980 96620 -72880
rect 98020 -72980 98120 -72880
rect 99520 -72980 99620 -72880
rect 101020 -72980 101120 -72880
rect 102520 -72980 102620 -72880
rect 104020 -72980 104120 -72880
rect 105520 -72980 105620 -72880
rect 107020 -72980 107120 -72880
rect 108520 -72980 108620 -72880
rect 110020 -72980 110120 -72880
rect 111520 -72980 111620 -72880
rect 113020 -72980 113120 -72880
rect 114520 -72980 114620 -72880
rect 116020 -72980 116120 -72880
rect 117520 -72980 117620 -72880
rect 119020 -72980 119120 -72880
rect 520 -74480 620 -74380
rect 2020 -74480 2120 -74380
rect 3520 -74480 3620 -74380
rect 5020 -74480 5120 -74380
rect 6520 -74480 6620 -74380
rect 8020 -74480 8120 -74380
rect 9520 -74480 9620 -74380
rect 11020 -74480 11120 -74380
rect 12520 -74480 12620 -74380
rect 14020 -74480 14120 -74380
rect 15520 -74480 15620 -74380
rect 17020 -74480 17120 -74380
rect 18520 -74480 18620 -74380
rect 20020 -74480 20120 -74380
rect 21520 -74480 21620 -74380
rect 23020 -74480 23120 -74380
rect 24520 -74480 24620 -74380
rect 26020 -74480 26120 -74380
rect 27520 -74480 27620 -74380
rect 29020 -74480 29120 -74380
rect 30520 -74480 30620 -74380
rect 32020 -74480 32120 -74380
rect 33520 -74480 33620 -74380
rect 35020 -74480 35120 -74380
rect 36520 -74480 36620 -74380
rect 38020 -74480 38120 -74380
rect 39520 -74480 39620 -74380
rect 41020 -74480 41120 -74380
rect 42520 -74480 42620 -74380
rect 44020 -74480 44120 -74380
rect 45520 -74480 45620 -74380
rect 47020 -74480 47120 -74380
rect 48520 -74480 48620 -74380
rect 50020 -74480 50120 -74380
rect 51520 -74480 51620 -74380
rect 53020 -74480 53120 -74380
rect 54520 -74480 54620 -74380
rect 56020 -74480 56120 -74380
rect 57520 -74480 57620 -74380
rect 59020 -74480 59120 -74380
rect 60520 -74480 60620 -74380
rect 62020 -74480 62120 -74380
rect 63520 -74480 63620 -74380
rect 65020 -74480 65120 -74380
rect 66520 -74480 66620 -74380
rect 68020 -74480 68120 -74380
rect 69520 -74480 69620 -74380
rect 71020 -74480 71120 -74380
rect 72520 -74480 72620 -74380
rect 74020 -74480 74120 -74380
rect 75520 -74480 75620 -74380
rect 77020 -74480 77120 -74380
rect 78520 -74480 78620 -74380
rect 80020 -74480 80120 -74380
rect 81520 -74480 81620 -74380
rect 83020 -74480 83120 -74380
rect 84520 -74480 84620 -74380
rect 86020 -74480 86120 -74380
rect 87520 -74480 87620 -74380
rect 89020 -74480 89120 -74380
rect 90520 -74480 90620 -74380
rect 92020 -74480 92120 -74380
rect 93520 -74480 93620 -74380
rect 95020 -74480 95120 -74380
rect 96520 -74480 96620 -74380
rect 98020 -74480 98120 -74380
rect 99520 -74480 99620 -74380
rect 101020 -74480 101120 -74380
rect 102520 -74480 102620 -74380
rect 104020 -74480 104120 -74380
rect 105520 -74480 105620 -74380
rect 107020 -74480 107120 -74380
rect 108520 -74480 108620 -74380
rect 110020 -74480 110120 -74380
rect 111520 -74480 111620 -74380
rect 113020 -74480 113120 -74380
rect 114520 -74480 114620 -74380
rect 116020 -74480 116120 -74380
rect 117520 -74480 117620 -74380
rect 119020 -74480 119120 -74380
rect 520 -75980 620 -75880
rect 2020 -75980 2120 -75880
rect 3520 -75980 3620 -75880
rect 5020 -75980 5120 -75880
rect 6520 -75980 6620 -75880
rect 8020 -75980 8120 -75880
rect 9520 -75980 9620 -75880
rect 11020 -75980 11120 -75880
rect 12520 -75980 12620 -75880
rect 14020 -75980 14120 -75880
rect 15520 -75980 15620 -75880
rect 17020 -75980 17120 -75880
rect 18520 -75980 18620 -75880
rect 20020 -75980 20120 -75880
rect 21520 -75980 21620 -75880
rect 23020 -75980 23120 -75880
rect 24520 -75980 24620 -75880
rect 26020 -75980 26120 -75880
rect 27520 -75980 27620 -75880
rect 29020 -75980 29120 -75880
rect 30520 -75980 30620 -75880
rect 32020 -75980 32120 -75880
rect 33520 -75980 33620 -75880
rect 35020 -75980 35120 -75880
rect 36520 -75980 36620 -75880
rect 38020 -75980 38120 -75880
rect 39520 -75980 39620 -75880
rect 41020 -75980 41120 -75880
rect 42520 -75980 42620 -75880
rect 44020 -75980 44120 -75880
rect 45520 -75980 45620 -75880
rect 47020 -75980 47120 -75880
rect 48520 -75980 48620 -75880
rect 50020 -75980 50120 -75880
rect 51520 -75980 51620 -75880
rect 53020 -75980 53120 -75880
rect 54520 -75980 54620 -75880
rect 56020 -75980 56120 -75880
rect 57520 -75980 57620 -75880
rect 59020 -75980 59120 -75880
rect 60520 -75980 60620 -75880
rect 62020 -75980 62120 -75880
rect 63520 -75980 63620 -75880
rect 65020 -75980 65120 -75880
rect 66520 -75980 66620 -75880
rect 68020 -75980 68120 -75880
rect 69520 -75980 69620 -75880
rect 71020 -75980 71120 -75880
rect 72520 -75980 72620 -75880
rect 74020 -75980 74120 -75880
rect 75520 -75980 75620 -75880
rect 77020 -75980 77120 -75880
rect 78520 -75980 78620 -75880
rect 80020 -75980 80120 -75880
rect 81520 -75980 81620 -75880
rect 83020 -75980 83120 -75880
rect 84520 -75980 84620 -75880
rect 86020 -75980 86120 -75880
rect 87520 -75980 87620 -75880
rect 89020 -75980 89120 -75880
rect 90520 -75980 90620 -75880
rect 92020 -75980 92120 -75880
rect 93520 -75980 93620 -75880
rect 95020 -75980 95120 -75880
rect 96520 -75980 96620 -75880
rect 98020 -75980 98120 -75880
rect 99520 -75980 99620 -75880
rect 101020 -75980 101120 -75880
rect 102520 -75980 102620 -75880
rect 104020 -75980 104120 -75880
rect 105520 -75980 105620 -75880
rect 107020 -75980 107120 -75880
rect 108520 -75980 108620 -75880
rect 110020 -75980 110120 -75880
rect 111520 -75980 111620 -75880
rect 113020 -75980 113120 -75880
rect 114520 -75980 114620 -75880
rect 116020 -75980 116120 -75880
rect 117520 -75980 117620 -75880
rect 119020 -75980 119120 -75880
rect 520 -77480 620 -77380
rect 2020 -77480 2120 -77380
rect 3520 -77480 3620 -77380
rect 5020 -77480 5120 -77380
rect 6520 -77480 6620 -77380
rect 8020 -77480 8120 -77380
rect 9520 -77480 9620 -77380
rect 11020 -77480 11120 -77380
rect 12520 -77480 12620 -77380
rect 14020 -77480 14120 -77380
rect 15520 -77480 15620 -77380
rect 17020 -77480 17120 -77380
rect 18520 -77480 18620 -77380
rect 20020 -77480 20120 -77380
rect 21520 -77480 21620 -77380
rect 23020 -77480 23120 -77380
rect 24520 -77480 24620 -77380
rect 26020 -77480 26120 -77380
rect 27520 -77480 27620 -77380
rect 29020 -77480 29120 -77380
rect 30520 -77480 30620 -77380
rect 32020 -77480 32120 -77380
rect 33520 -77480 33620 -77380
rect 35020 -77480 35120 -77380
rect 36520 -77480 36620 -77380
rect 38020 -77480 38120 -77380
rect 39520 -77480 39620 -77380
rect 41020 -77480 41120 -77380
rect 42520 -77480 42620 -77380
rect 44020 -77480 44120 -77380
rect 45520 -77480 45620 -77380
rect 47020 -77480 47120 -77380
rect 48520 -77480 48620 -77380
rect 50020 -77480 50120 -77380
rect 51520 -77480 51620 -77380
rect 53020 -77480 53120 -77380
rect 54520 -77480 54620 -77380
rect 56020 -77480 56120 -77380
rect 57520 -77480 57620 -77380
rect 59020 -77480 59120 -77380
rect 60520 -77480 60620 -77380
rect 62020 -77480 62120 -77380
rect 63520 -77480 63620 -77380
rect 65020 -77480 65120 -77380
rect 66520 -77480 66620 -77380
rect 68020 -77480 68120 -77380
rect 69520 -77480 69620 -77380
rect 71020 -77480 71120 -77380
rect 72520 -77480 72620 -77380
rect 74020 -77480 74120 -77380
rect 75520 -77480 75620 -77380
rect 77020 -77480 77120 -77380
rect 78520 -77480 78620 -77380
rect 80020 -77480 80120 -77380
rect 81520 -77480 81620 -77380
rect 83020 -77480 83120 -77380
rect 84520 -77480 84620 -77380
rect 86020 -77480 86120 -77380
rect 87520 -77480 87620 -77380
rect 89020 -77480 89120 -77380
rect 90520 -77480 90620 -77380
rect 92020 -77480 92120 -77380
rect 93520 -77480 93620 -77380
rect 95020 -77480 95120 -77380
rect 96520 -77480 96620 -77380
rect 98020 -77480 98120 -77380
rect 99520 -77480 99620 -77380
rect 101020 -77480 101120 -77380
rect 102520 -77480 102620 -77380
rect 104020 -77480 104120 -77380
rect 105520 -77480 105620 -77380
rect 107020 -77480 107120 -77380
rect 108520 -77480 108620 -77380
rect 110020 -77480 110120 -77380
rect 111520 -77480 111620 -77380
rect 113020 -77480 113120 -77380
rect 114520 -77480 114620 -77380
rect 116020 -77480 116120 -77380
rect 117520 -77480 117620 -77380
rect 119020 -77480 119120 -77380
rect 520 -78980 620 -78880
rect 2020 -78980 2120 -78880
rect 3520 -78980 3620 -78880
rect 5020 -78980 5120 -78880
rect 6520 -78980 6620 -78880
rect 8020 -78980 8120 -78880
rect 9520 -78980 9620 -78880
rect 11020 -78980 11120 -78880
rect 12520 -78980 12620 -78880
rect 14020 -78980 14120 -78880
rect 15520 -78980 15620 -78880
rect 17020 -78980 17120 -78880
rect 18520 -78980 18620 -78880
rect 20020 -78980 20120 -78880
rect 21520 -78980 21620 -78880
rect 23020 -78980 23120 -78880
rect 24520 -78980 24620 -78880
rect 26020 -78980 26120 -78880
rect 27520 -78980 27620 -78880
rect 29020 -78980 29120 -78880
rect 30520 -78980 30620 -78880
rect 32020 -78980 32120 -78880
rect 33520 -78980 33620 -78880
rect 35020 -78980 35120 -78880
rect 36520 -78980 36620 -78880
rect 38020 -78980 38120 -78880
rect 39520 -78980 39620 -78880
rect 41020 -78980 41120 -78880
rect 42520 -78980 42620 -78880
rect 44020 -78980 44120 -78880
rect 45520 -78980 45620 -78880
rect 47020 -78980 47120 -78880
rect 48520 -78980 48620 -78880
rect 50020 -78980 50120 -78880
rect 51520 -78980 51620 -78880
rect 53020 -78980 53120 -78880
rect 54520 -78980 54620 -78880
rect 56020 -78980 56120 -78880
rect 57520 -78980 57620 -78880
rect 59020 -78980 59120 -78880
rect 60520 -78980 60620 -78880
rect 62020 -78980 62120 -78880
rect 63520 -78980 63620 -78880
rect 65020 -78980 65120 -78880
rect 66520 -78980 66620 -78880
rect 68020 -78980 68120 -78880
rect 69520 -78980 69620 -78880
rect 71020 -78980 71120 -78880
rect 72520 -78980 72620 -78880
rect 74020 -78980 74120 -78880
rect 75520 -78980 75620 -78880
rect 77020 -78980 77120 -78880
rect 78520 -78980 78620 -78880
rect 80020 -78980 80120 -78880
rect 81520 -78980 81620 -78880
rect 83020 -78980 83120 -78880
rect 84520 -78980 84620 -78880
rect 86020 -78980 86120 -78880
rect 87520 -78980 87620 -78880
rect 89020 -78980 89120 -78880
rect 90520 -78980 90620 -78880
rect 92020 -78980 92120 -78880
rect 93520 -78980 93620 -78880
rect 95020 -78980 95120 -78880
rect 96520 -78980 96620 -78880
rect 98020 -78980 98120 -78880
rect 99520 -78980 99620 -78880
rect 101020 -78980 101120 -78880
rect 102520 -78980 102620 -78880
rect 104020 -78980 104120 -78880
rect 105520 -78980 105620 -78880
rect 107020 -78980 107120 -78880
rect 108520 -78980 108620 -78880
rect 110020 -78980 110120 -78880
rect 111520 -78980 111620 -78880
rect 113020 -78980 113120 -78880
rect 114520 -78980 114620 -78880
rect 116020 -78980 116120 -78880
rect 117520 -78980 117620 -78880
rect 119020 -78980 119120 -78880
rect 520 -80480 620 -80380
rect 2020 -80480 2120 -80380
rect 3520 -80480 3620 -80380
rect 5020 -80480 5120 -80380
rect 6520 -80480 6620 -80380
rect 8020 -80480 8120 -80380
rect 9520 -80480 9620 -80380
rect 11020 -80480 11120 -80380
rect 12520 -80480 12620 -80380
rect 14020 -80480 14120 -80380
rect 15520 -80480 15620 -80380
rect 17020 -80480 17120 -80380
rect 18520 -80480 18620 -80380
rect 20020 -80480 20120 -80380
rect 21520 -80480 21620 -80380
rect 23020 -80480 23120 -80380
rect 24520 -80480 24620 -80380
rect 26020 -80480 26120 -80380
rect 27520 -80480 27620 -80380
rect 29020 -80480 29120 -80380
rect 30520 -80480 30620 -80380
rect 32020 -80480 32120 -80380
rect 33520 -80480 33620 -80380
rect 35020 -80480 35120 -80380
rect 36520 -80480 36620 -80380
rect 38020 -80480 38120 -80380
rect 39520 -80480 39620 -80380
rect 41020 -80480 41120 -80380
rect 42520 -80480 42620 -80380
rect 44020 -80480 44120 -80380
rect 45520 -80480 45620 -80380
rect 47020 -80480 47120 -80380
rect 48520 -80480 48620 -80380
rect 50020 -80480 50120 -80380
rect 51520 -80480 51620 -80380
rect 53020 -80480 53120 -80380
rect 54520 -80480 54620 -80380
rect 56020 -80480 56120 -80380
rect 57520 -80480 57620 -80380
rect 59020 -80480 59120 -80380
rect 60520 -80480 60620 -80380
rect 62020 -80480 62120 -80380
rect 63520 -80480 63620 -80380
rect 65020 -80480 65120 -80380
rect 66520 -80480 66620 -80380
rect 68020 -80480 68120 -80380
rect 69520 -80480 69620 -80380
rect 71020 -80480 71120 -80380
rect 72520 -80480 72620 -80380
rect 74020 -80480 74120 -80380
rect 75520 -80480 75620 -80380
rect 77020 -80480 77120 -80380
rect 78520 -80480 78620 -80380
rect 80020 -80480 80120 -80380
rect 81520 -80480 81620 -80380
rect 83020 -80480 83120 -80380
rect 84520 -80480 84620 -80380
rect 86020 -80480 86120 -80380
rect 87520 -80480 87620 -80380
rect 89020 -80480 89120 -80380
rect 90520 -80480 90620 -80380
rect 92020 -80480 92120 -80380
rect 93520 -80480 93620 -80380
rect 95020 -80480 95120 -80380
rect 96520 -80480 96620 -80380
rect 98020 -80480 98120 -80380
rect 99520 -80480 99620 -80380
rect 101020 -80480 101120 -80380
rect 102520 -80480 102620 -80380
rect 104020 -80480 104120 -80380
rect 105520 -80480 105620 -80380
rect 107020 -80480 107120 -80380
rect 108520 -80480 108620 -80380
rect 110020 -80480 110120 -80380
rect 111520 -80480 111620 -80380
rect 113020 -80480 113120 -80380
rect 114520 -80480 114620 -80380
rect 116020 -80480 116120 -80380
rect 117520 -80480 117620 -80380
rect 119020 -80480 119120 -80380
rect 520 -81980 620 -81880
rect 2020 -81980 2120 -81880
rect 3520 -81980 3620 -81880
rect 5020 -81980 5120 -81880
rect 6520 -81980 6620 -81880
rect 8020 -81980 8120 -81880
rect 9520 -81980 9620 -81880
rect 11020 -81980 11120 -81880
rect 12520 -81980 12620 -81880
rect 14020 -81980 14120 -81880
rect 15520 -81980 15620 -81880
rect 17020 -81980 17120 -81880
rect 18520 -81980 18620 -81880
rect 20020 -81980 20120 -81880
rect 21520 -81980 21620 -81880
rect 23020 -81980 23120 -81880
rect 24520 -81980 24620 -81880
rect 26020 -81980 26120 -81880
rect 27520 -81980 27620 -81880
rect 29020 -81980 29120 -81880
rect 30520 -81980 30620 -81880
rect 32020 -81980 32120 -81880
rect 33520 -81980 33620 -81880
rect 35020 -81980 35120 -81880
rect 36520 -81980 36620 -81880
rect 38020 -81980 38120 -81880
rect 39520 -81980 39620 -81880
rect 41020 -81980 41120 -81880
rect 42520 -81980 42620 -81880
rect 44020 -81980 44120 -81880
rect 45520 -81980 45620 -81880
rect 47020 -81980 47120 -81880
rect 48520 -81980 48620 -81880
rect 50020 -81980 50120 -81880
rect 51520 -81980 51620 -81880
rect 53020 -81980 53120 -81880
rect 54520 -81980 54620 -81880
rect 56020 -81980 56120 -81880
rect 57520 -81980 57620 -81880
rect 59020 -81980 59120 -81880
rect 60520 -81980 60620 -81880
rect 62020 -81980 62120 -81880
rect 63520 -81980 63620 -81880
rect 65020 -81980 65120 -81880
rect 66520 -81980 66620 -81880
rect 68020 -81980 68120 -81880
rect 69520 -81980 69620 -81880
rect 71020 -81980 71120 -81880
rect 72520 -81980 72620 -81880
rect 74020 -81980 74120 -81880
rect 75520 -81980 75620 -81880
rect 77020 -81980 77120 -81880
rect 78520 -81980 78620 -81880
rect 80020 -81980 80120 -81880
rect 81520 -81980 81620 -81880
rect 83020 -81980 83120 -81880
rect 84520 -81980 84620 -81880
rect 86020 -81980 86120 -81880
rect 87520 -81980 87620 -81880
rect 89020 -81980 89120 -81880
rect 90520 -81980 90620 -81880
rect 92020 -81980 92120 -81880
rect 93520 -81980 93620 -81880
rect 95020 -81980 95120 -81880
rect 96520 -81980 96620 -81880
rect 98020 -81980 98120 -81880
rect 99520 -81980 99620 -81880
rect 101020 -81980 101120 -81880
rect 102520 -81980 102620 -81880
rect 104020 -81980 104120 -81880
rect 105520 -81980 105620 -81880
rect 107020 -81980 107120 -81880
rect 108520 -81980 108620 -81880
rect 110020 -81980 110120 -81880
rect 111520 -81980 111620 -81880
rect 113020 -81980 113120 -81880
rect 114520 -81980 114620 -81880
rect 116020 -81980 116120 -81880
rect 117520 -81980 117620 -81880
rect 119020 -81980 119120 -81880
rect 520 -83480 620 -83380
rect 2020 -83480 2120 -83380
rect 3520 -83480 3620 -83380
rect 5020 -83480 5120 -83380
rect 6520 -83480 6620 -83380
rect 8020 -83480 8120 -83380
rect 9520 -83480 9620 -83380
rect 11020 -83480 11120 -83380
rect 12520 -83480 12620 -83380
rect 14020 -83480 14120 -83380
rect 15520 -83480 15620 -83380
rect 17020 -83480 17120 -83380
rect 18520 -83480 18620 -83380
rect 20020 -83480 20120 -83380
rect 21520 -83480 21620 -83380
rect 23020 -83480 23120 -83380
rect 24520 -83480 24620 -83380
rect 26020 -83480 26120 -83380
rect 27520 -83480 27620 -83380
rect 29020 -83480 29120 -83380
rect 30520 -83480 30620 -83380
rect 32020 -83480 32120 -83380
rect 33520 -83480 33620 -83380
rect 35020 -83480 35120 -83380
rect 36520 -83480 36620 -83380
rect 38020 -83480 38120 -83380
rect 39520 -83480 39620 -83380
rect 41020 -83480 41120 -83380
rect 42520 -83480 42620 -83380
rect 44020 -83480 44120 -83380
rect 45520 -83480 45620 -83380
rect 47020 -83480 47120 -83380
rect 48520 -83480 48620 -83380
rect 50020 -83480 50120 -83380
rect 51520 -83480 51620 -83380
rect 53020 -83480 53120 -83380
rect 54520 -83480 54620 -83380
rect 56020 -83480 56120 -83380
rect 57520 -83480 57620 -83380
rect 59020 -83480 59120 -83380
rect 60520 -83480 60620 -83380
rect 62020 -83480 62120 -83380
rect 63520 -83480 63620 -83380
rect 65020 -83480 65120 -83380
rect 66520 -83480 66620 -83380
rect 68020 -83480 68120 -83380
rect 69520 -83480 69620 -83380
rect 71020 -83480 71120 -83380
rect 72520 -83480 72620 -83380
rect 74020 -83480 74120 -83380
rect 75520 -83480 75620 -83380
rect 77020 -83480 77120 -83380
rect 78520 -83480 78620 -83380
rect 80020 -83480 80120 -83380
rect 81520 -83480 81620 -83380
rect 83020 -83480 83120 -83380
rect 84520 -83480 84620 -83380
rect 86020 -83480 86120 -83380
rect 87520 -83480 87620 -83380
rect 89020 -83480 89120 -83380
rect 90520 -83480 90620 -83380
rect 92020 -83480 92120 -83380
rect 93520 -83480 93620 -83380
rect 95020 -83480 95120 -83380
rect 96520 -83480 96620 -83380
rect 98020 -83480 98120 -83380
rect 99520 -83480 99620 -83380
rect 101020 -83480 101120 -83380
rect 102520 -83480 102620 -83380
rect 104020 -83480 104120 -83380
rect 105520 -83480 105620 -83380
rect 107020 -83480 107120 -83380
rect 108520 -83480 108620 -83380
rect 110020 -83480 110120 -83380
rect 111520 -83480 111620 -83380
rect 113020 -83480 113120 -83380
rect 114520 -83480 114620 -83380
rect 116020 -83480 116120 -83380
rect 117520 -83480 117620 -83380
rect 119020 -83480 119120 -83380
rect 520 -84980 620 -84880
rect 2020 -84980 2120 -84880
rect 3520 -84980 3620 -84880
rect 5020 -84980 5120 -84880
rect 6520 -84980 6620 -84880
rect 8020 -84980 8120 -84880
rect 9520 -84980 9620 -84880
rect 11020 -84980 11120 -84880
rect 12520 -84980 12620 -84880
rect 14020 -84980 14120 -84880
rect 15520 -84980 15620 -84880
rect 17020 -84980 17120 -84880
rect 18520 -84980 18620 -84880
rect 20020 -84980 20120 -84880
rect 21520 -84980 21620 -84880
rect 23020 -84980 23120 -84880
rect 24520 -84980 24620 -84880
rect 26020 -84980 26120 -84880
rect 27520 -84980 27620 -84880
rect 29020 -84980 29120 -84880
rect 30520 -84980 30620 -84880
rect 32020 -84980 32120 -84880
rect 33520 -84980 33620 -84880
rect 35020 -84980 35120 -84880
rect 36520 -84980 36620 -84880
rect 38020 -84980 38120 -84880
rect 39520 -84980 39620 -84880
rect 41020 -84980 41120 -84880
rect 42520 -84980 42620 -84880
rect 44020 -84980 44120 -84880
rect 45520 -84980 45620 -84880
rect 47020 -84980 47120 -84880
rect 48520 -84980 48620 -84880
rect 50020 -84980 50120 -84880
rect 51520 -84980 51620 -84880
rect 53020 -84980 53120 -84880
rect 54520 -84980 54620 -84880
rect 56020 -84980 56120 -84880
rect 57520 -84980 57620 -84880
rect 59020 -84980 59120 -84880
rect 60520 -84980 60620 -84880
rect 62020 -84980 62120 -84880
rect 63520 -84980 63620 -84880
rect 65020 -84980 65120 -84880
rect 66520 -84980 66620 -84880
rect 68020 -84980 68120 -84880
rect 69520 -84980 69620 -84880
rect 71020 -84980 71120 -84880
rect 72520 -84980 72620 -84880
rect 74020 -84980 74120 -84880
rect 75520 -84980 75620 -84880
rect 77020 -84980 77120 -84880
rect 78520 -84980 78620 -84880
rect 80020 -84980 80120 -84880
rect 81520 -84980 81620 -84880
rect 83020 -84980 83120 -84880
rect 84520 -84980 84620 -84880
rect 86020 -84980 86120 -84880
rect 87520 -84980 87620 -84880
rect 89020 -84980 89120 -84880
rect 90520 -84980 90620 -84880
rect 92020 -84980 92120 -84880
rect 93520 -84980 93620 -84880
rect 95020 -84980 95120 -84880
rect 96520 -84980 96620 -84880
rect 98020 -84980 98120 -84880
rect 99520 -84980 99620 -84880
rect 101020 -84980 101120 -84880
rect 102520 -84980 102620 -84880
rect 104020 -84980 104120 -84880
rect 105520 -84980 105620 -84880
rect 107020 -84980 107120 -84880
rect 108520 -84980 108620 -84880
rect 110020 -84980 110120 -84880
rect 111520 -84980 111620 -84880
rect 113020 -84980 113120 -84880
rect 114520 -84980 114620 -84880
rect 116020 -84980 116120 -84880
rect 117520 -84980 117620 -84880
rect 119020 -84980 119120 -84880
rect 520 -86480 620 -86380
rect 2020 -86480 2120 -86380
rect 3520 -86480 3620 -86380
rect 5020 -86480 5120 -86380
rect 6520 -86480 6620 -86380
rect 8020 -86480 8120 -86380
rect 9520 -86480 9620 -86380
rect 11020 -86480 11120 -86380
rect 12520 -86480 12620 -86380
rect 14020 -86480 14120 -86380
rect 15520 -86480 15620 -86380
rect 17020 -86480 17120 -86380
rect 18520 -86480 18620 -86380
rect 20020 -86480 20120 -86380
rect 21520 -86480 21620 -86380
rect 23020 -86480 23120 -86380
rect 24520 -86480 24620 -86380
rect 26020 -86480 26120 -86380
rect 27520 -86480 27620 -86380
rect 29020 -86480 29120 -86380
rect 30520 -86480 30620 -86380
rect 32020 -86480 32120 -86380
rect 33520 -86480 33620 -86380
rect 35020 -86480 35120 -86380
rect 36520 -86480 36620 -86380
rect 38020 -86480 38120 -86380
rect 39520 -86480 39620 -86380
rect 41020 -86480 41120 -86380
rect 42520 -86480 42620 -86380
rect 44020 -86480 44120 -86380
rect 45520 -86480 45620 -86380
rect 47020 -86480 47120 -86380
rect 48520 -86480 48620 -86380
rect 50020 -86480 50120 -86380
rect 51520 -86480 51620 -86380
rect 53020 -86480 53120 -86380
rect 54520 -86480 54620 -86380
rect 56020 -86480 56120 -86380
rect 57520 -86480 57620 -86380
rect 59020 -86480 59120 -86380
rect 60520 -86480 60620 -86380
rect 62020 -86480 62120 -86380
rect 63520 -86480 63620 -86380
rect 65020 -86480 65120 -86380
rect 66520 -86480 66620 -86380
rect 68020 -86480 68120 -86380
rect 69520 -86480 69620 -86380
rect 71020 -86480 71120 -86380
rect 72520 -86480 72620 -86380
rect 74020 -86480 74120 -86380
rect 75520 -86480 75620 -86380
rect 77020 -86480 77120 -86380
rect 78520 -86480 78620 -86380
rect 80020 -86480 80120 -86380
rect 81520 -86480 81620 -86380
rect 83020 -86480 83120 -86380
rect 84520 -86480 84620 -86380
rect 86020 -86480 86120 -86380
rect 87520 -86480 87620 -86380
rect 89020 -86480 89120 -86380
rect 90520 -86480 90620 -86380
rect 92020 -86480 92120 -86380
rect 93520 -86480 93620 -86380
rect 95020 -86480 95120 -86380
rect 96520 -86480 96620 -86380
rect 98020 -86480 98120 -86380
rect 99520 -86480 99620 -86380
rect 101020 -86480 101120 -86380
rect 102520 -86480 102620 -86380
rect 104020 -86480 104120 -86380
rect 105520 -86480 105620 -86380
rect 107020 -86480 107120 -86380
rect 108520 -86480 108620 -86380
rect 110020 -86480 110120 -86380
rect 111520 -86480 111620 -86380
rect 113020 -86480 113120 -86380
rect 114520 -86480 114620 -86380
rect 116020 -86480 116120 -86380
rect 117520 -86480 117620 -86380
rect 119020 -86480 119120 -86380
rect 520 -87980 620 -87880
rect 2020 -87980 2120 -87880
rect 3520 -87980 3620 -87880
rect 5020 -87980 5120 -87880
rect 6520 -87980 6620 -87880
rect 8020 -87980 8120 -87880
rect 9520 -87980 9620 -87880
rect 11020 -87980 11120 -87880
rect 12520 -87980 12620 -87880
rect 14020 -87980 14120 -87880
rect 15520 -87980 15620 -87880
rect 17020 -87980 17120 -87880
rect 18520 -87980 18620 -87880
rect 20020 -87980 20120 -87880
rect 21520 -87980 21620 -87880
rect 23020 -87980 23120 -87880
rect 24520 -87980 24620 -87880
rect 26020 -87980 26120 -87880
rect 27520 -87980 27620 -87880
rect 29020 -87980 29120 -87880
rect 30520 -87980 30620 -87880
rect 32020 -87980 32120 -87880
rect 33520 -87980 33620 -87880
rect 35020 -87980 35120 -87880
rect 36520 -87980 36620 -87880
rect 38020 -87980 38120 -87880
rect 39520 -87980 39620 -87880
rect 41020 -87980 41120 -87880
rect 42520 -87980 42620 -87880
rect 44020 -87980 44120 -87880
rect 45520 -87980 45620 -87880
rect 47020 -87980 47120 -87880
rect 48520 -87980 48620 -87880
rect 50020 -87980 50120 -87880
rect 51520 -87980 51620 -87880
rect 53020 -87980 53120 -87880
rect 54520 -87980 54620 -87880
rect 56020 -87980 56120 -87880
rect 57520 -87980 57620 -87880
rect 59020 -87980 59120 -87880
rect 60520 -87980 60620 -87880
rect 62020 -87980 62120 -87880
rect 63520 -87980 63620 -87880
rect 65020 -87980 65120 -87880
rect 66520 -87980 66620 -87880
rect 68020 -87980 68120 -87880
rect 69520 -87980 69620 -87880
rect 71020 -87980 71120 -87880
rect 72520 -87980 72620 -87880
rect 74020 -87980 74120 -87880
rect 75520 -87980 75620 -87880
rect 77020 -87980 77120 -87880
rect 78520 -87980 78620 -87880
rect 80020 -87980 80120 -87880
rect 81520 -87980 81620 -87880
rect 83020 -87980 83120 -87880
rect 84520 -87980 84620 -87880
rect 86020 -87980 86120 -87880
rect 87520 -87980 87620 -87880
rect 89020 -87980 89120 -87880
rect 90520 -87980 90620 -87880
rect 92020 -87980 92120 -87880
rect 93520 -87980 93620 -87880
rect 95020 -87980 95120 -87880
rect 96520 -87980 96620 -87880
rect 98020 -87980 98120 -87880
rect 99520 -87980 99620 -87880
rect 101020 -87980 101120 -87880
rect 102520 -87980 102620 -87880
rect 104020 -87980 104120 -87880
rect 105520 -87980 105620 -87880
rect 107020 -87980 107120 -87880
rect 108520 -87980 108620 -87880
rect 110020 -87980 110120 -87880
rect 111520 -87980 111620 -87880
rect 113020 -87980 113120 -87880
rect 114520 -87980 114620 -87880
rect 116020 -87980 116120 -87880
rect 117520 -87980 117620 -87880
rect 119020 -87980 119120 -87880
rect 520 -89480 620 -89380
rect 2020 -89480 2120 -89380
rect 3520 -89480 3620 -89380
rect 5020 -89480 5120 -89380
rect 6520 -89480 6620 -89380
rect 8020 -89480 8120 -89380
rect 9520 -89480 9620 -89380
rect 11020 -89480 11120 -89380
rect 12520 -89480 12620 -89380
rect 14020 -89480 14120 -89380
rect 15520 -89480 15620 -89380
rect 17020 -89480 17120 -89380
rect 18520 -89480 18620 -89380
rect 20020 -89480 20120 -89380
rect 21520 -89480 21620 -89380
rect 23020 -89480 23120 -89380
rect 24520 -89480 24620 -89380
rect 26020 -89480 26120 -89380
rect 27520 -89480 27620 -89380
rect 29020 -89480 29120 -89380
rect 30520 -89480 30620 -89380
rect 32020 -89480 32120 -89380
rect 33520 -89480 33620 -89380
rect 35020 -89480 35120 -89380
rect 36520 -89480 36620 -89380
rect 38020 -89480 38120 -89380
rect 39520 -89480 39620 -89380
rect 41020 -89480 41120 -89380
rect 42520 -89480 42620 -89380
rect 44020 -89480 44120 -89380
rect 45520 -89480 45620 -89380
rect 47020 -89480 47120 -89380
rect 48520 -89480 48620 -89380
rect 50020 -89480 50120 -89380
rect 51520 -89480 51620 -89380
rect 53020 -89480 53120 -89380
rect 54520 -89480 54620 -89380
rect 56020 -89480 56120 -89380
rect 57520 -89480 57620 -89380
rect 59020 -89480 59120 -89380
rect 60520 -89480 60620 -89380
rect 62020 -89480 62120 -89380
rect 63520 -89480 63620 -89380
rect 65020 -89480 65120 -89380
rect 66520 -89480 66620 -89380
rect 68020 -89480 68120 -89380
rect 69520 -89480 69620 -89380
rect 71020 -89480 71120 -89380
rect 72520 -89480 72620 -89380
rect 74020 -89480 74120 -89380
rect 75520 -89480 75620 -89380
rect 77020 -89480 77120 -89380
rect 78520 -89480 78620 -89380
rect 80020 -89480 80120 -89380
rect 81520 -89480 81620 -89380
rect 83020 -89480 83120 -89380
rect 84520 -89480 84620 -89380
rect 86020 -89480 86120 -89380
rect 87520 -89480 87620 -89380
rect 89020 -89480 89120 -89380
rect 90520 -89480 90620 -89380
rect 92020 -89480 92120 -89380
rect 93520 -89480 93620 -89380
rect 95020 -89480 95120 -89380
rect 96520 -89480 96620 -89380
rect 98020 -89480 98120 -89380
rect 99520 -89480 99620 -89380
rect 101020 -89480 101120 -89380
rect 102520 -89480 102620 -89380
rect 104020 -89480 104120 -89380
rect 105520 -89480 105620 -89380
rect 107020 -89480 107120 -89380
rect 108520 -89480 108620 -89380
rect 110020 -89480 110120 -89380
rect 111520 -89480 111620 -89380
rect 113020 -89480 113120 -89380
rect 114520 -89480 114620 -89380
rect 116020 -89480 116120 -89380
rect 117520 -89480 117620 -89380
rect 119020 -89480 119120 -89380
rect 520 -90980 620 -90880
rect 2020 -90980 2120 -90880
rect 3520 -90980 3620 -90880
rect 5020 -90980 5120 -90880
rect 6520 -90980 6620 -90880
rect 8020 -90980 8120 -90880
rect 9520 -90980 9620 -90880
rect 11020 -90980 11120 -90880
rect 12520 -90980 12620 -90880
rect 14020 -90980 14120 -90880
rect 15520 -90980 15620 -90880
rect 17020 -90980 17120 -90880
rect 18520 -90980 18620 -90880
rect 20020 -90980 20120 -90880
rect 21520 -90980 21620 -90880
rect 23020 -90980 23120 -90880
rect 24520 -90980 24620 -90880
rect 26020 -90980 26120 -90880
rect 27520 -90980 27620 -90880
rect 29020 -90980 29120 -90880
rect 30520 -90980 30620 -90880
rect 32020 -90980 32120 -90880
rect 33520 -90980 33620 -90880
rect 35020 -90980 35120 -90880
rect 36520 -90980 36620 -90880
rect 38020 -90980 38120 -90880
rect 39520 -90980 39620 -90880
rect 41020 -90980 41120 -90880
rect 42520 -90980 42620 -90880
rect 44020 -90980 44120 -90880
rect 45520 -90980 45620 -90880
rect 47020 -90980 47120 -90880
rect 48520 -90980 48620 -90880
rect 50020 -90980 50120 -90880
rect 51520 -90980 51620 -90880
rect 53020 -90980 53120 -90880
rect 54520 -90980 54620 -90880
rect 56020 -90980 56120 -90880
rect 57520 -90980 57620 -90880
rect 59020 -90980 59120 -90880
rect 60520 -90980 60620 -90880
rect 62020 -90980 62120 -90880
rect 63520 -90980 63620 -90880
rect 65020 -90980 65120 -90880
rect 66520 -90980 66620 -90880
rect 68020 -90980 68120 -90880
rect 69520 -90980 69620 -90880
rect 71020 -90980 71120 -90880
rect 72520 -90980 72620 -90880
rect 74020 -90980 74120 -90880
rect 75520 -90980 75620 -90880
rect 77020 -90980 77120 -90880
rect 78520 -90980 78620 -90880
rect 80020 -90980 80120 -90880
rect 81520 -90980 81620 -90880
rect 83020 -90980 83120 -90880
rect 84520 -90980 84620 -90880
rect 86020 -90980 86120 -90880
rect 87520 -90980 87620 -90880
rect 89020 -90980 89120 -90880
rect 90520 -90980 90620 -90880
rect 92020 -90980 92120 -90880
rect 93520 -90980 93620 -90880
rect 95020 -90980 95120 -90880
rect 96520 -90980 96620 -90880
rect 98020 -90980 98120 -90880
rect 99520 -90980 99620 -90880
rect 101020 -90980 101120 -90880
rect 102520 -90980 102620 -90880
rect 104020 -90980 104120 -90880
rect 105520 -90980 105620 -90880
rect 107020 -90980 107120 -90880
rect 108520 -90980 108620 -90880
rect 110020 -90980 110120 -90880
rect 111520 -90980 111620 -90880
rect 113020 -90980 113120 -90880
rect 114520 -90980 114620 -90880
rect 116020 -90980 116120 -90880
rect 117520 -90980 117620 -90880
rect 119020 -90980 119120 -90880
rect 520 -92480 620 -92380
rect 2020 -92480 2120 -92380
rect 3520 -92480 3620 -92380
rect 5020 -92480 5120 -92380
rect 6520 -92480 6620 -92380
rect 8020 -92480 8120 -92380
rect 9520 -92480 9620 -92380
rect 11020 -92480 11120 -92380
rect 12520 -92480 12620 -92380
rect 14020 -92480 14120 -92380
rect 15520 -92480 15620 -92380
rect 17020 -92480 17120 -92380
rect 18520 -92480 18620 -92380
rect 20020 -92480 20120 -92380
rect 21520 -92480 21620 -92380
rect 23020 -92480 23120 -92380
rect 24520 -92480 24620 -92380
rect 26020 -92480 26120 -92380
rect 27520 -92480 27620 -92380
rect 29020 -92480 29120 -92380
rect 30520 -92480 30620 -92380
rect 32020 -92480 32120 -92380
rect 33520 -92480 33620 -92380
rect 35020 -92480 35120 -92380
rect 36520 -92480 36620 -92380
rect 38020 -92480 38120 -92380
rect 39520 -92480 39620 -92380
rect 41020 -92480 41120 -92380
rect 42520 -92480 42620 -92380
rect 44020 -92480 44120 -92380
rect 45520 -92480 45620 -92380
rect 47020 -92480 47120 -92380
rect 48520 -92480 48620 -92380
rect 50020 -92480 50120 -92380
rect 51520 -92480 51620 -92380
rect 53020 -92480 53120 -92380
rect 54520 -92480 54620 -92380
rect 56020 -92480 56120 -92380
rect 57520 -92480 57620 -92380
rect 59020 -92480 59120 -92380
rect 60520 -92480 60620 -92380
rect 62020 -92480 62120 -92380
rect 63520 -92480 63620 -92380
rect 65020 -92480 65120 -92380
rect 66520 -92480 66620 -92380
rect 68020 -92480 68120 -92380
rect 69520 -92480 69620 -92380
rect 71020 -92480 71120 -92380
rect 72520 -92480 72620 -92380
rect 74020 -92480 74120 -92380
rect 75520 -92480 75620 -92380
rect 77020 -92480 77120 -92380
rect 78520 -92480 78620 -92380
rect 80020 -92480 80120 -92380
rect 81520 -92480 81620 -92380
rect 83020 -92480 83120 -92380
rect 84520 -92480 84620 -92380
rect 86020 -92480 86120 -92380
rect 87520 -92480 87620 -92380
rect 89020 -92480 89120 -92380
rect 90520 -92480 90620 -92380
rect 92020 -92480 92120 -92380
rect 93520 -92480 93620 -92380
rect 95020 -92480 95120 -92380
rect 96520 -92480 96620 -92380
rect 98020 -92480 98120 -92380
rect 99520 -92480 99620 -92380
rect 101020 -92480 101120 -92380
rect 102520 -92480 102620 -92380
rect 104020 -92480 104120 -92380
rect 105520 -92480 105620 -92380
rect 107020 -92480 107120 -92380
rect 108520 -92480 108620 -92380
rect 110020 -92480 110120 -92380
rect 111520 -92480 111620 -92380
rect 113020 -92480 113120 -92380
rect 114520 -92480 114620 -92380
rect 116020 -92480 116120 -92380
rect 117520 -92480 117620 -92380
rect 119020 -92480 119120 -92380
rect 520 -93980 620 -93880
rect 2020 -93980 2120 -93880
rect 3520 -93980 3620 -93880
rect 5020 -93980 5120 -93880
rect 6520 -93980 6620 -93880
rect 8020 -93980 8120 -93880
rect 9520 -93980 9620 -93880
rect 11020 -93980 11120 -93880
rect 12520 -93980 12620 -93880
rect 14020 -93980 14120 -93880
rect 15520 -93980 15620 -93880
rect 17020 -93980 17120 -93880
rect 18520 -93980 18620 -93880
rect 20020 -93980 20120 -93880
rect 21520 -93980 21620 -93880
rect 23020 -93980 23120 -93880
rect 24520 -93980 24620 -93880
rect 26020 -93980 26120 -93880
rect 27520 -93980 27620 -93880
rect 29020 -93980 29120 -93880
rect 30520 -93980 30620 -93880
rect 32020 -93980 32120 -93880
rect 33520 -93980 33620 -93880
rect 35020 -93980 35120 -93880
rect 36520 -93980 36620 -93880
rect 38020 -93980 38120 -93880
rect 39520 -93980 39620 -93880
rect 41020 -93980 41120 -93880
rect 42520 -93980 42620 -93880
rect 44020 -93980 44120 -93880
rect 45520 -93980 45620 -93880
rect 47020 -93980 47120 -93880
rect 48520 -93980 48620 -93880
rect 50020 -93980 50120 -93880
rect 51520 -93980 51620 -93880
rect 53020 -93980 53120 -93880
rect 54520 -93980 54620 -93880
rect 56020 -93980 56120 -93880
rect 57520 -93980 57620 -93880
rect 59020 -93980 59120 -93880
rect 60520 -93980 60620 -93880
rect 62020 -93980 62120 -93880
rect 63520 -93980 63620 -93880
rect 65020 -93980 65120 -93880
rect 66520 -93980 66620 -93880
rect 68020 -93980 68120 -93880
rect 69520 -93980 69620 -93880
rect 71020 -93980 71120 -93880
rect 72520 -93980 72620 -93880
rect 74020 -93980 74120 -93880
rect 75520 -93980 75620 -93880
rect 77020 -93980 77120 -93880
rect 78520 -93980 78620 -93880
rect 80020 -93980 80120 -93880
rect 81520 -93980 81620 -93880
rect 83020 -93980 83120 -93880
rect 84520 -93980 84620 -93880
rect 86020 -93980 86120 -93880
rect 87520 -93980 87620 -93880
rect 89020 -93980 89120 -93880
rect 90520 -93980 90620 -93880
rect 92020 -93980 92120 -93880
rect 93520 -93980 93620 -93880
rect 95020 -93980 95120 -93880
rect 96520 -93980 96620 -93880
rect 98020 -93980 98120 -93880
rect 99520 -93980 99620 -93880
rect 101020 -93980 101120 -93880
rect 102520 -93980 102620 -93880
rect 104020 -93980 104120 -93880
rect 105520 -93980 105620 -93880
rect 107020 -93980 107120 -93880
rect 108520 -93980 108620 -93880
rect 110020 -93980 110120 -93880
rect 111520 -93980 111620 -93880
rect 113020 -93980 113120 -93880
rect 114520 -93980 114620 -93880
rect 116020 -93980 116120 -93880
rect 117520 -93980 117620 -93880
rect 119020 -93980 119120 -93880
rect 520 -95480 620 -95380
rect 2020 -95480 2120 -95380
rect 3520 -95480 3620 -95380
rect 5020 -95480 5120 -95380
rect 6520 -95480 6620 -95380
rect 8020 -95480 8120 -95380
rect 9520 -95480 9620 -95380
rect 11020 -95480 11120 -95380
rect 12520 -95480 12620 -95380
rect 14020 -95480 14120 -95380
rect 15520 -95480 15620 -95380
rect 17020 -95480 17120 -95380
rect 18520 -95480 18620 -95380
rect 20020 -95480 20120 -95380
rect 21520 -95480 21620 -95380
rect 23020 -95480 23120 -95380
rect 24520 -95480 24620 -95380
rect 26020 -95480 26120 -95380
rect 27520 -95480 27620 -95380
rect 29020 -95480 29120 -95380
rect 30520 -95480 30620 -95380
rect 32020 -95480 32120 -95380
rect 33520 -95480 33620 -95380
rect 35020 -95480 35120 -95380
rect 36520 -95480 36620 -95380
rect 38020 -95480 38120 -95380
rect 39520 -95480 39620 -95380
rect 41020 -95480 41120 -95380
rect 42520 -95480 42620 -95380
rect 44020 -95480 44120 -95380
rect 45520 -95480 45620 -95380
rect 47020 -95480 47120 -95380
rect 48520 -95480 48620 -95380
rect 50020 -95480 50120 -95380
rect 51520 -95480 51620 -95380
rect 53020 -95480 53120 -95380
rect 54520 -95480 54620 -95380
rect 56020 -95480 56120 -95380
rect 57520 -95480 57620 -95380
rect 59020 -95480 59120 -95380
rect 60520 -95480 60620 -95380
rect 62020 -95480 62120 -95380
rect 63520 -95480 63620 -95380
rect 65020 -95480 65120 -95380
rect 66520 -95480 66620 -95380
rect 68020 -95480 68120 -95380
rect 69520 -95480 69620 -95380
rect 71020 -95480 71120 -95380
rect 72520 -95480 72620 -95380
rect 74020 -95480 74120 -95380
rect 75520 -95480 75620 -95380
rect 77020 -95480 77120 -95380
rect 78520 -95480 78620 -95380
rect 80020 -95480 80120 -95380
rect 81520 -95480 81620 -95380
rect 83020 -95480 83120 -95380
rect 84520 -95480 84620 -95380
rect 86020 -95480 86120 -95380
rect 87520 -95480 87620 -95380
rect 89020 -95480 89120 -95380
rect 90520 -95480 90620 -95380
rect 92020 -95480 92120 -95380
rect 93520 -95480 93620 -95380
rect 95020 -95480 95120 -95380
rect 96520 -95480 96620 -95380
rect 98020 -95480 98120 -95380
rect 99520 -95480 99620 -95380
rect 101020 -95480 101120 -95380
rect 102520 -95480 102620 -95380
rect 104020 -95480 104120 -95380
rect 105520 -95480 105620 -95380
rect 107020 -95480 107120 -95380
rect 108520 -95480 108620 -95380
rect 110020 -95480 110120 -95380
rect 111520 -95480 111620 -95380
rect 113020 -95480 113120 -95380
rect 114520 -95480 114620 -95380
rect 116020 -95480 116120 -95380
rect 117520 -95480 117620 -95380
rect 119020 -95480 119120 -95380
rect 520 -96980 620 -96880
rect 2020 -96980 2120 -96880
rect 3520 -96980 3620 -96880
rect 5020 -96980 5120 -96880
rect 6520 -96980 6620 -96880
rect 8020 -96980 8120 -96880
rect 9520 -96980 9620 -96880
rect 11020 -96980 11120 -96880
rect 12520 -96980 12620 -96880
rect 14020 -96980 14120 -96880
rect 15520 -96980 15620 -96880
rect 17020 -96980 17120 -96880
rect 18520 -96980 18620 -96880
rect 20020 -96980 20120 -96880
rect 21520 -96980 21620 -96880
rect 23020 -96980 23120 -96880
rect 24520 -96980 24620 -96880
rect 26020 -96980 26120 -96880
rect 27520 -96980 27620 -96880
rect 29020 -96980 29120 -96880
rect 30520 -96980 30620 -96880
rect 32020 -96980 32120 -96880
rect 33520 -96980 33620 -96880
rect 35020 -96980 35120 -96880
rect 36520 -96980 36620 -96880
rect 38020 -96980 38120 -96880
rect 39520 -96980 39620 -96880
rect 41020 -96980 41120 -96880
rect 42520 -96980 42620 -96880
rect 44020 -96980 44120 -96880
rect 45520 -96980 45620 -96880
rect 47020 -96980 47120 -96880
rect 48520 -96980 48620 -96880
rect 50020 -96980 50120 -96880
rect 51520 -96980 51620 -96880
rect 53020 -96980 53120 -96880
rect 54520 -96980 54620 -96880
rect 56020 -96980 56120 -96880
rect 57520 -96980 57620 -96880
rect 59020 -96980 59120 -96880
rect 60520 -96980 60620 -96880
rect 62020 -96980 62120 -96880
rect 63520 -96980 63620 -96880
rect 65020 -96980 65120 -96880
rect 66520 -96980 66620 -96880
rect 68020 -96980 68120 -96880
rect 69520 -96980 69620 -96880
rect 71020 -96980 71120 -96880
rect 72520 -96980 72620 -96880
rect 74020 -96980 74120 -96880
rect 75520 -96980 75620 -96880
rect 77020 -96980 77120 -96880
rect 78520 -96980 78620 -96880
rect 80020 -96980 80120 -96880
rect 81520 -96980 81620 -96880
rect 83020 -96980 83120 -96880
rect 84520 -96980 84620 -96880
rect 86020 -96980 86120 -96880
rect 87520 -96980 87620 -96880
rect 89020 -96980 89120 -96880
rect 90520 -96980 90620 -96880
rect 92020 -96980 92120 -96880
rect 93520 -96980 93620 -96880
rect 95020 -96980 95120 -96880
rect 96520 -96980 96620 -96880
rect 98020 -96980 98120 -96880
rect 99520 -96980 99620 -96880
rect 101020 -96980 101120 -96880
rect 102520 -96980 102620 -96880
rect 104020 -96980 104120 -96880
rect 105520 -96980 105620 -96880
rect 107020 -96980 107120 -96880
rect 108520 -96980 108620 -96880
rect 110020 -96980 110120 -96880
rect 111520 -96980 111620 -96880
rect 113020 -96980 113120 -96880
rect 114520 -96980 114620 -96880
rect 116020 -96980 116120 -96880
rect 117520 -96980 117620 -96880
rect 119020 -96980 119120 -96880
rect 520 -98480 620 -98380
rect 2020 -98480 2120 -98380
rect 3520 -98480 3620 -98380
rect 5020 -98480 5120 -98380
rect 6520 -98480 6620 -98380
rect 8020 -98480 8120 -98380
rect 9520 -98480 9620 -98380
rect 11020 -98480 11120 -98380
rect 12520 -98480 12620 -98380
rect 14020 -98480 14120 -98380
rect 15520 -98480 15620 -98380
rect 17020 -98480 17120 -98380
rect 18520 -98480 18620 -98380
rect 20020 -98480 20120 -98380
rect 21520 -98480 21620 -98380
rect 23020 -98480 23120 -98380
rect 24520 -98480 24620 -98380
rect 26020 -98480 26120 -98380
rect 27520 -98480 27620 -98380
rect 29020 -98480 29120 -98380
rect 30520 -98480 30620 -98380
rect 32020 -98480 32120 -98380
rect 33520 -98480 33620 -98380
rect 35020 -98480 35120 -98380
rect 36520 -98480 36620 -98380
rect 38020 -98480 38120 -98380
rect 39520 -98480 39620 -98380
rect 41020 -98480 41120 -98380
rect 42520 -98480 42620 -98380
rect 44020 -98480 44120 -98380
rect 45520 -98480 45620 -98380
rect 47020 -98480 47120 -98380
rect 48520 -98480 48620 -98380
rect 50020 -98480 50120 -98380
rect 51520 -98480 51620 -98380
rect 53020 -98480 53120 -98380
rect 54520 -98480 54620 -98380
rect 56020 -98480 56120 -98380
rect 57520 -98480 57620 -98380
rect 59020 -98480 59120 -98380
rect 60520 -98480 60620 -98380
rect 62020 -98480 62120 -98380
rect 63520 -98480 63620 -98380
rect 65020 -98480 65120 -98380
rect 66520 -98480 66620 -98380
rect 68020 -98480 68120 -98380
rect 69520 -98480 69620 -98380
rect 71020 -98480 71120 -98380
rect 72520 -98480 72620 -98380
rect 74020 -98480 74120 -98380
rect 75520 -98480 75620 -98380
rect 77020 -98480 77120 -98380
rect 78520 -98480 78620 -98380
rect 80020 -98480 80120 -98380
rect 81520 -98480 81620 -98380
rect 83020 -98480 83120 -98380
rect 84520 -98480 84620 -98380
rect 86020 -98480 86120 -98380
rect 87520 -98480 87620 -98380
rect 89020 -98480 89120 -98380
rect 90520 -98480 90620 -98380
rect 92020 -98480 92120 -98380
rect 93520 -98480 93620 -98380
rect 95020 -98480 95120 -98380
rect 96520 -98480 96620 -98380
rect 98020 -98480 98120 -98380
rect 99520 -98480 99620 -98380
rect 101020 -98480 101120 -98380
rect 102520 -98480 102620 -98380
rect 104020 -98480 104120 -98380
rect 105520 -98480 105620 -98380
rect 107020 -98480 107120 -98380
rect 108520 -98480 108620 -98380
rect 110020 -98480 110120 -98380
rect 111520 -98480 111620 -98380
rect 113020 -98480 113120 -98380
rect 114520 -98480 114620 -98380
rect 116020 -98480 116120 -98380
rect 117520 -98480 117620 -98380
rect 119020 -98480 119120 -98380
rect 520 -99980 620 -99880
rect 2020 -99980 2120 -99880
rect 3520 -99980 3620 -99880
rect 5020 -99980 5120 -99880
rect 6520 -99980 6620 -99880
rect 8020 -99980 8120 -99880
rect 9520 -99980 9620 -99880
rect 11020 -99980 11120 -99880
rect 12520 -99980 12620 -99880
rect 14020 -99980 14120 -99880
rect 15520 -99980 15620 -99880
rect 17020 -99980 17120 -99880
rect 18520 -99980 18620 -99880
rect 20020 -99980 20120 -99880
rect 21520 -99980 21620 -99880
rect 23020 -99980 23120 -99880
rect 24520 -99980 24620 -99880
rect 26020 -99980 26120 -99880
rect 27520 -99980 27620 -99880
rect 29020 -99980 29120 -99880
rect 30520 -99980 30620 -99880
rect 32020 -99980 32120 -99880
rect 33520 -99980 33620 -99880
rect 35020 -99980 35120 -99880
rect 36520 -99980 36620 -99880
rect 38020 -99980 38120 -99880
rect 39520 -99980 39620 -99880
rect 41020 -99980 41120 -99880
rect 42520 -99980 42620 -99880
rect 44020 -99980 44120 -99880
rect 45520 -99980 45620 -99880
rect 47020 -99980 47120 -99880
rect 48520 -99980 48620 -99880
rect 50020 -99980 50120 -99880
rect 51520 -99980 51620 -99880
rect 53020 -99980 53120 -99880
rect 54520 -99980 54620 -99880
rect 56020 -99980 56120 -99880
rect 57520 -99980 57620 -99880
rect 59020 -99980 59120 -99880
rect 60520 -99980 60620 -99880
rect 62020 -99980 62120 -99880
rect 63520 -99980 63620 -99880
rect 65020 -99980 65120 -99880
rect 66520 -99980 66620 -99880
rect 68020 -99980 68120 -99880
rect 69520 -99980 69620 -99880
rect 71020 -99980 71120 -99880
rect 72520 -99980 72620 -99880
rect 74020 -99980 74120 -99880
rect 75520 -99980 75620 -99880
rect 77020 -99980 77120 -99880
rect 78520 -99980 78620 -99880
rect 80020 -99980 80120 -99880
rect 81520 -99980 81620 -99880
rect 83020 -99980 83120 -99880
rect 84520 -99980 84620 -99880
rect 86020 -99980 86120 -99880
rect 87520 -99980 87620 -99880
rect 89020 -99980 89120 -99880
rect 90520 -99980 90620 -99880
rect 92020 -99980 92120 -99880
rect 93520 -99980 93620 -99880
rect 95020 -99980 95120 -99880
rect 96520 -99980 96620 -99880
rect 98020 -99980 98120 -99880
rect 99520 -99980 99620 -99880
rect 101020 -99980 101120 -99880
rect 102520 -99980 102620 -99880
rect 104020 -99980 104120 -99880
rect 105520 -99980 105620 -99880
rect 107020 -99980 107120 -99880
rect 108520 -99980 108620 -99880
rect 110020 -99980 110120 -99880
rect 111520 -99980 111620 -99880
rect 113020 -99980 113120 -99880
rect 114520 -99980 114620 -99880
rect 116020 -99980 116120 -99880
rect 117520 -99980 117620 -99880
rect 119020 -99980 119120 -99880
rect 520 -101480 620 -101380
rect 2020 -101480 2120 -101380
rect 3520 -101480 3620 -101380
rect 5020 -101480 5120 -101380
rect 6520 -101480 6620 -101380
rect 8020 -101480 8120 -101380
rect 9520 -101480 9620 -101380
rect 11020 -101480 11120 -101380
rect 12520 -101480 12620 -101380
rect 14020 -101480 14120 -101380
rect 15520 -101480 15620 -101380
rect 17020 -101480 17120 -101380
rect 18520 -101480 18620 -101380
rect 20020 -101480 20120 -101380
rect 21520 -101480 21620 -101380
rect 23020 -101480 23120 -101380
rect 24520 -101480 24620 -101380
rect 26020 -101480 26120 -101380
rect 27520 -101480 27620 -101380
rect 29020 -101480 29120 -101380
rect 30520 -101480 30620 -101380
rect 32020 -101480 32120 -101380
rect 33520 -101480 33620 -101380
rect 35020 -101480 35120 -101380
rect 36520 -101480 36620 -101380
rect 38020 -101480 38120 -101380
rect 39520 -101480 39620 -101380
rect 41020 -101480 41120 -101380
rect 42520 -101480 42620 -101380
rect 44020 -101480 44120 -101380
rect 45520 -101480 45620 -101380
rect 47020 -101480 47120 -101380
rect 48520 -101480 48620 -101380
rect 50020 -101480 50120 -101380
rect 51520 -101480 51620 -101380
rect 53020 -101480 53120 -101380
rect 54520 -101480 54620 -101380
rect 56020 -101480 56120 -101380
rect 57520 -101480 57620 -101380
rect 59020 -101480 59120 -101380
rect 60520 -101480 60620 -101380
rect 62020 -101480 62120 -101380
rect 63520 -101480 63620 -101380
rect 65020 -101480 65120 -101380
rect 66520 -101480 66620 -101380
rect 68020 -101480 68120 -101380
rect 69520 -101480 69620 -101380
rect 71020 -101480 71120 -101380
rect 72520 -101480 72620 -101380
rect 74020 -101480 74120 -101380
rect 75520 -101480 75620 -101380
rect 77020 -101480 77120 -101380
rect 78520 -101480 78620 -101380
rect 80020 -101480 80120 -101380
rect 81520 -101480 81620 -101380
rect 83020 -101480 83120 -101380
rect 84520 -101480 84620 -101380
rect 86020 -101480 86120 -101380
rect 87520 -101480 87620 -101380
rect 89020 -101480 89120 -101380
rect 90520 -101480 90620 -101380
rect 92020 -101480 92120 -101380
rect 93520 -101480 93620 -101380
rect 95020 -101480 95120 -101380
rect 96520 -101480 96620 -101380
rect 98020 -101480 98120 -101380
rect 99520 -101480 99620 -101380
rect 101020 -101480 101120 -101380
rect 102520 -101480 102620 -101380
rect 104020 -101480 104120 -101380
rect 105520 -101480 105620 -101380
rect 107020 -101480 107120 -101380
rect 108520 -101480 108620 -101380
rect 110020 -101480 110120 -101380
rect 111520 -101480 111620 -101380
rect 113020 -101480 113120 -101380
rect 114520 -101480 114620 -101380
rect 116020 -101480 116120 -101380
rect 117520 -101480 117620 -101380
rect 119020 -101480 119120 -101380
rect 520 -102980 620 -102880
rect 2020 -102980 2120 -102880
rect 3520 -102980 3620 -102880
rect 5020 -102980 5120 -102880
rect 6520 -102980 6620 -102880
rect 8020 -102980 8120 -102880
rect 9520 -102980 9620 -102880
rect 11020 -102980 11120 -102880
rect 12520 -102980 12620 -102880
rect 14020 -102980 14120 -102880
rect 15520 -102980 15620 -102880
rect 17020 -102980 17120 -102880
rect 18520 -102980 18620 -102880
rect 20020 -102980 20120 -102880
rect 21520 -102980 21620 -102880
rect 23020 -102980 23120 -102880
rect 24520 -102980 24620 -102880
rect 26020 -102980 26120 -102880
rect 27520 -102980 27620 -102880
rect 29020 -102980 29120 -102880
rect 30520 -102980 30620 -102880
rect 32020 -102980 32120 -102880
rect 33520 -102980 33620 -102880
rect 35020 -102980 35120 -102880
rect 36520 -102980 36620 -102880
rect 38020 -102980 38120 -102880
rect 39520 -102980 39620 -102880
rect 41020 -102980 41120 -102880
rect 42520 -102980 42620 -102880
rect 44020 -102980 44120 -102880
rect 45520 -102980 45620 -102880
rect 47020 -102980 47120 -102880
rect 48520 -102980 48620 -102880
rect 50020 -102980 50120 -102880
rect 51520 -102980 51620 -102880
rect 53020 -102980 53120 -102880
rect 54520 -102980 54620 -102880
rect 56020 -102980 56120 -102880
rect 57520 -102980 57620 -102880
rect 59020 -102980 59120 -102880
rect 60520 -102980 60620 -102880
rect 62020 -102980 62120 -102880
rect 63520 -102980 63620 -102880
rect 65020 -102980 65120 -102880
rect 66520 -102980 66620 -102880
rect 68020 -102980 68120 -102880
rect 69520 -102980 69620 -102880
rect 71020 -102980 71120 -102880
rect 72520 -102980 72620 -102880
rect 74020 -102980 74120 -102880
rect 75520 -102980 75620 -102880
rect 77020 -102980 77120 -102880
rect 78520 -102980 78620 -102880
rect 80020 -102980 80120 -102880
rect 81520 -102980 81620 -102880
rect 83020 -102980 83120 -102880
rect 84520 -102980 84620 -102880
rect 86020 -102980 86120 -102880
rect 87520 -102980 87620 -102880
rect 89020 -102980 89120 -102880
rect 90520 -102980 90620 -102880
rect 92020 -102980 92120 -102880
rect 93520 -102980 93620 -102880
rect 95020 -102980 95120 -102880
rect 96520 -102980 96620 -102880
rect 98020 -102980 98120 -102880
rect 99520 -102980 99620 -102880
rect 101020 -102980 101120 -102880
rect 102520 -102980 102620 -102880
rect 104020 -102980 104120 -102880
rect 105520 -102980 105620 -102880
rect 107020 -102980 107120 -102880
rect 108520 -102980 108620 -102880
rect 110020 -102980 110120 -102880
rect 111520 -102980 111620 -102880
rect 113020 -102980 113120 -102880
rect 114520 -102980 114620 -102880
rect 116020 -102980 116120 -102880
rect 117520 -102980 117620 -102880
rect 119020 -102980 119120 -102880
rect 520 -104480 620 -104380
rect 2020 -104480 2120 -104380
rect 3520 -104480 3620 -104380
rect 5020 -104480 5120 -104380
rect 6520 -104480 6620 -104380
rect 8020 -104480 8120 -104380
rect 9520 -104480 9620 -104380
rect 11020 -104480 11120 -104380
rect 12520 -104480 12620 -104380
rect 14020 -104480 14120 -104380
rect 15520 -104480 15620 -104380
rect 17020 -104480 17120 -104380
rect 18520 -104480 18620 -104380
rect 20020 -104480 20120 -104380
rect 21520 -104480 21620 -104380
rect 23020 -104480 23120 -104380
rect 24520 -104480 24620 -104380
rect 26020 -104480 26120 -104380
rect 27520 -104480 27620 -104380
rect 29020 -104480 29120 -104380
rect 30520 -104480 30620 -104380
rect 32020 -104480 32120 -104380
rect 33520 -104480 33620 -104380
rect 35020 -104480 35120 -104380
rect 36520 -104480 36620 -104380
rect 38020 -104480 38120 -104380
rect 39520 -104480 39620 -104380
rect 41020 -104480 41120 -104380
rect 42520 -104480 42620 -104380
rect 44020 -104480 44120 -104380
rect 45520 -104480 45620 -104380
rect 47020 -104480 47120 -104380
rect 48520 -104480 48620 -104380
rect 50020 -104480 50120 -104380
rect 51520 -104480 51620 -104380
rect 53020 -104480 53120 -104380
rect 54520 -104480 54620 -104380
rect 56020 -104480 56120 -104380
rect 57520 -104480 57620 -104380
rect 59020 -104480 59120 -104380
rect 60520 -104480 60620 -104380
rect 62020 -104480 62120 -104380
rect 63520 -104480 63620 -104380
rect 65020 -104480 65120 -104380
rect 66520 -104480 66620 -104380
rect 68020 -104480 68120 -104380
rect 69520 -104480 69620 -104380
rect 71020 -104480 71120 -104380
rect 72520 -104480 72620 -104380
rect 74020 -104480 74120 -104380
rect 75520 -104480 75620 -104380
rect 77020 -104480 77120 -104380
rect 78520 -104480 78620 -104380
rect 80020 -104480 80120 -104380
rect 81520 -104480 81620 -104380
rect 83020 -104480 83120 -104380
rect 84520 -104480 84620 -104380
rect 86020 -104480 86120 -104380
rect 87520 -104480 87620 -104380
rect 89020 -104480 89120 -104380
rect 90520 -104480 90620 -104380
rect 92020 -104480 92120 -104380
rect 93520 -104480 93620 -104380
rect 95020 -104480 95120 -104380
rect 96520 -104480 96620 -104380
rect 98020 -104480 98120 -104380
rect 99520 -104480 99620 -104380
rect 101020 -104480 101120 -104380
rect 102520 -104480 102620 -104380
rect 104020 -104480 104120 -104380
rect 105520 -104480 105620 -104380
rect 107020 -104480 107120 -104380
rect 108520 -104480 108620 -104380
rect 110020 -104480 110120 -104380
rect 111520 -104480 111620 -104380
rect 113020 -104480 113120 -104380
rect 114520 -104480 114620 -104380
rect 116020 -104480 116120 -104380
rect 117520 -104480 117620 -104380
rect 119020 -104480 119120 -104380
rect 520 -105980 620 -105880
rect 2020 -105980 2120 -105880
rect 3520 -105980 3620 -105880
rect 5020 -105980 5120 -105880
rect 6520 -105980 6620 -105880
rect 8020 -105980 8120 -105880
rect 9520 -105980 9620 -105880
rect 11020 -105980 11120 -105880
rect 12520 -105980 12620 -105880
rect 14020 -105980 14120 -105880
rect 15520 -105980 15620 -105880
rect 17020 -105980 17120 -105880
rect 18520 -105980 18620 -105880
rect 20020 -105980 20120 -105880
rect 21520 -105980 21620 -105880
rect 23020 -105980 23120 -105880
rect 24520 -105980 24620 -105880
rect 26020 -105980 26120 -105880
rect 27520 -105980 27620 -105880
rect 29020 -105980 29120 -105880
rect 30520 -105980 30620 -105880
rect 32020 -105980 32120 -105880
rect 33520 -105980 33620 -105880
rect 35020 -105980 35120 -105880
rect 36520 -105980 36620 -105880
rect 38020 -105980 38120 -105880
rect 39520 -105980 39620 -105880
rect 41020 -105980 41120 -105880
rect 42520 -105980 42620 -105880
rect 44020 -105980 44120 -105880
rect 45520 -105980 45620 -105880
rect 47020 -105980 47120 -105880
rect 48520 -105980 48620 -105880
rect 50020 -105980 50120 -105880
rect 51520 -105980 51620 -105880
rect 53020 -105980 53120 -105880
rect 54520 -105980 54620 -105880
rect 56020 -105980 56120 -105880
rect 57520 -105980 57620 -105880
rect 59020 -105980 59120 -105880
rect 60520 -105980 60620 -105880
rect 62020 -105980 62120 -105880
rect 63520 -105980 63620 -105880
rect 65020 -105980 65120 -105880
rect 66520 -105980 66620 -105880
rect 68020 -105980 68120 -105880
rect 69520 -105980 69620 -105880
rect 71020 -105980 71120 -105880
rect 72520 -105980 72620 -105880
rect 74020 -105980 74120 -105880
rect 75520 -105980 75620 -105880
rect 77020 -105980 77120 -105880
rect 78520 -105980 78620 -105880
rect 80020 -105980 80120 -105880
rect 81520 -105980 81620 -105880
rect 83020 -105980 83120 -105880
rect 84520 -105980 84620 -105880
rect 86020 -105980 86120 -105880
rect 87520 -105980 87620 -105880
rect 89020 -105980 89120 -105880
rect 90520 -105980 90620 -105880
rect 92020 -105980 92120 -105880
rect 93520 -105980 93620 -105880
rect 95020 -105980 95120 -105880
rect 96520 -105980 96620 -105880
rect 98020 -105980 98120 -105880
rect 99520 -105980 99620 -105880
rect 101020 -105980 101120 -105880
rect 102520 -105980 102620 -105880
rect 104020 -105980 104120 -105880
rect 105520 -105980 105620 -105880
rect 107020 -105980 107120 -105880
rect 108520 -105980 108620 -105880
rect 110020 -105980 110120 -105880
rect 111520 -105980 111620 -105880
rect 113020 -105980 113120 -105880
rect 114520 -105980 114620 -105880
rect 116020 -105980 116120 -105880
rect 117520 -105980 117620 -105880
rect 119020 -105980 119120 -105880
rect 520 -107480 620 -107380
rect 2020 -107480 2120 -107380
rect 3520 -107480 3620 -107380
rect 5020 -107480 5120 -107380
rect 6520 -107480 6620 -107380
rect 8020 -107480 8120 -107380
rect 9520 -107480 9620 -107380
rect 11020 -107480 11120 -107380
rect 12520 -107480 12620 -107380
rect 14020 -107480 14120 -107380
rect 15520 -107480 15620 -107380
rect 17020 -107480 17120 -107380
rect 18520 -107480 18620 -107380
rect 20020 -107480 20120 -107380
rect 21520 -107480 21620 -107380
rect 23020 -107480 23120 -107380
rect 24520 -107480 24620 -107380
rect 26020 -107480 26120 -107380
rect 27520 -107480 27620 -107380
rect 29020 -107480 29120 -107380
rect 30520 -107480 30620 -107380
rect 32020 -107480 32120 -107380
rect 33520 -107480 33620 -107380
rect 35020 -107480 35120 -107380
rect 36520 -107480 36620 -107380
rect 38020 -107480 38120 -107380
rect 39520 -107480 39620 -107380
rect 41020 -107480 41120 -107380
rect 42520 -107480 42620 -107380
rect 44020 -107480 44120 -107380
rect 45520 -107480 45620 -107380
rect 47020 -107480 47120 -107380
rect 48520 -107480 48620 -107380
rect 50020 -107480 50120 -107380
rect 51520 -107480 51620 -107380
rect 53020 -107480 53120 -107380
rect 54520 -107480 54620 -107380
rect 56020 -107480 56120 -107380
rect 57520 -107480 57620 -107380
rect 59020 -107480 59120 -107380
rect 60520 -107480 60620 -107380
rect 62020 -107480 62120 -107380
rect 63520 -107480 63620 -107380
rect 65020 -107480 65120 -107380
rect 66520 -107480 66620 -107380
rect 68020 -107480 68120 -107380
rect 69520 -107480 69620 -107380
rect 71020 -107480 71120 -107380
rect 72520 -107480 72620 -107380
rect 74020 -107480 74120 -107380
rect 75520 -107480 75620 -107380
rect 77020 -107480 77120 -107380
rect 78520 -107480 78620 -107380
rect 80020 -107480 80120 -107380
rect 81520 -107480 81620 -107380
rect 83020 -107480 83120 -107380
rect 84520 -107480 84620 -107380
rect 86020 -107480 86120 -107380
rect 87520 -107480 87620 -107380
rect 89020 -107480 89120 -107380
rect 90520 -107480 90620 -107380
rect 92020 -107480 92120 -107380
rect 93520 -107480 93620 -107380
rect 95020 -107480 95120 -107380
rect 96520 -107480 96620 -107380
rect 98020 -107480 98120 -107380
rect 99520 -107480 99620 -107380
rect 101020 -107480 101120 -107380
rect 102520 -107480 102620 -107380
rect 104020 -107480 104120 -107380
rect 105520 -107480 105620 -107380
rect 107020 -107480 107120 -107380
rect 108520 -107480 108620 -107380
rect 110020 -107480 110120 -107380
rect 111520 -107480 111620 -107380
rect 113020 -107480 113120 -107380
rect 114520 -107480 114620 -107380
rect 116020 -107480 116120 -107380
rect 117520 -107480 117620 -107380
rect 119020 -107480 119120 -107380
rect 520 -108980 620 -108880
rect 2020 -108980 2120 -108880
rect 3520 -108980 3620 -108880
rect 5020 -108980 5120 -108880
rect 6520 -108980 6620 -108880
rect 8020 -108980 8120 -108880
rect 9520 -108980 9620 -108880
rect 11020 -108980 11120 -108880
rect 12520 -108980 12620 -108880
rect 14020 -108980 14120 -108880
rect 15520 -108980 15620 -108880
rect 17020 -108980 17120 -108880
rect 18520 -108980 18620 -108880
rect 20020 -108980 20120 -108880
rect 21520 -108980 21620 -108880
rect 23020 -108980 23120 -108880
rect 24520 -108980 24620 -108880
rect 26020 -108980 26120 -108880
rect 27520 -108980 27620 -108880
rect 29020 -108980 29120 -108880
rect 30520 -108980 30620 -108880
rect 32020 -108980 32120 -108880
rect 33520 -108980 33620 -108880
rect 35020 -108980 35120 -108880
rect 36520 -108980 36620 -108880
rect 38020 -108980 38120 -108880
rect 39520 -108980 39620 -108880
rect 41020 -108980 41120 -108880
rect 42520 -108980 42620 -108880
rect 44020 -108980 44120 -108880
rect 45520 -108980 45620 -108880
rect 47020 -108980 47120 -108880
rect 48520 -108980 48620 -108880
rect 50020 -108980 50120 -108880
rect 51520 -108980 51620 -108880
rect 53020 -108980 53120 -108880
rect 54520 -108980 54620 -108880
rect 56020 -108980 56120 -108880
rect 57520 -108980 57620 -108880
rect 59020 -108980 59120 -108880
rect 60520 -108980 60620 -108880
rect 62020 -108980 62120 -108880
rect 63520 -108980 63620 -108880
rect 65020 -108980 65120 -108880
rect 66520 -108980 66620 -108880
rect 68020 -108980 68120 -108880
rect 69520 -108980 69620 -108880
rect 71020 -108980 71120 -108880
rect 72520 -108980 72620 -108880
rect 74020 -108980 74120 -108880
rect 75520 -108980 75620 -108880
rect 77020 -108980 77120 -108880
rect 78520 -108980 78620 -108880
rect 80020 -108980 80120 -108880
rect 81520 -108980 81620 -108880
rect 83020 -108980 83120 -108880
rect 84520 -108980 84620 -108880
rect 86020 -108980 86120 -108880
rect 87520 -108980 87620 -108880
rect 89020 -108980 89120 -108880
rect 90520 -108980 90620 -108880
rect 92020 -108980 92120 -108880
rect 93520 -108980 93620 -108880
rect 95020 -108980 95120 -108880
rect 96520 -108980 96620 -108880
rect 98020 -108980 98120 -108880
rect 99520 -108980 99620 -108880
rect 101020 -108980 101120 -108880
rect 102520 -108980 102620 -108880
rect 104020 -108980 104120 -108880
rect 105520 -108980 105620 -108880
rect 107020 -108980 107120 -108880
rect 108520 -108980 108620 -108880
rect 110020 -108980 110120 -108880
rect 111520 -108980 111620 -108880
rect 113020 -108980 113120 -108880
rect 114520 -108980 114620 -108880
rect 116020 -108980 116120 -108880
rect 117520 -108980 117620 -108880
rect 119020 -108980 119120 -108880
rect 520 -110480 620 -110380
rect 2020 -110480 2120 -110380
rect 3520 -110480 3620 -110380
rect 5020 -110480 5120 -110380
rect 6520 -110480 6620 -110380
rect 8020 -110480 8120 -110380
rect 9520 -110480 9620 -110380
rect 11020 -110480 11120 -110380
rect 12520 -110480 12620 -110380
rect 14020 -110480 14120 -110380
rect 15520 -110480 15620 -110380
rect 17020 -110480 17120 -110380
rect 18520 -110480 18620 -110380
rect 20020 -110480 20120 -110380
rect 21520 -110480 21620 -110380
rect 23020 -110480 23120 -110380
rect 24520 -110480 24620 -110380
rect 26020 -110480 26120 -110380
rect 27520 -110480 27620 -110380
rect 29020 -110480 29120 -110380
rect 30520 -110480 30620 -110380
rect 32020 -110480 32120 -110380
rect 33520 -110480 33620 -110380
rect 35020 -110480 35120 -110380
rect 36520 -110480 36620 -110380
rect 38020 -110480 38120 -110380
rect 39520 -110480 39620 -110380
rect 41020 -110480 41120 -110380
rect 42520 -110480 42620 -110380
rect 44020 -110480 44120 -110380
rect 45520 -110480 45620 -110380
rect 47020 -110480 47120 -110380
rect 48520 -110480 48620 -110380
rect 50020 -110480 50120 -110380
rect 51520 -110480 51620 -110380
rect 53020 -110480 53120 -110380
rect 54520 -110480 54620 -110380
rect 56020 -110480 56120 -110380
rect 57520 -110480 57620 -110380
rect 59020 -110480 59120 -110380
rect 60520 -110480 60620 -110380
rect 62020 -110480 62120 -110380
rect 63520 -110480 63620 -110380
rect 65020 -110480 65120 -110380
rect 66520 -110480 66620 -110380
rect 68020 -110480 68120 -110380
rect 69520 -110480 69620 -110380
rect 71020 -110480 71120 -110380
rect 72520 -110480 72620 -110380
rect 74020 -110480 74120 -110380
rect 75520 -110480 75620 -110380
rect 77020 -110480 77120 -110380
rect 78520 -110480 78620 -110380
rect 80020 -110480 80120 -110380
rect 81520 -110480 81620 -110380
rect 83020 -110480 83120 -110380
rect 84520 -110480 84620 -110380
rect 86020 -110480 86120 -110380
rect 87520 -110480 87620 -110380
rect 89020 -110480 89120 -110380
rect 90520 -110480 90620 -110380
rect 92020 -110480 92120 -110380
rect 93520 -110480 93620 -110380
rect 95020 -110480 95120 -110380
rect 96520 -110480 96620 -110380
rect 98020 -110480 98120 -110380
rect 99520 -110480 99620 -110380
rect 101020 -110480 101120 -110380
rect 102520 -110480 102620 -110380
rect 104020 -110480 104120 -110380
rect 105520 -110480 105620 -110380
rect 107020 -110480 107120 -110380
rect 108520 -110480 108620 -110380
rect 110020 -110480 110120 -110380
rect 111520 -110480 111620 -110380
rect 113020 -110480 113120 -110380
rect 114520 -110480 114620 -110380
rect 116020 -110480 116120 -110380
rect 117520 -110480 117620 -110380
rect 119020 -110480 119120 -110380
rect 520 -111980 620 -111880
rect 2020 -111980 2120 -111880
rect 3520 -111980 3620 -111880
rect 5020 -111980 5120 -111880
rect 6520 -111980 6620 -111880
rect 8020 -111980 8120 -111880
rect 9520 -111980 9620 -111880
rect 11020 -111980 11120 -111880
rect 12520 -111980 12620 -111880
rect 14020 -111980 14120 -111880
rect 15520 -111980 15620 -111880
rect 17020 -111980 17120 -111880
rect 18520 -111980 18620 -111880
rect 20020 -111980 20120 -111880
rect 21520 -111980 21620 -111880
rect 23020 -111980 23120 -111880
rect 24520 -111980 24620 -111880
rect 26020 -111980 26120 -111880
rect 27520 -111980 27620 -111880
rect 29020 -111980 29120 -111880
rect 30520 -111980 30620 -111880
rect 32020 -111980 32120 -111880
rect 33520 -111980 33620 -111880
rect 35020 -111980 35120 -111880
rect 36520 -111980 36620 -111880
rect 38020 -111980 38120 -111880
rect 39520 -111980 39620 -111880
rect 41020 -111980 41120 -111880
rect 42520 -111980 42620 -111880
rect 44020 -111980 44120 -111880
rect 45520 -111980 45620 -111880
rect 47020 -111980 47120 -111880
rect 48520 -111980 48620 -111880
rect 50020 -111980 50120 -111880
rect 51520 -111980 51620 -111880
rect 53020 -111980 53120 -111880
rect 54520 -111980 54620 -111880
rect 56020 -111980 56120 -111880
rect 57520 -111980 57620 -111880
rect 59020 -111980 59120 -111880
rect 60520 -111980 60620 -111880
rect 62020 -111980 62120 -111880
rect 63520 -111980 63620 -111880
rect 65020 -111980 65120 -111880
rect 66520 -111980 66620 -111880
rect 68020 -111980 68120 -111880
rect 69520 -111980 69620 -111880
rect 71020 -111980 71120 -111880
rect 72520 -111980 72620 -111880
rect 74020 -111980 74120 -111880
rect 75520 -111980 75620 -111880
rect 77020 -111980 77120 -111880
rect 78520 -111980 78620 -111880
rect 80020 -111980 80120 -111880
rect 81520 -111980 81620 -111880
rect 83020 -111980 83120 -111880
rect 84520 -111980 84620 -111880
rect 86020 -111980 86120 -111880
rect 87520 -111980 87620 -111880
rect 89020 -111980 89120 -111880
rect 90520 -111980 90620 -111880
rect 92020 -111980 92120 -111880
rect 93520 -111980 93620 -111880
rect 95020 -111980 95120 -111880
rect 96520 -111980 96620 -111880
rect 98020 -111980 98120 -111880
rect 99520 -111980 99620 -111880
rect 101020 -111980 101120 -111880
rect 102520 -111980 102620 -111880
rect 104020 -111980 104120 -111880
rect 105520 -111980 105620 -111880
rect 107020 -111980 107120 -111880
rect 108520 -111980 108620 -111880
rect 110020 -111980 110120 -111880
rect 111520 -111980 111620 -111880
rect 113020 -111980 113120 -111880
rect 114520 -111980 114620 -111880
rect 116020 -111980 116120 -111880
rect 117520 -111980 117620 -111880
rect 119020 -111980 119120 -111880
rect 520 -113480 620 -113380
rect 2020 -113480 2120 -113380
rect 3520 -113480 3620 -113380
rect 5020 -113480 5120 -113380
rect 6520 -113480 6620 -113380
rect 8020 -113480 8120 -113380
rect 9520 -113480 9620 -113380
rect 11020 -113480 11120 -113380
rect 12520 -113480 12620 -113380
rect 14020 -113480 14120 -113380
rect 15520 -113480 15620 -113380
rect 17020 -113480 17120 -113380
rect 18520 -113480 18620 -113380
rect 20020 -113480 20120 -113380
rect 21520 -113480 21620 -113380
rect 23020 -113480 23120 -113380
rect 24520 -113480 24620 -113380
rect 26020 -113480 26120 -113380
rect 27520 -113480 27620 -113380
rect 29020 -113480 29120 -113380
rect 30520 -113480 30620 -113380
rect 32020 -113480 32120 -113380
rect 33520 -113480 33620 -113380
rect 35020 -113480 35120 -113380
rect 36520 -113480 36620 -113380
rect 38020 -113480 38120 -113380
rect 39520 -113480 39620 -113380
rect 41020 -113480 41120 -113380
rect 42520 -113480 42620 -113380
rect 44020 -113480 44120 -113380
rect 45520 -113480 45620 -113380
rect 47020 -113480 47120 -113380
rect 48520 -113480 48620 -113380
rect 50020 -113480 50120 -113380
rect 51520 -113480 51620 -113380
rect 53020 -113480 53120 -113380
rect 54520 -113480 54620 -113380
rect 56020 -113480 56120 -113380
rect 57520 -113480 57620 -113380
rect 59020 -113480 59120 -113380
rect 60520 -113480 60620 -113380
rect 62020 -113480 62120 -113380
rect 63520 -113480 63620 -113380
rect 65020 -113480 65120 -113380
rect 66520 -113480 66620 -113380
rect 68020 -113480 68120 -113380
rect 69520 -113480 69620 -113380
rect 71020 -113480 71120 -113380
rect 72520 -113480 72620 -113380
rect 74020 -113480 74120 -113380
rect 75520 -113480 75620 -113380
rect 77020 -113480 77120 -113380
rect 78520 -113480 78620 -113380
rect 80020 -113480 80120 -113380
rect 81520 -113480 81620 -113380
rect 83020 -113480 83120 -113380
rect 84520 -113480 84620 -113380
rect 86020 -113480 86120 -113380
rect 87520 -113480 87620 -113380
rect 89020 -113480 89120 -113380
rect 90520 -113480 90620 -113380
rect 92020 -113480 92120 -113380
rect 93520 -113480 93620 -113380
rect 95020 -113480 95120 -113380
rect 96520 -113480 96620 -113380
rect 98020 -113480 98120 -113380
rect 99520 -113480 99620 -113380
rect 101020 -113480 101120 -113380
rect 102520 -113480 102620 -113380
rect 104020 -113480 104120 -113380
rect 105520 -113480 105620 -113380
rect 107020 -113480 107120 -113380
rect 108520 -113480 108620 -113380
rect 110020 -113480 110120 -113380
rect 111520 -113480 111620 -113380
rect 113020 -113480 113120 -113380
rect 114520 -113480 114620 -113380
rect 116020 -113480 116120 -113380
rect 117520 -113480 117620 -113380
rect 119020 -113480 119120 -113380
rect 520 -114980 620 -114880
rect 2020 -114980 2120 -114880
rect 3520 -114980 3620 -114880
rect 5020 -114980 5120 -114880
rect 6520 -114980 6620 -114880
rect 8020 -114980 8120 -114880
rect 9520 -114980 9620 -114880
rect 11020 -114980 11120 -114880
rect 12520 -114980 12620 -114880
rect 14020 -114980 14120 -114880
rect 15520 -114980 15620 -114880
rect 17020 -114980 17120 -114880
rect 18520 -114980 18620 -114880
rect 20020 -114980 20120 -114880
rect 21520 -114980 21620 -114880
rect 23020 -114980 23120 -114880
rect 24520 -114980 24620 -114880
rect 26020 -114980 26120 -114880
rect 27520 -114980 27620 -114880
rect 29020 -114980 29120 -114880
rect 30520 -114980 30620 -114880
rect 32020 -114980 32120 -114880
rect 33520 -114980 33620 -114880
rect 35020 -114980 35120 -114880
rect 36520 -114980 36620 -114880
rect 38020 -114980 38120 -114880
rect 39520 -114980 39620 -114880
rect 41020 -114980 41120 -114880
rect 42520 -114980 42620 -114880
rect 44020 -114980 44120 -114880
rect 45520 -114980 45620 -114880
rect 47020 -114980 47120 -114880
rect 48520 -114980 48620 -114880
rect 50020 -114980 50120 -114880
rect 51520 -114980 51620 -114880
rect 53020 -114980 53120 -114880
rect 54520 -114980 54620 -114880
rect 56020 -114980 56120 -114880
rect 57520 -114980 57620 -114880
rect 59020 -114980 59120 -114880
rect 60520 -114980 60620 -114880
rect 62020 -114980 62120 -114880
rect 63520 -114980 63620 -114880
rect 65020 -114980 65120 -114880
rect 66520 -114980 66620 -114880
rect 68020 -114980 68120 -114880
rect 69520 -114980 69620 -114880
rect 71020 -114980 71120 -114880
rect 72520 -114980 72620 -114880
rect 74020 -114980 74120 -114880
rect 75520 -114980 75620 -114880
rect 77020 -114980 77120 -114880
rect 78520 -114980 78620 -114880
rect 80020 -114980 80120 -114880
rect 81520 -114980 81620 -114880
rect 83020 -114980 83120 -114880
rect 84520 -114980 84620 -114880
rect 86020 -114980 86120 -114880
rect 87520 -114980 87620 -114880
rect 89020 -114980 89120 -114880
rect 90520 -114980 90620 -114880
rect 92020 -114980 92120 -114880
rect 93520 -114980 93620 -114880
rect 95020 -114980 95120 -114880
rect 96520 -114980 96620 -114880
rect 98020 -114980 98120 -114880
rect 99520 -114980 99620 -114880
rect 101020 -114980 101120 -114880
rect 102520 -114980 102620 -114880
rect 104020 -114980 104120 -114880
rect 105520 -114980 105620 -114880
rect 107020 -114980 107120 -114880
rect 108520 -114980 108620 -114880
rect 110020 -114980 110120 -114880
rect 111520 -114980 111620 -114880
rect 113020 -114980 113120 -114880
rect 114520 -114980 114620 -114880
rect 116020 -114980 116120 -114880
rect 117520 -114980 117620 -114880
rect 119020 -114980 119120 -114880
rect 520 -116480 620 -116380
rect 2020 -116480 2120 -116380
rect 3520 -116480 3620 -116380
rect 5020 -116480 5120 -116380
rect 6520 -116480 6620 -116380
rect 8020 -116480 8120 -116380
rect 9520 -116480 9620 -116380
rect 11020 -116480 11120 -116380
rect 12520 -116480 12620 -116380
rect 14020 -116480 14120 -116380
rect 15520 -116480 15620 -116380
rect 17020 -116480 17120 -116380
rect 18520 -116480 18620 -116380
rect 20020 -116480 20120 -116380
rect 21520 -116480 21620 -116380
rect 23020 -116480 23120 -116380
rect 24520 -116480 24620 -116380
rect 26020 -116480 26120 -116380
rect 27520 -116480 27620 -116380
rect 29020 -116480 29120 -116380
rect 30520 -116480 30620 -116380
rect 32020 -116480 32120 -116380
rect 33520 -116480 33620 -116380
rect 35020 -116480 35120 -116380
rect 36520 -116480 36620 -116380
rect 38020 -116480 38120 -116380
rect 39520 -116480 39620 -116380
rect 41020 -116480 41120 -116380
rect 42520 -116480 42620 -116380
rect 44020 -116480 44120 -116380
rect 45520 -116480 45620 -116380
rect 47020 -116480 47120 -116380
rect 48520 -116480 48620 -116380
rect 50020 -116480 50120 -116380
rect 51520 -116480 51620 -116380
rect 53020 -116480 53120 -116380
rect 54520 -116480 54620 -116380
rect 56020 -116480 56120 -116380
rect 57520 -116480 57620 -116380
rect 59020 -116480 59120 -116380
rect 60520 -116480 60620 -116380
rect 62020 -116480 62120 -116380
rect 63520 -116480 63620 -116380
rect 65020 -116480 65120 -116380
rect 66520 -116480 66620 -116380
rect 68020 -116480 68120 -116380
rect 69520 -116480 69620 -116380
rect 71020 -116480 71120 -116380
rect 72520 -116480 72620 -116380
rect 74020 -116480 74120 -116380
rect 75520 -116480 75620 -116380
rect 77020 -116480 77120 -116380
rect 78520 -116480 78620 -116380
rect 80020 -116480 80120 -116380
rect 81520 -116480 81620 -116380
rect 83020 -116480 83120 -116380
rect 84520 -116480 84620 -116380
rect 86020 -116480 86120 -116380
rect 87520 -116480 87620 -116380
rect 89020 -116480 89120 -116380
rect 90520 -116480 90620 -116380
rect 92020 -116480 92120 -116380
rect 93520 -116480 93620 -116380
rect 95020 -116480 95120 -116380
rect 96520 -116480 96620 -116380
rect 98020 -116480 98120 -116380
rect 99520 -116480 99620 -116380
rect 101020 -116480 101120 -116380
rect 102520 -116480 102620 -116380
rect 104020 -116480 104120 -116380
rect 105520 -116480 105620 -116380
rect 107020 -116480 107120 -116380
rect 108520 -116480 108620 -116380
rect 110020 -116480 110120 -116380
rect 111520 -116480 111620 -116380
rect 113020 -116480 113120 -116380
rect 114520 -116480 114620 -116380
rect 116020 -116480 116120 -116380
rect 117520 -116480 117620 -116380
rect 119020 -116480 119120 -116380
rect 520 -117980 620 -117880
rect 2020 -117980 2120 -117880
rect 3520 -117980 3620 -117880
rect 5020 -117980 5120 -117880
rect 6520 -117980 6620 -117880
rect 8020 -117980 8120 -117880
rect 9520 -117980 9620 -117880
rect 11020 -117980 11120 -117880
rect 12520 -117980 12620 -117880
rect 14020 -117980 14120 -117880
rect 15520 -117980 15620 -117880
rect 17020 -117980 17120 -117880
rect 18520 -117980 18620 -117880
rect 20020 -117980 20120 -117880
rect 21520 -117980 21620 -117880
rect 23020 -117980 23120 -117880
rect 24520 -117980 24620 -117880
rect 26020 -117980 26120 -117880
rect 27520 -117980 27620 -117880
rect 29020 -117980 29120 -117880
rect 30520 -117980 30620 -117880
rect 32020 -117980 32120 -117880
rect 33520 -117980 33620 -117880
rect 35020 -117980 35120 -117880
rect 36520 -117980 36620 -117880
rect 38020 -117980 38120 -117880
rect 39520 -117980 39620 -117880
rect 41020 -117980 41120 -117880
rect 42520 -117980 42620 -117880
rect 44020 -117980 44120 -117880
rect 45520 -117980 45620 -117880
rect 47020 -117980 47120 -117880
rect 48520 -117980 48620 -117880
rect 50020 -117980 50120 -117880
rect 51520 -117980 51620 -117880
rect 53020 -117980 53120 -117880
rect 54520 -117980 54620 -117880
rect 56020 -117980 56120 -117880
rect 57520 -117980 57620 -117880
rect 59020 -117980 59120 -117880
rect 60520 -117980 60620 -117880
rect 62020 -117980 62120 -117880
rect 63520 -117980 63620 -117880
rect 65020 -117980 65120 -117880
rect 66520 -117980 66620 -117880
rect 68020 -117980 68120 -117880
rect 69520 -117980 69620 -117880
rect 71020 -117980 71120 -117880
rect 72520 -117980 72620 -117880
rect 74020 -117980 74120 -117880
rect 75520 -117980 75620 -117880
rect 77020 -117980 77120 -117880
rect 78520 -117980 78620 -117880
rect 80020 -117980 80120 -117880
rect 81520 -117980 81620 -117880
rect 83020 -117980 83120 -117880
rect 84520 -117980 84620 -117880
rect 86020 -117980 86120 -117880
rect 87520 -117980 87620 -117880
rect 89020 -117980 89120 -117880
rect 90520 -117980 90620 -117880
rect 92020 -117980 92120 -117880
rect 93520 -117980 93620 -117880
rect 95020 -117980 95120 -117880
rect 96520 -117980 96620 -117880
rect 98020 -117980 98120 -117880
rect 99520 -117980 99620 -117880
rect 101020 -117980 101120 -117880
rect 102520 -117980 102620 -117880
rect 104020 -117980 104120 -117880
rect 105520 -117980 105620 -117880
rect 107020 -117980 107120 -117880
rect 108520 -117980 108620 -117880
rect 110020 -117980 110120 -117880
rect 111520 -117980 111620 -117880
rect 113020 -117980 113120 -117880
rect 114520 -117980 114620 -117880
rect 116020 -117980 116120 -117880
rect 117520 -117980 117620 -117880
rect 119020 -117980 119120 -117880
use pixel  pixel_6320
timestamp 1654648307
transform 1 0 -1900 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6322
timestamp 1654648307
transform 1 0 1100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6321
timestamp 1654648307
transform 1 0 -400 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6324
timestamp 1654648307
transform 1 0 4100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6323
timestamp 1654648307
transform 1 0 2600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6326
timestamp 1654648307
transform 1 0 7100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6325
timestamp 1654648307
transform 1 0 5600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6328
timestamp 1654648307
transform 1 0 10100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6327
timestamp 1654648307
transform 1 0 8600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6330
timestamp 1654648307
transform 1 0 13100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6329
timestamp 1654648307
transform 1 0 11600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6332
timestamp 1654648307
transform 1 0 16100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6331
timestamp 1654648307
transform 1 0 14600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6334
timestamp 1654648307
transform 1 0 19100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6333
timestamp 1654648307
transform 1 0 17600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6336
timestamp 1654648307
transform 1 0 22100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6335
timestamp 1654648307
transform 1 0 20600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6338
timestamp 1654648307
transform 1 0 25100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6337
timestamp 1654648307
transform 1 0 23600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6340
timestamp 1654648307
transform 1 0 28100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6339
timestamp 1654648307
transform 1 0 26600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6342
timestamp 1654648307
transform 1 0 31100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6341
timestamp 1654648307
transform 1 0 29600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6344
timestamp 1654648307
transform 1 0 34100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6343
timestamp 1654648307
transform 1 0 32600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6346
timestamp 1654648307
transform 1 0 37100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6345
timestamp 1654648307
transform 1 0 35600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6348
timestamp 1654648307
transform 1 0 40100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6347
timestamp 1654648307
transform 1 0 38600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6350
timestamp 1654648307
transform 1 0 43100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6349
timestamp 1654648307
transform 1 0 41600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6352
timestamp 1654648307
transform 1 0 46100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6351
timestamp 1654648307
transform 1 0 44600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6354
timestamp 1654648307
transform 1 0 49100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6353
timestamp 1654648307
transform 1 0 47600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6356
timestamp 1654648307
transform 1 0 52100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6355
timestamp 1654648307
transform 1 0 50600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6358
timestamp 1654648307
transform 1 0 55100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6357
timestamp 1654648307
transform 1 0 53600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6360
timestamp 1654648307
transform 1 0 58100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6359
timestamp 1654648307
transform 1 0 56600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6362
timestamp 1654648307
transform 1 0 61100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6361
timestamp 1654648307
transform 1 0 59600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6364
timestamp 1654648307
transform 1 0 64100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6363
timestamp 1654648307
transform 1 0 62600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6366
timestamp 1654648307
transform 1 0 67100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6365
timestamp 1654648307
transform 1 0 65600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6368
timestamp 1654648307
transform 1 0 70100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6367
timestamp 1654648307
transform 1 0 68600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6370
timestamp 1654648307
transform 1 0 73100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6369
timestamp 1654648307
transform 1 0 71600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6372
timestamp 1654648307
transform 1 0 76100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6371
timestamp 1654648307
transform 1 0 74600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6374
timestamp 1654648307
transform 1 0 79100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6373
timestamp 1654648307
transform 1 0 77600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6376
timestamp 1654648307
transform 1 0 82100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6375
timestamp 1654648307
transform 1 0 80600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6378
timestamp 1654648307
transform 1 0 85100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6377
timestamp 1654648307
transform 1 0 83600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6380
timestamp 1654648307
transform 1 0 88100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6379
timestamp 1654648307
transform 1 0 86600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6382
timestamp 1654648307
transform 1 0 91100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6381
timestamp 1654648307
transform 1 0 89600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6384
timestamp 1654648307
transform 1 0 94100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6383
timestamp 1654648307
transform 1 0 92600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6386
timestamp 1654648307
transform 1 0 97100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6385
timestamp 1654648307
transform 1 0 95600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6388
timestamp 1654648307
transform 1 0 100100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6387
timestamp 1654648307
transform 1 0 98600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6390
timestamp 1654648307
transform 1 0 103100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6389
timestamp 1654648307
transform 1 0 101600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6392
timestamp 1654648307
transform 1 0 106100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6391
timestamp 1654648307
transform 1 0 104600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6394
timestamp 1654648307
transform 1 0 109100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6393
timestamp 1654648307
transform 1 0 107600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6396
timestamp 1654648307
transform 1 0 112100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6395
timestamp 1654648307
transform 1 0 110600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6398
timestamp 1654648307
transform 1 0 115100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6397
timestamp 1654648307
transform 1 0 113600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6399
timestamp 1654648307
transform 1 0 116600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_6240
timestamp 1654648307
transform 1 0 -1900 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6160
timestamp 1654648307
transform 1 0 -1900 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6242
timestamp 1654648307
transform 1 0 1100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6241
timestamp 1654648307
transform 1 0 -400 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6162
timestamp 1654648307
transform 1 0 1100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6161
timestamp 1654648307
transform 1 0 -400 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6244
timestamp 1654648307
transform 1 0 4100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6243
timestamp 1654648307
transform 1 0 2600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6164
timestamp 1654648307
transform 1 0 4100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6163
timestamp 1654648307
transform 1 0 2600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6246
timestamp 1654648307
transform 1 0 7100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6245
timestamp 1654648307
transform 1 0 5600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6166
timestamp 1654648307
transform 1 0 7100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6165
timestamp 1654648307
transform 1 0 5600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6248
timestamp 1654648307
transform 1 0 10100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6247
timestamp 1654648307
transform 1 0 8600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6168
timestamp 1654648307
transform 1 0 10100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6167
timestamp 1654648307
transform 1 0 8600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6250
timestamp 1654648307
transform 1 0 13100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6249
timestamp 1654648307
transform 1 0 11600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6170
timestamp 1654648307
transform 1 0 13100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6169
timestamp 1654648307
transform 1 0 11600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6252
timestamp 1654648307
transform 1 0 16100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6251
timestamp 1654648307
transform 1 0 14600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6172
timestamp 1654648307
transform 1 0 16100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6171
timestamp 1654648307
transform 1 0 14600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6254
timestamp 1654648307
transform 1 0 19100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6253
timestamp 1654648307
transform 1 0 17600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6174
timestamp 1654648307
transform 1 0 19100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6173
timestamp 1654648307
transform 1 0 17600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6256
timestamp 1654648307
transform 1 0 22100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6255
timestamp 1654648307
transform 1 0 20600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6176
timestamp 1654648307
transform 1 0 22100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6175
timestamp 1654648307
transform 1 0 20600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6258
timestamp 1654648307
transform 1 0 25100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6257
timestamp 1654648307
transform 1 0 23600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6178
timestamp 1654648307
transform 1 0 25100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6177
timestamp 1654648307
transform 1 0 23600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6260
timestamp 1654648307
transform 1 0 28100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6259
timestamp 1654648307
transform 1 0 26600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6180
timestamp 1654648307
transform 1 0 28100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6179
timestamp 1654648307
transform 1 0 26600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6262
timestamp 1654648307
transform 1 0 31100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6261
timestamp 1654648307
transform 1 0 29600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6182
timestamp 1654648307
transform 1 0 31100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6181
timestamp 1654648307
transform 1 0 29600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6264
timestamp 1654648307
transform 1 0 34100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6263
timestamp 1654648307
transform 1 0 32600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6184
timestamp 1654648307
transform 1 0 34100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6183
timestamp 1654648307
transform 1 0 32600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6266
timestamp 1654648307
transform 1 0 37100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6265
timestamp 1654648307
transform 1 0 35600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6186
timestamp 1654648307
transform 1 0 37100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6185
timestamp 1654648307
transform 1 0 35600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6268
timestamp 1654648307
transform 1 0 40100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6267
timestamp 1654648307
transform 1 0 38600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6188
timestamp 1654648307
transform 1 0 40100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6187
timestamp 1654648307
transform 1 0 38600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6270
timestamp 1654648307
transform 1 0 43100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6269
timestamp 1654648307
transform 1 0 41600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6190
timestamp 1654648307
transform 1 0 43100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6189
timestamp 1654648307
transform 1 0 41600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6272
timestamp 1654648307
transform 1 0 46100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6271
timestamp 1654648307
transform 1 0 44600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6192
timestamp 1654648307
transform 1 0 46100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6191
timestamp 1654648307
transform 1 0 44600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6274
timestamp 1654648307
transform 1 0 49100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6273
timestamp 1654648307
transform 1 0 47600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6194
timestamp 1654648307
transform 1 0 49100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6193
timestamp 1654648307
transform 1 0 47600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6276
timestamp 1654648307
transform 1 0 52100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6275
timestamp 1654648307
transform 1 0 50600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6196
timestamp 1654648307
transform 1 0 52100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6195
timestamp 1654648307
transform 1 0 50600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6278
timestamp 1654648307
transform 1 0 55100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6277
timestamp 1654648307
transform 1 0 53600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6198
timestamp 1654648307
transform 1 0 55100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6197
timestamp 1654648307
transform 1 0 53600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6280
timestamp 1654648307
transform 1 0 58100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6279
timestamp 1654648307
transform 1 0 56600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6200
timestamp 1654648307
transform 1 0 58100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6199
timestamp 1654648307
transform 1 0 56600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6282
timestamp 1654648307
transform 1 0 61100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6281
timestamp 1654648307
transform 1 0 59600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6202
timestamp 1654648307
transform 1 0 61100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6201
timestamp 1654648307
transform 1 0 59600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6284
timestamp 1654648307
transform 1 0 64100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6283
timestamp 1654648307
transform 1 0 62600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6204
timestamp 1654648307
transform 1 0 64100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6203
timestamp 1654648307
transform 1 0 62600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6286
timestamp 1654648307
transform 1 0 67100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6285
timestamp 1654648307
transform 1 0 65600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6206
timestamp 1654648307
transform 1 0 67100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6205
timestamp 1654648307
transform 1 0 65600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6288
timestamp 1654648307
transform 1 0 70100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6287
timestamp 1654648307
transform 1 0 68600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6208
timestamp 1654648307
transform 1 0 70100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6207
timestamp 1654648307
transform 1 0 68600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6290
timestamp 1654648307
transform 1 0 73100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6289
timestamp 1654648307
transform 1 0 71600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6210
timestamp 1654648307
transform 1 0 73100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6209
timestamp 1654648307
transform 1 0 71600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6292
timestamp 1654648307
transform 1 0 76100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6291
timestamp 1654648307
transform 1 0 74600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6212
timestamp 1654648307
transform 1 0 76100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6211
timestamp 1654648307
transform 1 0 74600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6294
timestamp 1654648307
transform 1 0 79100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6293
timestamp 1654648307
transform 1 0 77600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6214
timestamp 1654648307
transform 1 0 79100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6213
timestamp 1654648307
transform 1 0 77600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6296
timestamp 1654648307
transform 1 0 82100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6295
timestamp 1654648307
transform 1 0 80600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6216
timestamp 1654648307
transform 1 0 82100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6215
timestamp 1654648307
transform 1 0 80600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6298
timestamp 1654648307
transform 1 0 85100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6297
timestamp 1654648307
transform 1 0 83600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6218
timestamp 1654648307
transform 1 0 85100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6217
timestamp 1654648307
transform 1 0 83600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6300
timestamp 1654648307
transform 1 0 88100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6299
timestamp 1654648307
transform 1 0 86600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6220
timestamp 1654648307
transform 1 0 88100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6219
timestamp 1654648307
transform 1 0 86600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6302
timestamp 1654648307
transform 1 0 91100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6301
timestamp 1654648307
transform 1 0 89600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6222
timestamp 1654648307
transform 1 0 91100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6221
timestamp 1654648307
transform 1 0 89600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6304
timestamp 1654648307
transform 1 0 94100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6303
timestamp 1654648307
transform 1 0 92600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6224
timestamp 1654648307
transform 1 0 94100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6223
timestamp 1654648307
transform 1 0 92600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6306
timestamp 1654648307
transform 1 0 97100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6305
timestamp 1654648307
transform 1 0 95600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6226
timestamp 1654648307
transform 1 0 97100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6225
timestamp 1654648307
transform 1 0 95600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6308
timestamp 1654648307
transform 1 0 100100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6307
timestamp 1654648307
transform 1 0 98600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6228
timestamp 1654648307
transform 1 0 100100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6227
timestamp 1654648307
transform 1 0 98600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6310
timestamp 1654648307
transform 1 0 103100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6309
timestamp 1654648307
transform 1 0 101600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6230
timestamp 1654648307
transform 1 0 103100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6229
timestamp 1654648307
transform 1 0 101600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6312
timestamp 1654648307
transform 1 0 106100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6311
timestamp 1654648307
transform 1 0 104600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6232
timestamp 1654648307
transform 1 0 106100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6231
timestamp 1654648307
transform 1 0 104600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6314
timestamp 1654648307
transform 1 0 109100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6313
timestamp 1654648307
transform 1 0 107600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6234
timestamp 1654648307
transform 1 0 109100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6233
timestamp 1654648307
transform 1 0 107600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6316
timestamp 1654648307
transform 1 0 112100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6315
timestamp 1654648307
transform 1 0 110600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6236
timestamp 1654648307
transform 1 0 112100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6235
timestamp 1654648307
transform 1 0 110600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6318
timestamp 1654648307
transform 1 0 115100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6317
timestamp 1654648307
transform 1 0 113600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6238
timestamp 1654648307
transform 1 0 115100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6237
timestamp 1654648307
transform 1 0 113600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6319
timestamp 1654648307
transform 1 0 116600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_6239
timestamp 1654648307
transform 1 0 116600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_6080
timestamp 1654648307
transform 1 0 -1900 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6000
timestamp 1654648307
transform 1 0 -1900 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6082
timestamp 1654648307
transform 1 0 1100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6081
timestamp 1654648307
transform 1 0 -400 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6002
timestamp 1654648307
transform 1 0 1100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6001
timestamp 1654648307
transform 1 0 -400 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6084
timestamp 1654648307
transform 1 0 4100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6083
timestamp 1654648307
transform 1 0 2600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6004
timestamp 1654648307
transform 1 0 4100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6003
timestamp 1654648307
transform 1 0 2600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6086
timestamp 1654648307
transform 1 0 7100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6085
timestamp 1654648307
transform 1 0 5600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6006
timestamp 1654648307
transform 1 0 7100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6005
timestamp 1654648307
transform 1 0 5600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6088
timestamp 1654648307
transform 1 0 10100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6087
timestamp 1654648307
transform 1 0 8600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6008
timestamp 1654648307
transform 1 0 10100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6007
timestamp 1654648307
transform 1 0 8600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6090
timestamp 1654648307
transform 1 0 13100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6089
timestamp 1654648307
transform 1 0 11600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6010
timestamp 1654648307
transform 1 0 13100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6009
timestamp 1654648307
transform 1 0 11600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6092
timestamp 1654648307
transform 1 0 16100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6091
timestamp 1654648307
transform 1 0 14600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6012
timestamp 1654648307
transform 1 0 16100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6011
timestamp 1654648307
transform 1 0 14600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6094
timestamp 1654648307
transform 1 0 19100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6093
timestamp 1654648307
transform 1 0 17600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6014
timestamp 1654648307
transform 1 0 19100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6013
timestamp 1654648307
transform 1 0 17600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6096
timestamp 1654648307
transform 1 0 22100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6095
timestamp 1654648307
transform 1 0 20600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6016
timestamp 1654648307
transform 1 0 22100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6015
timestamp 1654648307
transform 1 0 20600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6098
timestamp 1654648307
transform 1 0 25100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6097
timestamp 1654648307
transform 1 0 23600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6018
timestamp 1654648307
transform 1 0 25100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6017
timestamp 1654648307
transform 1 0 23600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6100
timestamp 1654648307
transform 1 0 28100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6099
timestamp 1654648307
transform 1 0 26600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6020
timestamp 1654648307
transform 1 0 28100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6019
timestamp 1654648307
transform 1 0 26600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6102
timestamp 1654648307
transform 1 0 31100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6101
timestamp 1654648307
transform 1 0 29600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6022
timestamp 1654648307
transform 1 0 31100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6021
timestamp 1654648307
transform 1 0 29600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6104
timestamp 1654648307
transform 1 0 34100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6103
timestamp 1654648307
transform 1 0 32600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6024
timestamp 1654648307
transform 1 0 34100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6023
timestamp 1654648307
transform 1 0 32600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6106
timestamp 1654648307
transform 1 0 37100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6105
timestamp 1654648307
transform 1 0 35600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6026
timestamp 1654648307
transform 1 0 37100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6025
timestamp 1654648307
transform 1 0 35600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6108
timestamp 1654648307
transform 1 0 40100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6107
timestamp 1654648307
transform 1 0 38600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6028
timestamp 1654648307
transform 1 0 40100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6027
timestamp 1654648307
transform 1 0 38600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6110
timestamp 1654648307
transform 1 0 43100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6109
timestamp 1654648307
transform 1 0 41600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6030
timestamp 1654648307
transform 1 0 43100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6029
timestamp 1654648307
transform 1 0 41600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6112
timestamp 1654648307
transform 1 0 46100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6111
timestamp 1654648307
transform 1 0 44600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6032
timestamp 1654648307
transform 1 0 46100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6031
timestamp 1654648307
transform 1 0 44600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6114
timestamp 1654648307
transform 1 0 49100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6113
timestamp 1654648307
transform 1 0 47600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6034
timestamp 1654648307
transform 1 0 49100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6033
timestamp 1654648307
transform 1 0 47600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6116
timestamp 1654648307
transform 1 0 52100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6115
timestamp 1654648307
transform 1 0 50600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6036
timestamp 1654648307
transform 1 0 52100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6035
timestamp 1654648307
transform 1 0 50600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6118
timestamp 1654648307
transform 1 0 55100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6117
timestamp 1654648307
transform 1 0 53600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6038
timestamp 1654648307
transform 1 0 55100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6037
timestamp 1654648307
transform 1 0 53600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6120
timestamp 1654648307
transform 1 0 58100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6119
timestamp 1654648307
transform 1 0 56600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6040
timestamp 1654648307
transform 1 0 58100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6039
timestamp 1654648307
transform 1 0 56600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6122
timestamp 1654648307
transform 1 0 61100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6121
timestamp 1654648307
transform 1 0 59600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6042
timestamp 1654648307
transform 1 0 61100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6041
timestamp 1654648307
transform 1 0 59600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6124
timestamp 1654648307
transform 1 0 64100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6123
timestamp 1654648307
transform 1 0 62600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6044
timestamp 1654648307
transform 1 0 64100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6043
timestamp 1654648307
transform 1 0 62600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6126
timestamp 1654648307
transform 1 0 67100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6125
timestamp 1654648307
transform 1 0 65600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6046
timestamp 1654648307
transform 1 0 67100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6045
timestamp 1654648307
transform 1 0 65600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6128
timestamp 1654648307
transform 1 0 70100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6127
timestamp 1654648307
transform 1 0 68600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6048
timestamp 1654648307
transform 1 0 70100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6047
timestamp 1654648307
transform 1 0 68600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6130
timestamp 1654648307
transform 1 0 73100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6129
timestamp 1654648307
transform 1 0 71600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6050
timestamp 1654648307
transform 1 0 73100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6049
timestamp 1654648307
transform 1 0 71600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6132
timestamp 1654648307
transform 1 0 76100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6131
timestamp 1654648307
transform 1 0 74600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6052
timestamp 1654648307
transform 1 0 76100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6051
timestamp 1654648307
transform 1 0 74600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6134
timestamp 1654648307
transform 1 0 79100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6133
timestamp 1654648307
transform 1 0 77600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6054
timestamp 1654648307
transform 1 0 79100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6053
timestamp 1654648307
transform 1 0 77600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6136
timestamp 1654648307
transform 1 0 82100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6135
timestamp 1654648307
transform 1 0 80600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6056
timestamp 1654648307
transform 1 0 82100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6055
timestamp 1654648307
transform 1 0 80600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6138
timestamp 1654648307
transform 1 0 85100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6137
timestamp 1654648307
transform 1 0 83600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6058
timestamp 1654648307
transform 1 0 85100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6057
timestamp 1654648307
transform 1 0 83600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6140
timestamp 1654648307
transform 1 0 88100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6139
timestamp 1654648307
transform 1 0 86600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6060
timestamp 1654648307
transform 1 0 88100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6059
timestamp 1654648307
transform 1 0 86600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6142
timestamp 1654648307
transform 1 0 91100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6141
timestamp 1654648307
transform 1 0 89600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6062
timestamp 1654648307
transform 1 0 91100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6061
timestamp 1654648307
transform 1 0 89600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6144
timestamp 1654648307
transform 1 0 94100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6143
timestamp 1654648307
transform 1 0 92600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6064
timestamp 1654648307
transform 1 0 94100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6063
timestamp 1654648307
transform 1 0 92600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6146
timestamp 1654648307
transform 1 0 97100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6145
timestamp 1654648307
transform 1 0 95600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6066
timestamp 1654648307
transform 1 0 97100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6065
timestamp 1654648307
transform 1 0 95600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6148
timestamp 1654648307
transform 1 0 100100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6147
timestamp 1654648307
transform 1 0 98600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6068
timestamp 1654648307
transform 1 0 100100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6067
timestamp 1654648307
transform 1 0 98600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6150
timestamp 1654648307
transform 1 0 103100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6149
timestamp 1654648307
transform 1 0 101600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6070
timestamp 1654648307
transform 1 0 103100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6069
timestamp 1654648307
transform 1 0 101600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6152
timestamp 1654648307
transform 1 0 106100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6151
timestamp 1654648307
transform 1 0 104600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6072
timestamp 1654648307
transform 1 0 106100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6071
timestamp 1654648307
transform 1 0 104600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6154
timestamp 1654648307
transform 1 0 109100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6153
timestamp 1654648307
transform 1 0 107600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6074
timestamp 1654648307
transform 1 0 109100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6073
timestamp 1654648307
transform 1 0 107600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6156
timestamp 1654648307
transform 1 0 112100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6155
timestamp 1654648307
transform 1 0 110600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6076
timestamp 1654648307
transform 1 0 112100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6075
timestamp 1654648307
transform 1 0 110600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6158
timestamp 1654648307
transform 1 0 115100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6157
timestamp 1654648307
transform 1 0 113600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6078
timestamp 1654648307
transform 1 0 115100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6077
timestamp 1654648307
transform 1 0 113600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_6159
timestamp 1654648307
transform 1 0 116600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_6079
timestamp 1654648307
transform 1 0 116600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_5920
timestamp 1654648307
transform 1 0 -1900 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5840
timestamp 1654648307
transform 1 0 -1900 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5922
timestamp 1654648307
transform 1 0 1100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5921
timestamp 1654648307
transform 1 0 -400 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5842
timestamp 1654648307
transform 1 0 1100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5841
timestamp 1654648307
transform 1 0 -400 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5924
timestamp 1654648307
transform 1 0 4100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5923
timestamp 1654648307
transform 1 0 2600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5844
timestamp 1654648307
transform 1 0 4100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5843
timestamp 1654648307
transform 1 0 2600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5926
timestamp 1654648307
transform 1 0 7100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5925
timestamp 1654648307
transform 1 0 5600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5846
timestamp 1654648307
transform 1 0 7100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5845
timestamp 1654648307
transform 1 0 5600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5928
timestamp 1654648307
transform 1 0 10100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5927
timestamp 1654648307
transform 1 0 8600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5848
timestamp 1654648307
transform 1 0 10100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5847
timestamp 1654648307
transform 1 0 8600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5930
timestamp 1654648307
transform 1 0 13100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5929
timestamp 1654648307
transform 1 0 11600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5850
timestamp 1654648307
transform 1 0 13100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5849
timestamp 1654648307
transform 1 0 11600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5932
timestamp 1654648307
transform 1 0 16100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5931
timestamp 1654648307
transform 1 0 14600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5852
timestamp 1654648307
transform 1 0 16100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5851
timestamp 1654648307
transform 1 0 14600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5934
timestamp 1654648307
transform 1 0 19100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5933
timestamp 1654648307
transform 1 0 17600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5854
timestamp 1654648307
transform 1 0 19100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5853
timestamp 1654648307
transform 1 0 17600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5936
timestamp 1654648307
transform 1 0 22100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5935
timestamp 1654648307
transform 1 0 20600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5856
timestamp 1654648307
transform 1 0 22100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5855
timestamp 1654648307
transform 1 0 20600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5938
timestamp 1654648307
transform 1 0 25100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5937
timestamp 1654648307
transform 1 0 23600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5858
timestamp 1654648307
transform 1 0 25100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5857
timestamp 1654648307
transform 1 0 23600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5940
timestamp 1654648307
transform 1 0 28100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5939
timestamp 1654648307
transform 1 0 26600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5860
timestamp 1654648307
transform 1 0 28100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5859
timestamp 1654648307
transform 1 0 26600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5942
timestamp 1654648307
transform 1 0 31100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5941
timestamp 1654648307
transform 1 0 29600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5862
timestamp 1654648307
transform 1 0 31100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5861
timestamp 1654648307
transform 1 0 29600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5944
timestamp 1654648307
transform 1 0 34100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5943
timestamp 1654648307
transform 1 0 32600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5864
timestamp 1654648307
transform 1 0 34100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5863
timestamp 1654648307
transform 1 0 32600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5946
timestamp 1654648307
transform 1 0 37100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5945
timestamp 1654648307
transform 1 0 35600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5866
timestamp 1654648307
transform 1 0 37100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5865
timestamp 1654648307
transform 1 0 35600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5948
timestamp 1654648307
transform 1 0 40100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5947
timestamp 1654648307
transform 1 0 38600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5868
timestamp 1654648307
transform 1 0 40100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5867
timestamp 1654648307
transform 1 0 38600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5950
timestamp 1654648307
transform 1 0 43100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5949
timestamp 1654648307
transform 1 0 41600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5870
timestamp 1654648307
transform 1 0 43100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5869
timestamp 1654648307
transform 1 0 41600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5952
timestamp 1654648307
transform 1 0 46100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5951
timestamp 1654648307
transform 1 0 44600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5872
timestamp 1654648307
transform 1 0 46100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5871
timestamp 1654648307
transform 1 0 44600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5954
timestamp 1654648307
transform 1 0 49100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5953
timestamp 1654648307
transform 1 0 47600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5874
timestamp 1654648307
transform 1 0 49100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5873
timestamp 1654648307
transform 1 0 47600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5956
timestamp 1654648307
transform 1 0 52100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5955
timestamp 1654648307
transform 1 0 50600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5876
timestamp 1654648307
transform 1 0 52100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5875
timestamp 1654648307
transform 1 0 50600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5958
timestamp 1654648307
transform 1 0 55100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5957
timestamp 1654648307
transform 1 0 53600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5878
timestamp 1654648307
transform 1 0 55100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5877
timestamp 1654648307
transform 1 0 53600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5960
timestamp 1654648307
transform 1 0 58100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5959
timestamp 1654648307
transform 1 0 56600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5880
timestamp 1654648307
transform 1 0 58100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5879
timestamp 1654648307
transform 1 0 56600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5962
timestamp 1654648307
transform 1 0 61100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5961
timestamp 1654648307
transform 1 0 59600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5882
timestamp 1654648307
transform 1 0 61100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5881
timestamp 1654648307
transform 1 0 59600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5964
timestamp 1654648307
transform 1 0 64100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5963
timestamp 1654648307
transform 1 0 62600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5884
timestamp 1654648307
transform 1 0 64100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5883
timestamp 1654648307
transform 1 0 62600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5966
timestamp 1654648307
transform 1 0 67100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5965
timestamp 1654648307
transform 1 0 65600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5886
timestamp 1654648307
transform 1 0 67100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5885
timestamp 1654648307
transform 1 0 65600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5968
timestamp 1654648307
transform 1 0 70100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5967
timestamp 1654648307
transform 1 0 68600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5888
timestamp 1654648307
transform 1 0 70100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5887
timestamp 1654648307
transform 1 0 68600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5970
timestamp 1654648307
transform 1 0 73100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5969
timestamp 1654648307
transform 1 0 71600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5890
timestamp 1654648307
transform 1 0 73100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5889
timestamp 1654648307
transform 1 0 71600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5972
timestamp 1654648307
transform 1 0 76100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5971
timestamp 1654648307
transform 1 0 74600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5892
timestamp 1654648307
transform 1 0 76100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5891
timestamp 1654648307
transform 1 0 74600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5974
timestamp 1654648307
transform 1 0 79100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5973
timestamp 1654648307
transform 1 0 77600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5894
timestamp 1654648307
transform 1 0 79100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5893
timestamp 1654648307
transform 1 0 77600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5976
timestamp 1654648307
transform 1 0 82100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5975
timestamp 1654648307
transform 1 0 80600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5896
timestamp 1654648307
transform 1 0 82100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5895
timestamp 1654648307
transform 1 0 80600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5978
timestamp 1654648307
transform 1 0 85100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5977
timestamp 1654648307
transform 1 0 83600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5898
timestamp 1654648307
transform 1 0 85100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5897
timestamp 1654648307
transform 1 0 83600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5980
timestamp 1654648307
transform 1 0 88100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5979
timestamp 1654648307
transform 1 0 86600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5900
timestamp 1654648307
transform 1 0 88100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5899
timestamp 1654648307
transform 1 0 86600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5982
timestamp 1654648307
transform 1 0 91100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5981
timestamp 1654648307
transform 1 0 89600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5902
timestamp 1654648307
transform 1 0 91100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5901
timestamp 1654648307
transform 1 0 89600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5984
timestamp 1654648307
transform 1 0 94100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5983
timestamp 1654648307
transform 1 0 92600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5904
timestamp 1654648307
transform 1 0 94100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5903
timestamp 1654648307
transform 1 0 92600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5986
timestamp 1654648307
transform 1 0 97100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5985
timestamp 1654648307
transform 1 0 95600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5906
timestamp 1654648307
transform 1 0 97100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5905
timestamp 1654648307
transform 1 0 95600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5988
timestamp 1654648307
transform 1 0 100100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5987
timestamp 1654648307
transform 1 0 98600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5908
timestamp 1654648307
transform 1 0 100100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5907
timestamp 1654648307
transform 1 0 98600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5990
timestamp 1654648307
transform 1 0 103100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5989
timestamp 1654648307
transform 1 0 101600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5910
timestamp 1654648307
transform 1 0 103100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5909
timestamp 1654648307
transform 1 0 101600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5992
timestamp 1654648307
transform 1 0 106100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5991
timestamp 1654648307
transform 1 0 104600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5912
timestamp 1654648307
transform 1 0 106100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5911
timestamp 1654648307
transform 1 0 104600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5994
timestamp 1654648307
transform 1 0 109100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5993
timestamp 1654648307
transform 1 0 107600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5914
timestamp 1654648307
transform 1 0 109100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5913
timestamp 1654648307
transform 1 0 107600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5996
timestamp 1654648307
transform 1 0 112100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5995
timestamp 1654648307
transform 1 0 110600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5916
timestamp 1654648307
transform 1 0 112100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5915
timestamp 1654648307
transform 1 0 110600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5998
timestamp 1654648307
transform 1 0 115100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5997
timestamp 1654648307
transform 1 0 113600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5918
timestamp 1654648307
transform 1 0 115100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5917
timestamp 1654648307
transform 1 0 113600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5999
timestamp 1654648307
transform 1 0 116600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_5919
timestamp 1654648307
transform 1 0 116600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_5760
timestamp 1654648307
transform 1 0 -1900 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5680
timestamp 1654648307
transform 1 0 -1900 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5762
timestamp 1654648307
transform 1 0 1100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5761
timestamp 1654648307
transform 1 0 -400 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5682
timestamp 1654648307
transform 1 0 1100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5681
timestamp 1654648307
transform 1 0 -400 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5764
timestamp 1654648307
transform 1 0 4100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5763
timestamp 1654648307
transform 1 0 2600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5684
timestamp 1654648307
transform 1 0 4100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5683
timestamp 1654648307
transform 1 0 2600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5766
timestamp 1654648307
transform 1 0 7100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5765
timestamp 1654648307
transform 1 0 5600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5686
timestamp 1654648307
transform 1 0 7100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5685
timestamp 1654648307
transform 1 0 5600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5768
timestamp 1654648307
transform 1 0 10100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5767
timestamp 1654648307
transform 1 0 8600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5688
timestamp 1654648307
transform 1 0 10100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5687
timestamp 1654648307
transform 1 0 8600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5770
timestamp 1654648307
transform 1 0 13100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5769
timestamp 1654648307
transform 1 0 11600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5690
timestamp 1654648307
transform 1 0 13100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5689
timestamp 1654648307
transform 1 0 11600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5772
timestamp 1654648307
transform 1 0 16100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5771
timestamp 1654648307
transform 1 0 14600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5692
timestamp 1654648307
transform 1 0 16100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5691
timestamp 1654648307
transform 1 0 14600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5774
timestamp 1654648307
transform 1 0 19100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5773
timestamp 1654648307
transform 1 0 17600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5694
timestamp 1654648307
transform 1 0 19100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5693
timestamp 1654648307
transform 1 0 17600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5776
timestamp 1654648307
transform 1 0 22100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5775
timestamp 1654648307
transform 1 0 20600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5696
timestamp 1654648307
transform 1 0 22100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5695
timestamp 1654648307
transform 1 0 20600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5778
timestamp 1654648307
transform 1 0 25100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5777
timestamp 1654648307
transform 1 0 23600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5698
timestamp 1654648307
transform 1 0 25100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5697
timestamp 1654648307
transform 1 0 23600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5780
timestamp 1654648307
transform 1 0 28100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5779
timestamp 1654648307
transform 1 0 26600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5700
timestamp 1654648307
transform 1 0 28100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5699
timestamp 1654648307
transform 1 0 26600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5782
timestamp 1654648307
transform 1 0 31100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5781
timestamp 1654648307
transform 1 0 29600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5702
timestamp 1654648307
transform 1 0 31100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5701
timestamp 1654648307
transform 1 0 29600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5784
timestamp 1654648307
transform 1 0 34100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5783
timestamp 1654648307
transform 1 0 32600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5704
timestamp 1654648307
transform 1 0 34100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5703
timestamp 1654648307
transform 1 0 32600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5786
timestamp 1654648307
transform 1 0 37100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5785
timestamp 1654648307
transform 1 0 35600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5706
timestamp 1654648307
transform 1 0 37100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5705
timestamp 1654648307
transform 1 0 35600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5788
timestamp 1654648307
transform 1 0 40100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5787
timestamp 1654648307
transform 1 0 38600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5708
timestamp 1654648307
transform 1 0 40100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5707
timestamp 1654648307
transform 1 0 38600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5790
timestamp 1654648307
transform 1 0 43100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5789
timestamp 1654648307
transform 1 0 41600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5710
timestamp 1654648307
transform 1 0 43100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5709
timestamp 1654648307
transform 1 0 41600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5792
timestamp 1654648307
transform 1 0 46100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5791
timestamp 1654648307
transform 1 0 44600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5712
timestamp 1654648307
transform 1 0 46100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5711
timestamp 1654648307
transform 1 0 44600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5794
timestamp 1654648307
transform 1 0 49100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5793
timestamp 1654648307
transform 1 0 47600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5714
timestamp 1654648307
transform 1 0 49100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5713
timestamp 1654648307
transform 1 0 47600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5796
timestamp 1654648307
transform 1 0 52100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5795
timestamp 1654648307
transform 1 0 50600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5716
timestamp 1654648307
transform 1 0 52100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5715
timestamp 1654648307
transform 1 0 50600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5798
timestamp 1654648307
transform 1 0 55100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5797
timestamp 1654648307
transform 1 0 53600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5718
timestamp 1654648307
transform 1 0 55100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5717
timestamp 1654648307
transform 1 0 53600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5800
timestamp 1654648307
transform 1 0 58100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5799
timestamp 1654648307
transform 1 0 56600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5720
timestamp 1654648307
transform 1 0 58100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5719
timestamp 1654648307
transform 1 0 56600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5802
timestamp 1654648307
transform 1 0 61100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5801
timestamp 1654648307
transform 1 0 59600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5722
timestamp 1654648307
transform 1 0 61100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5721
timestamp 1654648307
transform 1 0 59600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5804
timestamp 1654648307
transform 1 0 64100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5803
timestamp 1654648307
transform 1 0 62600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5724
timestamp 1654648307
transform 1 0 64100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5723
timestamp 1654648307
transform 1 0 62600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5806
timestamp 1654648307
transform 1 0 67100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5805
timestamp 1654648307
transform 1 0 65600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5726
timestamp 1654648307
transform 1 0 67100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5725
timestamp 1654648307
transform 1 0 65600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5808
timestamp 1654648307
transform 1 0 70100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5807
timestamp 1654648307
transform 1 0 68600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5728
timestamp 1654648307
transform 1 0 70100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5727
timestamp 1654648307
transform 1 0 68600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5810
timestamp 1654648307
transform 1 0 73100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5809
timestamp 1654648307
transform 1 0 71600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5730
timestamp 1654648307
transform 1 0 73100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5729
timestamp 1654648307
transform 1 0 71600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5812
timestamp 1654648307
transform 1 0 76100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5811
timestamp 1654648307
transform 1 0 74600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5732
timestamp 1654648307
transform 1 0 76100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5731
timestamp 1654648307
transform 1 0 74600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5814
timestamp 1654648307
transform 1 0 79100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5813
timestamp 1654648307
transform 1 0 77600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5734
timestamp 1654648307
transform 1 0 79100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5733
timestamp 1654648307
transform 1 0 77600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5816
timestamp 1654648307
transform 1 0 82100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5815
timestamp 1654648307
transform 1 0 80600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5736
timestamp 1654648307
transform 1 0 82100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5735
timestamp 1654648307
transform 1 0 80600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5818
timestamp 1654648307
transform 1 0 85100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5817
timestamp 1654648307
transform 1 0 83600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5738
timestamp 1654648307
transform 1 0 85100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5737
timestamp 1654648307
transform 1 0 83600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5820
timestamp 1654648307
transform 1 0 88100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5819
timestamp 1654648307
transform 1 0 86600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5740
timestamp 1654648307
transform 1 0 88100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5739
timestamp 1654648307
transform 1 0 86600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5822
timestamp 1654648307
transform 1 0 91100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5821
timestamp 1654648307
transform 1 0 89600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5742
timestamp 1654648307
transform 1 0 91100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5741
timestamp 1654648307
transform 1 0 89600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5824
timestamp 1654648307
transform 1 0 94100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5823
timestamp 1654648307
transform 1 0 92600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5744
timestamp 1654648307
transform 1 0 94100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5743
timestamp 1654648307
transform 1 0 92600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5826
timestamp 1654648307
transform 1 0 97100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5825
timestamp 1654648307
transform 1 0 95600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5746
timestamp 1654648307
transform 1 0 97100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5745
timestamp 1654648307
transform 1 0 95600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5828
timestamp 1654648307
transform 1 0 100100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5827
timestamp 1654648307
transform 1 0 98600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5748
timestamp 1654648307
transform 1 0 100100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5747
timestamp 1654648307
transform 1 0 98600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5830
timestamp 1654648307
transform 1 0 103100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5829
timestamp 1654648307
transform 1 0 101600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5750
timestamp 1654648307
transform 1 0 103100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5749
timestamp 1654648307
transform 1 0 101600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5832
timestamp 1654648307
transform 1 0 106100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5831
timestamp 1654648307
transform 1 0 104600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5752
timestamp 1654648307
transform 1 0 106100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5751
timestamp 1654648307
transform 1 0 104600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5834
timestamp 1654648307
transform 1 0 109100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5833
timestamp 1654648307
transform 1 0 107600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5754
timestamp 1654648307
transform 1 0 109100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5753
timestamp 1654648307
transform 1 0 107600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5836
timestamp 1654648307
transform 1 0 112100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5835
timestamp 1654648307
transform 1 0 110600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5756
timestamp 1654648307
transform 1 0 112100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5755
timestamp 1654648307
transform 1 0 110600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5838
timestamp 1654648307
transform 1 0 115100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5837
timestamp 1654648307
transform 1 0 113600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5758
timestamp 1654648307
transform 1 0 115100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5757
timestamp 1654648307
transform 1 0 113600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5839
timestamp 1654648307
transform 1 0 116600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_5759
timestamp 1654648307
transform 1 0 116600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_5600
timestamp 1654648307
transform 1 0 -1900 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5520
timestamp 1654648307
transform 1 0 -1900 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5602
timestamp 1654648307
transform 1 0 1100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5601
timestamp 1654648307
transform 1 0 -400 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5522
timestamp 1654648307
transform 1 0 1100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5521
timestamp 1654648307
transform 1 0 -400 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5604
timestamp 1654648307
transform 1 0 4100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5603
timestamp 1654648307
transform 1 0 2600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5524
timestamp 1654648307
transform 1 0 4100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5523
timestamp 1654648307
transform 1 0 2600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5606
timestamp 1654648307
transform 1 0 7100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5605
timestamp 1654648307
transform 1 0 5600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5526
timestamp 1654648307
transform 1 0 7100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5525
timestamp 1654648307
transform 1 0 5600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5608
timestamp 1654648307
transform 1 0 10100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5607
timestamp 1654648307
transform 1 0 8600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5528
timestamp 1654648307
transform 1 0 10100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5527
timestamp 1654648307
transform 1 0 8600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5610
timestamp 1654648307
transform 1 0 13100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5609
timestamp 1654648307
transform 1 0 11600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5530
timestamp 1654648307
transform 1 0 13100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5529
timestamp 1654648307
transform 1 0 11600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5612
timestamp 1654648307
transform 1 0 16100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5611
timestamp 1654648307
transform 1 0 14600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5532
timestamp 1654648307
transform 1 0 16100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5531
timestamp 1654648307
transform 1 0 14600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5614
timestamp 1654648307
transform 1 0 19100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5613
timestamp 1654648307
transform 1 0 17600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5534
timestamp 1654648307
transform 1 0 19100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5533
timestamp 1654648307
transform 1 0 17600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5616
timestamp 1654648307
transform 1 0 22100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5615
timestamp 1654648307
transform 1 0 20600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5536
timestamp 1654648307
transform 1 0 22100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5535
timestamp 1654648307
transform 1 0 20600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5618
timestamp 1654648307
transform 1 0 25100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5617
timestamp 1654648307
transform 1 0 23600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5538
timestamp 1654648307
transform 1 0 25100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5537
timestamp 1654648307
transform 1 0 23600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5620
timestamp 1654648307
transform 1 0 28100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5619
timestamp 1654648307
transform 1 0 26600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5540
timestamp 1654648307
transform 1 0 28100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5539
timestamp 1654648307
transform 1 0 26600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5622
timestamp 1654648307
transform 1 0 31100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5621
timestamp 1654648307
transform 1 0 29600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5542
timestamp 1654648307
transform 1 0 31100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5541
timestamp 1654648307
transform 1 0 29600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5624
timestamp 1654648307
transform 1 0 34100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5623
timestamp 1654648307
transform 1 0 32600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5544
timestamp 1654648307
transform 1 0 34100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5543
timestamp 1654648307
transform 1 0 32600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5626
timestamp 1654648307
transform 1 0 37100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5625
timestamp 1654648307
transform 1 0 35600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5546
timestamp 1654648307
transform 1 0 37100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5545
timestamp 1654648307
transform 1 0 35600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5628
timestamp 1654648307
transform 1 0 40100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5627
timestamp 1654648307
transform 1 0 38600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5548
timestamp 1654648307
transform 1 0 40100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5547
timestamp 1654648307
transform 1 0 38600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5630
timestamp 1654648307
transform 1 0 43100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5629
timestamp 1654648307
transform 1 0 41600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5550
timestamp 1654648307
transform 1 0 43100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5549
timestamp 1654648307
transform 1 0 41600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5632
timestamp 1654648307
transform 1 0 46100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5631
timestamp 1654648307
transform 1 0 44600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5552
timestamp 1654648307
transform 1 0 46100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5551
timestamp 1654648307
transform 1 0 44600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5634
timestamp 1654648307
transform 1 0 49100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5633
timestamp 1654648307
transform 1 0 47600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5554
timestamp 1654648307
transform 1 0 49100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5553
timestamp 1654648307
transform 1 0 47600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5636
timestamp 1654648307
transform 1 0 52100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5635
timestamp 1654648307
transform 1 0 50600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5556
timestamp 1654648307
transform 1 0 52100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5555
timestamp 1654648307
transform 1 0 50600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5638
timestamp 1654648307
transform 1 0 55100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5637
timestamp 1654648307
transform 1 0 53600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5558
timestamp 1654648307
transform 1 0 55100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5557
timestamp 1654648307
transform 1 0 53600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5640
timestamp 1654648307
transform 1 0 58100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5639
timestamp 1654648307
transform 1 0 56600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5560
timestamp 1654648307
transform 1 0 58100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5559
timestamp 1654648307
transform 1 0 56600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5642
timestamp 1654648307
transform 1 0 61100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5641
timestamp 1654648307
transform 1 0 59600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5562
timestamp 1654648307
transform 1 0 61100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5561
timestamp 1654648307
transform 1 0 59600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5644
timestamp 1654648307
transform 1 0 64100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5643
timestamp 1654648307
transform 1 0 62600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5564
timestamp 1654648307
transform 1 0 64100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5563
timestamp 1654648307
transform 1 0 62600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5646
timestamp 1654648307
transform 1 0 67100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5645
timestamp 1654648307
transform 1 0 65600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5566
timestamp 1654648307
transform 1 0 67100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5565
timestamp 1654648307
transform 1 0 65600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5648
timestamp 1654648307
transform 1 0 70100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5647
timestamp 1654648307
transform 1 0 68600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5568
timestamp 1654648307
transform 1 0 70100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5567
timestamp 1654648307
transform 1 0 68600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5650
timestamp 1654648307
transform 1 0 73100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5649
timestamp 1654648307
transform 1 0 71600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5570
timestamp 1654648307
transform 1 0 73100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5569
timestamp 1654648307
transform 1 0 71600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5652
timestamp 1654648307
transform 1 0 76100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5651
timestamp 1654648307
transform 1 0 74600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5572
timestamp 1654648307
transform 1 0 76100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5571
timestamp 1654648307
transform 1 0 74600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5654
timestamp 1654648307
transform 1 0 79100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5653
timestamp 1654648307
transform 1 0 77600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5574
timestamp 1654648307
transform 1 0 79100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5573
timestamp 1654648307
transform 1 0 77600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5656
timestamp 1654648307
transform 1 0 82100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5655
timestamp 1654648307
transform 1 0 80600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5576
timestamp 1654648307
transform 1 0 82100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5575
timestamp 1654648307
transform 1 0 80600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5658
timestamp 1654648307
transform 1 0 85100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5657
timestamp 1654648307
transform 1 0 83600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5578
timestamp 1654648307
transform 1 0 85100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5577
timestamp 1654648307
transform 1 0 83600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5660
timestamp 1654648307
transform 1 0 88100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5659
timestamp 1654648307
transform 1 0 86600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5580
timestamp 1654648307
transform 1 0 88100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5579
timestamp 1654648307
transform 1 0 86600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5662
timestamp 1654648307
transform 1 0 91100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5661
timestamp 1654648307
transform 1 0 89600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5582
timestamp 1654648307
transform 1 0 91100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5581
timestamp 1654648307
transform 1 0 89600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5664
timestamp 1654648307
transform 1 0 94100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5663
timestamp 1654648307
transform 1 0 92600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5584
timestamp 1654648307
transform 1 0 94100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5583
timestamp 1654648307
transform 1 0 92600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5666
timestamp 1654648307
transform 1 0 97100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5665
timestamp 1654648307
transform 1 0 95600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5586
timestamp 1654648307
transform 1 0 97100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5585
timestamp 1654648307
transform 1 0 95600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5668
timestamp 1654648307
transform 1 0 100100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5667
timestamp 1654648307
transform 1 0 98600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5588
timestamp 1654648307
transform 1 0 100100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5587
timestamp 1654648307
transform 1 0 98600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5670
timestamp 1654648307
transform 1 0 103100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5669
timestamp 1654648307
transform 1 0 101600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5590
timestamp 1654648307
transform 1 0 103100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5589
timestamp 1654648307
transform 1 0 101600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5672
timestamp 1654648307
transform 1 0 106100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5671
timestamp 1654648307
transform 1 0 104600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5592
timestamp 1654648307
transform 1 0 106100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5591
timestamp 1654648307
transform 1 0 104600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5674
timestamp 1654648307
transform 1 0 109100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5673
timestamp 1654648307
transform 1 0 107600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5594
timestamp 1654648307
transform 1 0 109100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5593
timestamp 1654648307
transform 1 0 107600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5676
timestamp 1654648307
transform 1 0 112100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5675
timestamp 1654648307
transform 1 0 110600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5596
timestamp 1654648307
transform 1 0 112100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5595
timestamp 1654648307
transform 1 0 110600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5678
timestamp 1654648307
transform 1 0 115100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5677
timestamp 1654648307
transform 1 0 113600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5598
timestamp 1654648307
transform 1 0 115100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5597
timestamp 1654648307
transform 1 0 113600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5679
timestamp 1654648307
transform 1 0 116600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_5599
timestamp 1654648307
transform 1 0 116600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_5440
timestamp 1654648307
transform 1 0 -1900 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5360
timestamp 1654648307
transform 1 0 -1900 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5442
timestamp 1654648307
transform 1 0 1100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5441
timestamp 1654648307
transform 1 0 -400 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5362
timestamp 1654648307
transform 1 0 1100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5361
timestamp 1654648307
transform 1 0 -400 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5444
timestamp 1654648307
transform 1 0 4100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5443
timestamp 1654648307
transform 1 0 2600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5364
timestamp 1654648307
transform 1 0 4100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5363
timestamp 1654648307
transform 1 0 2600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5446
timestamp 1654648307
transform 1 0 7100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5445
timestamp 1654648307
transform 1 0 5600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5366
timestamp 1654648307
transform 1 0 7100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5365
timestamp 1654648307
transform 1 0 5600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5448
timestamp 1654648307
transform 1 0 10100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5447
timestamp 1654648307
transform 1 0 8600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5368
timestamp 1654648307
transform 1 0 10100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5367
timestamp 1654648307
transform 1 0 8600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5450
timestamp 1654648307
transform 1 0 13100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5449
timestamp 1654648307
transform 1 0 11600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5370
timestamp 1654648307
transform 1 0 13100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5369
timestamp 1654648307
transform 1 0 11600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5452
timestamp 1654648307
transform 1 0 16100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5451
timestamp 1654648307
transform 1 0 14600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5372
timestamp 1654648307
transform 1 0 16100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5371
timestamp 1654648307
transform 1 0 14600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5454
timestamp 1654648307
transform 1 0 19100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5453
timestamp 1654648307
transform 1 0 17600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5374
timestamp 1654648307
transform 1 0 19100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5373
timestamp 1654648307
transform 1 0 17600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5456
timestamp 1654648307
transform 1 0 22100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5455
timestamp 1654648307
transform 1 0 20600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5376
timestamp 1654648307
transform 1 0 22100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5375
timestamp 1654648307
transform 1 0 20600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5458
timestamp 1654648307
transform 1 0 25100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5457
timestamp 1654648307
transform 1 0 23600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5378
timestamp 1654648307
transform 1 0 25100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5377
timestamp 1654648307
transform 1 0 23600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5460
timestamp 1654648307
transform 1 0 28100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5459
timestamp 1654648307
transform 1 0 26600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5380
timestamp 1654648307
transform 1 0 28100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5379
timestamp 1654648307
transform 1 0 26600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5462
timestamp 1654648307
transform 1 0 31100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5461
timestamp 1654648307
transform 1 0 29600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5382
timestamp 1654648307
transform 1 0 31100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5381
timestamp 1654648307
transform 1 0 29600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5464
timestamp 1654648307
transform 1 0 34100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5463
timestamp 1654648307
transform 1 0 32600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5384
timestamp 1654648307
transform 1 0 34100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5383
timestamp 1654648307
transform 1 0 32600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5466
timestamp 1654648307
transform 1 0 37100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5465
timestamp 1654648307
transform 1 0 35600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5386
timestamp 1654648307
transform 1 0 37100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5385
timestamp 1654648307
transform 1 0 35600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5468
timestamp 1654648307
transform 1 0 40100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5467
timestamp 1654648307
transform 1 0 38600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5388
timestamp 1654648307
transform 1 0 40100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5387
timestamp 1654648307
transform 1 0 38600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5470
timestamp 1654648307
transform 1 0 43100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5469
timestamp 1654648307
transform 1 0 41600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5390
timestamp 1654648307
transform 1 0 43100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5389
timestamp 1654648307
transform 1 0 41600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5472
timestamp 1654648307
transform 1 0 46100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5471
timestamp 1654648307
transform 1 0 44600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5392
timestamp 1654648307
transform 1 0 46100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5391
timestamp 1654648307
transform 1 0 44600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5474
timestamp 1654648307
transform 1 0 49100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5473
timestamp 1654648307
transform 1 0 47600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5394
timestamp 1654648307
transform 1 0 49100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5393
timestamp 1654648307
transform 1 0 47600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5476
timestamp 1654648307
transform 1 0 52100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5475
timestamp 1654648307
transform 1 0 50600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5396
timestamp 1654648307
transform 1 0 52100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5395
timestamp 1654648307
transform 1 0 50600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5478
timestamp 1654648307
transform 1 0 55100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5477
timestamp 1654648307
transform 1 0 53600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5398
timestamp 1654648307
transform 1 0 55100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5397
timestamp 1654648307
transform 1 0 53600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5480
timestamp 1654648307
transform 1 0 58100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5479
timestamp 1654648307
transform 1 0 56600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5400
timestamp 1654648307
transform 1 0 58100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5399
timestamp 1654648307
transform 1 0 56600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5482
timestamp 1654648307
transform 1 0 61100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5481
timestamp 1654648307
transform 1 0 59600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5402
timestamp 1654648307
transform 1 0 61100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5401
timestamp 1654648307
transform 1 0 59600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5484
timestamp 1654648307
transform 1 0 64100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5483
timestamp 1654648307
transform 1 0 62600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5404
timestamp 1654648307
transform 1 0 64100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5403
timestamp 1654648307
transform 1 0 62600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5486
timestamp 1654648307
transform 1 0 67100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5485
timestamp 1654648307
transform 1 0 65600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5406
timestamp 1654648307
transform 1 0 67100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5405
timestamp 1654648307
transform 1 0 65600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5488
timestamp 1654648307
transform 1 0 70100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5487
timestamp 1654648307
transform 1 0 68600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5408
timestamp 1654648307
transform 1 0 70100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5407
timestamp 1654648307
transform 1 0 68600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5490
timestamp 1654648307
transform 1 0 73100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5489
timestamp 1654648307
transform 1 0 71600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5410
timestamp 1654648307
transform 1 0 73100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5409
timestamp 1654648307
transform 1 0 71600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5492
timestamp 1654648307
transform 1 0 76100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5491
timestamp 1654648307
transform 1 0 74600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5412
timestamp 1654648307
transform 1 0 76100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5411
timestamp 1654648307
transform 1 0 74600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5494
timestamp 1654648307
transform 1 0 79100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5493
timestamp 1654648307
transform 1 0 77600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5414
timestamp 1654648307
transform 1 0 79100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5413
timestamp 1654648307
transform 1 0 77600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5496
timestamp 1654648307
transform 1 0 82100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5495
timestamp 1654648307
transform 1 0 80600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5416
timestamp 1654648307
transform 1 0 82100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5415
timestamp 1654648307
transform 1 0 80600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5498
timestamp 1654648307
transform 1 0 85100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5497
timestamp 1654648307
transform 1 0 83600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5418
timestamp 1654648307
transform 1 0 85100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5417
timestamp 1654648307
transform 1 0 83600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5500
timestamp 1654648307
transform 1 0 88100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5499
timestamp 1654648307
transform 1 0 86600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5420
timestamp 1654648307
transform 1 0 88100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5419
timestamp 1654648307
transform 1 0 86600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5502
timestamp 1654648307
transform 1 0 91100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5501
timestamp 1654648307
transform 1 0 89600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5422
timestamp 1654648307
transform 1 0 91100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5421
timestamp 1654648307
transform 1 0 89600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5504
timestamp 1654648307
transform 1 0 94100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5503
timestamp 1654648307
transform 1 0 92600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5424
timestamp 1654648307
transform 1 0 94100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5423
timestamp 1654648307
transform 1 0 92600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5506
timestamp 1654648307
transform 1 0 97100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5505
timestamp 1654648307
transform 1 0 95600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5426
timestamp 1654648307
transform 1 0 97100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5425
timestamp 1654648307
transform 1 0 95600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5508
timestamp 1654648307
transform 1 0 100100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5507
timestamp 1654648307
transform 1 0 98600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5428
timestamp 1654648307
transform 1 0 100100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5427
timestamp 1654648307
transform 1 0 98600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5510
timestamp 1654648307
transform 1 0 103100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5509
timestamp 1654648307
transform 1 0 101600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5430
timestamp 1654648307
transform 1 0 103100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5429
timestamp 1654648307
transform 1 0 101600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5512
timestamp 1654648307
transform 1 0 106100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5511
timestamp 1654648307
transform 1 0 104600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5432
timestamp 1654648307
transform 1 0 106100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5431
timestamp 1654648307
transform 1 0 104600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5514
timestamp 1654648307
transform 1 0 109100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5513
timestamp 1654648307
transform 1 0 107600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5434
timestamp 1654648307
transform 1 0 109100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5433
timestamp 1654648307
transform 1 0 107600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5516
timestamp 1654648307
transform 1 0 112100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5515
timestamp 1654648307
transform 1 0 110600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5436
timestamp 1654648307
transform 1 0 112100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5435
timestamp 1654648307
transform 1 0 110600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5518
timestamp 1654648307
transform 1 0 115100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5517
timestamp 1654648307
transform 1 0 113600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5438
timestamp 1654648307
transform 1 0 115100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5437
timestamp 1654648307
transform 1 0 113600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5519
timestamp 1654648307
transform 1 0 116600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_5439
timestamp 1654648307
transform 1 0 116600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_5280
timestamp 1654648307
transform 1 0 -1900 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5200
timestamp 1654648307
transform 1 0 -1900 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5282
timestamp 1654648307
transform 1 0 1100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5281
timestamp 1654648307
transform 1 0 -400 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5202
timestamp 1654648307
transform 1 0 1100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5201
timestamp 1654648307
transform 1 0 -400 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5284
timestamp 1654648307
transform 1 0 4100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5283
timestamp 1654648307
transform 1 0 2600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5204
timestamp 1654648307
transform 1 0 4100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5203
timestamp 1654648307
transform 1 0 2600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5286
timestamp 1654648307
transform 1 0 7100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5285
timestamp 1654648307
transform 1 0 5600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5206
timestamp 1654648307
transform 1 0 7100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5205
timestamp 1654648307
transform 1 0 5600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5288
timestamp 1654648307
transform 1 0 10100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5287
timestamp 1654648307
transform 1 0 8600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5208
timestamp 1654648307
transform 1 0 10100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5207
timestamp 1654648307
transform 1 0 8600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5290
timestamp 1654648307
transform 1 0 13100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5289
timestamp 1654648307
transform 1 0 11600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5210
timestamp 1654648307
transform 1 0 13100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5209
timestamp 1654648307
transform 1 0 11600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5292
timestamp 1654648307
transform 1 0 16100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5291
timestamp 1654648307
transform 1 0 14600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5212
timestamp 1654648307
transform 1 0 16100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5211
timestamp 1654648307
transform 1 0 14600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5294
timestamp 1654648307
transform 1 0 19100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5293
timestamp 1654648307
transform 1 0 17600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5214
timestamp 1654648307
transform 1 0 19100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5213
timestamp 1654648307
transform 1 0 17600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5296
timestamp 1654648307
transform 1 0 22100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5295
timestamp 1654648307
transform 1 0 20600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5216
timestamp 1654648307
transform 1 0 22100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5215
timestamp 1654648307
transform 1 0 20600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5298
timestamp 1654648307
transform 1 0 25100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5297
timestamp 1654648307
transform 1 0 23600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5218
timestamp 1654648307
transform 1 0 25100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5217
timestamp 1654648307
transform 1 0 23600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5300
timestamp 1654648307
transform 1 0 28100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5299
timestamp 1654648307
transform 1 0 26600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5220
timestamp 1654648307
transform 1 0 28100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5219
timestamp 1654648307
transform 1 0 26600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5302
timestamp 1654648307
transform 1 0 31100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5301
timestamp 1654648307
transform 1 0 29600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5222
timestamp 1654648307
transform 1 0 31100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5221
timestamp 1654648307
transform 1 0 29600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5304
timestamp 1654648307
transform 1 0 34100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5303
timestamp 1654648307
transform 1 0 32600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5224
timestamp 1654648307
transform 1 0 34100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5223
timestamp 1654648307
transform 1 0 32600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5306
timestamp 1654648307
transform 1 0 37100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5305
timestamp 1654648307
transform 1 0 35600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5226
timestamp 1654648307
transform 1 0 37100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5225
timestamp 1654648307
transform 1 0 35600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5308
timestamp 1654648307
transform 1 0 40100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5307
timestamp 1654648307
transform 1 0 38600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5228
timestamp 1654648307
transform 1 0 40100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5227
timestamp 1654648307
transform 1 0 38600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5310
timestamp 1654648307
transform 1 0 43100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5309
timestamp 1654648307
transform 1 0 41600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5230
timestamp 1654648307
transform 1 0 43100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5229
timestamp 1654648307
transform 1 0 41600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5312
timestamp 1654648307
transform 1 0 46100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5311
timestamp 1654648307
transform 1 0 44600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5232
timestamp 1654648307
transform 1 0 46100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5231
timestamp 1654648307
transform 1 0 44600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5314
timestamp 1654648307
transform 1 0 49100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5313
timestamp 1654648307
transform 1 0 47600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5234
timestamp 1654648307
transform 1 0 49100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5233
timestamp 1654648307
transform 1 0 47600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5316
timestamp 1654648307
transform 1 0 52100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5315
timestamp 1654648307
transform 1 0 50600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5236
timestamp 1654648307
transform 1 0 52100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5235
timestamp 1654648307
transform 1 0 50600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5318
timestamp 1654648307
transform 1 0 55100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5317
timestamp 1654648307
transform 1 0 53600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5238
timestamp 1654648307
transform 1 0 55100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5237
timestamp 1654648307
transform 1 0 53600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5320
timestamp 1654648307
transform 1 0 58100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5319
timestamp 1654648307
transform 1 0 56600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5240
timestamp 1654648307
transform 1 0 58100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5239
timestamp 1654648307
transform 1 0 56600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5322
timestamp 1654648307
transform 1 0 61100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5321
timestamp 1654648307
transform 1 0 59600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5242
timestamp 1654648307
transform 1 0 61100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5241
timestamp 1654648307
transform 1 0 59600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5324
timestamp 1654648307
transform 1 0 64100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5323
timestamp 1654648307
transform 1 0 62600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5244
timestamp 1654648307
transform 1 0 64100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5243
timestamp 1654648307
transform 1 0 62600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5326
timestamp 1654648307
transform 1 0 67100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5325
timestamp 1654648307
transform 1 0 65600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5246
timestamp 1654648307
transform 1 0 67100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5245
timestamp 1654648307
transform 1 0 65600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5328
timestamp 1654648307
transform 1 0 70100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5327
timestamp 1654648307
transform 1 0 68600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5248
timestamp 1654648307
transform 1 0 70100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5247
timestamp 1654648307
transform 1 0 68600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5330
timestamp 1654648307
transform 1 0 73100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5329
timestamp 1654648307
transform 1 0 71600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5250
timestamp 1654648307
transform 1 0 73100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5249
timestamp 1654648307
transform 1 0 71600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5332
timestamp 1654648307
transform 1 0 76100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5331
timestamp 1654648307
transform 1 0 74600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5252
timestamp 1654648307
transform 1 0 76100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5251
timestamp 1654648307
transform 1 0 74600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5334
timestamp 1654648307
transform 1 0 79100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5333
timestamp 1654648307
transform 1 0 77600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5254
timestamp 1654648307
transform 1 0 79100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5253
timestamp 1654648307
transform 1 0 77600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5336
timestamp 1654648307
transform 1 0 82100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5335
timestamp 1654648307
transform 1 0 80600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5256
timestamp 1654648307
transform 1 0 82100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5255
timestamp 1654648307
transform 1 0 80600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5338
timestamp 1654648307
transform 1 0 85100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5337
timestamp 1654648307
transform 1 0 83600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5258
timestamp 1654648307
transform 1 0 85100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5257
timestamp 1654648307
transform 1 0 83600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5340
timestamp 1654648307
transform 1 0 88100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5339
timestamp 1654648307
transform 1 0 86600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5260
timestamp 1654648307
transform 1 0 88100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5259
timestamp 1654648307
transform 1 0 86600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5342
timestamp 1654648307
transform 1 0 91100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5341
timestamp 1654648307
transform 1 0 89600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5262
timestamp 1654648307
transform 1 0 91100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5261
timestamp 1654648307
transform 1 0 89600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5344
timestamp 1654648307
transform 1 0 94100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5343
timestamp 1654648307
transform 1 0 92600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5264
timestamp 1654648307
transform 1 0 94100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5263
timestamp 1654648307
transform 1 0 92600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5346
timestamp 1654648307
transform 1 0 97100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5345
timestamp 1654648307
transform 1 0 95600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5266
timestamp 1654648307
transform 1 0 97100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5265
timestamp 1654648307
transform 1 0 95600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5348
timestamp 1654648307
transform 1 0 100100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5347
timestamp 1654648307
transform 1 0 98600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5268
timestamp 1654648307
transform 1 0 100100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5267
timestamp 1654648307
transform 1 0 98600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5350
timestamp 1654648307
transform 1 0 103100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5349
timestamp 1654648307
transform 1 0 101600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5270
timestamp 1654648307
transform 1 0 103100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5269
timestamp 1654648307
transform 1 0 101600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5352
timestamp 1654648307
transform 1 0 106100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5351
timestamp 1654648307
transform 1 0 104600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5272
timestamp 1654648307
transform 1 0 106100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5271
timestamp 1654648307
transform 1 0 104600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5354
timestamp 1654648307
transform 1 0 109100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5353
timestamp 1654648307
transform 1 0 107600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5274
timestamp 1654648307
transform 1 0 109100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5273
timestamp 1654648307
transform 1 0 107600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5356
timestamp 1654648307
transform 1 0 112100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5355
timestamp 1654648307
transform 1 0 110600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5276
timestamp 1654648307
transform 1 0 112100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5275
timestamp 1654648307
transform 1 0 110600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5358
timestamp 1654648307
transform 1 0 115100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5357
timestamp 1654648307
transform 1 0 113600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5278
timestamp 1654648307
transform 1 0 115100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5277
timestamp 1654648307
transform 1 0 113600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5359
timestamp 1654648307
transform 1 0 116600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_5279
timestamp 1654648307
transform 1 0 116600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_5120
timestamp 1654648307
transform 1 0 -1900 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5040
timestamp 1654648307
transform 1 0 -1900 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5122
timestamp 1654648307
transform 1 0 1100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5121
timestamp 1654648307
transform 1 0 -400 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5042
timestamp 1654648307
transform 1 0 1100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5041
timestamp 1654648307
transform 1 0 -400 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5124
timestamp 1654648307
transform 1 0 4100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5123
timestamp 1654648307
transform 1 0 2600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5044
timestamp 1654648307
transform 1 0 4100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5043
timestamp 1654648307
transform 1 0 2600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5126
timestamp 1654648307
transform 1 0 7100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5125
timestamp 1654648307
transform 1 0 5600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5046
timestamp 1654648307
transform 1 0 7100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5045
timestamp 1654648307
transform 1 0 5600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5128
timestamp 1654648307
transform 1 0 10100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5127
timestamp 1654648307
transform 1 0 8600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5048
timestamp 1654648307
transform 1 0 10100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5047
timestamp 1654648307
transform 1 0 8600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5130
timestamp 1654648307
transform 1 0 13100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5129
timestamp 1654648307
transform 1 0 11600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5050
timestamp 1654648307
transform 1 0 13100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5049
timestamp 1654648307
transform 1 0 11600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5132
timestamp 1654648307
transform 1 0 16100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5131
timestamp 1654648307
transform 1 0 14600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5052
timestamp 1654648307
transform 1 0 16100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5051
timestamp 1654648307
transform 1 0 14600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5134
timestamp 1654648307
transform 1 0 19100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5133
timestamp 1654648307
transform 1 0 17600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5054
timestamp 1654648307
transform 1 0 19100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5053
timestamp 1654648307
transform 1 0 17600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5136
timestamp 1654648307
transform 1 0 22100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5135
timestamp 1654648307
transform 1 0 20600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5056
timestamp 1654648307
transform 1 0 22100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5055
timestamp 1654648307
transform 1 0 20600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5138
timestamp 1654648307
transform 1 0 25100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5137
timestamp 1654648307
transform 1 0 23600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5058
timestamp 1654648307
transform 1 0 25100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5057
timestamp 1654648307
transform 1 0 23600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5140
timestamp 1654648307
transform 1 0 28100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5139
timestamp 1654648307
transform 1 0 26600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5060
timestamp 1654648307
transform 1 0 28100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5059
timestamp 1654648307
transform 1 0 26600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5142
timestamp 1654648307
transform 1 0 31100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5141
timestamp 1654648307
transform 1 0 29600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5062
timestamp 1654648307
transform 1 0 31100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5061
timestamp 1654648307
transform 1 0 29600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5144
timestamp 1654648307
transform 1 0 34100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5143
timestamp 1654648307
transform 1 0 32600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5064
timestamp 1654648307
transform 1 0 34100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5063
timestamp 1654648307
transform 1 0 32600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5146
timestamp 1654648307
transform 1 0 37100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5145
timestamp 1654648307
transform 1 0 35600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5066
timestamp 1654648307
transform 1 0 37100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5065
timestamp 1654648307
transform 1 0 35600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5148
timestamp 1654648307
transform 1 0 40100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5147
timestamp 1654648307
transform 1 0 38600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5068
timestamp 1654648307
transform 1 0 40100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5067
timestamp 1654648307
transform 1 0 38600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5150
timestamp 1654648307
transform 1 0 43100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5149
timestamp 1654648307
transform 1 0 41600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5070
timestamp 1654648307
transform 1 0 43100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5069
timestamp 1654648307
transform 1 0 41600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5152
timestamp 1654648307
transform 1 0 46100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5151
timestamp 1654648307
transform 1 0 44600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5072
timestamp 1654648307
transform 1 0 46100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5071
timestamp 1654648307
transform 1 0 44600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5154
timestamp 1654648307
transform 1 0 49100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5153
timestamp 1654648307
transform 1 0 47600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5074
timestamp 1654648307
transform 1 0 49100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5073
timestamp 1654648307
transform 1 0 47600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5156
timestamp 1654648307
transform 1 0 52100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5155
timestamp 1654648307
transform 1 0 50600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5076
timestamp 1654648307
transform 1 0 52100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5075
timestamp 1654648307
transform 1 0 50600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5158
timestamp 1654648307
transform 1 0 55100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5157
timestamp 1654648307
transform 1 0 53600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5078
timestamp 1654648307
transform 1 0 55100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5077
timestamp 1654648307
transform 1 0 53600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5160
timestamp 1654648307
transform 1 0 58100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5159
timestamp 1654648307
transform 1 0 56600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5080
timestamp 1654648307
transform 1 0 58100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5079
timestamp 1654648307
transform 1 0 56600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5162
timestamp 1654648307
transform 1 0 61100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5161
timestamp 1654648307
transform 1 0 59600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5082
timestamp 1654648307
transform 1 0 61100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5081
timestamp 1654648307
transform 1 0 59600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5164
timestamp 1654648307
transform 1 0 64100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5163
timestamp 1654648307
transform 1 0 62600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5084
timestamp 1654648307
transform 1 0 64100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5083
timestamp 1654648307
transform 1 0 62600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5166
timestamp 1654648307
transform 1 0 67100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5165
timestamp 1654648307
transform 1 0 65600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5086
timestamp 1654648307
transform 1 0 67100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5085
timestamp 1654648307
transform 1 0 65600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5168
timestamp 1654648307
transform 1 0 70100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5167
timestamp 1654648307
transform 1 0 68600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5088
timestamp 1654648307
transform 1 0 70100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5087
timestamp 1654648307
transform 1 0 68600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5170
timestamp 1654648307
transform 1 0 73100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5169
timestamp 1654648307
transform 1 0 71600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5090
timestamp 1654648307
transform 1 0 73100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5089
timestamp 1654648307
transform 1 0 71600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5172
timestamp 1654648307
transform 1 0 76100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5171
timestamp 1654648307
transform 1 0 74600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5092
timestamp 1654648307
transform 1 0 76100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5091
timestamp 1654648307
transform 1 0 74600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5174
timestamp 1654648307
transform 1 0 79100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5173
timestamp 1654648307
transform 1 0 77600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5094
timestamp 1654648307
transform 1 0 79100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5093
timestamp 1654648307
transform 1 0 77600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5176
timestamp 1654648307
transform 1 0 82100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5175
timestamp 1654648307
transform 1 0 80600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5096
timestamp 1654648307
transform 1 0 82100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5095
timestamp 1654648307
transform 1 0 80600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5178
timestamp 1654648307
transform 1 0 85100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5177
timestamp 1654648307
transform 1 0 83600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5098
timestamp 1654648307
transform 1 0 85100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5097
timestamp 1654648307
transform 1 0 83600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5180
timestamp 1654648307
transform 1 0 88100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5179
timestamp 1654648307
transform 1 0 86600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5100
timestamp 1654648307
transform 1 0 88100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5099
timestamp 1654648307
transform 1 0 86600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5182
timestamp 1654648307
transform 1 0 91100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5181
timestamp 1654648307
transform 1 0 89600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5102
timestamp 1654648307
transform 1 0 91100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5101
timestamp 1654648307
transform 1 0 89600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5184
timestamp 1654648307
transform 1 0 94100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5183
timestamp 1654648307
transform 1 0 92600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5104
timestamp 1654648307
transform 1 0 94100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5103
timestamp 1654648307
transform 1 0 92600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5186
timestamp 1654648307
transform 1 0 97100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5185
timestamp 1654648307
transform 1 0 95600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5106
timestamp 1654648307
transform 1 0 97100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5105
timestamp 1654648307
transform 1 0 95600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5188
timestamp 1654648307
transform 1 0 100100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5187
timestamp 1654648307
transform 1 0 98600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5108
timestamp 1654648307
transform 1 0 100100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5107
timestamp 1654648307
transform 1 0 98600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5190
timestamp 1654648307
transform 1 0 103100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5189
timestamp 1654648307
transform 1 0 101600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5110
timestamp 1654648307
transform 1 0 103100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5109
timestamp 1654648307
transform 1 0 101600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5192
timestamp 1654648307
transform 1 0 106100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5191
timestamp 1654648307
transform 1 0 104600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5112
timestamp 1654648307
transform 1 0 106100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5111
timestamp 1654648307
transform 1 0 104600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5194
timestamp 1654648307
transform 1 0 109100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5193
timestamp 1654648307
transform 1 0 107600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5114
timestamp 1654648307
transform 1 0 109100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5113
timestamp 1654648307
transform 1 0 107600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5196
timestamp 1654648307
transform 1 0 112100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5195
timestamp 1654648307
transform 1 0 110600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5116
timestamp 1654648307
transform 1 0 112100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5115
timestamp 1654648307
transform 1 0 110600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5198
timestamp 1654648307
transform 1 0 115100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5197
timestamp 1654648307
transform 1 0 113600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5118
timestamp 1654648307
transform 1 0 115100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5117
timestamp 1654648307
transform 1 0 113600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_5199
timestamp 1654648307
transform 1 0 116600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_5119
timestamp 1654648307
transform 1 0 116600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_4960
timestamp 1654648307
transform 1 0 -1900 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4880
timestamp 1654648307
transform 1 0 -1900 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4962
timestamp 1654648307
transform 1 0 1100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4961
timestamp 1654648307
transform 1 0 -400 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4882
timestamp 1654648307
transform 1 0 1100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4881
timestamp 1654648307
transform 1 0 -400 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4964
timestamp 1654648307
transform 1 0 4100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4963
timestamp 1654648307
transform 1 0 2600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4884
timestamp 1654648307
transform 1 0 4100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4883
timestamp 1654648307
transform 1 0 2600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4966
timestamp 1654648307
transform 1 0 7100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4965
timestamp 1654648307
transform 1 0 5600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4886
timestamp 1654648307
transform 1 0 7100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4885
timestamp 1654648307
transform 1 0 5600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4968
timestamp 1654648307
transform 1 0 10100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4967
timestamp 1654648307
transform 1 0 8600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4888
timestamp 1654648307
transform 1 0 10100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4887
timestamp 1654648307
transform 1 0 8600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4970
timestamp 1654648307
transform 1 0 13100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4969
timestamp 1654648307
transform 1 0 11600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4890
timestamp 1654648307
transform 1 0 13100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4889
timestamp 1654648307
transform 1 0 11600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4972
timestamp 1654648307
transform 1 0 16100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4971
timestamp 1654648307
transform 1 0 14600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4892
timestamp 1654648307
transform 1 0 16100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4891
timestamp 1654648307
transform 1 0 14600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4974
timestamp 1654648307
transform 1 0 19100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4973
timestamp 1654648307
transform 1 0 17600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4894
timestamp 1654648307
transform 1 0 19100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4893
timestamp 1654648307
transform 1 0 17600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4976
timestamp 1654648307
transform 1 0 22100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4975
timestamp 1654648307
transform 1 0 20600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4896
timestamp 1654648307
transform 1 0 22100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4895
timestamp 1654648307
transform 1 0 20600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4978
timestamp 1654648307
transform 1 0 25100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4977
timestamp 1654648307
transform 1 0 23600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4898
timestamp 1654648307
transform 1 0 25100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4897
timestamp 1654648307
transform 1 0 23600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4980
timestamp 1654648307
transform 1 0 28100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4979
timestamp 1654648307
transform 1 0 26600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4900
timestamp 1654648307
transform 1 0 28100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4899
timestamp 1654648307
transform 1 0 26600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4982
timestamp 1654648307
transform 1 0 31100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4981
timestamp 1654648307
transform 1 0 29600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4902
timestamp 1654648307
transform 1 0 31100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4901
timestamp 1654648307
transform 1 0 29600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4984
timestamp 1654648307
transform 1 0 34100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4983
timestamp 1654648307
transform 1 0 32600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4904
timestamp 1654648307
transform 1 0 34100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4903
timestamp 1654648307
transform 1 0 32600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4986
timestamp 1654648307
transform 1 0 37100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4985
timestamp 1654648307
transform 1 0 35600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4906
timestamp 1654648307
transform 1 0 37100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4905
timestamp 1654648307
transform 1 0 35600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4988
timestamp 1654648307
transform 1 0 40100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4987
timestamp 1654648307
transform 1 0 38600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4908
timestamp 1654648307
transform 1 0 40100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4907
timestamp 1654648307
transform 1 0 38600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4990
timestamp 1654648307
transform 1 0 43100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4989
timestamp 1654648307
transform 1 0 41600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4910
timestamp 1654648307
transform 1 0 43100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4909
timestamp 1654648307
transform 1 0 41600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4992
timestamp 1654648307
transform 1 0 46100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4991
timestamp 1654648307
transform 1 0 44600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4912
timestamp 1654648307
transform 1 0 46100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4911
timestamp 1654648307
transform 1 0 44600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4994
timestamp 1654648307
transform 1 0 49100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4993
timestamp 1654648307
transform 1 0 47600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4914
timestamp 1654648307
transform 1 0 49100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4913
timestamp 1654648307
transform 1 0 47600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4996
timestamp 1654648307
transform 1 0 52100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4995
timestamp 1654648307
transform 1 0 50600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4916
timestamp 1654648307
transform 1 0 52100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4915
timestamp 1654648307
transform 1 0 50600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4998
timestamp 1654648307
transform 1 0 55100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4997
timestamp 1654648307
transform 1 0 53600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4918
timestamp 1654648307
transform 1 0 55100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4917
timestamp 1654648307
transform 1 0 53600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_5000
timestamp 1654648307
transform 1 0 58100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4999
timestamp 1654648307
transform 1 0 56600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4920
timestamp 1654648307
transform 1 0 58100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4919
timestamp 1654648307
transform 1 0 56600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_5002
timestamp 1654648307
transform 1 0 61100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_5001
timestamp 1654648307
transform 1 0 59600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4922
timestamp 1654648307
transform 1 0 61100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4921
timestamp 1654648307
transform 1 0 59600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_5004
timestamp 1654648307
transform 1 0 64100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_5003
timestamp 1654648307
transform 1 0 62600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4924
timestamp 1654648307
transform 1 0 64100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4923
timestamp 1654648307
transform 1 0 62600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_5006
timestamp 1654648307
transform 1 0 67100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_5005
timestamp 1654648307
transform 1 0 65600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4926
timestamp 1654648307
transform 1 0 67100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4925
timestamp 1654648307
transform 1 0 65600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_5008
timestamp 1654648307
transform 1 0 70100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_5007
timestamp 1654648307
transform 1 0 68600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4928
timestamp 1654648307
transform 1 0 70100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4927
timestamp 1654648307
transform 1 0 68600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_5010
timestamp 1654648307
transform 1 0 73100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_5009
timestamp 1654648307
transform 1 0 71600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4930
timestamp 1654648307
transform 1 0 73100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4929
timestamp 1654648307
transform 1 0 71600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_5012
timestamp 1654648307
transform 1 0 76100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_5011
timestamp 1654648307
transform 1 0 74600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4932
timestamp 1654648307
transform 1 0 76100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4931
timestamp 1654648307
transform 1 0 74600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_5014
timestamp 1654648307
transform 1 0 79100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_5013
timestamp 1654648307
transform 1 0 77600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4934
timestamp 1654648307
transform 1 0 79100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4933
timestamp 1654648307
transform 1 0 77600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_5016
timestamp 1654648307
transform 1 0 82100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_5015
timestamp 1654648307
transform 1 0 80600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4936
timestamp 1654648307
transform 1 0 82100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4935
timestamp 1654648307
transform 1 0 80600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_5018
timestamp 1654648307
transform 1 0 85100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_5017
timestamp 1654648307
transform 1 0 83600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4938
timestamp 1654648307
transform 1 0 85100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4937
timestamp 1654648307
transform 1 0 83600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_5020
timestamp 1654648307
transform 1 0 88100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_5019
timestamp 1654648307
transform 1 0 86600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4940
timestamp 1654648307
transform 1 0 88100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4939
timestamp 1654648307
transform 1 0 86600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_5022
timestamp 1654648307
transform 1 0 91100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_5021
timestamp 1654648307
transform 1 0 89600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4942
timestamp 1654648307
transform 1 0 91100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4941
timestamp 1654648307
transform 1 0 89600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_5024
timestamp 1654648307
transform 1 0 94100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_5023
timestamp 1654648307
transform 1 0 92600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4944
timestamp 1654648307
transform 1 0 94100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4943
timestamp 1654648307
transform 1 0 92600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_5026
timestamp 1654648307
transform 1 0 97100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_5025
timestamp 1654648307
transform 1 0 95600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4946
timestamp 1654648307
transform 1 0 97100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4945
timestamp 1654648307
transform 1 0 95600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_5028
timestamp 1654648307
transform 1 0 100100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_5027
timestamp 1654648307
transform 1 0 98600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4948
timestamp 1654648307
transform 1 0 100100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4947
timestamp 1654648307
transform 1 0 98600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_5030
timestamp 1654648307
transform 1 0 103100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_5029
timestamp 1654648307
transform 1 0 101600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4950
timestamp 1654648307
transform 1 0 103100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4949
timestamp 1654648307
transform 1 0 101600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_5032
timestamp 1654648307
transform 1 0 106100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_5031
timestamp 1654648307
transform 1 0 104600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4952
timestamp 1654648307
transform 1 0 106100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4951
timestamp 1654648307
transform 1 0 104600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_5034
timestamp 1654648307
transform 1 0 109100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_5033
timestamp 1654648307
transform 1 0 107600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4954
timestamp 1654648307
transform 1 0 109100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4953
timestamp 1654648307
transform 1 0 107600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_5036
timestamp 1654648307
transform 1 0 112100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_5035
timestamp 1654648307
transform 1 0 110600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4956
timestamp 1654648307
transform 1 0 112100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4955
timestamp 1654648307
transform 1 0 110600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_5038
timestamp 1654648307
transform 1 0 115100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_5037
timestamp 1654648307
transform 1 0 113600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4958
timestamp 1654648307
transform 1 0 115100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4957
timestamp 1654648307
transform 1 0 113600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_5039
timestamp 1654648307
transform 1 0 116600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_4959
timestamp 1654648307
transform 1 0 116600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_4720
timestamp 1654648307
transform 1 0 -1900 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4800
timestamp 1654648307
transform 1 0 -1900 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4722
timestamp 1654648307
transform 1 0 1100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4721
timestamp 1654648307
transform 1 0 -400 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4802
timestamp 1654648307
transform 1 0 1100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4801
timestamp 1654648307
transform 1 0 -400 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4724
timestamp 1654648307
transform 1 0 4100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4723
timestamp 1654648307
transform 1 0 2600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4804
timestamp 1654648307
transform 1 0 4100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4803
timestamp 1654648307
transform 1 0 2600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4726
timestamp 1654648307
transform 1 0 7100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4725
timestamp 1654648307
transform 1 0 5600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4806
timestamp 1654648307
transform 1 0 7100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4805
timestamp 1654648307
transform 1 0 5600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4728
timestamp 1654648307
transform 1 0 10100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4727
timestamp 1654648307
transform 1 0 8600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4808
timestamp 1654648307
transform 1 0 10100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4807
timestamp 1654648307
transform 1 0 8600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4810
timestamp 1654648307
transform 1 0 13100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4730
timestamp 1654648307
transform 1 0 13100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4729
timestamp 1654648307
transform 1 0 11600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4809
timestamp 1654648307
transform 1 0 11600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4812
timestamp 1654648307
transform 1 0 16100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4811
timestamp 1654648307
transform 1 0 14600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4732
timestamp 1654648307
transform 1 0 16100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4731
timestamp 1654648307
transform 1 0 14600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4814
timestamp 1654648307
transform 1 0 19100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4813
timestamp 1654648307
transform 1 0 17600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4734
timestamp 1654648307
transform 1 0 19100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4733
timestamp 1654648307
transform 1 0 17600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4816
timestamp 1654648307
transform 1 0 22100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4815
timestamp 1654648307
transform 1 0 20600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4736
timestamp 1654648307
transform 1 0 22100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4735
timestamp 1654648307
transform 1 0 20600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4818
timestamp 1654648307
transform 1 0 25100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4817
timestamp 1654648307
transform 1 0 23600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4738
timestamp 1654648307
transform 1 0 25100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4737
timestamp 1654648307
transform 1 0 23600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4820
timestamp 1654648307
transform 1 0 28100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4819
timestamp 1654648307
transform 1 0 26600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4740
timestamp 1654648307
transform 1 0 28100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4739
timestamp 1654648307
transform 1 0 26600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4822
timestamp 1654648307
transform 1 0 31100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4821
timestamp 1654648307
transform 1 0 29600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4742
timestamp 1654648307
transform 1 0 31100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4741
timestamp 1654648307
transform 1 0 29600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4824
timestamp 1654648307
transform 1 0 34100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4823
timestamp 1654648307
transform 1 0 32600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4744
timestamp 1654648307
transform 1 0 34100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4743
timestamp 1654648307
transform 1 0 32600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4826
timestamp 1654648307
transform 1 0 37100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4825
timestamp 1654648307
transform 1 0 35600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4746
timestamp 1654648307
transform 1 0 37100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4745
timestamp 1654648307
transform 1 0 35600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4828
timestamp 1654648307
transform 1 0 40100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4827
timestamp 1654648307
transform 1 0 38600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4748
timestamp 1654648307
transform 1 0 40100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4747
timestamp 1654648307
transform 1 0 38600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4830
timestamp 1654648307
transform 1 0 43100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4829
timestamp 1654648307
transform 1 0 41600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4750
timestamp 1654648307
transform 1 0 43100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4749
timestamp 1654648307
transform 1 0 41600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4832
timestamp 1654648307
transform 1 0 46100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4831
timestamp 1654648307
transform 1 0 44600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4752
timestamp 1654648307
transform 1 0 46100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4751
timestamp 1654648307
transform 1 0 44600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4834
timestamp 1654648307
transform 1 0 49100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4833
timestamp 1654648307
transform 1 0 47600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4754
timestamp 1654648307
transform 1 0 49100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4753
timestamp 1654648307
transform 1 0 47600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4836
timestamp 1654648307
transform 1 0 52100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4835
timestamp 1654648307
transform 1 0 50600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4756
timestamp 1654648307
transform 1 0 52100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4755
timestamp 1654648307
transform 1 0 50600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4838
timestamp 1654648307
transform 1 0 55100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4837
timestamp 1654648307
transform 1 0 53600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4758
timestamp 1654648307
transform 1 0 55100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4757
timestamp 1654648307
transform 1 0 53600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4840
timestamp 1654648307
transform 1 0 58100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4839
timestamp 1654648307
transform 1 0 56600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4760
timestamp 1654648307
transform 1 0 58100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4759
timestamp 1654648307
transform 1 0 56600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4842
timestamp 1654648307
transform 1 0 61100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4841
timestamp 1654648307
transform 1 0 59600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4762
timestamp 1654648307
transform 1 0 61100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4761
timestamp 1654648307
transform 1 0 59600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4844
timestamp 1654648307
transform 1 0 64100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4843
timestamp 1654648307
transform 1 0 62600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4763
timestamp 1654648307
transform 1 0 62600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4764
timestamp 1654648307
transform 1 0 64100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4846
timestamp 1654648307
transform 1 0 67100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4845
timestamp 1654648307
transform 1 0 65600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4765
timestamp 1654648307
transform 1 0 65600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4766
timestamp 1654648307
transform 1 0 67100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4848
timestamp 1654648307
transform 1 0 70100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4847
timestamp 1654648307
transform 1 0 68600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4767
timestamp 1654648307
transform 1 0 68600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4768
timestamp 1654648307
transform 1 0 70100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4850
timestamp 1654648307
transform 1 0 73100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4849
timestamp 1654648307
transform 1 0 71600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4769
timestamp 1654648307
transform 1 0 71600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4770
timestamp 1654648307
transform 1 0 73100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4852
timestamp 1654648307
transform 1 0 76100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4851
timestamp 1654648307
transform 1 0 74600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4771
timestamp 1654648307
transform 1 0 74600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4772
timestamp 1654648307
transform 1 0 76100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4854
timestamp 1654648307
transform 1 0 79100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4853
timestamp 1654648307
transform 1 0 77600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4773
timestamp 1654648307
transform 1 0 77600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4774
timestamp 1654648307
transform 1 0 79100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4856
timestamp 1654648307
transform 1 0 82100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4855
timestamp 1654648307
transform 1 0 80600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4775
timestamp 1654648307
transform 1 0 80600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4776
timestamp 1654648307
transform 1 0 82100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4858
timestamp 1654648307
transform 1 0 85100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4857
timestamp 1654648307
transform 1 0 83600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4777
timestamp 1654648307
transform 1 0 83600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4778
timestamp 1654648307
transform 1 0 85100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4860
timestamp 1654648307
transform 1 0 88100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4859
timestamp 1654648307
transform 1 0 86600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4779
timestamp 1654648307
transform 1 0 86600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4780
timestamp 1654648307
transform 1 0 88100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4862
timestamp 1654648307
transform 1 0 91100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4861
timestamp 1654648307
transform 1 0 89600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4781
timestamp 1654648307
transform 1 0 89600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4782
timestamp 1654648307
transform 1 0 91100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4864
timestamp 1654648307
transform 1 0 94100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4863
timestamp 1654648307
transform 1 0 92600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4783
timestamp 1654648307
transform 1 0 92600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4784
timestamp 1654648307
transform 1 0 94100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4866
timestamp 1654648307
transform 1 0 97100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4865
timestamp 1654648307
transform 1 0 95600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4785
timestamp 1654648307
transform 1 0 95600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4786
timestamp 1654648307
transform 1 0 97100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4868
timestamp 1654648307
transform 1 0 100100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4867
timestamp 1654648307
transform 1 0 98600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4787
timestamp 1654648307
transform 1 0 98600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4788
timestamp 1654648307
transform 1 0 100100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4870
timestamp 1654648307
transform 1 0 103100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4869
timestamp 1654648307
transform 1 0 101600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4789
timestamp 1654648307
transform 1 0 101600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4790
timestamp 1654648307
transform 1 0 103100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4872
timestamp 1654648307
transform 1 0 106100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4871
timestamp 1654648307
transform 1 0 104600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4791
timestamp 1654648307
transform 1 0 104600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4792
timestamp 1654648307
transform 1 0 106100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4874
timestamp 1654648307
transform 1 0 109100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4873
timestamp 1654648307
transform 1 0 107600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4793
timestamp 1654648307
transform 1 0 107600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4794
timestamp 1654648307
transform 1 0 109100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4876
timestamp 1654648307
transform 1 0 112100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4875
timestamp 1654648307
transform 1 0 110600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4795
timestamp 1654648307
transform 1 0 110600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4796
timestamp 1654648307
transform 1 0 112100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4878
timestamp 1654648307
transform 1 0 115100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4877
timestamp 1654648307
transform 1 0 113600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4797
timestamp 1654648307
transform 1 0 113600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4798
timestamp 1654648307
transform 1 0 115100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4879
timestamp 1654648307
transform 1 0 116600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_4799
timestamp 1654648307
transform 1 0 116600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_4640
timestamp 1654648307
transform 1 0 -1900 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4560
timestamp 1654648307
transform 1 0 -1900 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4642
timestamp 1654648307
transform 1 0 1100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4641
timestamp 1654648307
transform 1 0 -400 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4562
timestamp 1654648307
transform 1 0 1100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4561
timestamp 1654648307
transform 1 0 -400 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4644
timestamp 1654648307
transform 1 0 4100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4643
timestamp 1654648307
transform 1 0 2600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4564
timestamp 1654648307
transform 1 0 4100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4563
timestamp 1654648307
transform 1 0 2600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4646
timestamp 1654648307
transform 1 0 7100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4645
timestamp 1654648307
transform 1 0 5600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4566
timestamp 1654648307
transform 1 0 7100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4565
timestamp 1654648307
transform 1 0 5600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4648
timestamp 1654648307
transform 1 0 10100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4647
timestamp 1654648307
transform 1 0 8600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4568
timestamp 1654648307
transform 1 0 10100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4567
timestamp 1654648307
transform 1 0 8600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4650
timestamp 1654648307
transform 1 0 13100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4649
timestamp 1654648307
transform 1 0 11600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4570
timestamp 1654648307
transform 1 0 13100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4569
timestamp 1654648307
transform 1 0 11600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4652
timestamp 1654648307
transform 1 0 16100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4651
timestamp 1654648307
transform 1 0 14600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4572
timestamp 1654648307
transform 1 0 16100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4571
timestamp 1654648307
transform 1 0 14600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4654
timestamp 1654648307
transform 1 0 19100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4653
timestamp 1654648307
transform 1 0 17600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4574
timestamp 1654648307
transform 1 0 19100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4573
timestamp 1654648307
transform 1 0 17600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4656
timestamp 1654648307
transform 1 0 22100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4655
timestamp 1654648307
transform 1 0 20600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4576
timestamp 1654648307
transform 1 0 22100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4575
timestamp 1654648307
transform 1 0 20600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4658
timestamp 1654648307
transform 1 0 25100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4657
timestamp 1654648307
transform 1 0 23600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4578
timestamp 1654648307
transform 1 0 25100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4577
timestamp 1654648307
transform 1 0 23600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4660
timestamp 1654648307
transform 1 0 28100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4659
timestamp 1654648307
transform 1 0 26600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4580
timestamp 1654648307
transform 1 0 28100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4579
timestamp 1654648307
transform 1 0 26600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4662
timestamp 1654648307
transform 1 0 31100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4661
timestamp 1654648307
transform 1 0 29600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4582
timestamp 1654648307
transform 1 0 31100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4581
timestamp 1654648307
transform 1 0 29600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4664
timestamp 1654648307
transform 1 0 34100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4663
timestamp 1654648307
transform 1 0 32600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4584
timestamp 1654648307
transform 1 0 34100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4583
timestamp 1654648307
transform 1 0 32600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4666
timestamp 1654648307
transform 1 0 37100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4665
timestamp 1654648307
transform 1 0 35600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4586
timestamp 1654648307
transform 1 0 37100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4585
timestamp 1654648307
transform 1 0 35600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4668
timestamp 1654648307
transform 1 0 40100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4667
timestamp 1654648307
transform 1 0 38600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4588
timestamp 1654648307
transform 1 0 40100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4587
timestamp 1654648307
transform 1 0 38600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4670
timestamp 1654648307
transform 1 0 43100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4669
timestamp 1654648307
transform 1 0 41600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4590
timestamp 1654648307
transform 1 0 43100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4589
timestamp 1654648307
transform 1 0 41600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4672
timestamp 1654648307
transform 1 0 46100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4671
timestamp 1654648307
transform 1 0 44600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4592
timestamp 1654648307
transform 1 0 46100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4591
timestamp 1654648307
transform 1 0 44600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4674
timestamp 1654648307
transform 1 0 49100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4673
timestamp 1654648307
transform 1 0 47600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4594
timestamp 1654648307
transform 1 0 49100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4593
timestamp 1654648307
transform 1 0 47600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4676
timestamp 1654648307
transform 1 0 52100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4675
timestamp 1654648307
transform 1 0 50600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4596
timestamp 1654648307
transform 1 0 52100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4595
timestamp 1654648307
transform 1 0 50600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4678
timestamp 1654648307
transform 1 0 55100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4677
timestamp 1654648307
transform 1 0 53600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4598
timestamp 1654648307
transform 1 0 55100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4597
timestamp 1654648307
transform 1 0 53600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4680
timestamp 1654648307
transform 1 0 58100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4679
timestamp 1654648307
transform 1 0 56600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4600
timestamp 1654648307
transform 1 0 58100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4599
timestamp 1654648307
transform 1 0 56600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4682
timestamp 1654648307
transform 1 0 61100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4681
timestamp 1654648307
transform 1 0 59600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4602
timestamp 1654648307
transform 1 0 61100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4601
timestamp 1654648307
transform 1 0 59600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4683
timestamp 1654648307
transform 1 0 62600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4684
timestamp 1654648307
transform 1 0 64100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4603
timestamp 1654648307
transform 1 0 62600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4604
timestamp 1654648307
transform 1 0 64100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4685
timestamp 1654648307
transform 1 0 65600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4686
timestamp 1654648307
transform 1 0 67100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4605
timestamp 1654648307
transform 1 0 65600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4606
timestamp 1654648307
transform 1 0 67100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4687
timestamp 1654648307
transform 1 0 68600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4688
timestamp 1654648307
transform 1 0 70100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4607
timestamp 1654648307
transform 1 0 68600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4608
timestamp 1654648307
transform 1 0 70100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4689
timestamp 1654648307
transform 1 0 71600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4690
timestamp 1654648307
transform 1 0 73100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4609
timestamp 1654648307
transform 1 0 71600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4610
timestamp 1654648307
transform 1 0 73100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4691
timestamp 1654648307
transform 1 0 74600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4692
timestamp 1654648307
transform 1 0 76100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4611
timestamp 1654648307
transform 1 0 74600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4612
timestamp 1654648307
transform 1 0 76100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4693
timestamp 1654648307
transform 1 0 77600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4694
timestamp 1654648307
transform 1 0 79100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4613
timestamp 1654648307
transform 1 0 77600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4614
timestamp 1654648307
transform 1 0 79100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4695
timestamp 1654648307
transform 1 0 80600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4696
timestamp 1654648307
transform 1 0 82100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4615
timestamp 1654648307
transform 1 0 80600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4616
timestamp 1654648307
transform 1 0 82100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4697
timestamp 1654648307
transform 1 0 83600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4698
timestamp 1654648307
transform 1 0 85100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4617
timestamp 1654648307
transform 1 0 83600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4618
timestamp 1654648307
transform 1 0 85100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4699
timestamp 1654648307
transform 1 0 86600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4700
timestamp 1654648307
transform 1 0 88100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4619
timestamp 1654648307
transform 1 0 86600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4620
timestamp 1654648307
transform 1 0 88100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4701
timestamp 1654648307
transform 1 0 89600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4702
timestamp 1654648307
transform 1 0 91100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4621
timestamp 1654648307
transform 1 0 89600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4622
timestamp 1654648307
transform 1 0 91100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4703
timestamp 1654648307
transform 1 0 92600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4704
timestamp 1654648307
transform 1 0 94100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4623
timestamp 1654648307
transform 1 0 92600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4624
timestamp 1654648307
transform 1 0 94100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4705
timestamp 1654648307
transform 1 0 95600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4706
timestamp 1654648307
transform 1 0 97100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4625
timestamp 1654648307
transform 1 0 95600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4626
timestamp 1654648307
transform 1 0 97100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4707
timestamp 1654648307
transform 1 0 98600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4708
timestamp 1654648307
transform 1 0 100100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4627
timestamp 1654648307
transform 1 0 98600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4628
timestamp 1654648307
transform 1 0 100100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4709
timestamp 1654648307
transform 1 0 101600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4710
timestamp 1654648307
transform 1 0 103100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4629
timestamp 1654648307
transform 1 0 101600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4630
timestamp 1654648307
transform 1 0 103100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4711
timestamp 1654648307
transform 1 0 104600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4712
timestamp 1654648307
transform 1 0 106100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4631
timestamp 1654648307
transform 1 0 104600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4632
timestamp 1654648307
transform 1 0 106100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4713
timestamp 1654648307
transform 1 0 107600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4714
timestamp 1654648307
transform 1 0 109100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4633
timestamp 1654648307
transform 1 0 107600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4634
timestamp 1654648307
transform 1 0 109100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4715
timestamp 1654648307
transform 1 0 110600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4716
timestamp 1654648307
transform 1 0 112100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4635
timestamp 1654648307
transform 1 0 110600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4636
timestamp 1654648307
transform 1 0 112100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4717
timestamp 1654648307
transform 1 0 113600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4718
timestamp 1654648307
transform 1 0 115100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4637
timestamp 1654648307
transform 1 0 113600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4638
timestamp 1654648307
transform 1 0 115100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4719
timestamp 1654648307
transform 1 0 116600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_4639
timestamp 1654648307
transform 1 0 116600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_4480
timestamp 1654648307
transform 1 0 -1900 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4400
timestamp 1654648307
transform 1 0 -1900 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4482
timestamp 1654648307
transform 1 0 1100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4481
timestamp 1654648307
transform 1 0 -400 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4402
timestamp 1654648307
transform 1 0 1100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4401
timestamp 1654648307
transform 1 0 -400 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4484
timestamp 1654648307
transform 1 0 4100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4483
timestamp 1654648307
transform 1 0 2600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4404
timestamp 1654648307
transform 1 0 4100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4403
timestamp 1654648307
transform 1 0 2600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4486
timestamp 1654648307
transform 1 0 7100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4485
timestamp 1654648307
transform 1 0 5600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4406
timestamp 1654648307
transform 1 0 7100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4405
timestamp 1654648307
transform 1 0 5600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4488
timestamp 1654648307
transform 1 0 10100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4487
timestamp 1654648307
transform 1 0 8600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4408
timestamp 1654648307
transform 1 0 10100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4407
timestamp 1654648307
transform 1 0 8600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4490
timestamp 1654648307
transform 1 0 13100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4489
timestamp 1654648307
transform 1 0 11600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4410
timestamp 1654648307
transform 1 0 13100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4409
timestamp 1654648307
transform 1 0 11600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4492
timestamp 1654648307
transform 1 0 16100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4491
timestamp 1654648307
transform 1 0 14600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4412
timestamp 1654648307
transform 1 0 16100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4411
timestamp 1654648307
transform 1 0 14600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4494
timestamp 1654648307
transform 1 0 19100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4493
timestamp 1654648307
transform 1 0 17600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4414
timestamp 1654648307
transform 1 0 19100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4413
timestamp 1654648307
transform 1 0 17600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4496
timestamp 1654648307
transform 1 0 22100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4495
timestamp 1654648307
transform 1 0 20600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4416
timestamp 1654648307
transform 1 0 22100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4415
timestamp 1654648307
transform 1 0 20600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4498
timestamp 1654648307
transform 1 0 25100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4497
timestamp 1654648307
transform 1 0 23600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4418
timestamp 1654648307
transform 1 0 25100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4417
timestamp 1654648307
transform 1 0 23600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4500
timestamp 1654648307
transform 1 0 28100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4499
timestamp 1654648307
transform 1 0 26600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4420
timestamp 1654648307
transform 1 0 28100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4419
timestamp 1654648307
transform 1 0 26600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4502
timestamp 1654648307
transform 1 0 31100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4501
timestamp 1654648307
transform 1 0 29600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4422
timestamp 1654648307
transform 1 0 31100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4421
timestamp 1654648307
transform 1 0 29600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4504
timestamp 1654648307
transform 1 0 34100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4503
timestamp 1654648307
transform 1 0 32600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4424
timestamp 1654648307
transform 1 0 34100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4423
timestamp 1654648307
transform 1 0 32600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4506
timestamp 1654648307
transform 1 0 37100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4505
timestamp 1654648307
transform 1 0 35600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4426
timestamp 1654648307
transform 1 0 37100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4425
timestamp 1654648307
transform 1 0 35600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4508
timestamp 1654648307
transform 1 0 40100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4507
timestamp 1654648307
transform 1 0 38600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4428
timestamp 1654648307
transform 1 0 40100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4427
timestamp 1654648307
transform 1 0 38600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4510
timestamp 1654648307
transform 1 0 43100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4509
timestamp 1654648307
transform 1 0 41600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4430
timestamp 1654648307
transform 1 0 43100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4429
timestamp 1654648307
transform 1 0 41600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4512
timestamp 1654648307
transform 1 0 46100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4511
timestamp 1654648307
transform 1 0 44600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4432
timestamp 1654648307
transform 1 0 46100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4431
timestamp 1654648307
transform 1 0 44600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4514
timestamp 1654648307
transform 1 0 49100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4513
timestamp 1654648307
transform 1 0 47600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4434
timestamp 1654648307
transform 1 0 49100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4433
timestamp 1654648307
transform 1 0 47600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4516
timestamp 1654648307
transform 1 0 52100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4515
timestamp 1654648307
transform 1 0 50600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4436
timestamp 1654648307
transform 1 0 52100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4435
timestamp 1654648307
transform 1 0 50600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4518
timestamp 1654648307
transform 1 0 55100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4517
timestamp 1654648307
transform 1 0 53600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4438
timestamp 1654648307
transform 1 0 55100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4437
timestamp 1654648307
transform 1 0 53600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4520
timestamp 1654648307
transform 1 0 58100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4519
timestamp 1654648307
transform 1 0 56600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4440
timestamp 1654648307
transform 1 0 58100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4439
timestamp 1654648307
transform 1 0 56600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4522
timestamp 1654648307
transform 1 0 61100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4521
timestamp 1654648307
transform 1 0 59600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4442
timestamp 1654648307
transform 1 0 61100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4441
timestamp 1654648307
transform 1 0 59600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4523
timestamp 1654648307
transform 1 0 62600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4524
timestamp 1654648307
transform 1 0 64100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4443
timestamp 1654648307
transform 1 0 62600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4444
timestamp 1654648307
transform 1 0 64100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4525
timestamp 1654648307
transform 1 0 65600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4526
timestamp 1654648307
transform 1 0 67100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4445
timestamp 1654648307
transform 1 0 65600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4446
timestamp 1654648307
transform 1 0 67100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4527
timestamp 1654648307
transform 1 0 68600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4528
timestamp 1654648307
transform 1 0 70100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4447
timestamp 1654648307
transform 1 0 68600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4448
timestamp 1654648307
transform 1 0 70100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4529
timestamp 1654648307
transform 1 0 71600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4530
timestamp 1654648307
transform 1 0 73100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4449
timestamp 1654648307
transform 1 0 71600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4450
timestamp 1654648307
transform 1 0 73100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4531
timestamp 1654648307
transform 1 0 74600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4532
timestamp 1654648307
transform 1 0 76100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4451
timestamp 1654648307
transform 1 0 74600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4452
timestamp 1654648307
transform 1 0 76100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4533
timestamp 1654648307
transform 1 0 77600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4534
timestamp 1654648307
transform 1 0 79100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4453
timestamp 1654648307
transform 1 0 77600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4454
timestamp 1654648307
transform 1 0 79100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4535
timestamp 1654648307
transform 1 0 80600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4536
timestamp 1654648307
transform 1 0 82100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4455
timestamp 1654648307
transform 1 0 80600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4456
timestamp 1654648307
transform 1 0 82100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4537
timestamp 1654648307
transform 1 0 83600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4538
timestamp 1654648307
transform 1 0 85100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4457
timestamp 1654648307
transform 1 0 83600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4458
timestamp 1654648307
transform 1 0 85100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4539
timestamp 1654648307
transform 1 0 86600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4540
timestamp 1654648307
transform 1 0 88100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4459
timestamp 1654648307
transform 1 0 86600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4460
timestamp 1654648307
transform 1 0 88100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4541
timestamp 1654648307
transform 1 0 89600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4542
timestamp 1654648307
transform 1 0 91100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4461
timestamp 1654648307
transform 1 0 89600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4462
timestamp 1654648307
transform 1 0 91100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4543
timestamp 1654648307
transform 1 0 92600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4544
timestamp 1654648307
transform 1 0 94100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4463
timestamp 1654648307
transform 1 0 92600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4464
timestamp 1654648307
transform 1 0 94100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4545
timestamp 1654648307
transform 1 0 95600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4546
timestamp 1654648307
transform 1 0 97100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4465
timestamp 1654648307
transform 1 0 95600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4466
timestamp 1654648307
transform 1 0 97100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4547
timestamp 1654648307
transform 1 0 98600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4548
timestamp 1654648307
transform 1 0 100100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4467
timestamp 1654648307
transform 1 0 98600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4468
timestamp 1654648307
transform 1 0 100100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4549
timestamp 1654648307
transform 1 0 101600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4550
timestamp 1654648307
transform 1 0 103100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4469
timestamp 1654648307
transform 1 0 101600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4470
timestamp 1654648307
transform 1 0 103100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4551
timestamp 1654648307
transform 1 0 104600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4552
timestamp 1654648307
transform 1 0 106100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4471
timestamp 1654648307
transform 1 0 104600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4472
timestamp 1654648307
transform 1 0 106100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4553
timestamp 1654648307
transform 1 0 107600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4554
timestamp 1654648307
transform 1 0 109100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4473
timestamp 1654648307
transform 1 0 107600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4474
timestamp 1654648307
transform 1 0 109100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4555
timestamp 1654648307
transform 1 0 110600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4556
timestamp 1654648307
transform 1 0 112100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4475
timestamp 1654648307
transform 1 0 110600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4476
timestamp 1654648307
transform 1 0 112100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4557
timestamp 1654648307
transform 1 0 113600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4558
timestamp 1654648307
transform 1 0 115100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4477
timestamp 1654648307
transform 1 0 113600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4478
timestamp 1654648307
transform 1 0 115100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4559
timestamp 1654648307
transform 1 0 116600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_4479
timestamp 1654648307
transform 1 0 116600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_4320
timestamp 1654648307
transform 1 0 -1900 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4240
timestamp 1654648307
transform 1 0 -1900 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4322
timestamp 1654648307
transform 1 0 1100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4321
timestamp 1654648307
transform 1 0 -400 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4242
timestamp 1654648307
transform 1 0 1100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4241
timestamp 1654648307
transform 1 0 -400 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4324
timestamp 1654648307
transform 1 0 4100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4323
timestamp 1654648307
transform 1 0 2600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4244
timestamp 1654648307
transform 1 0 4100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4243
timestamp 1654648307
transform 1 0 2600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4326
timestamp 1654648307
transform 1 0 7100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4325
timestamp 1654648307
transform 1 0 5600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4246
timestamp 1654648307
transform 1 0 7100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4245
timestamp 1654648307
transform 1 0 5600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4328
timestamp 1654648307
transform 1 0 10100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4327
timestamp 1654648307
transform 1 0 8600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4248
timestamp 1654648307
transform 1 0 10100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4247
timestamp 1654648307
transform 1 0 8600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4330
timestamp 1654648307
transform 1 0 13100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4329
timestamp 1654648307
transform 1 0 11600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4250
timestamp 1654648307
transform 1 0 13100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4249
timestamp 1654648307
transform 1 0 11600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4332
timestamp 1654648307
transform 1 0 16100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4331
timestamp 1654648307
transform 1 0 14600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4252
timestamp 1654648307
transform 1 0 16100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4251
timestamp 1654648307
transform 1 0 14600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4334
timestamp 1654648307
transform 1 0 19100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4333
timestamp 1654648307
transform 1 0 17600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4254
timestamp 1654648307
transform 1 0 19100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4253
timestamp 1654648307
transform 1 0 17600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4336
timestamp 1654648307
transform 1 0 22100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4335
timestamp 1654648307
transform 1 0 20600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4256
timestamp 1654648307
transform 1 0 22100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4255
timestamp 1654648307
transform 1 0 20600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4338
timestamp 1654648307
transform 1 0 25100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4337
timestamp 1654648307
transform 1 0 23600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4258
timestamp 1654648307
transform 1 0 25100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4257
timestamp 1654648307
transform 1 0 23600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4340
timestamp 1654648307
transform 1 0 28100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4339
timestamp 1654648307
transform 1 0 26600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4260
timestamp 1654648307
transform 1 0 28100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4259
timestamp 1654648307
transform 1 0 26600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4342
timestamp 1654648307
transform 1 0 31100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4341
timestamp 1654648307
transform 1 0 29600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4262
timestamp 1654648307
transform 1 0 31100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4261
timestamp 1654648307
transform 1 0 29600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4344
timestamp 1654648307
transform 1 0 34100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4343
timestamp 1654648307
transform 1 0 32600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4264
timestamp 1654648307
transform 1 0 34100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4263
timestamp 1654648307
transform 1 0 32600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4346
timestamp 1654648307
transform 1 0 37100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4345
timestamp 1654648307
transform 1 0 35600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4266
timestamp 1654648307
transform 1 0 37100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4265
timestamp 1654648307
transform 1 0 35600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4348
timestamp 1654648307
transform 1 0 40100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4347
timestamp 1654648307
transform 1 0 38600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4268
timestamp 1654648307
transform 1 0 40100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4267
timestamp 1654648307
transform 1 0 38600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4350
timestamp 1654648307
transform 1 0 43100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4349
timestamp 1654648307
transform 1 0 41600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4270
timestamp 1654648307
transform 1 0 43100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4269
timestamp 1654648307
transform 1 0 41600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4352
timestamp 1654648307
transform 1 0 46100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4351
timestamp 1654648307
transform 1 0 44600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4272
timestamp 1654648307
transform 1 0 46100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4271
timestamp 1654648307
transform 1 0 44600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4354
timestamp 1654648307
transform 1 0 49100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4353
timestamp 1654648307
transform 1 0 47600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4274
timestamp 1654648307
transform 1 0 49100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4273
timestamp 1654648307
transform 1 0 47600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4356
timestamp 1654648307
transform 1 0 52100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4355
timestamp 1654648307
transform 1 0 50600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4276
timestamp 1654648307
transform 1 0 52100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4275
timestamp 1654648307
transform 1 0 50600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4358
timestamp 1654648307
transform 1 0 55100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4357
timestamp 1654648307
transform 1 0 53600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4278
timestamp 1654648307
transform 1 0 55100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4277
timestamp 1654648307
transform 1 0 53600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4360
timestamp 1654648307
transform 1 0 58100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4359
timestamp 1654648307
transform 1 0 56600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4280
timestamp 1654648307
transform 1 0 58100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4279
timestamp 1654648307
transform 1 0 56600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4362
timestamp 1654648307
transform 1 0 61100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4361
timestamp 1654648307
transform 1 0 59600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4282
timestamp 1654648307
transform 1 0 61100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4281
timestamp 1654648307
transform 1 0 59600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4363
timestamp 1654648307
transform 1 0 62600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4283
timestamp 1654648307
transform 1 0 62600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4364
timestamp 1654648307
transform 1 0 64100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4284
timestamp 1654648307
transform 1 0 64100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4365
timestamp 1654648307
transform 1 0 65600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4285
timestamp 1654648307
transform 1 0 65600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4366
timestamp 1654648307
transform 1 0 67100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4286
timestamp 1654648307
transform 1 0 67100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4367
timestamp 1654648307
transform 1 0 68600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4287
timestamp 1654648307
transform 1 0 68600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4368
timestamp 1654648307
transform 1 0 70100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4288
timestamp 1654648307
transform 1 0 70100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4369
timestamp 1654648307
transform 1 0 71600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4289
timestamp 1654648307
transform 1 0 71600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4370
timestamp 1654648307
transform 1 0 73100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4290
timestamp 1654648307
transform 1 0 73100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4371
timestamp 1654648307
transform 1 0 74600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4291
timestamp 1654648307
transform 1 0 74600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4372
timestamp 1654648307
transform 1 0 76100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4292
timestamp 1654648307
transform 1 0 76100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4373
timestamp 1654648307
transform 1 0 77600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4293
timestamp 1654648307
transform 1 0 77600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4374
timestamp 1654648307
transform 1 0 79100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4294
timestamp 1654648307
transform 1 0 79100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4375
timestamp 1654648307
transform 1 0 80600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4295
timestamp 1654648307
transform 1 0 80600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4376
timestamp 1654648307
transform 1 0 82100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4296
timestamp 1654648307
transform 1 0 82100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4377
timestamp 1654648307
transform 1 0 83600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4297
timestamp 1654648307
transform 1 0 83600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4378
timestamp 1654648307
transform 1 0 85100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4298
timestamp 1654648307
transform 1 0 85100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4379
timestamp 1654648307
transform 1 0 86600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4299
timestamp 1654648307
transform 1 0 86600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4380
timestamp 1654648307
transform 1 0 88100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4300
timestamp 1654648307
transform 1 0 88100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4381
timestamp 1654648307
transform 1 0 89600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4301
timestamp 1654648307
transform 1 0 89600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4382
timestamp 1654648307
transform 1 0 91100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4302
timestamp 1654648307
transform 1 0 91100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4383
timestamp 1654648307
transform 1 0 92600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4303
timestamp 1654648307
transform 1 0 92600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4384
timestamp 1654648307
transform 1 0 94100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4304
timestamp 1654648307
transform 1 0 94100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4385
timestamp 1654648307
transform 1 0 95600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4305
timestamp 1654648307
transform 1 0 95600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4386
timestamp 1654648307
transform 1 0 97100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4306
timestamp 1654648307
transform 1 0 97100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4387
timestamp 1654648307
transform 1 0 98600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4307
timestamp 1654648307
transform 1 0 98600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4388
timestamp 1654648307
transform 1 0 100100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4308
timestamp 1654648307
transform 1 0 100100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4389
timestamp 1654648307
transform 1 0 101600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4309
timestamp 1654648307
transform 1 0 101600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4390
timestamp 1654648307
transform 1 0 103100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4310
timestamp 1654648307
transform 1 0 103100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4391
timestamp 1654648307
transform 1 0 104600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4311
timestamp 1654648307
transform 1 0 104600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4392
timestamp 1654648307
transform 1 0 106100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4312
timestamp 1654648307
transform 1 0 106100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4393
timestamp 1654648307
transform 1 0 107600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4313
timestamp 1654648307
transform 1 0 107600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4394
timestamp 1654648307
transform 1 0 109100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4314
timestamp 1654648307
transform 1 0 109100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4395
timestamp 1654648307
transform 1 0 110600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4315
timestamp 1654648307
transform 1 0 110600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4396
timestamp 1654648307
transform 1 0 112100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4316
timestamp 1654648307
transform 1 0 112100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4397
timestamp 1654648307
transform 1 0 113600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4317
timestamp 1654648307
transform 1 0 113600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4398
timestamp 1654648307
transform 1 0 115100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4318
timestamp 1654648307
transform 1 0 115100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4399
timestamp 1654648307
transform 1 0 116600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_4319
timestamp 1654648307
transform 1 0 116600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_4160
timestamp 1654648307
transform 1 0 -1900 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4080
timestamp 1654648307
transform 1 0 -1900 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4162
timestamp 1654648307
transform 1 0 1100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4161
timestamp 1654648307
transform 1 0 -400 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4082
timestamp 1654648307
transform 1 0 1100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4081
timestamp 1654648307
transform 1 0 -400 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4164
timestamp 1654648307
transform 1 0 4100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4163
timestamp 1654648307
transform 1 0 2600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4084
timestamp 1654648307
transform 1 0 4100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4083
timestamp 1654648307
transform 1 0 2600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4166
timestamp 1654648307
transform 1 0 7100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4165
timestamp 1654648307
transform 1 0 5600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4086
timestamp 1654648307
transform 1 0 7100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4085
timestamp 1654648307
transform 1 0 5600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4168
timestamp 1654648307
transform 1 0 10100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4167
timestamp 1654648307
transform 1 0 8600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4088
timestamp 1654648307
transform 1 0 10100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4087
timestamp 1654648307
transform 1 0 8600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4170
timestamp 1654648307
transform 1 0 13100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4169
timestamp 1654648307
transform 1 0 11600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4090
timestamp 1654648307
transform 1 0 13100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4089
timestamp 1654648307
transform 1 0 11600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4172
timestamp 1654648307
transform 1 0 16100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4171
timestamp 1654648307
transform 1 0 14600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4092
timestamp 1654648307
transform 1 0 16100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4091
timestamp 1654648307
transform 1 0 14600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4174
timestamp 1654648307
transform 1 0 19100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4173
timestamp 1654648307
transform 1 0 17600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4094
timestamp 1654648307
transform 1 0 19100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4093
timestamp 1654648307
transform 1 0 17600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4176
timestamp 1654648307
transform 1 0 22100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4175
timestamp 1654648307
transform 1 0 20600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4096
timestamp 1654648307
transform 1 0 22100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4095
timestamp 1654648307
transform 1 0 20600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4178
timestamp 1654648307
transform 1 0 25100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4177
timestamp 1654648307
transform 1 0 23600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4098
timestamp 1654648307
transform 1 0 25100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4097
timestamp 1654648307
transform 1 0 23600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4180
timestamp 1654648307
transform 1 0 28100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4179
timestamp 1654648307
transform 1 0 26600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4100
timestamp 1654648307
transform 1 0 28100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4099
timestamp 1654648307
transform 1 0 26600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4182
timestamp 1654648307
transform 1 0 31100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4181
timestamp 1654648307
transform 1 0 29600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4102
timestamp 1654648307
transform 1 0 31100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4101
timestamp 1654648307
transform 1 0 29600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4184
timestamp 1654648307
transform 1 0 34100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4183
timestamp 1654648307
transform 1 0 32600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4104
timestamp 1654648307
transform 1 0 34100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4103
timestamp 1654648307
transform 1 0 32600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4186
timestamp 1654648307
transform 1 0 37100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4185
timestamp 1654648307
transform 1 0 35600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4106
timestamp 1654648307
transform 1 0 37100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4105
timestamp 1654648307
transform 1 0 35600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4188
timestamp 1654648307
transform 1 0 40100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4187
timestamp 1654648307
transform 1 0 38600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4108
timestamp 1654648307
transform 1 0 40100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4107
timestamp 1654648307
transform 1 0 38600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4190
timestamp 1654648307
transform 1 0 43100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4189
timestamp 1654648307
transform 1 0 41600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4110
timestamp 1654648307
transform 1 0 43100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4109
timestamp 1654648307
transform 1 0 41600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4192
timestamp 1654648307
transform 1 0 46100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4191
timestamp 1654648307
transform 1 0 44600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4112
timestamp 1654648307
transform 1 0 46100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4111
timestamp 1654648307
transform 1 0 44600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4194
timestamp 1654648307
transform 1 0 49100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4193
timestamp 1654648307
transform 1 0 47600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4114
timestamp 1654648307
transform 1 0 49100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4113
timestamp 1654648307
transform 1 0 47600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4196
timestamp 1654648307
transform 1 0 52100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4195
timestamp 1654648307
transform 1 0 50600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4116
timestamp 1654648307
transform 1 0 52100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4115
timestamp 1654648307
transform 1 0 50600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4198
timestamp 1654648307
transform 1 0 55100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4197
timestamp 1654648307
transform 1 0 53600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4118
timestamp 1654648307
transform 1 0 55100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4117
timestamp 1654648307
transform 1 0 53600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4200
timestamp 1654648307
transform 1 0 58100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4199
timestamp 1654648307
transform 1 0 56600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4120
timestamp 1654648307
transform 1 0 58100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4119
timestamp 1654648307
transform 1 0 56600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4202
timestamp 1654648307
transform 1 0 61100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4201
timestamp 1654648307
transform 1 0 59600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4122
timestamp 1654648307
transform 1 0 61100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4121
timestamp 1654648307
transform 1 0 59600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4203
timestamp 1654648307
transform 1 0 62600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4123
timestamp 1654648307
transform 1 0 62600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4204
timestamp 1654648307
transform 1 0 64100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4124
timestamp 1654648307
transform 1 0 64100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4205
timestamp 1654648307
transform 1 0 65600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4125
timestamp 1654648307
transform 1 0 65600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4206
timestamp 1654648307
transform 1 0 67100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4126
timestamp 1654648307
transform 1 0 67100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4207
timestamp 1654648307
transform 1 0 68600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4127
timestamp 1654648307
transform 1 0 68600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4208
timestamp 1654648307
transform 1 0 70100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4128
timestamp 1654648307
transform 1 0 70100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4209
timestamp 1654648307
transform 1 0 71600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4129
timestamp 1654648307
transform 1 0 71600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4210
timestamp 1654648307
transform 1 0 73100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4130
timestamp 1654648307
transform 1 0 73100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4211
timestamp 1654648307
transform 1 0 74600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4131
timestamp 1654648307
transform 1 0 74600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4212
timestamp 1654648307
transform 1 0 76100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4132
timestamp 1654648307
transform 1 0 76100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4213
timestamp 1654648307
transform 1 0 77600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4133
timestamp 1654648307
transform 1 0 77600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4214
timestamp 1654648307
transform 1 0 79100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4134
timestamp 1654648307
transform 1 0 79100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4215
timestamp 1654648307
transform 1 0 80600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4135
timestamp 1654648307
transform 1 0 80600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4216
timestamp 1654648307
transform 1 0 82100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4136
timestamp 1654648307
transform 1 0 82100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4217
timestamp 1654648307
transform 1 0 83600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4137
timestamp 1654648307
transform 1 0 83600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4218
timestamp 1654648307
transform 1 0 85100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4138
timestamp 1654648307
transform 1 0 85100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4219
timestamp 1654648307
transform 1 0 86600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4139
timestamp 1654648307
transform 1 0 86600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4220
timestamp 1654648307
transform 1 0 88100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4140
timestamp 1654648307
transform 1 0 88100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4221
timestamp 1654648307
transform 1 0 89600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4141
timestamp 1654648307
transform 1 0 89600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4222
timestamp 1654648307
transform 1 0 91100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4142
timestamp 1654648307
transform 1 0 91100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4223
timestamp 1654648307
transform 1 0 92600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4143
timestamp 1654648307
transform 1 0 92600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4224
timestamp 1654648307
transform 1 0 94100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4144
timestamp 1654648307
transform 1 0 94100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4225
timestamp 1654648307
transform 1 0 95600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4145
timestamp 1654648307
transform 1 0 95600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4226
timestamp 1654648307
transform 1 0 97100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4146
timestamp 1654648307
transform 1 0 97100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4227
timestamp 1654648307
transform 1 0 98600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4147
timestamp 1654648307
transform 1 0 98600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4228
timestamp 1654648307
transform 1 0 100100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4148
timestamp 1654648307
transform 1 0 100100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4229
timestamp 1654648307
transform 1 0 101600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4149
timestamp 1654648307
transform 1 0 101600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4230
timestamp 1654648307
transform 1 0 103100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4150
timestamp 1654648307
transform 1 0 103100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4231
timestamp 1654648307
transform 1 0 104600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4151
timestamp 1654648307
transform 1 0 104600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4232
timestamp 1654648307
transform 1 0 106100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4152
timestamp 1654648307
transform 1 0 106100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4233
timestamp 1654648307
transform 1 0 107600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4153
timestamp 1654648307
transform 1 0 107600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4234
timestamp 1654648307
transform 1 0 109100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4154
timestamp 1654648307
transform 1 0 109100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4235
timestamp 1654648307
transform 1 0 110600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4155
timestamp 1654648307
transform 1 0 110600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4236
timestamp 1654648307
transform 1 0 112100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4156
timestamp 1654648307
transform 1 0 112100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4237
timestamp 1654648307
transform 1 0 113600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4157
timestamp 1654648307
transform 1 0 113600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4238
timestamp 1654648307
transform 1 0 115100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4158
timestamp 1654648307
transform 1 0 115100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4239
timestamp 1654648307
transform 1 0 116600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_4159
timestamp 1654648307
transform 1 0 116600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_4000
timestamp 1654648307
transform 1 0 -1900 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3920
timestamp 1654648307
transform 1 0 -1900 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4002
timestamp 1654648307
transform 1 0 1100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_4001
timestamp 1654648307
transform 1 0 -400 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3922
timestamp 1654648307
transform 1 0 1100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_3921
timestamp 1654648307
transform 1 0 -400 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4004
timestamp 1654648307
transform 1 0 4100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_4003
timestamp 1654648307
transform 1 0 2600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3924
timestamp 1654648307
transform 1 0 4100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_3923
timestamp 1654648307
transform 1 0 2600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4006
timestamp 1654648307
transform 1 0 7100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_4005
timestamp 1654648307
transform 1 0 5600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3926
timestamp 1654648307
transform 1 0 7100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_3925
timestamp 1654648307
transform 1 0 5600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4008
timestamp 1654648307
transform 1 0 10100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_4007
timestamp 1654648307
transform 1 0 8600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3928
timestamp 1654648307
transform 1 0 10100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_3927
timestamp 1654648307
transform 1 0 8600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4010
timestamp 1654648307
transform 1 0 13100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_4009
timestamp 1654648307
transform 1 0 11600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3930
timestamp 1654648307
transform 1 0 13100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_3929
timestamp 1654648307
transform 1 0 11600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4012
timestamp 1654648307
transform 1 0 16100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_4011
timestamp 1654648307
transform 1 0 14600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3932
timestamp 1654648307
transform 1 0 16100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_3931
timestamp 1654648307
transform 1 0 14600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4014
timestamp 1654648307
transform 1 0 19100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_4013
timestamp 1654648307
transform 1 0 17600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3934
timestamp 1654648307
transform 1 0 19100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_3933
timestamp 1654648307
transform 1 0 17600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4016
timestamp 1654648307
transform 1 0 22100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_4015
timestamp 1654648307
transform 1 0 20600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3936
timestamp 1654648307
transform 1 0 22100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_3935
timestamp 1654648307
transform 1 0 20600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4018
timestamp 1654648307
transform 1 0 25100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_4017
timestamp 1654648307
transform 1 0 23600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3938
timestamp 1654648307
transform 1 0 25100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_3937
timestamp 1654648307
transform 1 0 23600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4020
timestamp 1654648307
transform 1 0 28100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_4019
timestamp 1654648307
transform 1 0 26600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3940
timestamp 1654648307
transform 1 0 28100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_3939
timestamp 1654648307
transform 1 0 26600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4022
timestamp 1654648307
transform 1 0 31100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_4021
timestamp 1654648307
transform 1 0 29600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3942
timestamp 1654648307
transform 1 0 31100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_3941
timestamp 1654648307
transform 1 0 29600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4024
timestamp 1654648307
transform 1 0 34100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_4023
timestamp 1654648307
transform 1 0 32600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3944
timestamp 1654648307
transform 1 0 34100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_3943
timestamp 1654648307
transform 1 0 32600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4026
timestamp 1654648307
transform 1 0 37100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_4025
timestamp 1654648307
transform 1 0 35600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3946
timestamp 1654648307
transform 1 0 37100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_3945
timestamp 1654648307
transform 1 0 35600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4028
timestamp 1654648307
transform 1 0 40100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_4027
timestamp 1654648307
transform 1 0 38600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3948
timestamp 1654648307
transform 1 0 40100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_3947
timestamp 1654648307
transform 1 0 38600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4030
timestamp 1654648307
transform 1 0 43100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_4029
timestamp 1654648307
transform 1 0 41600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3950
timestamp 1654648307
transform 1 0 43100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_3949
timestamp 1654648307
transform 1 0 41600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4032
timestamp 1654648307
transform 1 0 46100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_4031
timestamp 1654648307
transform 1 0 44600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3952
timestamp 1654648307
transform 1 0 46100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_3951
timestamp 1654648307
transform 1 0 44600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4034
timestamp 1654648307
transform 1 0 49100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_4033
timestamp 1654648307
transform 1 0 47600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3954
timestamp 1654648307
transform 1 0 49100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_3953
timestamp 1654648307
transform 1 0 47600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4036
timestamp 1654648307
transform 1 0 52100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_4035
timestamp 1654648307
transform 1 0 50600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3956
timestamp 1654648307
transform 1 0 52100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_3955
timestamp 1654648307
transform 1 0 50600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4038
timestamp 1654648307
transform 1 0 55100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_4037
timestamp 1654648307
transform 1 0 53600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3958
timestamp 1654648307
transform 1 0 55100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_3957
timestamp 1654648307
transform 1 0 53600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4040
timestamp 1654648307
transform 1 0 58100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_4039
timestamp 1654648307
transform 1 0 56600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3960
timestamp 1654648307
transform 1 0 58100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_3959
timestamp 1654648307
transform 1 0 56600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4042
timestamp 1654648307
transform 1 0 61100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_4041
timestamp 1654648307
transform 1 0 59600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3962
timestamp 1654648307
transform 1 0 61100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_3961
timestamp 1654648307
transform 1 0 59600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4043
timestamp 1654648307
transform 1 0 62600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3963
timestamp 1654648307
transform 1 0 62600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4044
timestamp 1654648307
transform 1 0 64100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3964
timestamp 1654648307
transform 1 0 64100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4045
timestamp 1654648307
transform 1 0 65600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3965
timestamp 1654648307
transform 1 0 65600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4046
timestamp 1654648307
transform 1 0 67100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3966
timestamp 1654648307
transform 1 0 67100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4047
timestamp 1654648307
transform 1 0 68600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3967
timestamp 1654648307
transform 1 0 68600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4048
timestamp 1654648307
transform 1 0 70100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3968
timestamp 1654648307
transform 1 0 70100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4049
timestamp 1654648307
transform 1 0 71600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3969
timestamp 1654648307
transform 1 0 71600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4050
timestamp 1654648307
transform 1 0 73100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3970
timestamp 1654648307
transform 1 0 73100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4051
timestamp 1654648307
transform 1 0 74600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3971
timestamp 1654648307
transform 1 0 74600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4052
timestamp 1654648307
transform 1 0 76100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3972
timestamp 1654648307
transform 1 0 76100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4053
timestamp 1654648307
transform 1 0 77600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3973
timestamp 1654648307
transform 1 0 77600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4054
timestamp 1654648307
transform 1 0 79100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3974
timestamp 1654648307
transform 1 0 79100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4055
timestamp 1654648307
transform 1 0 80600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3975
timestamp 1654648307
transform 1 0 80600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4056
timestamp 1654648307
transform 1 0 82100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3976
timestamp 1654648307
transform 1 0 82100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4057
timestamp 1654648307
transform 1 0 83600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3977
timestamp 1654648307
transform 1 0 83600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4058
timestamp 1654648307
transform 1 0 85100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3978
timestamp 1654648307
transform 1 0 85100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4059
timestamp 1654648307
transform 1 0 86600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3979
timestamp 1654648307
transform 1 0 86600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4060
timestamp 1654648307
transform 1 0 88100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3980
timestamp 1654648307
transform 1 0 88100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4061
timestamp 1654648307
transform 1 0 89600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3981
timestamp 1654648307
transform 1 0 89600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4062
timestamp 1654648307
transform 1 0 91100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3982
timestamp 1654648307
transform 1 0 91100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4063
timestamp 1654648307
transform 1 0 92600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3983
timestamp 1654648307
transform 1 0 92600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4064
timestamp 1654648307
transform 1 0 94100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3984
timestamp 1654648307
transform 1 0 94100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4065
timestamp 1654648307
transform 1 0 95600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3985
timestamp 1654648307
transform 1 0 95600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4066
timestamp 1654648307
transform 1 0 97100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3986
timestamp 1654648307
transform 1 0 97100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4067
timestamp 1654648307
transform 1 0 98600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3987
timestamp 1654648307
transform 1 0 98600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4068
timestamp 1654648307
transform 1 0 100100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3988
timestamp 1654648307
transform 1 0 100100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4069
timestamp 1654648307
transform 1 0 101600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3989
timestamp 1654648307
transform 1 0 101600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4070
timestamp 1654648307
transform 1 0 103100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3990
timestamp 1654648307
transform 1 0 103100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4071
timestamp 1654648307
transform 1 0 104600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3991
timestamp 1654648307
transform 1 0 104600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4072
timestamp 1654648307
transform 1 0 106100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3992
timestamp 1654648307
transform 1 0 106100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4073
timestamp 1654648307
transform 1 0 107600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3993
timestamp 1654648307
transform 1 0 107600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4074
timestamp 1654648307
transform 1 0 109100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3994
timestamp 1654648307
transform 1 0 109100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4075
timestamp 1654648307
transform 1 0 110600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3995
timestamp 1654648307
transform 1 0 110600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4076
timestamp 1654648307
transform 1 0 112100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3996
timestamp 1654648307
transform 1 0 112100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4077
timestamp 1654648307
transform 1 0 113600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3997
timestamp 1654648307
transform 1 0 113600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4078
timestamp 1654648307
transform 1 0 115100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3998
timestamp 1654648307
transform 1 0 115100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4079
timestamp 1654648307
transform 1 0 116600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_3999
timestamp 1654648307
transform 1 0 116600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_3840
timestamp 1654648307
transform 1 0 -1900 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3760
timestamp 1654648307
transform 1 0 -1900 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3842
timestamp 1654648307
transform 1 0 1100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3841
timestamp 1654648307
transform 1 0 -400 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3762
timestamp 1654648307
transform 1 0 1100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3761
timestamp 1654648307
transform 1 0 -400 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3844
timestamp 1654648307
transform 1 0 4100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3843
timestamp 1654648307
transform 1 0 2600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3764
timestamp 1654648307
transform 1 0 4100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3763
timestamp 1654648307
transform 1 0 2600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3846
timestamp 1654648307
transform 1 0 7100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3845
timestamp 1654648307
transform 1 0 5600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3766
timestamp 1654648307
transform 1 0 7100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3765
timestamp 1654648307
transform 1 0 5600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3848
timestamp 1654648307
transform 1 0 10100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3847
timestamp 1654648307
transform 1 0 8600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3768
timestamp 1654648307
transform 1 0 10100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3767
timestamp 1654648307
transform 1 0 8600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3850
timestamp 1654648307
transform 1 0 13100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3849
timestamp 1654648307
transform 1 0 11600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3770
timestamp 1654648307
transform 1 0 13100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3769
timestamp 1654648307
transform 1 0 11600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3852
timestamp 1654648307
transform 1 0 16100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3851
timestamp 1654648307
transform 1 0 14600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3772
timestamp 1654648307
transform 1 0 16100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3771
timestamp 1654648307
transform 1 0 14600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3854
timestamp 1654648307
transform 1 0 19100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3853
timestamp 1654648307
transform 1 0 17600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3774
timestamp 1654648307
transform 1 0 19100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3773
timestamp 1654648307
transform 1 0 17600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3856
timestamp 1654648307
transform 1 0 22100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3855
timestamp 1654648307
transform 1 0 20600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3776
timestamp 1654648307
transform 1 0 22100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3775
timestamp 1654648307
transform 1 0 20600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3858
timestamp 1654648307
transform 1 0 25100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3857
timestamp 1654648307
transform 1 0 23600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3778
timestamp 1654648307
transform 1 0 25100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3777
timestamp 1654648307
transform 1 0 23600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3860
timestamp 1654648307
transform 1 0 28100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3859
timestamp 1654648307
transform 1 0 26600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3780
timestamp 1654648307
transform 1 0 28100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3779
timestamp 1654648307
transform 1 0 26600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3862
timestamp 1654648307
transform 1 0 31100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3861
timestamp 1654648307
transform 1 0 29600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3782
timestamp 1654648307
transform 1 0 31100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3781
timestamp 1654648307
transform 1 0 29600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3864
timestamp 1654648307
transform 1 0 34100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3863
timestamp 1654648307
transform 1 0 32600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3784
timestamp 1654648307
transform 1 0 34100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3783
timestamp 1654648307
transform 1 0 32600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3866
timestamp 1654648307
transform 1 0 37100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3865
timestamp 1654648307
transform 1 0 35600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3786
timestamp 1654648307
transform 1 0 37100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3785
timestamp 1654648307
transform 1 0 35600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3868
timestamp 1654648307
transform 1 0 40100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3867
timestamp 1654648307
transform 1 0 38600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3788
timestamp 1654648307
transform 1 0 40100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3787
timestamp 1654648307
transform 1 0 38600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3870
timestamp 1654648307
transform 1 0 43100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3869
timestamp 1654648307
transform 1 0 41600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3790
timestamp 1654648307
transform 1 0 43100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3789
timestamp 1654648307
transform 1 0 41600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3872
timestamp 1654648307
transform 1 0 46100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3871
timestamp 1654648307
transform 1 0 44600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3792
timestamp 1654648307
transform 1 0 46100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3791
timestamp 1654648307
transform 1 0 44600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3874
timestamp 1654648307
transform 1 0 49100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3873
timestamp 1654648307
transform 1 0 47600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3794
timestamp 1654648307
transform 1 0 49100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3793
timestamp 1654648307
transform 1 0 47600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3876
timestamp 1654648307
transform 1 0 52100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3875
timestamp 1654648307
transform 1 0 50600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3796
timestamp 1654648307
transform 1 0 52100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3795
timestamp 1654648307
transform 1 0 50600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3878
timestamp 1654648307
transform 1 0 55100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3877
timestamp 1654648307
transform 1 0 53600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3798
timestamp 1654648307
transform 1 0 55100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3797
timestamp 1654648307
transform 1 0 53600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3880
timestamp 1654648307
transform 1 0 58100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3879
timestamp 1654648307
transform 1 0 56600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3800
timestamp 1654648307
transform 1 0 58100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3799
timestamp 1654648307
transform 1 0 56600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3882
timestamp 1654648307
transform 1 0 61100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3881
timestamp 1654648307
transform 1 0 59600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3802
timestamp 1654648307
transform 1 0 61100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3801
timestamp 1654648307
transform 1 0 59600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3883
timestamp 1654648307
transform 1 0 62600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3803
timestamp 1654648307
transform 1 0 62600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3884
timestamp 1654648307
transform 1 0 64100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3804
timestamp 1654648307
transform 1 0 64100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3885
timestamp 1654648307
transform 1 0 65600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3805
timestamp 1654648307
transform 1 0 65600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3886
timestamp 1654648307
transform 1 0 67100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3806
timestamp 1654648307
transform 1 0 67100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3887
timestamp 1654648307
transform 1 0 68600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3807
timestamp 1654648307
transform 1 0 68600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3888
timestamp 1654648307
transform 1 0 70100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3808
timestamp 1654648307
transform 1 0 70100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3889
timestamp 1654648307
transform 1 0 71600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3809
timestamp 1654648307
transform 1 0 71600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3890
timestamp 1654648307
transform 1 0 73100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3810
timestamp 1654648307
transform 1 0 73100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3891
timestamp 1654648307
transform 1 0 74600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3811
timestamp 1654648307
transform 1 0 74600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3892
timestamp 1654648307
transform 1 0 76100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3812
timestamp 1654648307
transform 1 0 76100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3893
timestamp 1654648307
transform 1 0 77600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3813
timestamp 1654648307
transform 1 0 77600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3894
timestamp 1654648307
transform 1 0 79100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3814
timestamp 1654648307
transform 1 0 79100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3895
timestamp 1654648307
transform 1 0 80600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3815
timestamp 1654648307
transform 1 0 80600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3896
timestamp 1654648307
transform 1 0 82100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3816
timestamp 1654648307
transform 1 0 82100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3897
timestamp 1654648307
transform 1 0 83600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3817
timestamp 1654648307
transform 1 0 83600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3898
timestamp 1654648307
transform 1 0 85100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3818
timestamp 1654648307
transform 1 0 85100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3899
timestamp 1654648307
transform 1 0 86600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3819
timestamp 1654648307
transform 1 0 86600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3900
timestamp 1654648307
transform 1 0 88100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3820
timestamp 1654648307
transform 1 0 88100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3901
timestamp 1654648307
transform 1 0 89600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3821
timestamp 1654648307
transform 1 0 89600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3902
timestamp 1654648307
transform 1 0 91100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3822
timestamp 1654648307
transform 1 0 91100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3903
timestamp 1654648307
transform 1 0 92600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3823
timestamp 1654648307
transform 1 0 92600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3904
timestamp 1654648307
transform 1 0 94100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3824
timestamp 1654648307
transform 1 0 94100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3905
timestamp 1654648307
transform 1 0 95600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3825
timestamp 1654648307
transform 1 0 95600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3906
timestamp 1654648307
transform 1 0 97100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3826
timestamp 1654648307
transform 1 0 97100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3907
timestamp 1654648307
transform 1 0 98600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3827
timestamp 1654648307
transform 1 0 98600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3908
timestamp 1654648307
transform 1 0 100100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3828
timestamp 1654648307
transform 1 0 100100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3909
timestamp 1654648307
transform 1 0 101600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3829
timestamp 1654648307
transform 1 0 101600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3910
timestamp 1654648307
transform 1 0 103100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3830
timestamp 1654648307
transform 1 0 103100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3911
timestamp 1654648307
transform 1 0 104600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3831
timestamp 1654648307
transform 1 0 104600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3912
timestamp 1654648307
transform 1 0 106100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3832
timestamp 1654648307
transform 1 0 106100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3913
timestamp 1654648307
transform 1 0 107600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3833
timestamp 1654648307
transform 1 0 107600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3914
timestamp 1654648307
transform 1 0 109100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3834
timestamp 1654648307
transform 1 0 109100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3915
timestamp 1654648307
transform 1 0 110600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3835
timestamp 1654648307
transform 1 0 110600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3916
timestamp 1654648307
transform 1 0 112100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3836
timestamp 1654648307
transform 1 0 112100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3917
timestamp 1654648307
transform 1 0 113600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3837
timestamp 1654648307
transform 1 0 113600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3918
timestamp 1654648307
transform 1 0 115100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3838
timestamp 1654648307
transform 1 0 115100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3919
timestamp 1654648307
transform 1 0 116600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_3839
timestamp 1654648307
transform 1 0 116600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_3680
timestamp 1654648307
transform 1 0 -1900 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3600
timestamp 1654648307
transform 1 0 -1900 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3682
timestamp 1654648307
transform 1 0 1100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3681
timestamp 1654648307
transform 1 0 -400 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3602
timestamp 1654648307
transform 1 0 1100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3601
timestamp 1654648307
transform 1 0 -400 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3684
timestamp 1654648307
transform 1 0 4100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3683
timestamp 1654648307
transform 1 0 2600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3604
timestamp 1654648307
transform 1 0 4100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3603
timestamp 1654648307
transform 1 0 2600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3686
timestamp 1654648307
transform 1 0 7100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3685
timestamp 1654648307
transform 1 0 5600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3606
timestamp 1654648307
transform 1 0 7100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3605
timestamp 1654648307
transform 1 0 5600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3688
timestamp 1654648307
transform 1 0 10100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3687
timestamp 1654648307
transform 1 0 8600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3608
timestamp 1654648307
transform 1 0 10100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3607
timestamp 1654648307
transform 1 0 8600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3690
timestamp 1654648307
transform 1 0 13100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3689
timestamp 1654648307
transform 1 0 11600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3610
timestamp 1654648307
transform 1 0 13100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3609
timestamp 1654648307
transform 1 0 11600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3692
timestamp 1654648307
transform 1 0 16100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3691
timestamp 1654648307
transform 1 0 14600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3612
timestamp 1654648307
transform 1 0 16100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3611
timestamp 1654648307
transform 1 0 14600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3694
timestamp 1654648307
transform 1 0 19100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3693
timestamp 1654648307
transform 1 0 17600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3614
timestamp 1654648307
transform 1 0 19100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3613
timestamp 1654648307
transform 1 0 17600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3696
timestamp 1654648307
transform 1 0 22100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3695
timestamp 1654648307
transform 1 0 20600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3616
timestamp 1654648307
transform 1 0 22100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3615
timestamp 1654648307
transform 1 0 20600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3698
timestamp 1654648307
transform 1 0 25100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3697
timestamp 1654648307
transform 1 0 23600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3618
timestamp 1654648307
transform 1 0 25100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3617
timestamp 1654648307
transform 1 0 23600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3700
timestamp 1654648307
transform 1 0 28100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3699
timestamp 1654648307
transform 1 0 26600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3620
timestamp 1654648307
transform 1 0 28100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3619
timestamp 1654648307
transform 1 0 26600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3702
timestamp 1654648307
transform 1 0 31100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3701
timestamp 1654648307
transform 1 0 29600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3622
timestamp 1654648307
transform 1 0 31100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3621
timestamp 1654648307
transform 1 0 29600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3704
timestamp 1654648307
transform 1 0 34100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3703
timestamp 1654648307
transform 1 0 32600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3624
timestamp 1654648307
transform 1 0 34100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3623
timestamp 1654648307
transform 1 0 32600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3706
timestamp 1654648307
transform 1 0 37100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3705
timestamp 1654648307
transform 1 0 35600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3626
timestamp 1654648307
transform 1 0 37100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3625
timestamp 1654648307
transform 1 0 35600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3708
timestamp 1654648307
transform 1 0 40100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3707
timestamp 1654648307
transform 1 0 38600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3628
timestamp 1654648307
transform 1 0 40100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3627
timestamp 1654648307
transform 1 0 38600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3710
timestamp 1654648307
transform 1 0 43100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3709
timestamp 1654648307
transform 1 0 41600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3630
timestamp 1654648307
transform 1 0 43100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3629
timestamp 1654648307
transform 1 0 41600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3712
timestamp 1654648307
transform 1 0 46100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3711
timestamp 1654648307
transform 1 0 44600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3632
timestamp 1654648307
transform 1 0 46100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3631
timestamp 1654648307
transform 1 0 44600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3714
timestamp 1654648307
transform 1 0 49100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3713
timestamp 1654648307
transform 1 0 47600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3634
timestamp 1654648307
transform 1 0 49100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3633
timestamp 1654648307
transform 1 0 47600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3716
timestamp 1654648307
transform 1 0 52100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3715
timestamp 1654648307
transform 1 0 50600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3636
timestamp 1654648307
transform 1 0 52100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3635
timestamp 1654648307
transform 1 0 50600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3718
timestamp 1654648307
transform 1 0 55100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3717
timestamp 1654648307
transform 1 0 53600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3638
timestamp 1654648307
transform 1 0 55100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3637
timestamp 1654648307
transform 1 0 53600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3720
timestamp 1654648307
transform 1 0 58100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3719
timestamp 1654648307
transform 1 0 56600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3640
timestamp 1654648307
transform 1 0 58100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3639
timestamp 1654648307
transform 1 0 56600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3722
timestamp 1654648307
transform 1 0 61100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3721
timestamp 1654648307
transform 1 0 59600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3642
timestamp 1654648307
transform 1 0 61100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3641
timestamp 1654648307
transform 1 0 59600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3723
timestamp 1654648307
transform 1 0 62600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3643
timestamp 1654648307
transform 1 0 62600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3724
timestamp 1654648307
transform 1 0 64100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3644
timestamp 1654648307
transform 1 0 64100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3725
timestamp 1654648307
transform 1 0 65600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3645
timestamp 1654648307
transform 1 0 65600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3726
timestamp 1654648307
transform 1 0 67100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3646
timestamp 1654648307
transform 1 0 67100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3727
timestamp 1654648307
transform 1 0 68600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3647
timestamp 1654648307
transform 1 0 68600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3728
timestamp 1654648307
transform 1 0 70100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3648
timestamp 1654648307
transform 1 0 70100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3729
timestamp 1654648307
transform 1 0 71600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3649
timestamp 1654648307
transform 1 0 71600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3730
timestamp 1654648307
transform 1 0 73100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3650
timestamp 1654648307
transform 1 0 73100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3731
timestamp 1654648307
transform 1 0 74600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3651
timestamp 1654648307
transform 1 0 74600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3732
timestamp 1654648307
transform 1 0 76100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3652
timestamp 1654648307
transform 1 0 76100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3733
timestamp 1654648307
transform 1 0 77600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3653
timestamp 1654648307
transform 1 0 77600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3734
timestamp 1654648307
transform 1 0 79100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3654
timestamp 1654648307
transform 1 0 79100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3735
timestamp 1654648307
transform 1 0 80600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3655
timestamp 1654648307
transform 1 0 80600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3736
timestamp 1654648307
transform 1 0 82100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3656
timestamp 1654648307
transform 1 0 82100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3737
timestamp 1654648307
transform 1 0 83600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3657
timestamp 1654648307
transform 1 0 83600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3738
timestamp 1654648307
transform 1 0 85100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3658
timestamp 1654648307
transform 1 0 85100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3739
timestamp 1654648307
transform 1 0 86600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3659
timestamp 1654648307
transform 1 0 86600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3740
timestamp 1654648307
transform 1 0 88100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3660
timestamp 1654648307
transform 1 0 88100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3741
timestamp 1654648307
transform 1 0 89600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3661
timestamp 1654648307
transform 1 0 89600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3742
timestamp 1654648307
transform 1 0 91100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3662
timestamp 1654648307
transform 1 0 91100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3743
timestamp 1654648307
transform 1 0 92600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3663
timestamp 1654648307
transform 1 0 92600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3744
timestamp 1654648307
transform 1 0 94100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3664
timestamp 1654648307
transform 1 0 94100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3745
timestamp 1654648307
transform 1 0 95600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3665
timestamp 1654648307
transform 1 0 95600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3746
timestamp 1654648307
transform 1 0 97100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3666
timestamp 1654648307
transform 1 0 97100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3747
timestamp 1654648307
transform 1 0 98600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3667
timestamp 1654648307
transform 1 0 98600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3748
timestamp 1654648307
transform 1 0 100100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3668
timestamp 1654648307
transform 1 0 100100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3749
timestamp 1654648307
transform 1 0 101600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3669
timestamp 1654648307
transform 1 0 101600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3750
timestamp 1654648307
transform 1 0 103100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3670
timestamp 1654648307
transform 1 0 103100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3751
timestamp 1654648307
transform 1 0 104600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3671
timestamp 1654648307
transform 1 0 104600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3752
timestamp 1654648307
transform 1 0 106100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3672
timestamp 1654648307
transform 1 0 106100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3753
timestamp 1654648307
transform 1 0 107600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3673
timestamp 1654648307
transform 1 0 107600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3754
timestamp 1654648307
transform 1 0 109100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3674
timestamp 1654648307
transform 1 0 109100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3755
timestamp 1654648307
transform 1 0 110600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3675
timestamp 1654648307
transform 1 0 110600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3756
timestamp 1654648307
transform 1 0 112100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3676
timestamp 1654648307
transform 1 0 112100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3757
timestamp 1654648307
transform 1 0 113600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3677
timestamp 1654648307
transform 1 0 113600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3758
timestamp 1654648307
transform 1 0 115100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3678
timestamp 1654648307
transform 1 0 115100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3759
timestamp 1654648307
transform 1 0 116600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_3679
timestamp 1654648307
transform 1 0 116600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_3520
timestamp 1654648307
transform 1 0 -1900 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3440
timestamp 1654648307
transform 1 0 -1900 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3522
timestamp 1654648307
transform 1 0 1100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3521
timestamp 1654648307
transform 1 0 -400 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3442
timestamp 1654648307
transform 1 0 1100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3441
timestamp 1654648307
transform 1 0 -400 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3524
timestamp 1654648307
transform 1 0 4100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3523
timestamp 1654648307
transform 1 0 2600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3444
timestamp 1654648307
transform 1 0 4100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3443
timestamp 1654648307
transform 1 0 2600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3526
timestamp 1654648307
transform 1 0 7100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3525
timestamp 1654648307
transform 1 0 5600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3446
timestamp 1654648307
transform 1 0 7100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3445
timestamp 1654648307
transform 1 0 5600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3528
timestamp 1654648307
transform 1 0 10100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3527
timestamp 1654648307
transform 1 0 8600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3448
timestamp 1654648307
transform 1 0 10100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3447
timestamp 1654648307
transform 1 0 8600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3530
timestamp 1654648307
transform 1 0 13100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3529
timestamp 1654648307
transform 1 0 11600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3450
timestamp 1654648307
transform 1 0 13100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3449
timestamp 1654648307
transform 1 0 11600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3532
timestamp 1654648307
transform 1 0 16100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3531
timestamp 1654648307
transform 1 0 14600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3452
timestamp 1654648307
transform 1 0 16100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3451
timestamp 1654648307
transform 1 0 14600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3534
timestamp 1654648307
transform 1 0 19100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3533
timestamp 1654648307
transform 1 0 17600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3454
timestamp 1654648307
transform 1 0 19100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3453
timestamp 1654648307
transform 1 0 17600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3536
timestamp 1654648307
transform 1 0 22100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3535
timestamp 1654648307
transform 1 0 20600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3456
timestamp 1654648307
transform 1 0 22100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3455
timestamp 1654648307
transform 1 0 20600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3538
timestamp 1654648307
transform 1 0 25100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3537
timestamp 1654648307
transform 1 0 23600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3458
timestamp 1654648307
transform 1 0 25100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3457
timestamp 1654648307
transform 1 0 23600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3540
timestamp 1654648307
transform 1 0 28100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3539
timestamp 1654648307
transform 1 0 26600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3460
timestamp 1654648307
transform 1 0 28100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3459
timestamp 1654648307
transform 1 0 26600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3542
timestamp 1654648307
transform 1 0 31100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3541
timestamp 1654648307
transform 1 0 29600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3462
timestamp 1654648307
transform 1 0 31100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3461
timestamp 1654648307
transform 1 0 29600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3544
timestamp 1654648307
transform 1 0 34100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3543
timestamp 1654648307
transform 1 0 32600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3464
timestamp 1654648307
transform 1 0 34100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3463
timestamp 1654648307
transform 1 0 32600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3546
timestamp 1654648307
transform 1 0 37100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3545
timestamp 1654648307
transform 1 0 35600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3466
timestamp 1654648307
transform 1 0 37100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3465
timestamp 1654648307
transform 1 0 35600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3548
timestamp 1654648307
transform 1 0 40100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3547
timestamp 1654648307
transform 1 0 38600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3468
timestamp 1654648307
transform 1 0 40100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3467
timestamp 1654648307
transform 1 0 38600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3550
timestamp 1654648307
transform 1 0 43100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3549
timestamp 1654648307
transform 1 0 41600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3470
timestamp 1654648307
transform 1 0 43100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3469
timestamp 1654648307
transform 1 0 41600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3552
timestamp 1654648307
transform 1 0 46100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3551
timestamp 1654648307
transform 1 0 44600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3472
timestamp 1654648307
transform 1 0 46100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3471
timestamp 1654648307
transform 1 0 44600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3554
timestamp 1654648307
transform 1 0 49100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3553
timestamp 1654648307
transform 1 0 47600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3474
timestamp 1654648307
transform 1 0 49100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3473
timestamp 1654648307
transform 1 0 47600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3556
timestamp 1654648307
transform 1 0 52100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3555
timestamp 1654648307
transform 1 0 50600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3476
timestamp 1654648307
transform 1 0 52100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3475
timestamp 1654648307
transform 1 0 50600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3558
timestamp 1654648307
transform 1 0 55100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3557
timestamp 1654648307
transform 1 0 53600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3478
timestamp 1654648307
transform 1 0 55100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3477
timestamp 1654648307
transform 1 0 53600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3560
timestamp 1654648307
transform 1 0 58100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3559
timestamp 1654648307
transform 1 0 56600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3480
timestamp 1654648307
transform 1 0 58100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3479
timestamp 1654648307
transform 1 0 56600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3562
timestamp 1654648307
transform 1 0 61100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3561
timestamp 1654648307
transform 1 0 59600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3482
timestamp 1654648307
transform 1 0 61100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3481
timestamp 1654648307
transform 1 0 59600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3563
timestamp 1654648307
transform 1 0 62600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3483
timestamp 1654648307
transform 1 0 62600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3564
timestamp 1654648307
transform 1 0 64100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3484
timestamp 1654648307
transform 1 0 64100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3565
timestamp 1654648307
transform 1 0 65600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3485
timestamp 1654648307
transform 1 0 65600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3566
timestamp 1654648307
transform 1 0 67100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3486
timestamp 1654648307
transform 1 0 67100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3567
timestamp 1654648307
transform 1 0 68600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3487
timestamp 1654648307
transform 1 0 68600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3568
timestamp 1654648307
transform 1 0 70100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3488
timestamp 1654648307
transform 1 0 70100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3569
timestamp 1654648307
transform 1 0 71600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3489
timestamp 1654648307
transform 1 0 71600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3570
timestamp 1654648307
transform 1 0 73100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3490
timestamp 1654648307
transform 1 0 73100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3571
timestamp 1654648307
transform 1 0 74600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3491
timestamp 1654648307
transform 1 0 74600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3572
timestamp 1654648307
transform 1 0 76100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3492
timestamp 1654648307
transform 1 0 76100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3573
timestamp 1654648307
transform 1 0 77600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3493
timestamp 1654648307
transform 1 0 77600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3574
timestamp 1654648307
transform 1 0 79100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3494
timestamp 1654648307
transform 1 0 79100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3575
timestamp 1654648307
transform 1 0 80600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3495
timestamp 1654648307
transform 1 0 80600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3576
timestamp 1654648307
transform 1 0 82100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3496
timestamp 1654648307
transform 1 0 82100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3577
timestamp 1654648307
transform 1 0 83600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3497
timestamp 1654648307
transform 1 0 83600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3578
timestamp 1654648307
transform 1 0 85100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3498
timestamp 1654648307
transform 1 0 85100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3579
timestamp 1654648307
transform 1 0 86600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3499
timestamp 1654648307
transform 1 0 86600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3580
timestamp 1654648307
transform 1 0 88100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3500
timestamp 1654648307
transform 1 0 88100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3581
timestamp 1654648307
transform 1 0 89600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3501
timestamp 1654648307
transform 1 0 89600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3582
timestamp 1654648307
transform 1 0 91100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3502
timestamp 1654648307
transform 1 0 91100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3583
timestamp 1654648307
transform 1 0 92600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3503
timestamp 1654648307
transform 1 0 92600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3584
timestamp 1654648307
transform 1 0 94100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3504
timestamp 1654648307
transform 1 0 94100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3585
timestamp 1654648307
transform 1 0 95600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3505
timestamp 1654648307
transform 1 0 95600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3586
timestamp 1654648307
transform 1 0 97100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3506
timestamp 1654648307
transform 1 0 97100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3587
timestamp 1654648307
transform 1 0 98600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3507
timestamp 1654648307
transform 1 0 98600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3588
timestamp 1654648307
transform 1 0 100100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3508
timestamp 1654648307
transform 1 0 100100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3589
timestamp 1654648307
transform 1 0 101600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3509
timestamp 1654648307
transform 1 0 101600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3590
timestamp 1654648307
transform 1 0 103100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3510
timestamp 1654648307
transform 1 0 103100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3591
timestamp 1654648307
transform 1 0 104600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3511
timestamp 1654648307
transform 1 0 104600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3592
timestamp 1654648307
transform 1 0 106100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3512
timestamp 1654648307
transform 1 0 106100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3593
timestamp 1654648307
transform 1 0 107600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3513
timestamp 1654648307
transform 1 0 107600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3594
timestamp 1654648307
transform 1 0 109100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3514
timestamp 1654648307
transform 1 0 109100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3595
timestamp 1654648307
transform 1 0 110600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3515
timestamp 1654648307
transform 1 0 110600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3596
timestamp 1654648307
transform 1 0 112100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3516
timestamp 1654648307
transform 1 0 112100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3597
timestamp 1654648307
transform 1 0 113600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3517
timestamp 1654648307
transform 1 0 113600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3598
timestamp 1654648307
transform 1 0 115100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3518
timestamp 1654648307
transform 1 0 115100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3599
timestamp 1654648307
transform 1 0 116600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_3519
timestamp 1654648307
transform 1 0 116600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_3360
timestamp 1654648307
transform 1 0 -1900 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3280
timestamp 1654648307
transform 1 0 -1900 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3362
timestamp 1654648307
transform 1 0 1100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3361
timestamp 1654648307
transform 1 0 -400 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3282
timestamp 1654648307
transform 1 0 1100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3281
timestamp 1654648307
transform 1 0 -400 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3364
timestamp 1654648307
transform 1 0 4100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3363
timestamp 1654648307
transform 1 0 2600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3284
timestamp 1654648307
transform 1 0 4100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3283
timestamp 1654648307
transform 1 0 2600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3366
timestamp 1654648307
transform 1 0 7100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3365
timestamp 1654648307
transform 1 0 5600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3286
timestamp 1654648307
transform 1 0 7100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3285
timestamp 1654648307
transform 1 0 5600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3368
timestamp 1654648307
transform 1 0 10100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3367
timestamp 1654648307
transform 1 0 8600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3288
timestamp 1654648307
transform 1 0 10100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3287
timestamp 1654648307
transform 1 0 8600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3370
timestamp 1654648307
transform 1 0 13100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3369
timestamp 1654648307
transform 1 0 11600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3290
timestamp 1654648307
transform 1 0 13100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3289
timestamp 1654648307
transform 1 0 11600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3372
timestamp 1654648307
transform 1 0 16100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3371
timestamp 1654648307
transform 1 0 14600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3292
timestamp 1654648307
transform 1 0 16100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3291
timestamp 1654648307
transform 1 0 14600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3374
timestamp 1654648307
transform 1 0 19100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3373
timestamp 1654648307
transform 1 0 17600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3294
timestamp 1654648307
transform 1 0 19100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3293
timestamp 1654648307
transform 1 0 17600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3376
timestamp 1654648307
transform 1 0 22100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3375
timestamp 1654648307
transform 1 0 20600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3296
timestamp 1654648307
transform 1 0 22100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3295
timestamp 1654648307
transform 1 0 20600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3378
timestamp 1654648307
transform 1 0 25100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3377
timestamp 1654648307
transform 1 0 23600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3298
timestamp 1654648307
transform 1 0 25100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3297
timestamp 1654648307
transform 1 0 23600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3380
timestamp 1654648307
transform 1 0 28100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3379
timestamp 1654648307
transform 1 0 26600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3300
timestamp 1654648307
transform 1 0 28100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3299
timestamp 1654648307
transform 1 0 26600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3382
timestamp 1654648307
transform 1 0 31100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3381
timestamp 1654648307
transform 1 0 29600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3302
timestamp 1654648307
transform 1 0 31100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3301
timestamp 1654648307
transform 1 0 29600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3384
timestamp 1654648307
transform 1 0 34100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3383
timestamp 1654648307
transform 1 0 32600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3304
timestamp 1654648307
transform 1 0 34100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3303
timestamp 1654648307
transform 1 0 32600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3386
timestamp 1654648307
transform 1 0 37100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3385
timestamp 1654648307
transform 1 0 35600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3306
timestamp 1654648307
transform 1 0 37100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3305
timestamp 1654648307
transform 1 0 35600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3388
timestamp 1654648307
transform 1 0 40100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3387
timestamp 1654648307
transform 1 0 38600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3308
timestamp 1654648307
transform 1 0 40100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3307
timestamp 1654648307
transform 1 0 38600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3390
timestamp 1654648307
transform 1 0 43100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3389
timestamp 1654648307
transform 1 0 41600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3310
timestamp 1654648307
transform 1 0 43100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3309
timestamp 1654648307
transform 1 0 41600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3392
timestamp 1654648307
transform 1 0 46100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3391
timestamp 1654648307
transform 1 0 44600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3312
timestamp 1654648307
transform 1 0 46100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3311
timestamp 1654648307
transform 1 0 44600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3394
timestamp 1654648307
transform 1 0 49100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3393
timestamp 1654648307
transform 1 0 47600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3314
timestamp 1654648307
transform 1 0 49100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3313
timestamp 1654648307
transform 1 0 47600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3396
timestamp 1654648307
transform 1 0 52100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3395
timestamp 1654648307
transform 1 0 50600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3316
timestamp 1654648307
transform 1 0 52100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3315
timestamp 1654648307
transform 1 0 50600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3398
timestamp 1654648307
transform 1 0 55100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3397
timestamp 1654648307
transform 1 0 53600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3318
timestamp 1654648307
transform 1 0 55100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3317
timestamp 1654648307
transform 1 0 53600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3400
timestamp 1654648307
transform 1 0 58100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3399
timestamp 1654648307
transform 1 0 56600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3320
timestamp 1654648307
transform 1 0 58100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3319
timestamp 1654648307
transform 1 0 56600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3402
timestamp 1654648307
transform 1 0 61100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3401
timestamp 1654648307
transform 1 0 59600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3322
timestamp 1654648307
transform 1 0 61100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3321
timestamp 1654648307
transform 1 0 59600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3403
timestamp 1654648307
transform 1 0 62600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3323
timestamp 1654648307
transform 1 0 62600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3404
timestamp 1654648307
transform 1 0 64100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3324
timestamp 1654648307
transform 1 0 64100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3405
timestamp 1654648307
transform 1 0 65600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3325
timestamp 1654648307
transform 1 0 65600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3406
timestamp 1654648307
transform 1 0 67100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3326
timestamp 1654648307
transform 1 0 67100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3407
timestamp 1654648307
transform 1 0 68600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3327
timestamp 1654648307
transform 1 0 68600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3408
timestamp 1654648307
transform 1 0 70100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3328
timestamp 1654648307
transform 1 0 70100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3409
timestamp 1654648307
transform 1 0 71600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3329
timestamp 1654648307
transform 1 0 71600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3410
timestamp 1654648307
transform 1 0 73100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3330
timestamp 1654648307
transform 1 0 73100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3411
timestamp 1654648307
transform 1 0 74600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3331
timestamp 1654648307
transform 1 0 74600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3412
timestamp 1654648307
transform 1 0 76100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3332
timestamp 1654648307
transform 1 0 76100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3413
timestamp 1654648307
transform 1 0 77600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3333
timestamp 1654648307
transform 1 0 77600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3414
timestamp 1654648307
transform 1 0 79100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3334
timestamp 1654648307
transform 1 0 79100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3415
timestamp 1654648307
transform 1 0 80600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3335
timestamp 1654648307
transform 1 0 80600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3416
timestamp 1654648307
transform 1 0 82100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3336
timestamp 1654648307
transform 1 0 82100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3417
timestamp 1654648307
transform 1 0 83600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3337
timestamp 1654648307
transform 1 0 83600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3418
timestamp 1654648307
transform 1 0 85100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3338
timestamp 1654648307
transform 1 0 85100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3419
timestamp 1654648307
transform 1 0 86600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3339
timestamp 1654648307
transform 1 0 86600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3420
timestamp 1654648307
transform 1 0 88100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3340
timestamp 1654648307
transform 1 0 88100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3421
timestamp 1654648307
transform 1 0 89600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3341
timestamp 1654648307
transform 1 0 89600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3422
timestamp 1654648307
transform 1 0 91100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3342
timestamp 1654648307
transform 1 0 91100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3423
timestamp 1654648307
transform 1 0 92600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3343
timestamp 1654648307
transform 1 0 92600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3424
timestamp 1654648307
transform 1 0 94100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3344
timestamp 1654648307
transform 1 0 94100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3425
timestamp 1654648307
transform 1 0 95600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3345
timestamp 1654648307
transform 1 0 95600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3426
timestamp 1654648307
transform 1 0 97100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3346
timestamp 1654648307
transform 1 0 97100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3427
timestamp 1654648307
transform 1 0 98600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3347
timestamp 1654648307
transform 1 0 98600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3428
timestamp 1654648307
transform 1 0 100100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3348
timestamp 1654648307
transform 1 0 100100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3429
timestamp 1654648307
transform 1 0 101600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3349
timestamp 1654648307
transform 1 0 101600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3430
timestamp 1654648307
transform 1 0 103100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3350
timestamp 1654648307
transform 1 0 103100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3431
timestamp 1654648307
transform 1 0 104600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3351
timestamp 1654648307
transform 1 0 104600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3432
timestamp 1654648307
transform 1 0 106100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3352
timestamp 1654648307
transform 1 0 106100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3433
timestamp 1654648307
transform 1 0 107600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3353
timestamp 1654648307
transform 1 0 107600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3434
timestamp 1654648307
transform 1 0 109100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3354
timestamp 1654648307
transform 1 0 109100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3435
timestamp 1654648307
transform 1 0 110600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3355
timestamp 1654648307
transform 1 0 110600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3436
timestamp 1654648307
transform 1 0 112100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3356
timestamp 1654648307
transform 1 0 112100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3437
timestamp 1654648307
transform 1 0 113600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3357
timestamp 1654648307
transform 1 0 113600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3438
timestamp 1654648307
transform 1 0 115100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3358
timestamp 1654648307
transform 1 0 115100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3439
timestamp 1654648307
transform 1 0 116600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_3359
timestamp 1654648307
transform 1 0 116600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_3200
timestamp 1654648307
transform 1 0 -1900 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3120
timestamp 1654648307
transform 1 0 -1900 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3202
timestamp 1654648307
transform 1 0 1100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3201
timestamp 1654648307
transform 1 0 -400 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3122
timestamp 1654648307
transform 1 0 1100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3121
timestamp 1654648307
transform 1 0 -400 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3204
timestamp 1654648307
transform 1 0 4100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3203
timestamp 1654648307
transform 1 0 2600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3124
timestamp 1654648307
transform 1 0 4100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3123
timestamp 1654648307
transform 1 0 2600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3206
timestamp 1654648307
transform 1 0 7100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3205
timestamp 1654648307
transform 1 0 5600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3126
timestamp 1654648307
transform 1 0 7100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3125
timestamp 1654648307
transform 1 0 5600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3208
timestamp 1654648307
transform 1 0 10100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3207
timestamp 1654648307
transform 1 0 8600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3128
timestamp 1654648307
transform 1 0 10100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3127
timestamp 1654648307
transform 1 0 8600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3210
timestamp 1654648307
transform 1 0 13100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3209
timestamp 1654648307
transform 1 0 11600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3130
timestamp 1654648307
transform 1 0 13100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3129
timestamp 1654648307
transform 1 0 11600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3212
timestamp 1654648307
transform 1 0 16100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3211
timestamp 1654648307
transform 1 0 14600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3132
timestamp 1654648307
transform 1 0 16100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3131
timestamp 1654648307
transform 1 0 14600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3214
timestamp 1654648307
transform 1 0 19100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3213
timestamp 1654648307
transform 1 0 17600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3134
timestamp 1654648307
transform 1 0 19100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3133
timestamp 1654648307
transform 1 0 17600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3216
timestamp 1654648307
transform 1 0 22100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3215
timestamp 1654648307
transform 1 0 20600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3136
timestamp 1654648307
transform 1 0 22100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3135
timestamp 1654648307
transform 1 0 20600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3218
timestamp 1654648307
transform 1 0 25100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3217
timestamp 1654648307
transform 1 0 23600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3138
timestamp 1654648307
transform 1 0 25100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3137
timestamp 1654648307
transform 1 0 23600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3220
timestamp 1654648307
transform 1 0 28100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3219
timestamp 1654648307
transform 1 0 26600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3140
timestamp 1654648307
transform 1 0 28100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3139
timestamp 1654648307
transform 1 0 26600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3222
timestamp 1654648307
transform 1 0 31100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3221
timestamp 1654648307
transform 1 0 29600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3142
timestamp 1654648307
transform 1 0 31100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3141
timestamp 1654648307
transform 1 0 29600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3224
timestamp 1654648307
transform 1 0 34100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3223
timestamp 1654648307
transform 1 0 32600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3144
timestamp 1654648307
transform 1 0 34100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3143
timestamp 1654648307
transform 1 0 32600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3226
timestamp 1654648307
transform 1 0 37100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3225
timestamp 1654648307
transform 1 0 35600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3146
timestamp 1654648307
transform 1 0 37100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3145
timestamp 1654648307
transform 1 0 35600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3228
timestamp 1654648307
transform 1 0 40100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3227
timestamp 1654648307
transform 1 0 38600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3148
timestamp 1654648307
transform 1 0 40100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3147
timestamp 1654648307
transform 1 0 38600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3230
timestamp 1654648307
transform 1 0 43100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3229
timestamp 1654648307
transform 1 0 41600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3150
timestamp 1654648307
transform 1 0 43100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3149
timestamp 1654648307
transform 1 0 41600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3232
timestamp 1654648307
transform 1 0 46100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3231
timestamp 1654648307
transform 1 0 44600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3152
timestamp 1654648307
transform 1 0 46100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3151
timestamp 1654648307
transform 1 0 44600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3234
timestamp 1654648307
transform 1 0 49100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3233
timestamp 1654648307
transform 1 0 47600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3154
timestamp 1654648307
transform 1 0 49100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3153
timestamp 1654648307
transform 1 0 47600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3236
timestamp 1654648307
transform 1 0 52100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3235
timestamp 1654648307
transform 1 0 50600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3156
timestamp 1654648307
transform 1 0 52100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3155
timestamp 1654648307
transform 1 0 50600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3238
timestamp 1654648307
transform 1 0 55100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3237
timestamp 1654648307
transform 1 0 53600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3158
timestamp 1654648307
transform 1 0 55100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3157
timestamp 1654648307
transform 1 0 53600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3240
timestamp 1654648307
transform 1 0 58100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3239
timestamp 1654648307
transform 1 0 56600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3160
timestamp 1654648307
transform 1 0 58100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3159
timestamp 1654648307
transform 1 0 56600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3242
timestamp 1654648307
transform 1 0 61100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3241
timestamp 1654648307
transform 1 0 59600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3162
timestamp 1654648307
transform 1 0 61100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3161
timestamp 1654648307
transform 1 0 59600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3243
timestamp 1654648307
transform 1 0 62600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3163
timestamp 1654648307
transform 1 0 62600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3244
timestamp 1654648307
transform 1 0 64100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3164
timestamp 1654648307
transform 1 0 64100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3245
timestamp 1654648307
transform 1 0 65600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3165
timestamp 1654648307
transform 1 0 65600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3246
timestamp 1654648307
transform 1 0 67100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3166
timestamp 1654648307
transform 1 0 67100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3247
timestamp 1654648307
transform 1 0 68600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3167
timestamp 1654648307
transform 1 0 68600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3248
timestamp 1654648307
transform 1 0 70100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3168
timestamp 1654648307
transform 1 0 70100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3249
timestamp 1654648307
transform 1 0 71600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3169
timestamp 1654648307
transform 1 0 71600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3250
timestamp 1654648307
transform 1 0 73100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3170
timestamp 1654648307
transform 1 0 73100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3251
timestamp 1654648307
transform 1 0 74600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3171
timestamp 1654648307
transform 1 0 74600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3252
timestamp 1654648307
transform 1 0 76100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3172
timestamp 1654648307
transform 1 0 76100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3253
timestamp 1654648307
transform 1 0 77600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3173
timestamp 1654648307
transform 1 0 77600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3254
timestamp 1654648307
transform 1 0 79100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3174
timestamp 1654648307
transform 1 0 79100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3255
timestamp 1654648307
transform 1 0 80600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3175
timestamp 1654648307
transform 1 0 80600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3256
timestamp 1654648307
transform 1 0 82100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3176
timestamp 1654648307
transform 1 0 82100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3257
timestamp 1654648307
transform 1 0 83600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3177
timestamp 1654648307
transform 1 0 83600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3258
timestamp 1654648307
transform 1 0 85100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3178
timestamp 1654648307
transform 1 0 85100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3259
timestamp 1654648307
transform 1 0 86600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3179
timestamp 1654648307
transform 1 0 86600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3260
timestamp 1654648307
transform 1 0 88100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3180
timestamp 1654648307
transform 1 0 88100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3261
timestamp 1654648307
transform 1 0 89600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3181
timestamp 1654648307
transform 1 0 89600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3262
timestamp 1654648307
transform 1 0 91100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3182
timestamp 1654648307
transform 1 0 91100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3263
timestamp 1654648307
transform 1 0 92600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3183
timestamp 1654648307
transform 1 0 92600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3264
timestamp 1654648307
transform 1 0 94100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3184
timestamp 1654648307
transform 1 0 94100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3265
timestamp 1654648307
transform 1 0 95600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3185
timestamp 1654648307
transform 1 0 95600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3266
timestamp 1654648307
transform 1 0 97100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3186
timestamp 1654648307
transform 1 0 97100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3267
timestamp 1654648307
transform 1 0 98600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3187
timestamp 1654648307
transform 1 0 98600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3268
timestamp 1654648307
transform 1 0 100100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3188
timestamp 1654648307
transform 1 0 100100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3269
timestamp 1654648307
transform 1 0 101600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3189
timestamp 1654648307
transform 1 0 101600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3270
timestamp 1654648307
transform 1 0 103100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3190
timestamp 1654648307
transform 1 0 103100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3271
timestamp 1654648307
transform 1 0 104600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3191
timestamp 1654648307
transform 1 0 104600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3272
timestamp 1654648307
transform 1 0 106100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3192
timestamp 1654648307
transform 1 0 106100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3273
timestamp 1654648307
transform 1 0 107600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3193
timestamp 1654648307
transform 1 0 107600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3274
timestamp 1654648307
transform 1 0 109100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3194
timestamp 1654648307
transform 1 0 109100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3275
timestamp 1654648307
transform 1 0 110600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3195
timestamp 1654648307
transform 1 0 110600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3276
timestamp 1654648307
transform 1 0 112100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3196
timestamp 1654648307
transform 1 0 112100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3277
timestamp 1654648307
transform 1 0 113600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3197
timestamp 1654648307
transform 1 0 113600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3278
timestamp 1654648307
transform 1 0 115100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3198
timestamp 1654648307
transform 1 0 115100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3279
timestamp 1654648307
transform 1 0 116600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_3199
timestamp 1654648307
transform 1 0 116600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3040
timestamp 1654648307
transform 1 0 -1900 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2960
timestamp 1654648307
transform 1 0 -1900 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3042
timestamp 1654648307
transform 1 0 1100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3041
timestamp 1654648307
transform 1 0 -400 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2962
timestamp 1654648307
transform 1 0 1100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_2961
timestamp 1654648307
transform 1 0 -400 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3044
timestamp 1654648307
transform 1 0 4100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3043
timestamp 1654648307
transform 1 0 2600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2964
timestamp 1654648307
transform 1 0 4100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_2963
timestamp 1654648307
transform 1 0 2600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3046
timestamp 1654648307
transform 1 0 7100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3045
timestamp 1654648307
transform 1 0 5600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2966
timestamp 1654648307
transform 1 0 7100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_2965
timestamp 1654648307
transform 1 0 5600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3048
timestamp 1654648307
transform 1 0 10100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3047
timestamp 1654648307
transform 1 0 8600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2968
timestamp 1654648307
transform 1 0 10100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_2967
timestamp 1654648307
transform 1 0 8600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3050
timestamp 1654648307
transform 1 0 13100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3049
timestamp 1654648307
transform 1 0 11600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2970
timestamp 1654648307
transform 1 0 13100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_2969
timestamp 1654648307
transform 1 0 11600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3052
timestamp 1654648307
transform 1 0 16100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3051
timestamp 1654648307
transform 1 0 14600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2972
timestamp 1654648307
transform 1 0 16100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_2971
timestamp 1654648307
transform 1 0 14600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3054
timestamp 1654648307
transform 1 0 19100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3053
timestamp 1654648307
transform 1 0 17600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2974
timestamp 1654648307
transform 1 0 19100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_2973
timestamp 1654648307
transform 1 0 17600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3055
timestamp 1654648307
transform 1 0 20600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2975
timestamp 1654648307
transform 1 0 20600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3056
timestamp 1654648307
transform 1 0 22100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2976
timestamp 1654648307
transform 1 0 22100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3057
timestamp 1654648307
transform 1 0 23600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2977
timestamp 1654648307
transform 1 0 23600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3058
timestamp 1654648307
transform 1 0 25100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2978
timestamp 1654648307
transform 1 0 25100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3059
timestamp 1654648307
transform 1 0 26600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2979
timestamp 1654648307
transform 1 0 26600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3060
timestamp 1654648307
transform 1 0 28100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2980
timestamp 1654648307
transform 1 0 28100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3061
timestamp 1654648307
transform 1 0 29600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2981
timestamp 1654648307
transform 1 0 29600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3062
timestamp 1654648307
transform 1 0 31100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2982
timestamp 1654648307
transform 1 0 31100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3063
timestamp 1654648307
transform 1 0 32600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2983
timestamp 1654648307
transform 1 0 32600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3064
timestamp 1654648307
transform 1 0 34100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2984
timestamp 1654648307
transform 1 0 34100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3065
timestamp 1654648307
transform 1 0 35600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2985
timestamp 1654648307
transform 1 0 35600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3066
timestamp 1654648307
transform 1 0 37100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2986
timestamp 1654648307
transform 1 0 37100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3067
timestamp 1654648307
transform 1 0 38600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2987
timestamp 1654648307
transform 1 0 38600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3068
timestamp 1654648307
transform 1 0 40100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2988
timestamp 1654648307
transform 1 0 40100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3069
timestamp 1654648307
transform 1 0 41600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2989
timestamp 1654648307
transform 1 0 41600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3070
timestamp 1654648307
transform 1 0 43100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2990
timestamp 1654648307
transform 1 0 43100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3071
timestamp 1654648307
transform 1 0 44600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2991
timestamp 1654648307
transform 1 0 44600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3072
timestamp 1654648307
transform 1 0 46100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2992
timestamp 1654648307
transform 1 0 46100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3073
timestamp 1654648307
transform 1 0 47600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2993
timestamp 1654648307
transform 1 0 47600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3074
timestamp 1654648307
transform 1 0 49100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2994
timestamp 1654648307
transform 1 0 49100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3075
timestamp 1654648307
transform 1 0 50600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2995
timestamp 1654648307
transform 1 0 50600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3076
timestamp 1654648307
transform 1 0 52100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2996
timestamp 1654648307
transform 1 0 52100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3077
timestamp 1654648307
transform 1 0 53600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2997
timestamp 1654648307
transform 1 0 53600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3078
timestamp 1654648307
transform 1 0 55100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2998
timestamp 1654648307
transform 1 0 55100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3079
timestamp 1654648307
transform 1 0 56600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_2999
timestamp 1654648307
transform 1 0 56600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3080
timestamp 1654648307
transform 1 0 58100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3000
timestamp 1654648307
transform 1 0 58100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3081
timestamp 1654648307
transform 1 0 59600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3001
timestamp 1654648307
transform 1 0 59600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3082
timestamp 1654648307
transform 1 0 61100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3002
timestamp 1654648307
transform 1 0 61100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3083
timestamp 1654648307
transform 1 0 62600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3003
timestamp 1654648307
transform 1 0 62600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3084
timestamp 1654648307
transform 1 0 64100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3004
timestamp 1654648307
transform 1 0 64100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3085
timestamp 1654648307
transform 1 0 65600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3005
timestamp 1654648307
transform 1 0 65600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3086
timestamp 1654648307
transform 1 0 67100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3006
timestamp 1654648307
transform 1 0 67100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3087
timestamp 1654648307
transform 1 0 68600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3007
timestamp 1654648307
transform 1 0 68600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3088
timestamp 1654648307
transform 1 0 70100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3008
timestamp 1654648307
transform 1 0 70100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3089
timestamp 1654648307
transform 1 0 71600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3009
timestamp 1654648307
transform 1 0 71600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3090
timestamp 1654648307
transform 1 0 73100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3010
timestamp 1654648307
transform 1 0 73100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3091
timestamp 1654648307
transform 1 0 74600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3011
timestamp 1654648307
transform 1 0 74600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3092
timestamp 1654648307
transform 1 0 76100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3012
timestamp 1654648307
transform 1 0 76100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3093
timestamp 1654648307
transform 1 0 77600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3013
timestamp 1654648307
transform 1 0 77600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3094
timestamp 1654648307
transform 1 0 79100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3014
timestamp 1654648307
transform 1 0 79100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3095
timestamp 1654648307
transform 1 0 80600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3015
timestamp 1654648307
transform 1 0 80600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3096
timestamp 1654648307
transform 1 0 82100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3016
timestamp 1654648307
transform 1 0 82100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3097
timestamp 1654648307
transform 1 0 83600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3017
timestamp 1654648307
transform 1 0 83600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3098
timestamp 1654648307
transform 1 0 85100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3018
timestamp 1654648307
transform 1 0 85100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3099
timestamp 1654648307
transform 1 0 86600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3019
timestamp 1654648307
transform 1 0 86600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3100
timestamp 1654648307
transform 1 0 88100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3020
timestamp 1654648307
transform 1 0 88100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3101
timestamp 1654648307
transform 1 0 89600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3021
timestamp 1654648307
transform 1 0 89600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3102
timestamp 1654648307
transform 1 0 91100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3022
timestamp 1654648307
transform 1 0 91100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3103
timestamp 1654648307
transform 1 0 92600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3023
timestamp 1654648307
transform 1 0 92600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3104
timestamp 1654648307
transform 1 0 94100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3024
timestamp 1654648307
transform 1 0 94100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3105
timestamp 1654648307
transform 1 0 95600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3025
timestamp 1654648307
transform 1 0 95600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3106
timestamp 1654648307
transform 1 0 97100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3026
timestamp 1654648307
transform 1 0 97100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3107
timestamp 1654648307
transform 1 0 98600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3027
timestamp 1654648307
transform 1 0 98600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3108
timestamp 1654648307
transform 1 0 100100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3028
timestamp 1654648307
transform 1 0 100100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3109
timestamp 1654648307
transform 1 0 101600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3029
timestamp 1654648307
transform 1 0 101600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3110
timestamp 1654648307
transform 1 0 103100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3030
timestamp 1654648307
transform 1 0 103100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3111
timestamp 1654648307
transform 1 0 104600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3031
timestamp 1654648307
transform 1 0 104600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3112
timestamp 1654648307
transform 1 0 106100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3032
timestamp 1654648307
transform 1 0 106100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3113
timestamp 1654648307
transform 1 0 107600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3033
timestamp 1654648307
transform 1 0 107600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3114
timestamp 1654648307
transform 1 0 109100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3034
timestamp 1654648307
transform 1 0 109100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3115
timestamp 1654648307
transform 1 0 110600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3035
timestamp 1654648307
transform 1 0 110600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3116
timestamp 1654648307
transform 1 0 112100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3036
timestamp 1654648307
transform 1 0 112100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3117
timestamp 1654648307
transform 1 0 113600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3037
timestamp 1654648307
transform 1 0 113600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3118
timestamp 1654648307
transform 1 0 115100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3038
timestamp 1654648307
transform 1 0 115100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3119
timestamp 1654648307
transform 1 0 116600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3039
timestamp 1654648307
transform 1 0 116600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_2880
timestamp 1654648307
transform 1 0 -1900 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2800
timestamp 1654648307
transform 1 0 -1900 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2882
timestamp 1654648307
transform 1 0 1100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2881
timestamp 1654648307
transform 1 0 -400 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2802
timestamp 1654648307
transform 1 0 1100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2801
timestamp 1654648307
transform 1 0 -400 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2884
timestamp 1654648307
transform 1 0 4100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2883
timestamp 1654648307
transform 1 0 2600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2804
timestamp 1654648307
transform 1 0 4100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2803
timestamp 1654648307
transform 1 0 2600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2886
timestamp 1654648307
transform 1 0 7100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2885
timestamp 1654648307
transform 1 0 5600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2806
timestamp 1654648307
transform 1 0 7100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2805
timestamp 1654648307
transform 1 0 5600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2888
timestamp 1654648307
transform 1 0 10100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2887
timestamp 1654648307
transform 1 0 8600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2808
timestamp 1654648307
transform 1 0 10100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2807
timestamp 1654648307
transform 1 0 8600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2890
timestamp 1654648307
transform 1 0 13100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2889
timestamp 1654648307
transform 1 0 11600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2810
timestamp 1654648307
transform 1 0 13100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2809
timestamp 1654648307
transform 1 0 11600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2892
timestamp 1654648307
transform 1 0 16100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2891
timestamp 1654648307
transform 1 0 14600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2812
timestamp 1654648307
transform 1 0 16100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2811
timestamp 1654648307
transform 1 0 14600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2894
timestamp 1654648307
transform 1 0 19100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2893
timestamp 1654648307
transform 1 0 17600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2814
timestamp 1654648307
transform 1 0 19100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2813
timestamp 1654648307
transform 1 0 17600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2895
timestamp 1654648307
transform 1 0 20600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2815
timestamp 1654648307
transform 1 0 20600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2896
timestamp 1654648307
transform 1 0 22100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2816
timestamp 1654648307
transform 1 0 22100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2897
timestamp 1654648307
transform 1 0 23600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2817
timestamp 1654648307
transform 1 0 23600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2898
timestamp 1654648307
transform 1 0 25100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2818
timestamp 1654648307
transform 1 0 25100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2899
timestamp 1654648307
transform 1 0 26600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2819
timestamp 1654648307
transform 1 0 26600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2900
timestamp 1654648307
transform 1 0 28100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2820
timestamp 1654648307
transform 1 0 28100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2901
timestamp 1654648307
transform 1 0 29600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2821
timestamp 1654648307
transform 1 0 29600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2902
timestamp 1654648307
transform 1 0 31100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2822
timestamp 1654648307
transform 1 0 31100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2903
timestamp 1654648307
transform 1 0 32600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2823
timestamp 1654648307
transform 1 0 32600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2904
timestamp 1654648307
transform 1 0 34100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2824
timestamp 1654648307
transform 1 0 34100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2905
timestamp 1654648307
transform 1 0 35600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2825
timestamp 1654648307
transform 1 0 35600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2906
timestamp 1654648307
transform 1 0 37100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2826
timestamp 1654648307
transform 1 0 37100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2907
timestamp 1654648307
transform 1 0 38600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2827
timestamp 1654648307
transform 1 0 38600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2908
timestamp 1654648307
transform 1 0 40100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2828
timestamp 1654648307
transform 1 0 40100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2909
timestamp 1654648307
transform 1 0 41600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2829
timestamp 1654648307
transform 1 0 41600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2910
timestamp 1654648307
transform 1 0 43100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2830
timestamp 1654648307
transform 1 0 43100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2911
timestamp 1654648307
transform 1 0 44600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2831
timestamp 1654648307
transform 1 0 44600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2912
timestamp 1654648307
transform 1 0 46100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2832
timestamp 1654648307
transform 1 0 46100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2913
timestamp 1654648307
transform 1 0 47600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2833
timestamp 1654648307
transform 1 0 47600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2914
timestamp 1654648307
transform 1 0 49100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2834
timestamp 1654648307
transform 1 0 49100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2915
timestamp 1654648307
transform 1 0 50600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2835
timestamp 1654648307
transform 1 0 50600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2916
timestamp 1654648307
transform 1 0 52100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2836
timestamp 1654648307
transform 1 0 52100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2917
timestamp 1654648307
transform 1 0 53600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2837
timestamp 1654648307
transform 1 0 53600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2918
timestamp 1654648307
transform 1 0 55100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2838
timestamp 1654648307
transform 1 0 55100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2919
timestamp 1654648307
transform 1 0 56600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2839
timestamp 1654648307
transform 1 0 56600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2920
timestamp 1654648307
transform 1 0 58100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2840
timestamp 1654648307
transform 1 0 58100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2921
timestamp 1654648307
transform 1 0 59600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2841
timestamp 1654648307
transform 1 0 59600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2922
timestamp 1654648307
transform 1 0 61100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2842
timestamp 1654648307
transform 1 0 61100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2923
timestamp 1654648307
transform 1 0 62600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2843
timestamp 1654648307
transform 1 0 62600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2924
timestamp 1654648307
transform 1 0 64100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2844
timestamp 1654648307
transform 1 0 64100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2925
timestamp 1654648307
transform 1 0 65600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2845
timestamp 1654648307
transform 1 0 65600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2926
timestamp 1654648307
transform 1 0 67100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2846
timestamp 1654648307
transform 1 0 67100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2927
timestamp 1654648307
transform 1 0 68600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2847
timestamp 1654648307
transform 1 0 68600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2928
timestamp 1654648307
transform 1 0 70100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2848
timestamp 1654648307
transform 1 0 70100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2929
timestamp 1654648307
transform 1 0 71600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2849
timestamp 1654648307
transform 1 0 71600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2930
timestamp 1654648307
transform 1 0 73100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2850
timestamp 1654648307
transform 1 0 73100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2931
timestamp 1654648307
transform 1 0 74600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2851
timestamp 1654648307
transform 1 0 74600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2932
timestamp 1654648307
transform 1 0 76100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2852
timestamp 1654648307
transform 1 0 76100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2933
timestamp 1654648307
transform 1 0 77600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2853
timestamp 1654648307
transform 1 0 77600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2934
timestamp 1654648307
transform 1 0 79100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2854
timestamp 1654648307
transform 1 0 79100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2935
timestamp 1654648307
transform 1 0 80600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2855
timestamp 1654648307
transform 1 0 80600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2936
timestamp 1654648307
transform 1 0 82100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2856
timestamp 1654648307
transform 1 0 82100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2937
timestamp 1654648307
transform 1 0 83600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2857
timestamp 1654648307
transform 1 0 83600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2938
timestamp 1654648307
transform 1 0 85100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2858
timestamp 1654648307
transform 1 0 85100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2939
timestamp 1654648307
transform 1 0 86600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2859
timestamp 1654648307
transform 1 0 86600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2940
timestamp 1654648307
transform 1 0 88100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2860
timestamp 1654648307
transform 1 0 88100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2941
timestamp 1654648307
transform 1 0 89600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2861
timestamp 1654648307
transform 1 0 89600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2942
timestamp 1654648307
transform 1 0 91100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2862
timestamp 1654648307
transform 1 0 91100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2943
timestamp 1654648307
transform 1 0 92600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2863
timestamp 1654648307
transform 1 0 92600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2944
timestamp 1654648307
transform 1 0 94100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2864
timestamp 1654648307
transform 1 0 94100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2945
timestamp 1654648307
transform 1 0 95600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2865
timestamp 1654648307
transform 1 0 95600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2946
timestamp 1654648307
transform 1 0 97100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2866
timestamp 1654648307
transform 1 0 97100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2947
timestamp 1654648307
transform 1 0 98600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2867
timestamp 1654648307
transform 1 0 98600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2948
timestamp 1654648307
transform 1 0 100100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2868
timestamp 1654648307
transform 1 0 100100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2949
timestamp 1654648307
transform 1 0 101600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2869
timestamp 1654648307
transform 1 0 101600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2950
timestamp 1654648307
transform 1 0 103100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2870
timestamp 1654648307
transform 1 0 103100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2951
timestamp 1654648307
transform 1 0 104600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2871
timestamp 1654648307
transform 1 0 104600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2952
timestamp 1654648307
transform 1 0 106100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2872
timestamp 1654648307
transform 1 0 106100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2953
timestamp 1654648307
transform 1 0 107600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2873
timestamp 1654648307
transform 1 0 107600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2954
timestamp 1654648307
transform 1 0 109100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2874
timestamp 1654648307
transform 1 0 109100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2955
timestamp 1654648307
transform 1 0 110600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2875
timestamp 1654648307
transform 1 0 110600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2956
timestamp 1654648307
transform 1 0 112100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2876
timestamp 1654648307
transform 1 0 112100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2957
timestamp 1654648307
transform 1 0 113600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2877
timestamp 1654648307
transform 1 0 113600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2958
timestamp 1654648307
transform 1 0 115100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2878
timestamp 1654648307
transform 1 0 115100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2959
timestamp 1654648307
transform 1 0 116600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_2879
timestamp 1654648307
transform 1 0 116600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_2720
timestamp 1654648307
transform 1 0 -1900 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2640
timestamp 1654648307
transform 1 0 -1900 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2722
timestamp 1654648307
transform 1 0 1100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2721
timestamp 1654648307
transform 1 0 -400 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2642
timestamp 1654648307
transform 1 0 1100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2641
timestamp 1654648307
transform 1 0 -400 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2724
timestamp 1654648307
transform 1 0 4100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2723
timestamp 1654648307
transform 1 0 2600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2644
timestamp 1654648307
transform 1 0 4100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2643
timestamp 1654648307
transform 1 0 2600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2726
timestamp 1654648307
transform 1 0 7100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2725
timestamp 1654648307
transform 1 0 5600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2646
timestamp 1654648307
transform 1 0 7100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2645
timestamp 1654648307
transform 1 0 5600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2728
timestamp 1654648307
transform 1 0 10100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2727
timestamp 1654648307
transform 1 0 8600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2648
timestamp 1654648307
transform 1 0 10100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2647
timestamp 1654648307
transform 1 0 8600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2730
timestamp 1654648307
transform 1 0 13100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2729
timestamp 1654648307
transform 1 0 11600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2650
timestamp 1654648307
transform 1 0 13100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2649
timestamp 1654648307
transform 1 0 11600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2732
timestamp 1654648307
transform 1 0 16100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2731
timestamp 1654648307
transform 1 0 14600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2652
timestamp 1654648307
transform 1 0 16100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2651
timestamp 1654648307
transform 1 0 14600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2734
timestamp 1654648307
transform 1 0 19100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2733
timestamp 1654648307
transform 1 0 17600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2654
timestamp 1654648307
transform 1 0 19100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2653
timestamp 1654648307
transform 1 0 17600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2735
timestamp 1654648307
transform 1 0 20600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2736
timestamp 1654648307
transform 1 0 22100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2655
timestamp 1654648307
transform 1 0 20600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2656
timestamp 1654648307
transform 1 0 22100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2737
timestamp 1654648307
transform 1 0 23600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2738
timestamp 1654648307
transform 1 0 25100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2657
timestamp 1654648307
transform 1 0 23600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2658
timestamp 1654648307
transform 1 0 25100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2739
timestamp 1654648307
transform 1 0 26600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2740
timestamp 1654648307
transform 1 0 28100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2659
timestamp 1654648307
transform 1 0 26600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2660
timestamp 1654648307
transform 1 0 28100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2741
timestamp 1654648307
transform 1 0 29600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2742
timestamp 1654648307
transform 1 0 31100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2661
timestamp 1654648307
transform 1 0 29600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2662
timestamp 1654648307
transform 1 0 31100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2743
timestamp 1654648307
transform 1 0 32600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2744
timestamp 1654648307
transform 1 0 34100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2663
timestamp 1654648307
transform 1 0 32600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2664
timestamp 1654648307
transform 1 0 34100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2745
timestamp 1654648307
transform 1 0 35600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2746
timestamp 1654648307
transform 1 0 37100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2665
timestamp 1654648307
transform 1 0 35600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2666
timestamp 1654648307
transform 1 0 37100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2747
timestamp 1654648307
transform 1 0 38600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2748
timestamp 1654648307
transform 1 0 40100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2667
timestamp 1654648307
transform 1 0 38600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2668
timestamp 1654648307
transform 1 0 40100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2749
timestamp 1654648307
transform 1 0 41600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2750
timestamp 1654648307
transform 1 0 43100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2669
timestamp 1654648307
transform 1 0 41600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2670
timestamp 1654648307
transform 1 0 43100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2751
timestamp 1654648307
transform 1 0 44600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2752
timestamp 1654648307
transform 1 0 46100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2671
timestamp 1654648307
transform 1 0 44600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2672
timestamp 1654648307
transform 1 0 46100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2753
timestamp 1654648307
transform 1 0 47600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2754
timestamp 1654648307
transform 1 0 49100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2673
timestamp 1654648307
transform 1 0 47600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2674
timestamp 1654648307
transform 1 0 49100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2755
timestamp 1654648307
transform 1 0 50600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2756
timestamp 1654648307
transform 1 0 52100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2675
timestamp 1654648307
transform 1 0 50600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2676
timestamp 1654648307
transform 1 0 52100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2757
timestamp 1654648307
transform 1 0 53600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2758
timestamp 1654648307
transform 1 0 55100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2677
timestamp 1654648307
transform 1 0 53600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2678
timestamp 1654648307
transform 1 0 55100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2759
timestamp 1654648307
transform 1 0 56600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2760
timestamp 1654648307
transform 1 0 58100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2679
timestamp 1654648307
transform 1 0 56600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2680
timestamp 1654648307
transform 1 0 58100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2761
timestamp 1654648307
transform 1 0 59600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2762
timestamp 1654648307
transform 1 0 61100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2681
timestamp 1654648307
transform 1 0 59600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2682
timestamp 1654648307
transform 1 0 61100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2763
timestamp 1654648307
transform 1 0 62600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2683
timestamp 1654648307
transform 1 0 62600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2764
timestamp 1654648307
transform 1 0 64100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2684
timestamp 1654648307
transform 1 0 64100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2765
timestamp 1654648307
transform 1 0 65600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2685
timestamp 1654648307
transform 1 0 65600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2766
timestamp 1654648307
transform 1 0 67100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2686
timestamp 1654648307
transform 1 0 67100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2767
timestamp 1654648307
transform 1 0 68600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2687
timestamp 1654648307
transform 1 0 68600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2768
timestamp 1654648307
transform 1 0 70100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2688
timestamp 1654648307
transform 1 0 70100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2769
timestamp 1654648307
transform 1 0 71600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2689
timestamp 1654648307
transform 1 0 71600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2770
timestamp 1654648307
transform 1 0 73100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2690
timestamp 1654648307
transform 1 0 73100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2771
timestamp 1654648307
transform 1 0 74600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2691
timestamp 1654648307
transform 1 0 74600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2772
timestamp 1654648307
transform 1 0 76100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2692
timestamp 1654648307
transform 1 0 76100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2773
timestamp 1654648307
transform 1 0 77600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2693
timestamp 1654648307
transform 1 0 77600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2774
timestamp 1654648307
transform 1 0 79100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2694
timestamp 1654648307
transform 1 0 79100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2775
timestamp 1654648307
transform 1 0 80600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2695
timestamp 1654648307
transform 1 0 80600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2776
timestamp 1654648307
transform 1 0 82100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2696
timestamp 1654648307
transform 1 0 82100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2777
timestamp 1654648307
transform 1 0 83600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2697
timestamp 1654648307
transform 1 0 83600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2778
timestamp 1654648307
transform 1 0 85100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2698
timestamp 1654648307
transform 1 0 85100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2779
timestamp 1654648307
transform 1 0 86600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2699
timestamp 1654648307
transform 1 0 86600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2780
timestamp 1654648307
transform 1 0 88100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2700
timestamp 1654648307
transform 1 0 88100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2781
timestamp 1654648307
transform 1 0 89600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2701
timestamp 1654648307
transform 1 0 89600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2782
timestamp 1654648307
transform 1 0 91100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2702
timestamp 1654648307
transform 1 0 91100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2783
timestamp 1654648307
transform 1 0 92600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2703
timestamp 1654648307
transform 1 0 92600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2784
timestamp 1654648307
transform 1 0 94100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2704
timestamp 1654648307
transform 1 0 94100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2785
timestamp 1654648307
transform 1 0 95600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2705
timestamp 1654648307
transform 1 0 95600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2786
timestamp 1654648307
transform 1 0 97100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2706
timestamp 1654648307
transform 1 0 97100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2787
timestamp 1654648307
transform 1 0 98600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2707
timestamp 1654648307
transform 1 0 98600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2788
timestamp 1654648307
transform 1 0 100100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2708
timestamp 1654648307
transform 1 0 100100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2789
timestamp 1654648307
transform 1 0 101600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2709
timestamp 1654648307
transform 1 0 101600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2790
timestamp 1654648307
transform 1 0 103100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2710
timestamp 1654648307
transform 1 0 103100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2791
timestamp 1654648307
transform 1 0 104600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2711
timestamp 1654648307
transform 1 0 104600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2792
timestamp 1654648307
transform 1 0 106100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2712
timestamp 1654648307
transform 1 0 106100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2793
timestamp 1654648307
transform 1 0 107600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2713
timestamp 1654648307
transform 1 0 107600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2794
timestamp 1654648307
transform 1 0 109100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2714
timestamp 1654648307
transform 1 0 109100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2795
timestamp 1654648307
transform 1 0 110600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2715
timestamp 1654648307
transform 1 0 110600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2796
timestamp 1654648307
transform 1 0 112100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2716
timestamp 1654648307
transform 1 0 112100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2797
timestamp 1654648307
transform 1 0 113600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2717
timestamp 1654648307
transform 1 0 113600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2798
timestamp 1654648307
transform 1 0 115100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2718
timestamp 1654648307
transform 1 0 115100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2799
timestamp 1654648307
transform 1 0 116600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_2719
timestamp 1654648307
transform 1 0 116600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_2560
timestamp 1654648307
transform 1 0 -1900 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2480
timestamp 1654648307
transform 1 0 -1900 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2562
timestamp 1654648307
transform 1 0 1100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2561
timestamp 1654648307
transform 1 0 -400 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2482
timestamp 1654648307
transform 1 0 1100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2481
timestamp 1654648307
transform 1 0 -400 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2564
timestamp 1654648307
transform 1 0 4100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2563
timestamp 1654648307
transform 1 0 2600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2484
timestamp 1654648307
transform 1 0 4100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2483
timestamp 1654648307
transform 1 0 2600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2566
timestamp 1654648307
transform 1 0 7100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2565
timestamp 1654648307
transform 1 0 5600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2486
timestamp 1654648307
transform 1 0 7100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2485
timestamp 1654648307
transform 1 0 5600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2568
timestamp 1654648307
transform 1 0 10100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2567
timestamp 1654648307
transform 1 0 8600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2488
timestamp 1654648307
transform 1 0 10100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2487
timestamp 1654648307
transform 1 0 8600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2570
timestamp 1654648307
transform 1 0 13100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2569
timestamp 1654648307
transform 1 0 11600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2490
timestamp 1654648307
transform 1 0 13100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2489
timestamp 1654648307
transform 1 0 11600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2572
timestamp 1654648307
transform 1 0 16100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2571
timestamp 1654648307
transform 1 0 14600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2492
timestamp 1654648307
transform 1 0 16100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2491
timestamp 1654648307
transform 1 0 14600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2574
timestamp 1654648307
transform 1 0 19100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2573
timestamp 1654648307
transform 1 0 17600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2494
timestamp 1654648307
transform 1 0 19100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2493
timestamp 1654648307
transform 1 0 17600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2575
timestamp 1654648307
transform 1 0 20600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2576
timestamp 1654648307
transform 1 0 22100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2495
timestamp 1654648307
transform 1 0 20600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2496
timestamp 1654648307
transform 1 0 22100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2577
timestamp 1654648307
transform 1 0 23600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2578
timestamp 1654648307
transform 1 0 25100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2497
timestamp 1654648307
transform 1 0 23600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2498
timestamp 1654648307
transform 1 0 25100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2579
timestamp 1654648307
transform 1 0 26600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2580
timestamp 1654648307
transform 1 0 28100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2499
timestamp 1654648307
transform 1 0 26600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2500
timestamp 1654648307
transform 1 0 28100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2581
timestamp 1654648307
transform 1 0 29600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2582
timestamp 1654648307
transform 1 0 31100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2501
timestamp 1654648307
transform 1 0 29600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2502
timestamp 1654648307
transform 1 0 31100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2583
timestamp 1654648307
transform 1 0 32600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2584
timestamp 1654648307
transform 1 0 34100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2503
timestamp 1654648307
transform 1 0 32600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2504
timestamp 1654648307
transform 1 0 34100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2585
timestamp 1654648307
transform 1 0 35600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2586
timestamp 1654648307
transform 1 0 37100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2505
timestamp 1654648307
transform 1 0 35600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2506
timestamp 1654648307
transform 1 0 37100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2587
timestamp 1654648307
transform 1 0 38600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2588
timestamp 1654648307
transform 1 0 40100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2507
timestamp 1654648307
transform 1 0 38600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2508
timestamp 1654648307
transform 1 0 40100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2589
timestamp 1654648307
transform 1 0 41600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2590
timestamp 1654648307
transform 1 0 43100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2509
timestamp 1654648307
transform 1 0 41600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2510
timestamp 1654648307
transform 1 0 43100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2591
timestamp 1654648307
transform 1 0 44600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2592
timestamp 1654648307
transform 1 0 46100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2511
timestamp 1654648307
transform 1 0 44600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2512
timestamp 1654648307
transform 1 0 46100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2593
timestamp 1654648307
transform 1 0 47600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2594
timestamp 1654648307
transform 1 0 49100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2513
timestamp 1654648307
transform 1 0 47600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2514
timestamp 1654648307
transform 1 0 49100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2595
timestamp 1654648307
transform 1 0 50600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2596
timestamp 1654648307
transform 1 0 52100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2515
timestamp 1654648307
transform 1 0 50600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2516
timestamp 1654648307
transform 1 0 52100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2597
timestamp 1654648307
transform 1 0 53600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2598
timestamp 1654648307
transform 1 0 55100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2517
timestamp 1654648307
transform 1 0 53600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2518
timestamp 1654648307
transform 1 0 55100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2599
timestamp 1654648307
transform 1 0 56600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2600
timestamp 1654648307
transform 1 0 58100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2519
timestamp 1654648307
transform 1 0 56600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2520
timestamp 1654648307
transform 1 0 58100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2601
timestamp 1654648307
transform 1 0 59600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2602
timestamp 1654648307
transform 1 0 61100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2521
timestamp 1654648307
transform 1 0 59600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2522
timestamp 1654648307
transform 1 0 61100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2603
timestamp 1654648307
transform 1 0 62600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2523
timestamp 1654648307
transform 1 0 62600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2604
timestamp 1654648307
transform 1 0 64100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2524
timestamp 1654648307
transform 1 0 64100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2605
timestamp 1654648307
transform 1 0 65600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2525
timestamp 1654648307
transform 1 0 65600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2606
timestamp 1654648307
transform 1 0 67100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2526
timestamp 1654648307
transform 1 0 67100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2607
timestamp 1654648307
transform 1 0 68600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2527
timestamp 1654648307
transform 1 0 68600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2608
timestamp 1654648307
transform 1 0 70100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2528
timestamp 1654648307
transform 1 0 70100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2609
timestamp 1654648307
transform 1 0 71600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2529
timestamp 1654648307
transform 1 0 71600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2610
timestamp 1654648307
transform 1 0 73100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2530
timestamp 1654648307
transform 1 0 73100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2611
timestamp 1654648307
transform 1 0 74600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2531
timestamp 1654648307
transform 1 0 74600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2612
timestamp 1654648307
transform 1 0 76100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2532
timestamp 1654648307
transform 1 0 76100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2613
timestamp 1654648307
transform 1 0 77600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2533
timestamp 1654648307
transform 1 0 77600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2614
timestamp 1654648307
transform 1 0 79100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2534
timestamp 1654648307
transform 1 0 79100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2615
timestamp 1654648307
transform 1 0 80600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2535
timestamp 1654648307
transform 1 0 80600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2616
timestamp 1654648307
transform 1 0 82100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2536
timestamp 1654648307
transform 1 0 82100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2617
timestamp 1654648307
transform 1 0 83600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2537
timestamp 1654648307
transform 1 0 83600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2618
timestamp 1654648307
transform 1 0 85100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2538
timestamp 1654648307
transform 1 0 85100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2619
timestamp 1654648307
transform 1 0 86600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2539
timestamp 1654648307
transform 1 0 86600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2620
timestamp 1654648307
transform 1 0 88100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2540
timestamp 1654648307
transform 1 0 88100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2621
timestamp 1654648307
transform 1 0 89600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2541
timestamp 1654648307
transform 1 0 89600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2622
timestamp 1654648307
transform 1 0 91100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2542
timestamp 1654648307
transform 1 0 91100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2623
timestamp 1654648307
transform 1 0 92600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2543
timestamp 1654648307
transform 1 0 92600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2624
timestamp 1654648307
transform 1 0 94100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2544
timestamp 1654648307
transform 1 0 94100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2625
timestamp 1654648307
transform 1 0 95600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2545
timestamp 1654648307
transform 1 0 95600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2626
timestamp 1654648307
transform 1 0 97100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2546
timestamp 1654648307
transform 1 0 97100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2627
timestamp 1654648307
transform 1 0 98600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2547
timestamp 1654648307
transform 1 0 98600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2628
timestamp 1654648307
transform 1 0 100100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2548
timestamp 1654648307
transform 1 0 100100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2629
timestamp 1654648307
transform 1 0 101600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2549
timestamp 1654648307
transform 1 0 101600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2630
timestamp 1654648307
transform 1 0 103100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2550
timestamp 1654648307
transform 1 0 103100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2631
timestamp 1654648307
transform 1 0 104600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2551
timestamp 1654648307
transform 1 0 104600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2632
timestamp 1654648307
transform 1 0 106100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2552
timestamp 1654648307
transform 1 0 106100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2633
timestamp 1654648307
transform 1 0 107600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2553
timestamp 1654648307
transform 1 0 107600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2634
timestamp 1654648307
transform 1 0 109100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2554
timestamp 1654648307
transform 1 0 109100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2635
timestamp 1654648307
transform 1 0 110600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2555
timestamp 1654648307
transform 1 0 110600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2636
timestamp 1654648307
transform 1 0 112100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2556
timestamp 1654648307
transform 1 0 112100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2637
timestamp 1654648307
transform 1 0 113600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2557
timestamp 1654648307
transform 1 0 113600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2638
timestamp 1654648307
transform 1 0 115100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2558
timestamp 1654648307
transform 1 0 115100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2639
timestamp 1654648307
transform 1 0 116600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_2559
timestamp 1654648307
transform 1 0 116600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_2400
timestamp 1654648307
transform 1 0 -1900 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2320
timestamp 1654648307
transform 1 0 -1900 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2402
timestamp 1654648307
transform 1 0 1100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2401
timestamp 1654648307
transform 1 0 -400 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2322
timestamp 1654648307
transform 1 0 1100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2321
timestamp 1654648307
transform 1 0 -400 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2404
timestamp 1654648307
transform 1 0 4100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2403
timestamp 1654648307
transform 1 0 2600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2324
timestamp 1654648307
transform 1 0 4100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2323
timestamp 1654648307
transform 1 0 2600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2406
timestamp 1654648307
transform 1 0 7100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2405
timestamp 1654648307
transform 1 0 5600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2326
timestamp 1654648307
transform 1 0 7100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2325
timestamp 1654648307
transform 1 0 5600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2408
timestamp 1654648307
transform 1 0 10100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2407
timestamp 1654648307
transform 1 0 8600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2328
timestamp 1654648307
transform 1 0 10100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2327
timestamp 1654648307
transform 1 0 8600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2410
timestamp 1654648307
transform 1 0 13100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2409
timestamp 1654648307
transform 1 0 11600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2330
timestamp 1654648307
transform 1 0 13100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2329
timestamp 1654648307
transform 1 0 11600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2412
timestamp 1654648307
transform 1 0 16100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2411
timestamp 1654648307
transform 1 0 14600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2332
timestamp 1654648307
transform 1 0 16100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2331
timestamp 1654648307
transform 1 0 14600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2414
timestamp 1654648307
transform 1 0 19100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2413
timestamp 1654648307
transform 1 0 17600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2334
timestamp 1654648307
transform 1 0 19100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2333
timestamp 1654648307
transform 1 0 17600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2415
timestamp 1654648307
transform 1 0 20600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2416
timestamp 1654648307
transform 1 0 22100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2335
timestamp 1654648307
transform 1 0 20600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2336
timestamp 1654648307
transform 1 0 22100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2417
timestamp 1654648307
transform 1 0 23600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2418
timestamp 1654648307
transform 1 0 25100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2337
timestamp 1654648307
transform 1 0 23600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2338
timestamp 1654648307
transform 1 0 25100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2419
timestamp 1654648307
transform 1 0 26600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2420
timestamp 1654648307
transform 1 0 28100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2339
timestamp 1654648307
transform 1 0 26600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2340
timestamp 1654648307
transform 1 0 28100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2421
timestamp 1654648307
transform 1 0 29600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2422
timestamp 1654648307
transform 1 0 31100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2341
timestamp 1654648307
transform 1 0 29600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2342
timestamp 1654648307
transform 1 0 31100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2423
timestamp 1654648307
transform 1 0 32600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2424
timestamp 1654648307
transform 1 0 34100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2343
timestamp 1654648307
transform 1 0 32600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2344
timestamp 1654648307
transform 1 0 34100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2425
timestamp 1654648307
transform 1 0 35600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2426
timestamp 1654648307
transform 1 0 37100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2345
timestamp 1654648307
transform 1 0 35600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2346
timestamp 1654648307
transform 1 0 37100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2427
timestamp 1654648307
transform 1 0 38600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2428
timestamp 1654648307
transform 1 0 40100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2347
timestamp 1654648307
transform 1 0 38600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2348
timestamp 1654648307
transform 1 0 40100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2429
timestamp 1654648307
transform 1 0 41600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2430
timestamp 1654648307
transform 1 0 43100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2349
timestamp 1654648307
transform 1 0 41600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2350
timestamp 1654648307
transform 1 0 43100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2431
timestamp 1654648307
transform 1 0 44600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2432
timestamp 1654648307
transform 1 0 46100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2351
timestamp 1654648307
transform 1 0 44600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2352
timestamp 1654648307
transform 1 0 46100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2433
timestamp 1654648307
transform 1 0 47600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2434
timestamp 1654648307
transform 1 0 49100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2353
timestamp 1654648307
transform 1 0 47600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2354
timestamp 1654648307
transform 1 0 49100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2435
timestamp 1654648307
transform 1 0 50600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2436
timestamp 1654648307
transform 1 0 52100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2355
timestamp 1654648307
transform 1 0 50600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2356
timestamp 1654648307
transform 1 0 52100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2437
timestamp 1654648307
transform 1 0 53600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2438
timestamp 1654648307
transform 1 0 55100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2357
timestamp 1654648307
transform 1 0 53600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2358
timestamp 1654648307
transform 1 0 55100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2439
timestamp 1654648307
transform 1 0 56600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2440
timestamp 1654648307
transform 1 0 58100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2359
timestamp 1654648307
transform 1 0 56600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2360
timestamp 1654648307
transform 1 0 58100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2441
timestamp 1654648307
transform 1 0 59600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2442
timestamp 1654648307
transform 1 0 61100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2361
timestamp 1654648307
transform 1 0 59600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2362
timestamp 1654648307
transform 1 0 61100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2443
timestamp 1654648307
transform 1 0 62600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2363
timestamp 1654648307
transform 1 0 62600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2444
timestamp 1654648307
transform 1 0 64100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2364
timestamp 1654648307
transform 1 0 64100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2445
timestamp 1654648307
transform 1 0 65600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2365
timestamp 1654648307
transform 1 0 65600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2446
timestamp 1654648307
transform 1 0 67100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2366
timestamp 1654648307
transform 1 0 67100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2447
timestamp 1654648307
transform 1 0 68600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2367
timestamp 1654648307
transform 1 0 68600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2448
timestamp 1654648307
transform 1 0 70100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2368
timestamp 1654648307
transform 1 0 70100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2449
timestamp 1654648307
transform 1 0 71600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2369
timestamp 1654648307
transform 1 0 71600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2450
timestamp 1654648307
transform 1 0 73100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2370
timestamp 1654648307
transform 1 0 73100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2451
timestamp 1654648307
transform 1 0 74600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2371
timestamp 1654648307
transform 1 0 74600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2452
timestamp 1654648307
transform 1 0 76100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2372
timestamp 1654648307
transform 1 0 76100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2453
timestamp 1654648307
transform 1 0 77600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2373
timestamp 1654648307
transform 1 0 77600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2454
timestamp 1654648307
transform 1 0 79100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2374
timestamp 1654648307
transform 1 0 79100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2455
timestamp 1654648307
transform 1 0 80600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2375
timestamp 1654648307
transform 1 0 80600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2456
timestamp 1654648307
transform 1 0 82100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2376
timestamp 1654648307
transform 1 0 82100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2457
timestamp 1654648307
transform 1 0 83600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2377
timestamp 1654648307
transform 1 0 83600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2458
timestamp 1654648307
transform 1 0 85100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2378
timestamp 1654648307
transform 1 0 85100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2459
timestamp 1654648307
transform 1 0 86600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2379
timestamp 1654648307
transform 1 0 86600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2460
timestamp 1654648307
transform 1 0 88100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2380
timestamp 1654648307
transform 1 0 88100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2461
timestamp 1654648307
transform 1 0 89600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2381
timestamp 1654648307
transform 1 0 89600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2462
timestamp 1654648307
transform 1 0 91100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2382
timestamp 1654648307
transform 1 0 91100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2463
timestamp 1654648307
transform 1 0 92600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2383
timestamp 1654648307
transform 1 0 92600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2464
timestamp 1654648307
transform 1 0 94100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2384
timestamp 1654648307
transform 1 0 94100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2465
timestamp 1654648307
transform 1 0 95600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2385
timestamp 1654648307
transform 1 0 95600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2466
timestamp 1654648307
transform 1 0 97100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2386
timestamp 1654648307
transform 1 0 97100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2467
timestamp 1654648307
transform 1 0 98600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2387
timestamp 1654648307
transform 1 0 98600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2468
timestamp 1654648307
transform 1 0 100100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2388
timestamp 1654648307
transform 1 0 100100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2469
timestamp 1654648307
transform 1 0 101600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2389
timestamp 1654648307
transform 1 0 101600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2470
timestamp 1654648307
transform 1 0 103100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2390
timestamp 1654648307
transform 1 0 103100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2471
timestamp 1654648307
transform 1 0 104600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2391
timestamp 1654648307
transform 1 0 104600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2472
timestamp 1654648307
transform 1 0 106100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2392
timestamp 1654648307
transform 1 0 106100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2473
timestamp 1654648307
transform 1 0 107600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2393
timestamp 1654648307
transform 1 0 107600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2474
timestamp 1654648307
transform 1 0 109100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2394
timestamp 1654648307
transform 1 0 109100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2475
timestamp 1654648307
transform 1 0 110600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2395
timestamp 1654648307
transform 1 0 110600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2476
timestamp 1654648307
transform 1 0 112100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2396
timestamp 1654648307
transform 1 0 112100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2477
timestamp 1654648307
transform 1 0 113600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2397
timestamp 1654648307
transform 1 0 113600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2478
timestamp 1654648307
transform 1 0 115100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2398
timestamp 1654648307
transform 1 0 115100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2479
timestamp 1654648307
transform 1 0 116600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_2399
timestamp 1654648307
transform 1 0 116600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2240
timestamp 1654648307
transform 1 0 -1900 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2160
timestamp 1654648307
transform 1 0 -1900 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2080
timestamp 1654648307
transform 1 0 -1900 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2242
timestamp 1654648307
transform 1 0 1100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2241
timestamp 1654648307
transform 1 0 -400 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2162
timestamp 1654648307
transform 1 0 1100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2161
timestamp 1654648307
transform 1 0 -400 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2082
timestamp 1654648307
transform 1 0 1100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2081
timestamp 1654648307
transform 1 0 -400 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2244
timestamp 1654648307
transform 1 0 4100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2243
timestamp 1654648307
transform 1 0 2600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2164
timestamp 1654648307
transform 1 0 4100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2163
timestamp 1654648307
transform 1 0 2600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2084
timestamp 1654648307
transform 1 0 4100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2083
timestamp 1654648307
transform 1 0 2600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2246
timestamp 1654648307
transform 1 0 7100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2245
timestamp 1654648307
transform 1 0 5600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2166
timestamp 1654648307
transform 1 0 7100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2165
timestamp 1654648307
transform 1 0 5600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2086
timestamp 1654648307
transform 1 0 7100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2085
timestamp 1654648307
transform 1 0 5600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2248
timestamp 1654648307
transform 1 0 10100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2247
timestamp 1654648307
transform 1 0 8600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2168
timestamp 1654648307
transform 1 0 10100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2167
timestamp 1654648307
transform 1 0 8600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2088
timestamp 1654648307
transform 1 0 10100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2087
timestamp 1654648307
transform 1 0 8600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2250
timestamp 1654648307
transform 1 0 13100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2249
timestamp 1654648307
transform 1 0 11600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2170
timestamp 1654648307
transform 1 0 13100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2169
timestamp 1654648307
transform 1 0 11600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2090
timestamp 1654648307
transform 1 0 13100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2089
timestamp 1654648307
transform 1 0 11600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2252
timestamp 1654648307
transform 1 0 16100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2251
timestamp 1654648307
transform 1 0 14600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2172
timestamp 1654648307
transform 1 0 16100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2171
timestamp 1654648307
transform 1 0 14600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2092
timestamp 1654648307
transform 1 0 16100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2091
timestamp 1654648307
transform 1 0 14600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2254
timestamp 1654648307
transform 1 0 19100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2253
timestamp 1654648307
transform 1 0 17600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2174
timestamp 1654648307
transform 1 0 19100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2173
timestamp 1654648307
transform 1 0 17600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2094
timestamp 1654648307
transform 1 0 19100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2093
timestamp 1654648307
transform 1 0 17600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2255
timestamp 1654648307
transform 1 0 20600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2256
timestamp 1654648307
transform 1 0 22100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2175
timestamp 1654648307
transform 1 0 20600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2176
timestamp 1654648307
transform 1 0 22100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2095
timestamp 1654648307
transform 1 0 20600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2096
timestamp 1654648307
transform 1 0 22100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2257
timestamp 1654648307
transform 1 0 23600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2258
timestamp 1654648307
transform 1 0 25100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2177
timestamp 1654648307
transform 1 0 23600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2178
timestamp 1654648307
transform 1 0 25100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2097
timestamp 1654648307
transform 1 0 23600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2098
timestamp 1654648307
transform 1 0 25100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2259
timestamp 1654648307
transform 1 0 26600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2260
timestamp 1654648307
transform 1 0 28100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2179
timestamp 1654648307
transform 1 0 26600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2180
timestamp 1654648307
transform 1 0 28100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2099
timestamp 1654648307
transform 1 0 26600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2100
timestamp 1654648307
transform 1 0 28100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2261
timestamp 1654648307
transform 1 0 29600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2262
timestamp 1654648307
transform 1 0 31100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2181
timestamp 1654648307
transform 1 0 29600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2182
timestamp 1654648307
transform 1 0 31100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2101
timestamp 1654648307
transform 1 0 29600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2102
timestamp 1654648307
transform 1 0 31100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2263
timestamp 1654648307
transform 1 0 32600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2264
timestamp 1654648307
transform 1 0 34100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2183
timestamp 1654648307
transform 1 0 32600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2184
timestamp 1654648307
transform 1 0 34100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2103
timestamp 1654648307
transform 1 0 32600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2104
timestamp 1654648307
transform 1 0 34100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2265
timestamp 1654648307
transform 1 0 35600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2266
timestamp 1654648307
transform 1 0 37100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2185
timestamp 1654648307
transform 1 0 35600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2186
timestamp 1654648307
transform 1 0 37100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2105
timestamp 1654648307
transform 1 0 35600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2106
timestamp 1654648307
transform 1 0 37100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2267
timestamp 1654648307
transform 1 0 38600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2268
timestamp 1654648307
transform 1 0 40100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2187
timestamp 1654648307
transform 1 0 38600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2188
timestamp 1654648307
transform 1 0 40100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2107
timestamp 1654648307
transform 1 0 38600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2108
timestamp 1654648307
transform 1 0 40100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2269
timestamp 1654648307
transform 1 0 41600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2270
timestamp 1654648307
transform 1 0 43100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2189
timestamp 1654648307
transform 1 0 41600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2190
timestamp 1654648307
transform 1 0 43100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2109
timestamp 1654648307
transform 1 0 41600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2110
timestamp 1654648307
transform 1 0 43100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2271
timestamp 1654648307
transform 1 0 44600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2272
timestamp 1654648307
transform 1 0 46100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2191
timestamp 1654648307
transform 1 0 44600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2192
timestamp 1654648307
transform 1 0 46100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2111
timestamp 1654648307
transform 1 0 44600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2112
timestamp 1654648307
transform 1 0 46100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2273
timestamp 1654648307
transform 1 0 47600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2274
timestamp 1654648307
transform 1 0 49100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2193
timestamp 1654648307
transform 1 0 47600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2194
timestamp 1654648307
transform 1 0 49100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2113
timestamp 1654648307
transform 1 0 47600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2114
timestamp 1654648307
transform 1 0 49100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2275
timestamp 1654648307
transform 1 0 50600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2276
timestamp 1654648307
transform 1 0 52100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2195
timestamp 1654648307
transform 1 0 50600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2196
timestamp 1654648307
transform 1 0 52100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2115
timestamp 1654648307
transform 1 0 50600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2116
timestamp 1654648307
transform 1 0 52100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2277
timestamp 1654648307
transform 1 0 53600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2278
timestamp 1654648307
transform 1 0 55100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2197
timestamp 1654648307
transform 1 0 53600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2198
timestamp 1654648307
transform 1 0 55100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2117
timestamp 1654648307
transform 1 0 53600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2118
timestamp 1654648307
transform 1 0 55100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2279
timestamp 1654648307
transform 1 0 56600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2280
timestamp 1654648307
transform 1 0 58100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2199
timestamp 1654648307
transform 1 0 56600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2200
timestamp 1654648307
transform 1 0 58100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2119
timestamp 1654648307
transform 1 0 56600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2120
timestamp 1654648307
transform 1 0 58100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2281
timestamp 1654648307
transform 1 0 59600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2282
timestamp 1654648307
transform 1 0 61100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2201
timestamp 1654648307
transform 1 0 59600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2202
timestamp 1654648307
transform 1 0 61100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2121
timestamp 1654648307
transform 1 0 59600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2122
timestamp 1654648307
transform 1 0 61100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2283
timestamp 1654648307
transform 1 0 62600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2203
timestamp 1654648307
transform 1 0 62600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2284
timestamp 1654648307
transform 1 0 64100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2204
timestamp 1654648307
transform 1 0 64100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2123
timestamp 1654648307
transform 1 0 62600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2124
timestamp 1654648307
transform 1 0 64100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2285
timestamp 1654648307
transform 1 0 65600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2205
timestamp 1654648307
transform 1 0 65600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2286
timestamp 1654648307
transform 1 0 67100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2206
timestamp 1654648307
transform 1 0 67100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2125
timestamp 1654648307
transform 1 0 65600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2126
timestamp 1654648307
transform 1 0 67100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2287
timestamp 1654648307
transform 1 0 68600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2207
timestamp 1654648307
transform 1 0 68600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2288
timestamp 1654648307
transform 1 0 70100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2208
timestamp 1654648307
transform 1 0 70100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2127
timestamp 1654648307
transform 1 0 68600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2128
timestamp 1654648307
transform 1 0 70100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2289
timestamp 1654648307
transform 1 0 71600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2209
timestamp 1654648307
transform 1 0 71600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2290
timestamp 1654648307
transform 1 0 73100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2210
timestamp 1654648307
transform 1 0 73100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2129
timestamp 1654648307
transform 1 0 71600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2130
timestamp 1654648307
transform 1 0 73100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2291
timestamp 1654648307
transform 1 0 74600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2211
timestamp 1654648307
transform 1 0 74600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2292
timestamp 1654648307
transform 1 0 76100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2212
timestamp 1654648307
transform 1 0 76100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2131
timestamp 1654648307
transform 1 0 74600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2132
timestamp 1654648307
transform 1 0 76100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2293
timestamp 1654648307
transform 1 0 77600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2213
timestamp 1654648307
transform 1 0 77600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2294
timestamp 1654648307
transform 1 0 79100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2214
timestamp 1654648307
transform 1 0 79100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2133
timestamp 1654648307
transform 1 0 77600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2134
timestamp 1654648307
transform 1 0 79100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2295
timestamp 1654648307
transform 1 0 80600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2215
timestamp 1654648307
transform 1 0 80600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2296
timestamp 1654648307
transform 1 0 82100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2216
timestamp 1654648307
transform 1 0 82100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2135
timestamp 1654648307
transform 1 0 80600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2136
timestamp 1654648307
transform 1 0 82100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2297
timestamp 1654648307
transform 1 0 83600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2217
timestamp 1654648307
transform 1 0 83600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2298
timestamp 1654648307
transform 1 0 85100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2218
timestamp 1654648307
transform 1 0 85100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2137
timestamp 1654648307
transform 1 0 83600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2138
timestamp 1654648307
transform 1 0 85100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2299
timestamp 1654648307
transform 1 0 86600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2219
timestamp 1654648307
transform 1 0 86600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2300
timestamp 1654648307
transform 1 0 88100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2220
timestamp 1654648307
transform 1 0 88100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2139
timestamp 1654648307
transform 1 0 86600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2140
timestamp 1654648307
transform 1 0 88100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2301
timestamp 1654648307
transform 1 0 89600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2221
timestamp 1654648307
transform 1 0 89600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2302
timestamp 1654648307
transform 1 0 91100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2222
timestamp 1654648307
transform 1 0 91100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2141
timestamp 1654648307
transform 1 0 89600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2142
timestamp 1654648307
transform 1 0 91100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2303
timestamp 1654648307
transform 1 0 92600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2223
timestamp 1654648307
transform 1 0 92600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2304
timestamp 1654648307
transform 1 0 94100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2224
timestamp 1654648307
transform 1 0 94100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2143
timestamp 1654648307
transform 1 0 92600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2144
timestamp 1654648307
transform 1 0 94100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2305
timestamp 1654648307
transform 1 0 95600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2225
timestamp 1654648307
transform 1 0 95600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2306
timestamp 1654648307
transform 1 0 97100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2226
timestamp 1654648307
transform 1 0 97100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2145
timestamp 1654648307
transform 1 0 95600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2146
timestamp 1654648307
transform 1 0 97100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2307
timestamp 1654648307
transform 1 0 98600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2227
timestamp 1654648307
transform 1 0 98600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2308
timestamp 1654648307
transform 1 0 100100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2228
timestamp 1654648307
transform 1 0 100100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2147
timestamp 1654648307
transform 1 0 98600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2148
timestamp 1654648307
transform 1 0 100100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2309
timestamp 1654648307
transform 1 0 101600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2229
timestamp 1654648307
transform 1 0 101600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2310
timestamp 1654648307
transform 1 0 103100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2230
timestamp 1654648307
transform 1 0 103100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2149
timestamp 1654648307
transform 1 0 101600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2150
timestamp 1654648307
transform 1 0 103100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2311
timestamp 1654648307
transform 1 0 104600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2231
timestamp 1654648307
transform 1 0 104600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2312
timestamp 1654648307
transform 1 0 106100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2232
timestamp 1654648307
transform 1 0 106100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2151
timestamp 1654648307
transform 1 0 104600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2152
timestamp 1654648307
transform 1 0 106100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2313
timestamp 1654648307
transform 1 0 107600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2233
timestamp 1654648307
transform 1 0 107600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2314
timestamp 1654648307
transform 1 0 109100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2234
timestamp 1654648307
transform 1 0 109100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2153
timestamp 1654648307
transform 1 0 107600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2154
timestamp 1654648307
transform 1 0 109100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2315
timestamp 1654648307
transform 1 0 110600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2235
timestamp 1654648307
transform 1 0 110600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2316
timestamp 1654648307
transform 1 0 112100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2236
timestamp 1654648307
transform 1 0 112100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2155
timestamp 1654648307
transform 1 0 110600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2156
timestamp 1654648307
transform 1 0 112100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2317
timestamp 1654648307
transform 1 0 113600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2237
timestamp 1654648307
transform 1 0 113600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2318
timestamp 1654648307
transform 1 0 115100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2238
timestamp 1654648307
transform 1 0 115100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2157
timestamp 1654648307
transform 1 0 113600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2158
timestamp 1654648307
transform 1 0 115100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2319
timestamp 1654648307
transform 1 0 116600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2239
timestamp 1654648307
transform 1 0 116600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2159
timestamp 1654648307
transform 1 0 116600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2000
timestamp 1654648307
transform 1 0 -1900 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1920
timestamp 1654648307
transform 1 0 -1900 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2002
timestamp 1654648307
transform 1 0 1100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2001
timestamp 1654648307
transform 1 0 -400 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1921
timestamp 1654648307
transform 1 0 -400 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1922
timestamp 1654648307
transform 1 0 1100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2004
timestamp 1654648307
transform 1 0 4100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2003
timestamp 1654648307
transform 1 0 2600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1923
timestamp 1654648307
transform 1 0 2600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1924
timestamp 1654648307
transform 1 0 4100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2006
timestamp 1654648307
transform 1 0 7100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2005
timestamp 1654648307
transform 1 0 5600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1925
timestamp 1654648307
transform 1 0 5600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1926
timestamp 1654648307
transform 1 0 7100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2008
timestamp 1654648307
transform 1 0 10100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2007
timestamp 1654648307
transform 1 0 8600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1927
timestamp 1654648307
transform 1 0 8600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1928
timestamp 1654648307
transform 1 0 10100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2010
timestamp 1654648307
transform 1 0 13100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2009
timestamp 1654648307
transform 1 0 11600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1929
timestamp 1654648307
transform 1 0 11600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1930
timestamp 1654648307
transform 1 0 13100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2012
timestamp 1654648307
transform 1 0 16100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2011
timestamp 1654648307
transform 1 0 14600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1931
timestamp 1654648307
transform 1 0 14600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1932
timestamp 1654648307
transform 1 0 16100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2014
timestamp 1654648307
transform 1 0 19100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2013
timestamp 1654648307
transform 1 0 17600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1933
timestamp 1654648307
transform 1 0 17600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1934
timestamp 1654648307
transform 1 0 19100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2015
timestamp 1654648307
transform 1 0 20600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2016
timestamp 1654648307
transform 1 0 22100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1935
timestamp 1654648307
transform 1 0 20600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1936
timestamp 1654648307
transform 1 0 22100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2017
timestamp 1654648307
transform 1 0 23600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2018
timestamp 1654648307
transform 1 0 25100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1937
timestamp 1654648307
transform 1 0 23600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1938
timestamp 1654648307
transform 1 0 25100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2019
timestamp 1654648307
transform 1 0 26600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2020
timestamp 1654648307
transform 1 0 28100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1939
timestamp 1654648307
transform 1 0 26600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1940
timestamp 1654648307
transform 1 0 28100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2021
timestamp 1654648307
transform 1 0 29600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2022
timestamp 1654648307
transform 1 0 31100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1941
timestamp 1654648307
transform 1 0 29600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1942
timestamp 1654648307
transform 1 0 31100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2023
timestamp 1654648307
transform 1 0 32600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2024
timestamp 1654648307
transform 1 0 34100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1943
timestamp 1654648307
transform 1 0 32600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1944
timestamp 1654648307
transform 1 0 34100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2025
timestamp 1654648307
transform 1 0 35600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2026
timestamp 1654648307
transform 1 0 37100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1945
timestamp 1654648307
transform 1 0 35600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1946
timestamp 1654648307
transform 1 0 37100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2027
timestamp 1654648307
transform 1 0 38600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2028
timestamp 1654648307
transform 1 0 40100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1947
timestamp 1654648307
transform 1 0 38600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1948
timestamp 1654648307
transform 1 0 40100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2029
timestamp 1654648307
transform 1 0 41600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2030
timestamp 1654648307
transform 1 0 43100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1949
timestamp 1654648307
transform 1 0 41600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1950
timestamp 1654648307
transform 1 0 43100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2031
timestamp 1654648307
transform 1 0 44600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2032
timestamp 1654648307
transform 1 0 46100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1951
timestamp 1654648307
transform 1 0 44600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1952
timestamp 1654648307
transform 1 0 46100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2033
timestamp 1654648307
transform 1 0 47600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2034
timestamp 1654648307
transform 1 0 49100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1953
timestamp 1654648307
transform 1 0 47600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1954
timestamp 1654648307
transform 1 0 49100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2035
timestamp 1654648307
transform 1 0 50600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2036
timestamp 1654648307
transform 1 0 52100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1955
timestamp 1654648307
transform 1 0 50600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1956
timestamp 1654648307
transform 1 0 52100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2037
timestamp 1654648307
transform 1 0 53600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2038
timestamp 1654648307
transform 1 0 55100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1957
timestamp 1654648307
transform 1 0 53600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1958
timestamp 1654648307
transform 1 0 55100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2039
timestamp 1654648307
transform 1 0 56600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2040
timestamp 1654648307
transform 1 0 58100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1959
timestamp 1654648307
transform 1 0 56600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1960
timestamp 1654648307
transform 1 0 58100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2041
timestamp 1654648307
transform 1 0 59600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2042
timestamp 1654648307
transform 1 0 61100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1961
timestamp 1654648307
transform 1 0 59600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1962
timestamp 1654648307
transform 1 0 61100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2043
timestamp 1654648307
transform 1 0 62600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2044
timestamp 1654648307
transform 1 0 64100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1963
timestamp 1654648307
transform 1 0 62600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1964
timestamp 1654648307
transform 1 0 64100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2045
timestamp 1654648307
transform 1 0 65600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2046
timestamp 1654648307
transform 1 0 67100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1965
timestamp 1654648307
transform 1 0 65600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1966
timestamp 1654648307
transform 1 0 67100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2047
timestamp 1654648307
transform 1 0 68600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2048
timestamp 1654648307
transform 1 0 70100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1967
timestamp 1654648307
transform 1 0 68600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1968
timestamp 1654648307
transform 1 0 70100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2049
timestamp 1654648307
transform 1 0 71600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2050
timestamp 1654648307
transform 1 0 73100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1969
timestamp 1654648307
transform 1 0 71600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1970
timestamp 1654648307
transform 1 0 73100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2051
timestamp 1654648307
transform 1 0 74600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2052
timestamp 1654648307
transform 1 0 76100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1971
timestamp 1654648307
transform 1 0 74600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1972
timestamp 1654648307
transform 1 0 76100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2053
timestamp 1654648307
transform 1 0 77600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2054
timestamp 1654648307
transform 1 0 79100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1973
timestamp 1654648307
transform 1 0 77600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1974
timestamp 1654648307
transform 1 0 79100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2055
timestamp 1654648307
transform 1 0 80600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2056
timestamp 1654648307
transform 1 0 82100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1975
timestamp 1654648307
transform 1 0 80600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1976
timestamp 1654648307
transform 1 0 82100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2057
timestamp 1654648307
transform 1 0 83600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2058
timestamp 1654648307
transform 1 0 85100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1977
timestamp 1654648307
transform 1 0 83600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1978
timestamp 1654648307
transform 1 0 85100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2059
timestamp 1654648307
transform 1 0 86600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2060
timestamp 1654648307
transform 1 0 88100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1979
timestamp 1654648307
transform 1 0 86600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1980
timestamp 1654648307
transform 1 0 88100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2061
timestamp 1654648307
transform 1 0 89600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2062
timestamp 1654648307
transform 1 0 91100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1981
timestamp 1654648307
transform 1 0 89600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1982
timestamp 1654648307
transform 1 0 91100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2063
timestamp 1654648307
transform 1 0 92600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2064
timestamp 1654648307
transform 1 0 94100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1983
timestamp 1654648307
transform 1 0 92600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1984
timestamp 1654648307
transform 1 0 94100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2065
timestamp 1654648307
transform 1 0 95600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2066
timestamp 1654648307
transform 1 0 97100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1985
timestamp 1654648307
transform 1 0 95600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1986
timestamp 1654648307
transform 1 0 97100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2067
timestamp 1654648307
transform 1 0 98600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2068
timestamp 1654648307
transform 1 0 100100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1987
timestamp 1654648307
transform 1 0 98600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1988
timestamp 1654648307
transform 1 0 100100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2069
timestamp 1654648307
transform 1 0 101600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2070
timestamp 1654648307
transform 1 0 103100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1989
timestamp 1654648307
transform 1 0 101600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1990
timestamp 1654648307
transform 1 0 103100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2071
timestamp 1654648307
transform 1 0 104600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2072
timestamp 1654648307
transform 1 0 106100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1991
timestamp 1654648307
transform 1 0 104600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1992
timestamp 1654648307
transform 1 0 106100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2073
timestamp 1654648307
transform 1 0 107600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2074
timestamp 1654648307
transform 1 0 109100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1993
timestamp 1654648307
transform 1 0 107600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1994
timestamp 1654648307
transform 1 0 109100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2075
timestamp 1654648307
transform 1 0 110600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2076
timestamp 1654648307
transform 1 0 112100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1995
timestamp 1654648307
transform 1 0 110600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1996
timestamp 1654648307
transform 1 0 112100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2077
timestamp 1654648307
transform 1 0 113600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2078
timestamp 1654648307
transform 1 0 115100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1997
timestamp 1654648307
transform 1 0 113600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1998
timestamp 1654648307
transform 1 0 115100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2079
timestamp 1654648307
transform 1 0 116600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_1999
timestamp 1654648307
transform 1 0 116600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_1840
timestamp 1654648307
transform 1 0 -1900 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1760
timestamp 1654648307
transform 1 0 -1900 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1841
timestamp 1654648307
transform 1 0 -400 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1842
timestamp 1654648307
transform 1 0 1100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1761
timestamp 1654648307
transform 1 0 -400 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1762
timestamp 1654648307
transform 1 0 1100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1843
timestamp 1654648307
transform 1 0 2600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1844
timestamp 1654648307
transform 1 0 4100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1763
timestamp 1654648307
transform 1 0 2600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1764
timestamp 1654648307
transform 1 0 4100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1845
timestamp 1654648307
transform 1 0 5600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1846
timestamp 1654648307
transform 1 0 7100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1765
timestamp 1654648307
transform 1 0 5600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1766
timestamp 1654648307
transform 1 0 7100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1847
timestamp 1654648307
transform 1 0 8600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1848
timestamp 1654648307
transform 1 0 10100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1767
timestamp 1654648307
transform 1 0 8600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1768
timestamp 1654648307
transform 1 0 10100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1849
timestamp 1654648307
transform 1 0 11600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1850
timestamp 1654648307
transform 1 0 13100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1769
timestamp 1654648307
transform 1 0 11600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1770
timestamp 1654648307
transform 1 0 13100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1851
timestamp 1654648307
transform 1 0 14600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1852
timestamp 1654648307
transform 1 0 16100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1771
timestamp 1654648307
transform 1 0 14600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1772
timestamp 1654648307
transform 1 0 16100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1853
timestamp 1654648307
transform 1 0 17600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1854
timestamp 1654648307
transform 1 0 19100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1773
timestamp 1654648307
transform 1 0 17600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1774
timestamp 1654648307
transform 1 0 19100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1855
timestamp 1654648307
transform 1 0 20600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1856
timestamp 1654648307
transform 1 0 22100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1775
timestamp 1654648307
transform 1 0 20600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1776
timestamp 1654648307
transform 1 0 22100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1857
timestamp 1654648307
transform 1 0 23600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1858
timestamp 1654648307
transform 1 0 25100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1777
timestamp 1654648307
transform 1 0 23600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1778
timestamp 1654648307
transform 1 0 25100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1859
timestamp 1654648307
transform 1 0 26600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1860
timestamp 1654648307
transform 1 0 28100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1779
timestamp 1654648307
transform 1 0 26600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1780
timestamp 1654648307
transform 1 0 28100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1861
timestamp 1654648307
transform 1 0 29600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1862
timestamp 1654648307
transform 1 0 31100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1781
timestamp 1654648307
transform 1 0 29600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1782
timestamp 1654648307
transform 1 0 31100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1863
timestamp 1654648307
transform 1 0 32600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1864
timestamp 1654648307
transform 1 0 34100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1783
timestamp 1654648307
transform 1 0 32600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1784
timestamp 1654648307
transform 1 0 34100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1865
timestamp 1654648307
transform 1 0 35600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1866
timestamp 1654648307
transform 1 0 37100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1785
timestamp 1654648307
transform 1 0 35600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1786
timestamp 1654648307
transform 1 0 37100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1867
timestamp 1654648307
transform 1 0 38600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1868
timestamp 1654648307
transform 1 0 40100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1787
timestamp 1654648307
transform 1 0 38600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1788
timestamp 1654648307
transform 1 0 40100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1869
timestamp 1654648307
transform 1 0 41600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1870
timestamp 1654648307
transform 1 0 43100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1789
timestamp 1654648307
transform 1 0 41600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1790
timestamp 1654648307
transform 1 0 43100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1871
timestamp 1654648307
transform 1 0 44600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1872
timestamp 1654648307
transform 1 0 46100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1791
timestamp 1654648307
transform 1 0 44600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1792
timestamp 1654648307
transform 1 0 46100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1873
timestamp 1654648307
transform 1 0 47600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1874
timestamp 1654648307
transform 1 0 49100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1793
timestamp 1654648307
transform 1 0 47600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1794
timestamp 1654648307
transform 1 0 49100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1875
timestamp 1654648307
transform 1 0 50600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1876
timestamp 1654648307
transform 1 0 52100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1795
timestamp 1654648307
transform 1 0 50600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1796
timestamp 1654648307
transform 1 0 52100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1877
timestamp 1654648307
transform 1 0 53600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1878
timestamp 1654648307
transform 1 0 55100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1797
timestamp 1654648307
transform 1 0 53600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1798
timestamp 1654648307
transform 1 0 55100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1879
timestamp 1654648307
transform 1 0 56600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1880
timestamp 1654648307
transform 1 0 58100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1799
timestamp 1654648307
transform 1 0 56600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1800
timestamp 1654648307
transform 1 0 58100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1881
timestamp 1654648307
transform 1 0 59600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1882
timestamp 1654648307
transform 1 0 61100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1801
timestamp 1654648307
transform 1 0 59600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1802
timestamp 1654648307
transform 1 0 61100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1883
timestamp 1654648307
transform 1 0 62600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1884
timestamp 1654648307
transform 1 0 64100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1803
timestamp 1654648307
transform 1 0 62600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1804
timestamp 1654648307
transform 1 0 64100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1885
timestamp 1654648307
transform 1 0 65600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1886
timestamp 1654648307
transform 1 0 67100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1805
timestamp 1654648307
transform 1 0 65600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1806
timestamp 1654648307
transform 1 0 67100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1887
timestamp 1654648307
transform 1 0 68600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1888
timestamp 1654648307
transform 1 0 70100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1807
timestamp 1654648307
transform 1 0 68600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1808
timestamp 1654648307
transform 1 0 70100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1889
timestamp 1654648307
transform 1 0 71600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1890
timestamp 1654648307
transform 1 0 73100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1809
timestamp 1654648307
transform 1 0 71600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1810
timestamp 1654648307
transform 1 0 73100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1891
timestamp 1654648307
transform 1 0 74600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1892
timestamp 1654648307
transform 1 0 76100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1811
timestamp 1654648307
transform 1 0 74600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1812
timestamp 1654648307
transform 1 0 76100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1893
timestamp 1654648307
transform 1 0 77600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1894
timestamp 1654648307
transform 1 0 79100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1813
timestamp 1654648307
transform 1 0 77600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1814
timestamp 1654648307
transform 1 0 79100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1895
timestamp 1654648307
transform 1 0 80600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1896
timestamp 1654648307
transform 1 0 82100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1815
timestamp 1654648307
transform 1 0 80600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1816
timestamp 1654648307
transform 1 0 82100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1897
timestamp 1654648307
transform 1 0 83600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1898
timestamp 1654648307
transform 1 0 85100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1817
timestamp 1654648307
transform 1 0 83600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1818
timestamp 1654648307
transform 1 0 85100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1899
timestamp 1654648307
transform 1 0 86600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1900
timestamp 1654648307
transform 1 0 88100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1819
timestamp 1654648307
transform 1 0 86600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1820
timestamp 1654648307
transform 1 0 88100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1901
timestamp 1654648307
transform 1 0 89600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1902
timestamp 1654648307
transform 1 0 91100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1821
timestamp 1654648307
transform 1 0 89600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1822
timestamp 1654648307
transform 1 0 91100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1903
timestamp 1654648307
transform 1 0 92600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1904
timestamp 1654648307
transform 1 0 94100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1823
timestamp 1654648307
transform 1 0 92600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1824
timestamp 1654648307
transform 1 0 94100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1905
timestamp 1654648307
transform 1 0 95600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1906
timestamp 1654648307
transform 1 0 97100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1825
timestamp 1654648307
transform 1 0 95600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1826
timestamp 1654648307
transform 1 0 97100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1907
timestamp 1654648307
transform 1 0 98600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1908
timestamp 1654648307
transform 1 0 100100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1827
timestamp 1654648307
transform 1 0 98600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1828
timestamp 1654648307
transform 1 0 100100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1909
timestamp 1654648307
transform 1 0 101600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1910
timestamp 1654648307
transform 1 0 103100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1829
timestamp 1654648307
transform 1 0 101600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1830
timestamp 1654648307
transform 1 0 103100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1911
timestamp 1654648307
transform 1 0 104600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1912
timestamp 1654648307
transform 1 0 106100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1831
timestamp 1654648307
transform 1 0 104600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1832
timestamp 1654648307
transform 1 0 106100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1913
timestamp 1654648307
transform 1 0 107600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1914
timestamp 1654648307
transform 1 0 109100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1833
timestamp 1654648307
transform 1 0 107600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1834
timestamp 1654648307
transform 1 0 109100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1915
timestamp 1654648307
transform 1 0 110600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1916
timestamp 1654648307
transform 1 0 112100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1835
timestamp 1654648307
transform 1 0 110600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1836
timestamp 1654648307
transform 1 0 112100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1917
timestamp 1654648307
transform 1 0 113600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1918
timestamp 1654648307
transform 1 0 115100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1837
timestamp 1654648307
transform 1 0 113600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1838
timestamp 1654648307
transform 1 0 115100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1919
timestamp 1654648307
transform 1 0 116600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_1839
timestamp 1654648307
transform 1 0 116600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_1680
timestamp 1654648307
transform 1 0 -1900 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1600
timestamp 1654648307
transform 1 0 -1900 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1681
timestamp 1654648307
transform 1 0 -400 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1682
timestamp 1654648307
transform 1 0 1100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1601
timestamp 1654648307
transform 1 0 -400 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1602
timestamp 1654648307
transform 1 0 1100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1683
timestamp 1654648307
transform 1 0 2600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1684
timestamp 1654648307
transform 1 0 4100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1603
timestamp 1654648307
transform 1 0 2600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1604
timestamp 1654648307
transform 1 0 4100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1685
timestamp 1654648307
transform 1 0 5600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1686
timestamp 1654648307
transform 1 0 7100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1605
timestamp 1654648307
transform 1 0 5600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1606
timestamp 1654648307
transform 1 0 7100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1687
timestamp 1654648307
transform 1 0 8600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1688
timestamp 1654648307
transform 1 0 10100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1607
timestamp 1654648307
transform 1 0 8600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1608
timestamp 1654648307
transform 1 0 10100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1689
timestamp 1654648307
transform 1 0 11600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1690
timestamp 1654648307
transform 1 0 13100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1609
timestamp 1654648307
transform 1 0 11600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1610
timestamp 1654648307
transform 1 0 13100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1691
timestamp 1654648307
transform 1 0 14600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1692
timestamp 1654648307
transform 1 0 16100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1611
timestamp 1654648307
transform 1 0 14600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1612
timestamp 1654648307
transform 1 0 16100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1693
timestamp 1654648307
transform 1 0 17600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1694
timestamp 1654648307
transform 1 0 19100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1613
timestamp 1654648307
transform 1 0 17600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1614
timestamp 1654648307
transform 1 0 19100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1695
timestamp 1654648307
transform 1 0 20600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1696
timestamp 1654648307
transform 1 0 22100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1615
timestamp 1654648307
transform 1 0 20600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1616
timestamp 1654648307
transform 1 0 22100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1697
timestamp 1654648307
transform 1 0 23600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1698
timestamp 1654648307
transform 1 0 25100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1617
timestamp 1654648307
transform 1 0 23600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1618
timestamp 1654648307
transform 1 0 25100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1699
timestamp 1654648307
transform 1 0 26600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1700
timestamp 1654648307
transform 1 0 28100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1619
timestamp 1654648307
transform 1 0 26600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1620
timestamp 1654648307
transform 1 0 28100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1701
timestamp 1654648307
transform 1 0 29600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1702
timestamp 1654648307
transform 1 0 31100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1621
timestamp 1654648307
transform 1 0 29600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1622
timestamp 1654648307
transform 1 0 31100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1703
timestamp 1654648307
transform 1 0 32600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1704
timestamp 1654648307
transform 1 0 34100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1623
timestamp 1654648307
transform 1 0 32600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1624
timestamp 1654648307
transform 1 0 34100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1705
timestamp 1654648307
transform 1 0 35600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1706
timestamp 1654648307
transform 1 0 37100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1625
timestamp 1654648307
transform 1 0 35600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1626
timestamp 1654648307
transform 1 0 37100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1707
timestamp 1654648307
transform 1 0 38600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1708
timestamp 1654648307
transform 1 0 40100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1627
timestamp 1654648307
transform 1 0 38600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1628
timestamp 1654648307
transform 1 0 40100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1709
timestamp 1654648307
transform 1 0 41600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1710
timestamp 1654648307
transform 1 0 43100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1629
timestamp 1654648307
transform 1 0 41600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1630
timestamp 1654648307
transform 1 0 43100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1711
timestamp 1654648307
transform 1 0 44600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1712
timestamp 1654648307
transform 1 0 46100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1631
timestamp 1654648307
transform 1 0 44600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1632
timestamp 1654648307
transform 1 0 46100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1713
timestamp 1654648307
transform 1 0 47600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1714
timestamp 1654648307
transform 1 0 49100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1633
timestamp 1654648307
transform 1 0 47600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1634
timestamp 1654648307
transform 1 0 49100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1715
timestamp 1654648307
transform 1 0 50600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1716
timestamp 1654648307
transform 1 0 52100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1635
timestamp 1654648307
transform 1 0 50600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1636
timestamp 1654648307
transform 1 0 52100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1717
timestamp 1654648307
transform 1 0 53600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1718
timestamp 1654648307
transform 1 0 55100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1637
timestamp 1654648307
transform 1 0 53600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1638
timestamp 1654648307
transform 1 0 55100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1719
timestamp 1654648307
transform 1 0 56600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1720
timestamp 1654648307
transform 1 0 58100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1639
timestamp 1654648307
transform 1 0 56600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1640
timestamp 1654648307
transform 1 0 58100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1721
timestamp 1654648307
transform 1 0 59600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1722
timestamp 1654648307
transform 1 0 61100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1641
timestamp 1654648307
transform 1 0 59600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1642
timestamp 1654648307
transform 1 0 61100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1723
timestamp 1654648307
transform 1 0 62600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1724
timestamp 1654648307
transform 1 0 64100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1643
timestamp 1654648307
transform 1 0 62600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1644
timestamp 1654648307
transform 1 0 64100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1725
timestamp 1654648307
transform 1 0 65600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1726
timestamp 1654648307
transform 1 0 67100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1645
timestamp 1654648307
transform 1 0 65600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1646
timestamp 1654648307
transform 1 0 67100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1727
timestamp 1654648307
transform 1 0 68600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1728
timestamp 1654648307
transform 1 0 70100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1647
timestamp 1654648307
transform 1 0 68600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1648
timestamp 1654648307
transform 1 0 70100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1729
timestamp 1654648307
transform 1 0 71600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1730
timestamp 1654648307
transform 1 0 73100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1649
timestamp 1654648307
transform 1 0 71600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1650
timestamp 1654648307
transform 1 0 73100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1731
timestamp 1654648307
transform 1 0 74600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1732
timestamp 1654648307
transform 1 0 76100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1651
timestamp 1654648307
transform 1 0 74600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1652
timestamp 1654648307
transform 1 0 76100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1733
timestamp 1654648307
transform 1 0 77600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1734
timestamp 1654648307
transform 1 0 79100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1653
timestamp 1654648307
transform 1 0 77600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1654
timestamp 1654648307
transform 1 0 79100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1735
timestamp 1654648307
transform 1 0 80600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1736
timestamp 1654648307
transform 1 0 82100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1655
timestamp 1654648307
transform 1 0 80600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1656
timestamp 1654648307
transform 1 0 82100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1737
timestamp 1654648307
transform 1 0 83600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1738
timestamp 1654648307
transform 1 0 85100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1657
timestamp 1654648307
transform 1 0 83600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1658
timestamp 1654648307
transform 1 0 85100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1739
timestamp 1654648307
transform 1 0 86600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1740
timestamp 1654648307
transform 1 0 88100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1659
timestamp 1654648307
transform 1 0 86600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1660
timestamp 1654648307
transform 1 0 88100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1741
timestamp 1654648307
transform 1 0 89600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1742
timestamp 1654648307
transform 1 0 91100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1661
timestamp 1654648307
transform 1 0 89600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1662
timestamp 1654648307
transform 1 0 91100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1743
timestamp 1654648307
transform 1 0 92600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1744
timestamp 1654648307
transform 1 0 94100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1663
timestamp 1654648307
transform 1 0 92600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1664
timestamp 1654648307
transform 1 0 94100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1745
timestamp 1654648307
transform 1 0 95600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1746
timestamp 1654648307
transform 1 0 97100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1665
timestamp 1654648307
transform 1 0 95600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1666
timestamp 1654648307
transform 1 0 97100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1747
timestamp 1654648307
transform 1 0 98600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1748
timestamp 1654648307
transform 1 0 100100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1667
timestamp 1654648307
transform 1 0 98600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1668
timestamp 1654648307
transform 1 0 100100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1749
timestamp 1654648307
transform 1 0 101600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1750
timestamp 1654648307
transform 1 0 103100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1669
timestamp 1654648307
transform 1 0 101600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1670
timestamp 1654648307
transform 1 0 103100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1751
timestamp 1654648307
transform 1 0 104600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1752
timestamp 1654648307
transform 1 0 106100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1671
timestamp 1654648307
transform 1 0 104600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1672
timestamp 1654648307
transform 1 0 106100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1753
timestamp 1654648307
transform 1 0 107600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1754
timestamp 1654648307
transform 1 0 109100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1673
timestamp 1654648307
transform 1 0 107600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1674
timestamp 1654648307
transform 1 0 109100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1755
timestamp 1654648307
transform 1 0 110600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1756
timestamp 1654648307
transform 1 0 112100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1675
timestamp 1654648307
transform 1 0 110600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1676
timestamp 1654648307
transform 1 0 112100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1757
timestamp 1654648307
transform 1 0 113600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1758
timestamp 1654648307
transform 1 0 115100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1677
timestamp 1654648307
transform 1 0 113600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1678
timestamp 1654648307
transform 1 0 115100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1759
timestamp 1654648307
transform 1 0 116600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_1679
timestamp 1654648307
transform 1 0 116600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_1520
timestamp 1654648307
transform 1 0 -1900 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1440
timestamp 1654648307
transform 1 0 -1900 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1521
timestamp 1654648307
transform 1 0 -400 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1522
timestamp 1654648307
transform 1 0 1100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1441
timestamp 1654648307
transform 1 0 -400 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1442
timestamp 1654648307
transform 1 0 1100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1523
timestamp 1654648307
transform 1 0 2600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1524
timestamp 1654648307
transform 1 0 4100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1443
timestamp 1654648307
transform 1 0 2600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1444
timestamp 1654648307
transform 1 0 4100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1525
timestamp 1654648307
transform 1 0 5600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1526
timestamp 1654648307
transform 1 0 7100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1445
timestamp 1654648307
transform 1 0 5600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1446
timestamp 1654648307
transform 1 0 7100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1527
timestamp 1654648307
transform 1 0 8600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1528
timestamp 1654648307
transform 1 0 10100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1447
timestamp 1654648307
transform 1 0 8600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1448
timestamp 1654648307
transform 1 0 10100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1529
timestamp 1654648307
transform 1 0 11600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1530
timestamp 1654648307
transform 1 0 13100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1449
timestamp 1654648307
transform 1 0 11600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1450
timestamp 1654648307
transform 1 0 13100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1531
timestamp 1654648307
transform 1 0 14600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1532
timestamp 1654648307
transform 1 0 16100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1451
timestamp 1654648307
transform 1 0 14600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1452
timestamp 1654648307
transform 1 0 16100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1533
timestamp 1654648307
transform 1 0 17600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1534
timestamp 1654648307
transform 1 0 19100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1453
timestamp 1654648307
transform 1 0 17600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1454
timestamp 1654648307
transform 1 0 19100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1535
timestamp 1654648307
transform 1 0 20600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1536
timestamp 1654648307
transform 1 0 22100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1455
timestamp 1654648307
transform 1 0 20600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1456
timestamp 1654648307
transform 1 0 22100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1537
timestamp 1654648307
transform 1 0 23600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1538
timestamp 1654648307
transform 1 0 25100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1457
timestamp 1654648307
transform 1 0 23600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1458
timestamp 1654648307
transform 1 0 25100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1539
timestamp 1654648307
transform 1 0 26600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1540
timestamp 1654648307
transform 1 0 28100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1459
timestamp 1654648307
transform 1 0 26600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1460
timestamp 1654648307
transform 1 0 28100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1541
timestamp 1654648307
transform 1 0 29600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1542
timestamp 1654648307
transform 1 0 31100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1461
timestamp 1654648307
transform 1 0 29600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1462
timestamp 1654648307
transform 1 0 31100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1543
timestamp 1654648307
transform 1 0 32600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1544
timestamp 1654648307
transform 1 0 34100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1463
timestamp 1654648307
transform 1 0 32600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1464
timestamp 1654648307
transform 1 0 34100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1545
timestamp 1654648307
transform 1 0 35600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1546
timestamp 1654648307
transform 1 0 37100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1465
timestamp 1654648307
transform 1 0 35600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1466
timestamp 1654648307
transform 1 0 37100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1547
timestamp 1654648307
transform 1 0 38600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1548
timestamp 1654648307
transform 1 0 40100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1467
timestamp 1654648307
transform 1 0 38600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1468
timestamp 1654648307
transform 1 0 40100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1549
timestamp 1654648307
transform 1 0 41600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1550
timestamp 1654648307
transform 1 0 43100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1469
timestamp 1654648307
transform 1 0 41600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1470
timestamp 1654648307
transform 1 0 43100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1551
timestamp 1654648307
transform 1 0 44600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1552
timestamp 1654648307
transform 1 0 46100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1471
timestamp 1654648307
transform 1 0 44600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1472
timestamp 1654648307
transform 1 0 46100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1553
timestamp 1654648307
transform 1 0 47600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1554
timestamp 1654648307
transform 1 0 49100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1473
timestamp 1654648307
transform 1 0 47600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1474
timestamp 1654648307
transform 1 0 49100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1555
timestamp 1654648307
transform 1 0 50600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1556
timestamp 1654648307
transform 1 0 52100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1475
timestamp 1654648307
transform 1 0 50600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1476
timestamp 1654648307
transform 1 0 52100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1557
timestamp 1654648307
transform 1 0 53600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1558
timestamp 1654648307
transform 1 0 55100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1477
timestamp 1654648307
transform 1 0 53600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1478
timestamp 1654648307
transform 1 0 55100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1559
timestamp 1654648307
transform 1 0 56600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1560
timestamp 1654648307
transform 1 0 58100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1479
timestamp 1654648307
transform 1 0 56600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1480
timestamp 1654648307
transform 1 0 58100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1561
timestamp 1654648307
transform 1 0 59600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1562
timestamp 1654648307
transform 1 0 61100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1481
timestamp 1654648307
transform 1 0 59600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1482
timestamp 1654648307
transform 1 0 61100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1563
timestamp 1654648307
transform 1 0 62600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1564
timestamp 1654648307
transform 1 0 64100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1483
timestamp 1654648307
transform 1 0 62600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1484
timestamp 1654648307
transform 1 0 64100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1565
timestamp 1654648307
transform 1 0 65600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1566
timestamp 1654648307
transform 1 0 67100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1485
timestamp 1654648307
transform 1 0 65600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1486
timestamp 1654648307
transform 1 0 67100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1567
timestamp 1654648307
transform 1 0 68600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1568
timestamp 1654648307
transform 1 0 70100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1487
timestamp 1654648307
transform 1 0 68600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1488
timestamp 1654648307
transform 1 0 70100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1569
timestamp 1654648307
transform 1 0 71600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1570
timestamp 1654648307
transform 1 0 73100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1489
timestamp 1654648307
transform 1 0 71600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1490
timestamp 1654648307
transform 1 0 73100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1571
timestamp 1654648307
transform 1 0 74600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1572
timestamp 1654648307
transform 1 0 76100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1491
timestamp 1654648307
transform 1 0 74600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1492
timestamp 1654648307
transform 1 0 76100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1573
timestamp 1654648307
transform 1 0 77600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1574
timestamp 1654648307
transform 1 0 79100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1493
timestamp 1654648307
transform 1 0 77600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1494
timestamp 1654648307
transform 1 0 79100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1575
timestamp 1654648307
transform 1 0 80600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1576
timestamp 1654648307
transform 1 0 82100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1495
timestamp 1654648307
transform 1 0 80600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1496
timestamp 1654648307
transform 1 0 82100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1577
timestamp 1654648307
transform 1 0 83600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1578
timestamp 1654648307
transform 1 0 85100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1497
timestamp 1654648307
transform 1 0 83600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1498
timestamp 1654648307
transform 1 0 85100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1579
timestamp 1654648307
transform 1 0 86600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1580
timestamp 1654648307
transform 1 0 88100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1499
timestamp 1654648307
transform 1 0 86600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1500
timestamp 1654648307
transform 1 0 88100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1581
timestamp 1654648307
transform 1 0 89600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1582
timestamp 1654648307
transform 1 0 91100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1501
timestamp 1654648307
transform 1 0 89600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1502
timestamp 1654648307
transform 1 0 91100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1583
timestamp 1654648307
transform 1 0 92600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1584
timestamp 1654648307
transform 1 0 94100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1503
timestamp 1654648307
transform 1 0 92600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1504
timestamp 1654648307
transform 1 0 94100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1585
timestamp 1654648307
transform 1 0 95600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1586
timestamp 1654648307
transform 1 0 97100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1505
timestamp 1654648307
transform 1 0 95600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1506
timestamp 1654648307
transform 1 0 97100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1587
timestamp 1654648307
transform 1 0 98600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1588
timestamp 1654648307
transform 1 0 100100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1507
timestamp 1654648307
transform 1 0 98600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1508
timestamp 1654648307
transform 1 0 100100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1589
timestamp 1654648307
transform 1 0 101600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1590
timestamp 1654648307
transform 1 0 103100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1509
timestamp 1654648307
transform 1 0 101600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1510
timestamp 1654648307
transform 1 0 103100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1591
timestamp 1654648307
transform 1 0 104600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1592
timestamp 1654648307
transform 1 0 106100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1511
timestamp 1654648307
transform 1 0 104600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1512
timestamp 1654648307
transform 1 0 106100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1593
timestamp 1654648307
transform 1 0 107600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1594
timestamp 1654648307
transform 1 0 109100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1513
timestamp 1654648307
transform 1 0 107600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1514
timestamp 1654648307
transform 1 0 109100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1595
timestamp 1654648307
transform 1 0 110600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1596
timestamp 1654648307
transform 1 0 112100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1515
timestamp 1654648307
transform 1 0 110600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1516
timestamp 1654648307
transform 1 0 112100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1597
timestamp 1654648307
transform 1 0 113600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1598
timestamp 1654648307
transform 1 0 115100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1517
timestamp 1654648307
transform 1 0 113600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1518
timestamp 1654648307
transform 1 0 115100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1599
timestamp 1654648307
transform 1 0 116600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1519
timestamp 1654648307
transform 1 0 116600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1360
timestamp 1654648307
transform 1 0 -1900 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1280
timestamp 1654648307
transform 1 0 -1900 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1361
timestamp 1654648307
transform 1 0 -400 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1362
timestamp 1654648307
transform 1 0 1100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1281
timestamp 1654648307
transform 1 0 -400 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1282
timestamp 1654648307
transform 1 0 1100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1363
timestamp 1654648307
transform 1 0 2600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1364
timestamp 1654648307
transform 1 0 4100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1283
timestamp 1654648307
transform 1 0 2600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1284
timestamp 1654648307
transform 1 0 4100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1365
timestamp 1654648307
transform 1 0 5600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1366
timestamp 1654648307
transform 1 0 7100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1285
timestamp 1654648307
transform 1 0 5600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1286
timestamp 1654648307
transform 1 0 7100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1367
timestamp 1654648307
transform 1 0 8600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1368
timestamp 1654648307
transform 1 0 10100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1287
timestamp 1654648307
transform 1 0 8600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1288
timestamp 1654648307
transform 1 0 10100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1369
timestamp 1654648307
transform 1 0 11600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1370
timestamp 1654648307
transform 1 0 13100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1289
timestamp 1654648307
transform 1 0 11600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1290
timestamp 1654648307
transform 1 0 13100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1371
timestamp 1654648307
transform 1 0 14600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1372
timestamp 1654648307
transform 1 0 16100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1291
timestamp 1654648307
transform 1 0 14600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1292
timestamp 1654648307
transform 1 0 16100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1373
timestamp 1654648307
transform 1 0 17600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1374
timestamp 1654648307
transform 1 0 19100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1293
timestamp 1654648307
transform 1 0 17600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1294
timestamp 1654648307
transform 1 0 19100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1375
timestamp 1654648307
transform 1 0 20600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1376
timestamp 1654648307
transform 1 0 22100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1295
timestamp 1654648307
transform 1 0 20600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1296
timestamp 1654648307
transform 1 0 22100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1377
timestamp 1654648307
transform 1 0 23600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1378
timestamp 1654648307
transform 1 0 25100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1297
timestamp 1654648307
transform 1 0 23600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1298
timestamp 1654648307
transform 1 0 25100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1379
timestamp 1654648307
transform 1 0 26600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1380
timestamp 1654648307
transform 1 0 28100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1299
timestamp 1654648307
transform 1 0 26600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1300
timestamp 1654648307
transform 1 0 28100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1381
timestamp 1654648307
transform 1 0 29600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1382
timestamp 1654648307
transform 1 0 31100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1301
timestamp 1654648307
transform 1 0 29600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1302
timestamp 1654648307
transform 1 0 31100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1383
timestamp 1654648307
transform 1 0 32600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1384
timestamp 1654648307
transform 1 0 34100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1303
timestamp 1654648307
transform 1 0 32600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1304
timestamp 1654648307
transform 1 0 34100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1385
timestamp 1654648307
transform 1 0 35600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1386
timestamp 1654648307
transform 1 0 37100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1305
timestamp 1654648307
transform 1 0 35600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1306
timestamp 1654648307
transform 1 0 37100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1387
timestamp 1654648307
transform 1 0 38600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1388
timestamp 1654648307
transform 1 0 40100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1307
timestamp 1654648307
transform 1 0 38600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1308
timestamp 1654648307
transform 1 0 40100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1389
timestamp 1654648307
transform 1 0 41600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1390
timestamp 1654648307
transform 1 0 43100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1309
timestamp 1654648307
transform 1 0 41600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1310
timestamp 1654648307
transform 1 0 43100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1391
timestamp 1654648307
transform 1 0 44600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1392
timestamp 1654648307
transform 1 0 46100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1311
timestamp 1654648307
transform 1 0 44600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1312
timestamp 1654648307
transform 1 0 46100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1393
timestamp 1654648307
transform 1 0 47600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1394
timestamp 1654648307
transform 1 0 49100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1313
timestamp 1654648307
transform 1 0 47600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1314
timestamp 1654648307
transform 1 0 49100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1395
timestamp 1654648307
transform 1 0 50600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1396
timestamp 1654648307
transform 1 0 52100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1315
timestamp 1654648307
transform 1 0 50600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1316
timestamp 1654648307
transform 1 0 52100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1397
timestamp 1654648307
transform 1 0 53600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1398
timestamp 1654648307
transform 1 0 55100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1317
timestamp 1654648307
transform 1 0 53600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1318
timestamp 1654648307
transform 1 0 55100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1399
timestamp 1654648307
transform 1 0 56600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1400
timestamp 1654648307
transform 1 0 58100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1319
timestamp 1654648307
transform 1 0 56600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1320
timestamp 1654648307
transform 1 0 58100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1401
timestamp 1654648307
transform 1 0 59600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1402
timestamp 1654648307
transform 1 0 61100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1321
timestamp 1654648307
transform 1 0 59600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1322
timestamp 1654648307
transform 1 0 61100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1403
timestamp 1654648307
transform 1 0 62600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1404
timestamp 1654648307
transform 1 0 64100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1323
timestamp 1654648307
transform 1 0 62600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1324
timestamp 1654648307
transform 1 0 64100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1405
timestamp 1654648307
transform 1 0 65600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1406
timestamp 1654648307
transform 1 0 67100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1325
timestamp 1654648307
transform 1 0 65600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1326
timestamp 1654648307
transform 1 0 67100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1407
timestamp 1654648307
transform 1 0 68600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1408
timestamp 1654648307
transform 1 0 70100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1327
timestamp 1654648307
transform 1 0 68600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1328
timestamp 1654648307
transform 1 0 70100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1409
timestamp 1654648307
transform 1 0 71600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1410
timestamp 1654648307
transform 1 0 73100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1329
timestamp 1654648307
transform 1 0 71600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1330
timestamp 1654648307
transform 1 0 73100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1411
timestamp 1654648307
transform 1 0 74600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1412
timestamp 1654648307
transform 1 0 76100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1331
timestamp 1654648307
transform 1 0 74600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1332
timestamp 1654648307
transform 1 0 76100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1413
timestamp 1654648307
transform 1 0 77600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1414
timestamp 1654648307
transform 1 0 79100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1333
timestamp 1654648307
transform 1 0 77600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1334
timestamp 1654648307
transform 1 0 79100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1415
timestamp 1654648307
transform 1 0 80600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1416
timestamp 1654648307
transform 1 0 82100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1335
timestamp 1654648307
transform 1 0 80600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1336
timestamp 1654648307
transform 1 0 82100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1417
timestamp 1654648307
transform 1 0 83600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1418
timestamp 1654648307
transform 1 0 85100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1337
timestamp 1654648307
transform 1 0 83600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1338
timestamp 1654648307
transform 1 0 85100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1419
timestamp 1654648307
transform 1 0 86600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1420
timestamp 1654648307
transform 1 0 88100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1339
timestamp 1654648307
transform 1 0 86600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1340
timestamp 1654648307
transform 1 0 88100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1421
timestamp 1654648307
transform 1 0 89600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1422
timestamp 1654648307
transform 1 0 91100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1341
timestamp 1654648307
transform 1 0 89600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1342
timestamp 1654648307
transform 1 0 91100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1423
timestamp 1654648307
transform 1 0 92600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1424
timestamp 1654648307
transform 1 0 94100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1343
timestamp 1654648307
transform 1 0 92600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1344
timestamp 1654648307
transform 1 0 94100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1425
timestamp 1654648307
transform 1 0 95600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1426
timestamp 1654648307
transform 1 0 97100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1345
timestamp 1654648307
transform 1 0 95600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1346
timestamp 1654648307
transform 1 0 97100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1427
timestamp 1654648307
transform 1 0 98600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1428
timestamp 1654648307
transform 1 0 100100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1347
timestamp 1654648307
transform 1 0 98600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1348
timestamp 1654648307
transform 1 0 100100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1429
timestamp 1654648307
transform 1 0 101600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1430
timestamp 1654648307
transform 1 0 103100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1349
timestamp 1654648307
transform 1 0 101600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1350
timestamp 1654648307
transform 1 0 103100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1431
timestamp 1654648307
transform 1 0 104600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1432
timestamp 1654648307
transform 1 0 106100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1351
timestamp 1654648307
transform 1 0 104600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1352
timestamp 1654648307
transform 1 0 106100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1433
timestamp 1654648307
transform 1 0 107600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1434
timestamp 1654648307
transform 1 0 109100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1353
timestamp 1654648307
transform 1 0 107600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1354
timestamp 1654648307
transform 1 0 109100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1435
timestamp 1654648307
transform 1 0 110600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1436
timestamp 1654648307
transform 1 0 112100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1355
timestamp 1654648307
transform 1 0 110600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1356
timestamp 1654648307
transform 1 0 112100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1437
timestamp 1654648307
transform 1 0 113600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1438
timestamp 1654648307
transform 1 0 115100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1357
timestamp 1654648307
transform 1 0 113600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1358
timestamp 1654648307
transform 1 0 115100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1439
timestamp 1654648307
transform 1 0 116600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1359
timestamp 1654648307
transform 1 0 116600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1200
timestamp 1654648307
transform 1 0 -1900 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1120
timestamp 1654648307
transform 1 0 -1900 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1201
timestamp 1654648307
transform 1 0 -400 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1202
timestamp 1654648307
transform 1 0 1100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1121
timestamp 1654648307
transform 1 0 -400 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1122
timestamp 1654648307
transform 1 0 1100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1203
timestamp 1654648307
transform 1 0 2600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1204
timestamp 1654648307
transform 1 0 4100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1123
timestamp 1654648307
transform 1 0 2600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1124
timestamp 1654648307
transform 1 0 4100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1205
timestamp 1654648307
transform 1 0 5600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1206
timestamp 1654648307
transform 1 0 7100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1125
timestamp 1654648307
transform 1 0 5600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1126
timestamp 1654648307
transform 1 0 7100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1207
timestamp 1654648307
transform 1 0 8600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1208
timestamp 1654648307
transform 1 0 10100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1127
timestamp 1654648307
transform 1 0 8600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1128
timestamp 1654648307
transform 1 0 10100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1209
timestamp 1654648307
transform 1 0 11600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1210
timestamp 1654648307
transform 1 0 13100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1129
timestamp 1654648307
transform 1 0 11600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1130
timestamp 1654648307
transform 1 0 13100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1211
timestamp 1654648307
transform 1 0 14600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1212
timestamp 1654648307
transform 1 0 16100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1131
timestamp 1654648307
transform 1 0 14600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1132
timestamp 1654648307
transform 1 0 16100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1213
timestamp 1654648307
transform 1 0 17600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1214
timestamp 1654648307
transform 1 0 19100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1133
timestamp 1654648307
transform 1 0 17600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1134
timestamp 1654648307
transform 1 0 19100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1215
timestamp 1654648307
transform 1 0 20600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1216
timestamp 1654648307
transform 1 0 22100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1135
timestamp 1654648307
transform 1 0 20600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1136
timestamp 1654648307
transform 1 0 22100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1217
timestamp 1654648307
transform 1 0 23600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1218
timestamp 1654648307
transform 1 0 25100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1137
timestamp 1654648307
transform 1 0 23600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1138
timestamp 1654648307
transform 1 0 25100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1219
timestamp 1654648307
transform 1 0 26600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1220
timestamp 1654648307
transform 1 0 28100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1139
timestamp 1654648307
transform 1 0 26600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1140
timestamp 1654648307
transform 1 0 28100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1221
timestamp 1654648307
transform 1 0 29600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1222
timestamp 1654648307
transform 1 0 31100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1141
timestamp 1654648307
transform 1 0 29600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1142
timestamp 1654648307
transform 1 0 31100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1223
timestamp 1654648307
transform 1 0 32600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1224
timestamp 1654648307
transform 1 0 34100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1143
timestamp 1654648307
transform 1 0 32600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1144
timestamp 1654648307
transform 1 0 34100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1225
timestamp 1654648307
transform 1 0 35600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1226
timestamp 1654648307
transform 1 0 37100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1145
timestamp 1654648307
transform 1 0 35600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1146
timestamp 1654648307
transform 1 0 37100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1227
timestamp 1654648307
transform 1 0 38600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1228
timestamp 1654648307
transform 1 0 40100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1147
timestamp 1654648307
transform 1 0 38600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1148
timestamp 1654648307
transform 1 0 40100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1229
timestamp 1654648307
transform 1 0 41600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1230
timestamp 1654648307
transform 1 0 43100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1149
timestamp 1654648307
transform 1 0 41600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1150
timestamp 1654648307
transform 1 0 43100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1231
timestamp 1654648307
transform 1 0 44600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1232
timestamp 1654648307
transform 1 0 46100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1151
timestamp 1654648307
transform 1 0 44600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1152
timestamp 1654648307
transform 1 0 46100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1233
timestamp 1654648307
transform 1 0 47600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1234
timestamp 1654648307
transform 1 0 49100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1153
timestamp 1654648307
transform 1 0 47600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1154
timestamp 1654648307
transform 1 0 49100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1235
timestamp 1654648307
transform 1 0 50600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1236
timestamp 1654648307
transform 1 0 52100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1155
timestamp 1654648307
transform 1 0 50600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1156
timestamp 1654648307
transform 1 0 52100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1237
timestamp 1654648307
transform 1 0 53600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1238
timestamp 1654648307
transform 1 0 55100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1157
timestamp 1654648307
transform 1 0 53600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1158
timestamp 1654648307
transform 1 0 55100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1239
timestamp 1654648307
transform 1 0 56600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1240
timestamp 1654648307
transform 1 0 58100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1159
timestamp 1654648307
transform 1 0 56600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1160
timestamp 1654648307
transform 1 0 58100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1241
timestamp 1654648307
transform 1 0 59600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1242
timestamp 1654648307
transform 1 0 61100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1161
timestamp 1654648307
transform 1 0 59600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1162
timestamp 1654648307
transform 1 0 61100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1243
timestamp 1654648307
transform 1 0 62600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1244
timestamp 1654648307
transform 1 0 64100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1163
timestamp 1654648307
transform 1 0 62600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1164
timestamp 1654648307
transform 1 0 64100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1245
timestamp 1654648307
transform 1 0 65600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1246
timestamp 1654648307
transform 1 0 67100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1165
timestamp 1654648307
transform 1 0 65600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1166
timestamp 1654648307
transform 1 0 67100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1247
timestamp 1654648307
transform 1 0 68600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1248
timestamp 1654648307
transform 1 0 70100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1167
timestamp 1654648307
transform 1 0 68600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1168
timestamp 1654648307
transform 1 0 70100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1249
timestamp 1654648307
transform 1 0 71600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1250
timestamp 1654648307
transform 1 0 73100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1169
timestamp 1654648307
transform 1 0 71600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1170
timestamp 1654648307
transform 1 0 73100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1251
timestamp 1654648307
transform 1 0 74600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1252
timestamp 1654648307
transform 1 0 76100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1171
timestamp 1654648307
transform 1 0 74600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1172
timestamp 1654648307
transform 1 0 76100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1253
timestamp 1654648307
transform 1 0 77600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1254
timestamp 1654648307
transform 1 0 79100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1173
timestamp 1654648307
transform 1 0 77600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1174
timestamp 1654648307
transform 1 0 79100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1255
timestamp 1654648307
transform 1 0 80600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1256
timestamp 1654648307
transform 1 0 82100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1175
timestamp 1654648307
transform 1 0 80600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1176
timestamp 1654648307
transform 1 0 82100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1257
timestamp 1654648307
transform 1 0 83600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1258
timestamp 1654648307
transform 1 0 85100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1177
timestamp 1654648307
transform 1 0 83600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1178
timestamp 1654648307
transform 1 0 85100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1259
timestamp 1654648307
transform 1 0 86600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1260
timestamp 1654648307
transform 1 0 88100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1179
timestamp 1654648307
transform 1 0 86600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1180
timestamp 1654648307
transform 1 0 88100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1261
timestamp 1654648307
transform 1 0 89600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1262
timestamp 1654648307
transform 1 0 91100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1181
timestamp 1654648307
transform 1 0 89600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1182
timestamp 1654648307
transform 1 0 91100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1263
timestamp 1654648307
transform 1 0 92600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1264
timestamp 1654648307
transform 1 0 94100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1183
timestamp 1654648307
transform 1 0 92600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1184
timestamp 1654648307
transform 1 0 94100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1265
timestamp 1654648307
transform 1 0 95600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1266
timestamp 1654648307
transform 1 0 97100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1185
timestamp 1654648307
transform 1 0 95600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1186
timestamp 1654648307
transform 1 0 97100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1267
timestamp 1654648307
transform 1 0 98600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1268
timestamp 1654648307
transform 1 0 100100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1187
timestamp 1654648307
transform 1 0 98600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1188
timestamp 1654648307
transform 1 0 100100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1269
timestamp 1654648307
transform 1 0 101600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1270
timestamp 1654648307
transform 1 0 103100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1189
timestamp 1654648307
transform 1 0 101600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1190
timestamp 1654648307
transform 1 0 103100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1271
timestamp 1654648307
transform 1 0 104600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1272
timestamp 1654648307
transform 1 0 106100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1191
timestamp 1654648307
transform 1 0 104600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1192
timestamp 1654648307
transform 1 0 106100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1273
timestamp 1654648307
transform 1 0 107600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1274
timestamp 1654648307
transform 1 0 109100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1193
timestamp 1654648307
transform 1 0 107600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1194
timestamp 1654648307
transform 1 0 109100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1275
timestamp 1654648307
transform 1 0 110600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1276
timestamp 1654648307
transform 1 0 112100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1195
timestamp 1654648307
transform 1 0 110600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1196
timestamp 1654648307
transform 1 0 112100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1277
timestamp 1654648307
transform 1 0 113600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1278
timestamp 1654648307
transform 1 0 115100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1197
timestamp 1654648307
transform 1 0 113600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1198
timestamp 1654648307
transform 1 0 115100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1279
timestamp 1654648307
transform 1 0 116600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1199
timestamp 1654648307
transform 1 0 116600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1040
timestamp 1654648307
transform 1 0 -1900 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_960
timestamp 1654648307
transform 1 0 -1900 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1041
timestamp 1654648307
transform 1 0 -400 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1042
timestamp 1654648307
transform 1 0 1100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_961
timestamp 1654648307
transform 1 0 -400 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_962
timestamp 1654648307
transform 1 0 1100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1043
timestamp 1654648307
transform 1 0 2600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1044
timestamp 1654648307
transform 1 0 4100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_963
timestamp 1654648307
transform 1 0 2600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_964
timestamp 1654648307
transform 1 0 4100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1045
timestamp 1654648307
transform 1 0 5600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1046
timestamp 1654648307
transform 1 0 7100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_965
timestamp 1654648307
transform 1 0 5600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_966
timestamp 1654648307
transform 1 0 7100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1047
timestamp 1654648307
transform 1 0 8600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1048
timestamp 1654648307
transform 1 0 10100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_967
timestamp 1654648307
transform 1 0 8600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_968
timestamp 1654648307
transform 1 0 10100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1049
timestamp 1654648307
transform 1 0 11600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1050
timestamp 1654648307
transform 1 0 13100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_969
timestamp 1654648307
transform 1 0 11600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_970
timestamp 1654648307
transform 1 0 13100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1051
timestamp 1654648307
transform 1 0 14600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1052
timestamp 1654648307
transform 1 0 16100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_971
timestamp 1654648307
transform 1 0 14600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_972
timestamp 1654648307
transform 1 0 16100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1053
timestamp 1654648307
transform 1 0 17600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1054
timestamp 1654648307
transform 1 0 19100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_973
timestamp 1654648307
transform 1 0 17600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_974
timestamp 1654648307
transform 1 0 19100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1055
timestamp 1654648307
transform 1 0 20600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1056
timestamp 1654648307
transform 1 0 22100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_975
timestamp 1654648307
transform 1 0 20600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_976
timestamp 1654648307
transform 1 0 22100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1057
timestamp 1654648307
transform 1 0 23600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1058
timestamp 1654648307
transform 1 0 25100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_977
timestamp 1654648307
transform 1 0 23600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_978
timestamp 1654648307
transform 1 0 25100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1059
timestamp 1654648307
transform 1 0 26600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1060
timestamp 1654648307
transform 1 0 28100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_979
timestamp 1654648307
transform 1 0 26600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_980
timestamp 1654648307
transform 1 0 28100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1061
timestamp 1654648307
transform 1 0 29600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1062
timestamp 1654648307
transform 1 0 31100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_981
timestamp 1654648307
transform 1 0 29600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_982
timestamp 1654648307
transform 1 0 31100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1063
timestamp 1654648307
transform 1 0 32600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1064
timestamp 1654648307
transform 1 0 34100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_983
timestamp 1654648307
transform 1 0 32600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_984
timestamp 1654648307
transform 1 0 34100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1065
timestamp 1654648307
transform 1 0 35600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1066
timestamp 1654648307
transform 1 0 37100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_985
timestamp 1654648307
transform 1 0 35600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_986
timestamp 1654648307
transform 1 0 37100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1067
timestamp 1654648307
transform 1 0 38600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1068
timestamp 1654648307
transform 1 0 40100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_987
timestamp 1654648307
transform 1 0 38600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_988
timestamp 1654648307
transform 1 0 40100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1069
timestamp 1654648307
transform 1 0 41600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1070
timestamp 1654648307
transform 1 0 43100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_989
timestamp 1654648307
transform 1 0 41600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_990
timestamp 1654648307
transform 1 0 43100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1071
timestamp 1654648307
transform 1 0 44600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1072
timestamp 1654648307
transform 1 0 46100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_991
timestamp 1654648307
transform 1 0 44600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_992
timestamp 1654648307
transform 1 0 46100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1073
timestamp 1654648307
transform 1 0 47600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1074
timestamp 1654648307
transform 1 0 49100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_993
timestamp 1654648307
transform 1 0 47600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_994
timestamp 1654648307
transform 1 0 49100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1075
timestamp 1654648307
transform 1 0 50600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1076
timestamp 1654648307
transform 1 0 52100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_995
timestamp 1654648307
transform 1 0 50600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_996
timestamp 1654648307
transform 1 0 52100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1077
timestamp 1654648307
transform 1 0 53600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1078
timestamp 1654648307
transform 1 0 55100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_997
timestamp 1654648307
transform 1 0 53600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_998
timestamp 1654648307
transform 1 0 55100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1079
timestamp 1654648307
transform 1 0 56600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1080
timestamp 1654648307
transform 1 0 58100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_999
timestamp 1654648307
transform 1 0 56600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1000
timestamp 1654648307
transform 1 0 58100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1081
timestamp 1654648307
transform 1 0 59600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1082
timestamp 1654648307
transform 1 0 61100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1001
timestamp 1654648307
transform 1 0 59600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1002
timestamp 1654648307
transform 1 0 61100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1083
timestamp 1654648307
transform 1 0 62600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1084
timestamp 1654648307
transform 1 0 64100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1003
timestamp 1654648307
transform 1 0 62600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1004
timestamp 1654648307
transform 1 0 64100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1085
timestamp 1654648307
transform 1 0 65600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1086
timestamp 1654648307
transform 1 0 67100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1005
timestamp 1654648307
transform 1 0 65600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1006
timestamp 1654648307
transform 1 0 67100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1087
timestamp 1654648307
transform 1 0 68600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1088
timestamp 1654648307
transform 1 0 70100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1007
timestamp 1654648307
transform 1 0 68600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1008
timestamp 1654648307
transform 1 0 70100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1089
timestamp 1654648307
transform 1 0 71600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1090
timestamp 1654648307
transform 1 0 73100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1009
timestamp 1654648307
transform 1 0 71600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1010
timestamp 1654648307
transform 1 0 73100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1091
timestamp 1654648307
transform 1 0 74600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1092
timestamp 1654648307
transform 1 0 76100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1011
timestamp 1654648307
transform 1 0 74600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1012
timestamp 1654648307
transform 1 0 76100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1093
timestamp 1654648307
transform 1 0 77600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1094
timestamp 1654648307
transform 1 0 79100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1013
timestamp 1654648307
transform 1 0 77600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1014
timestamp 1654648307
transform 1 0 79100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1095
timestamp 1654648307
transform 1 0 80600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1096
timestamp 1654648307
transform 1 0 82100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1015
timestamp 1654648307
transform 1 0 80600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1016
timestamp 1654648307
transform 1 0 82100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1097
timestamp 1654648307
transform 1 0 83600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1098
timestamp 1654648307
transform 1 0 85100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1017
timestamp 1654648307
transform 1 0 83600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1018
timestamp 1654648307
transform 1 0 85100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1099
timestamp 1654648307
transform 1 0 86600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1100
timestamp 1654648307
transform 1 0 88100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1019
timestamp 1654648307
transform 1 0 86600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1020
timestamp 1654648307
transform 1 0 88100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1101
timestamp 1654648307
transform 1 0 89600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1102
timestamp 1654648307
transform 1 0 91100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1021
timestamp 1654648307
transform 1 0 89600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1022
timestamp 1654648307
transform 1 0 91100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1103
timestamp 1654648307
transform 1 0 92600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1104
timestamp 1654648307
transform 1 0 94100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1023
timestamp 1654648307
transform 1 0 92600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1024
timestamp 1654648307
transform 1 0 94100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1105
timestamp 1654648307
transform 1 0 95600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1106
timestamp 1654648307
transform 1 0 97100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1025
timestamp 1654648307
transform 1 0 95600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1026
timestamp 1654648307
transform 1 0 97100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1107
timestamp 1654648307
transform 1 0 98600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1108
timestamp 1654648307
transform 1 0 100100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1027
timestamp 1654648307
transform 1 0 98600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1028
timestamp 1654648307
transform 1 0 100100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1109
timestamp 1654648307
transform 1 0 101600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1110
timestamp 1654648307
transform 1 0 103100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1029
timestamp 1654648307
transform 1 0 101600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1030
timestamp 1654648307
transform 1 0 103100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1111
timestamp 1654648307
transform 1 0 104600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1112
timestamp 1654648307
transform 1 0 106100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1031
timestamp 1654648307
transform 1 0 104600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1032
timestamp 1654648307
transform 1 0 106100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1113
timestamp 1654648307
transform 1 0 107600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1114
timestamp 1654648307
transform 1 0 109100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1033
timestamp 1654648307
transform 1 0 107600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1034
timestamp 1654648307
transform 1 0 109100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1115
timestamp 1654648307
transform 1 0 110600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1116
timestamp 1654648307
transform 1 0 112100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1035
timestamp 1654648307
transform 1 0 110600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1036
timestamp 1654648307
transform 1 0 112100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1117
timestamp 1654648307
transform 1 0 113600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1118
timestamp 1654648307
transform 1 0 115100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1037
timestamp 1654648307
transform 1 0 113600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1038
timestamp 1654648307
transform 1 0 115100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1119
timestamp 1654648307
transform 1 0 116600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1039
timestamp 1654648307
transform 1 0 116600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_880
timestamp 1654648307
transform 1 0 -1900 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_800
timestamp 1654648307
transform 1 0 -1900 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_881
timestamp 1654648307
transform 1 0 -400 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_882
timestamp 1654648307
transform 1 0 1100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_801
timestamp 1654648307
transform 1 0 -400 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_802
timestamp 1654648307
transform 1 0 1100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_883
timestamp 1654648307
transform 1 0 2600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_884
timestamp 1654648307
transform 1 0 4100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_803
timestamp 1654648307
transform 1 0 2600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_804
timestamp 1654648307
transform 1 0 4100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_885
timestamp 1654648307
transform 1 0 5600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_886
timestamp 1654648307
transform 1 0 7100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_805
timestamp 1654648307
transform 1 0 5600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_806
timestamp 1654648307
transform 1 0 7100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_887
timestamp 1654648307
transform 1 0 8600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_888
timestamp 1654648307
transform 1 0 10100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_807
timestamp 1654648307
transform 1 0 8600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_808
timestamp 1654648307
transform 1 0 10100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_889
timestamp 1654648307
transform 1 0 11600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_890
timestamp 1654648307
transform 1 0 13100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_809
timestamp 1654648307
transform 1 0 11600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_810
timestamp 1654648307
transform 1 0 13100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_891
timestamp 1654648307
transform 1 0 14600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_892
timestamp 1654648307
transform 1 0 16100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_811
timestamp 1654648307
transform 1 0 14600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_812
timestamp 1654648307
transform 1 0 16100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_893
timestamp 1654648307
transform 1 0 17600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_894
timestamp 1654648307
transform 1 0 19100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_813
timestamp 1654648307
transform 1 0 17600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_814
timestamp 1654648307
transform 1 0 19100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_895
timestamp 1654648307
transform 1 0 20600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_896
timestamp 1654648307
transform 1 0 22100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_815
timestamp 1654648307
transform 1 0 20600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_816
timestamp 1654648307
transform 1 0 22100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_897
timestamp 1654648307
transform 1 0 23600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_898
timestamp 1654648307
transform 1 0 25100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_817
timestamp 1654648307
transform 1 0 23600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_818
timestamp 1654648307
transform 1 0 25100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_899
timestamp 1654648307
transform 1 0 26600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_900
timestamp 1654648307
transform 1 0 28100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_819
timestamp 1654648307
transform 1 0 26600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_820
timestamp 1654648307
transform 1 0 28100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_901
timestamp 1654648307
transform 1 0 29600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_902
timestamp 1654648307
transform 1 0 31100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_821
timestamp 1654648307
transform 1 0 29600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_822
timestamp 1654648307
transform 1 0 31100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_903
timestamp 1654648307
transform 1 0 32600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_904
timestamp 1654648307
transform 1 0 34100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_823
timestamp 1654648307
transform 1 0 32600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_824
timestamp 1654648307
transform 1 0 34100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_905
timestamp 1654648307
transform 1 0 35600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_906
timestamp 1654648307
transform 1 0 37100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_825
timestamp 1654648307
transform 1 0 35600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_826
timestamp 1654648307
transform 1 0 37100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_907
timestamp 1654648307
transform 1 0 38600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_908
timestamp 1654648307
transform 1 0 40100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_827
timestamp 1654648307
transform 1 0 38600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_828
timestamp 1654648307
transform 1 0 40100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_909
timestamp 1654648307
transform 1 0 41600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_910
timestamp 1654648307
transform 1 0 43100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_829
timestamp 1654648307
transform 1 0 41600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_830
timestamp 1654648307
transform 1 0 43100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_911
timestamp 1654648307
transform 1 0 44600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_912
timestamp 1654648307
transform 1 0 46100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_831
timestamp 1654648307
transform 1 0 44600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_832
timestamp 1654648307
transform 1 0 46100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_913
timestamp 1654648307
transform 1 0 47600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_914
timestamp 1654648307
transform 1 0 49100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_833
timestamp 1654648307
transform 1 0 47600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_834
timestamp 1654648307
transform 1 0 49100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_915
timestamp 1654648307
transform 1 0 50600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_916
timestamp 1654648307
transform 1 0 52100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_835
timestamp 1654648307
transform 1 0 50600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_836
timestamp 1654648307
transform 1 0 52100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_917
timestamp 1654648307
transform 1 0 53600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_918
timestamp 1654648307
transform 1 0 55100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_837
timestamp 1654648307
transform 1 0 53600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_838
timestamp 1654648307
transform 1 0 55100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_919
timestamp 1654648307
transform 1 0 56600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_920
timestamp 1654648307
transform 1 0 58100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_839
timestamp 1654648307
transform 1 0 56600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_840
timestamp 1654648307
transform 1 0 58100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_921
timestamp 1654648307
transform 1 0 59600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_922
timestamp 1654648307
transform 1 0 61100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_841
timestamp 1654648307
transform 1 0 59600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_842
timestamp 1654648307
transform 1 0 61100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_923
timestamp 1654648307
transform 1 0 62600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_924
timestamp 1654648307
transform 1 0 64100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_843
timestamp 1654648307
transform 1 0 62600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_844
timestamp 1654648307
transform 1 0 64100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_925
timestamp 1654648307
transform 1 0 65600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_926
timestamp 1654648307
transform 1 0 67100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_845
timestamp 1654648307
transform 1 0 65600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_846
timestamp 1654648307
transform 1 0 67100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_927
timestamp 1654648307
transform 1 0 68600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_928
timestamp 1654648307
transform 1 0 70100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_847
timestamp 1654648307
transform 1 0 68600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_848
timestamp 1654648307
transform 1 0 70100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_929
timestamp 1654648307
transform 1 0 71600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_930
timestamp 1654648307
transform 1 0 73100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_849
timestamp 1654648307
transform 1 0 71600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_850
timestamp 1654648307
transform 1 0 73100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_931
timestamp 1654648307
transform 1 0 74600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_932
timestamp 1654648307
transform 1 0 76100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_851
timestamp 1654648307
transform 1 0 74600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_852
timestamp 1654648307
transform 1 0 76100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_933
timestamp 1654648307
transform 1 0 77600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_934
timestamp 1654648307
transform 1 0 79100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_853
timestamp 1654648307
transform 1 0 77600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_854
timestamp 1654648307
transform 1 0 79100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_935
timestamp 1654648307
transform 1 0 80600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_936
timestamp 1654648307
transform 1 0 82100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_855
timestamp 1654648307
transform 1 0 80600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_856
timestamp 1654648307
transform 1 0 82100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_937
timestamp 1654648307
transform 1 0 83600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_938
timestamp 1654648307
transform 1 0 85100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_857
timestamp 1654648307
transform 1 0 83600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_858
timestamp 1654648307
transform 1 0 85100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_939
timestamp 1654648307
transform 1 0 86600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_940
timestamp 1654648307
transform 1 0 88100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_859
timestamp 1654648307
transform 1 0 86600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_860
timestamp 1654648307
transform 1 0 88100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_941
timestamp 1654648307
transform 1 0 89600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_942
timestamp 1654648307
transform 1 0 91100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_861
timestamp 1654648307
transform 1 0 89600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_862
timestamp 1654648307
transform 1 0 91100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_943
timestamp 1654648307
transform 1 0 92600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_944
timestamp 1654648307
transform 1 0 94100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_863
timestamp 1654648307
transform 1 0 92600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_864
timestamp 1654648307
transform 1 0 94100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_945
timestamp 1654648307
transform 1 0 95600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_946
timestamp 1654648307
transform 1 0 97100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_865
timestamp 1654648307
transform 1 0 95600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_866
timestamp 1654648307
transform 1 0 97100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_947
timestamp 1654648307
transform 1 0 98600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_948
timestamp 1654648307
transform 1 0 100100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_867
timestamp 1654648307
transform 1 0 98600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_868
timestamp 1654648307
transform 1 0 100100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_949
timestamp 1654648307
transform 1 0 101600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_950
timestamp 1654648307
transform 1 0 103100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_869
timestamp 1654648307
transform 1 0 101600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_870
timestamp 1654648307
transform 1 0 103100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_951
timestamp 1654648307
transform 1 0 104600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_952
timestamp 1654648307
transform 1 0 106100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_871
timestamp 1654648307
transform 1 0 104600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_872
timestamp 1654648307
transform 1 0 106100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_953
timestamp 1654648307
transform 1 0 107600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_954
timestamp 1654648307
transform 1 0 109100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_873
timestamp 1654648307
transform 1 0 107600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_874
timestamp 1654648307
transform 1 0 109100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_955
timestamp 1654648307
transform 1 0 110600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_956
timestamp 1654648307
transform 1 0 112100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_875
timestamp 1654648307
transform 1 0 110600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_876
timestamp 1654648307
transform 1 0 112100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_957
timestamp 1654648307
transform 1 0 113600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_958
timestamp 1654648307
transform 1 0 115100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_877
timestamp 1654648307
transform 1 0 113600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_878
timestamp 1654648307
transform 1 0 115100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_959
timestamp 1654648307
transform 1 0 116600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_879
timestamp 1654648307
transform 1 0 116600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_720
timestamp 1654648307
transform 1 0 -1900 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_640
timestamp 1654648307
transform 1 0 -1900 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_721
timestamp 1654648307
transform 1 0 -400 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_722
timestamp 1654648307
transform 1 0 1100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_641
timestamp 1654648307
transform 1 0 -400 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_642
timestamp 1654648307
transform 1 0 1100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_723
timestamp 1654648307
transform 1 0 2600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_724
timestamp 1654648307
transform 1 0 4100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_643
timestamp 1654648307
transform 1 0 2600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_644
timestamp 1654648307
transform 1 0 4100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_725
timestamp 1654648307
transform 1 0 5600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_726
timestamp 1654648307
transform 1 0 7100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_645
timestamp 1654648307
transform 1 0 5600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_646
timestamp 1654648307
transform 1 0 7100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_727
timestamp 1654648307
transform 1 0 8600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_728
timestamp 1654648307
transform 1 0 10100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_647
timestamp 1654648307
transform 1 0 8600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_648
timestamp 1654648307
transform 1 0 10100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_729
timestamp 1654648307
transform 1 0 11600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_730
timestamp 1654648307
transform 1 0 13100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_649
timestamp 1654648307
transform 1 0 11600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_650
timestamp 1654648307
transform 1 0 13100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_731
timestamp 1654648307
transform 1 0 14600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_732
timestamp 1654648307
transform 1 0 16100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_651
timestamp 1654648307
transform 1 0 14600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_652
timestamp 1654648307
transform 1 0 16100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_733
timestamp 1654648307
transform 1 0 17600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_734
timestamp 1654648307
transform 1 0 19100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_653
timestamp 1654648307
transform 1 0 17600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_654
timestamp 1654648307
transform 1 0 19100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_735
timestamp 1654648307
transform 1 0 20600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_736
timestamp 1654648307
transform 1 0 22100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_655
timestamp 1654648307
transform 1 0 20600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_656
timestamp 1654648307
transform 1 0 22100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_737
timestamp 1654648307
transform 1 0 23600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_738
timestamp 1654648307
transform 1 0 25100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_657
timestamp 1654648307
transform 1 0 23600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_658
timestamp 1654648307
transform 1 0 25100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_739
timestamp 1654648307
transform 1 0 26600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_740
timestamp 1654648307
transform 1 0 28100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_659
timestamp 1654648307
transform 1 0 26600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_660
timestamp 1654648307
transform 1 0 28100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_741
timestamp 1654648307
transform 1 0 29600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_742
timestamp 1654648307
transform 1 0 31100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_661
timestamp 1654648307
transform 1 0 29600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_662
timestamp 1654648307
transform 1 0 31100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_743
timestamp 1654648307
transform 1 0 32600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_744
timestamp 1654648307
transform 1 0 34100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_663
timestamp 1654648307
transform 1 0 32600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_664
timestamp 1654648307
transform 1 0 34100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_745
timestamp 1654648307
transform 1 0 35600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_746
timestamp 1654648307
transform 1 0 37100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_665
timestamp 1654648307
transform 1 0 35600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_666
timestamp 1654648307
transform 1 0 37100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_747
timestamp 1654648307
transform 1 0 38600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_748
timestamp 1654648307
transform 1 0 40100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_667
timestamp 1654648307
transform 1 0 38600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_668
timestamp 1654648307
transform 1 0 40100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_749
timestamp 1654648307
transform 1 0 41600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_750
timestamp 1654648307
transform 1 0 43100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_669
timestamp 1654648307
transform 1 0 41600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_670
timestamp 1654648307
transform 1 0 43100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_751
timestamp 1654648307
transform 1 0 44600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_752
timestamp 1654648307
transform 1 0 46100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_671
timestamp 1654648307
transform 1 0 44600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_672
timestamp 1654648307
transform 1 0 46100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_753
timestamp 1654648307
transform 1 0 47600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_754
timestamp 1654648307
transform 1 0 49100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_673
timestamp 1654648307
transform 1 0 47600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_674
timestamp 1654648307
transform 1 0 49100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_755
timestamp 1654648307
transform 1 0 50600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_756
timestamp 1654648307
transform 1 0 52100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_675
timestamp 1654648307
transform 1 0 50600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_676
timestamp 1654648307
transform 1 0 52100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_757
timestamp 1654648307
transform 1 0 53600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_758
timestamp 1654648307
transform 1 0 55100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_677
timestamp 1654648307
transform 1 0 53600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_678
timestamp 1654648307
transform 1 0 55100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_759
timestamp 1654648307
transform 1 0 56600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_760
timestamp 1654648307
transform 1 0 58100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_679
timestamp 1654648307
transform 1 0 56600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_680
timestamp 1654648307
transform 1 0 58100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_761
timestamp 1654648307
transform 1 0 59600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_762
timestamp 1654648307
transform 1 0 61100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_681
timestamp 1654648307
transform 1 0 59600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_682
timestamp 1654648307
transform 1 0 61100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_763
timestamp 1654648307
transform 1 0 62600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_764
timestamp 1654648307
transform 1 0 64100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_683
timestamp 1654648307
transform 1 0 62600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_684
timestamp 1654648307
transform 1 0 64100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_765
timestamp 1654648307
transform 1 0 65600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_766
timestamp 1654648307
transform 1 0 67100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_685
timestamp 1654648307
transform 1 0 65600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_686
timestamp 1654648307
transform 1 0 67100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_767
timestamp 1654648307
transform 1 0 68600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_768
timestamp 1654648307
transform 1 0 70100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_687
timestamp 1654648307
transform 1 0 68600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_688
timestamp 1654648307
transform 1 0 70100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_769
timestamp 1654648307
transform 1 0 71600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_770
timestamp 1654648307
transform 1 0 73100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_689
timestamp 1654648307
transform 1 0 71600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_690
timestamp 1654648307
transform 1 0 73100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_771
timestamp 1654648307
transform 1 0 74600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_772
timestamp 1654648307
transform 1 0 76100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_691
timestamp 1654648307
transform 1 0 74600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_692
timestamp 1654648307
transform 1 0 76100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_773
timestamp 1654648307
transform 1 0 77600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_774
timestamp 1654648307
transform 1 0 79100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_693
timestamp 1654648307
transform 1 0 77600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_694
timestamp 1654648307
transform 1 0 79100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_775
timestamp 1654648307
transform 1 0 80600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_776
timestamp 1654648307
transform 1 0 82100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_695
timestamp 1654648307
transform 1 0 80600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_696
timestamp 1654648307
transform 1 0 82100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_777
timestamp 1654648307
transform 1 0 83600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_778
timestamp 1654648307
transform 1 0 85100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_697
timestamp 1654648307
transform 1 0 83600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_698
timestamp 1654648307
transform 1 0 85100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_779
timestamp 1654648307
transform 1 0 86600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_780
timestamp 1654648307
transform 1 0 88100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_699
timestamp 1654648307
transform 1 0 86600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_700
timestamp 1654648307
transform 1 0 88100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_781
timestamp 1654648307
transform 1 0 89600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_782
timestamp 1654648307
transform 1 0 91100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_701
timestamp 1654648307
transform 1 0 89600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_702
timestamp 1654648307
transform 1 0 91100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_783
timestamp 1654648307
transform 1 0 92600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_784
timestamp 1654648307
transform 1 0 94100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_703
timestamp 1654648307
transform 1 0 92600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_704
timestamp 1654648307
transform 1 0 94100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_785
timestamp 1654648307
transform 1 0 95600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_786
timestamp 1654648307
transform 1 0 97100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_705
timestamp 1654648307
transform 1 0 95600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_706
timestamp 1654648307
transform 1 0 97100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_787
timestamp 1654648307
transform 1 0 98600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_788
timestamp 1654648307
transform 1 0 100100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_707
timestamp 1654648307
transform 1 0 98600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_708
timestamp 1654648307
transform 1 0 100100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_789
timestamp 1654648307
transform 1 0 101600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_790
timestamp 1654648307
transform 1 0 103100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_709
timestamp 1654648307
transform 1 0 101600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_710
timestamp 1654648307
transform 1 0 103100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_791
timestamp 1654648307
transform 1 0 104600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_792
timestamp 1654648307
transform 1 0 106100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_711
timestamp 1654648307
transform 1 0 104600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_712
timestamp 1654648307
transform 1 0 106100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_793
timestamp 1654648307
transform 1 0 107600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_794
timestamp 1654648307
transform 1 0 109100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_713
timestamp 1654648307
transform 1 0 107600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_714
timestamp 1654648307
transform 1 0 109100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_795
timestamp 1654648307
transform 1 0 110600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_796
timestamp 1654648307
transform 1 0 112100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_715
timestamp 1654648307
transform 1 0 110600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_716
timestamp 1654648307
transform 1 0 112100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_797
timestamp 1654648307
transform 1 0 113600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_798
timestamp 1654648307
transform 1 0 115100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_717
timestamp 1654648307
transform 1 0 113600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_718
timestamp 1654648307
transform 1 0 115100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_799
timestamp 1654648307
transform 1 0 116600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_719
timestamp 1654648307
transform 1 0 116600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_560
timestamp 1654648307
transform 1 0 -1900 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_480
timestamp 1654648307
transform 1 0 -1900 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_561
timestamp 1654648307
transform 1 0 -400 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_562
timestamp 1654648307
transform 1 0 1100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_481
timestamp 1654648307
transform 1 0 -400 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_482
timestamp 1654648307
transform 1 0 1100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_563
timestamp 1654648307
transform 1 0 2600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_564
timestamp 1654648307
transform 1 0 4100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_483
timestamp 1654648307
transform 1 0 2600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_484
timestamp 1654648307
transform 1 0 4100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_565
timestamp 1654648307
transform 1 0 5600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_566
timestamp 1654648307
transform 1 0 7100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_485
timestamp 1654648307
transform 1 0 5600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_486
timestamp 1654648307
transform 1 0 7100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_567
timestamp 1654648307
transform 1 0 8600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_568
timestamp 1654648307
transform 1 0 10100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_487
timestamp 1654648307
transform 1 0 8600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_488
timestamp 1654648307
transform 1 0 10100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_569
timestamp 1654648307
transform 1 0 11600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_570
timestamp 1654648307
transform 1 0 13100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_489
timestamp 1654648307
transform 1 0 11600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_490
timestamp 1654648307
transform 1 0 13100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_571
timestamp 1654648307
transform 1 0 14600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_572
timestamp 1654648307
transform 1 0 16100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_491
timestamp 1654648307
transform 1 0 14600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_492
timestamp 1654648307
transform 1 0 16100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_573
timestamp 1654648307
transform 1 0 17600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_574
timestamp 1654648307
transform 1 0 19100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_493
timestamp 1654648307
transform 1 0 17600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_494
timestamp 1654648307
transform 1 0 19100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_575
timestamp 1654648307
transform 1 0 20600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_576
timestamp 1654648307
transform 1 0 22100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_495
timestamp 1654648307
transform 1 0 20600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_496
timestamp 1654648307
transform 1 0 22100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_577
timestamp 1654648307
transform 1 0 23600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_578
timestamp 1654648307
transform 1 0 25100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_497
timestamp 1654648307
transform 1 0 23600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_498
timestamp 1654648307
transform 1 0 25100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_579
timestamp 1654648307
transform 1 0 26600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_580
timestamp 1654648307
transform 1 0 28100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_499
timestamp 1654648307
transform 1 0 26600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_500
timestamp 1654648307
transform 1 0 28100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_581
timestamp 1654648307
transform 1 0 29600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_582
timestamp 1654648307
transform 1 0 31100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_501
timestamp 1654648307
transform 1 0 29600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_502
timestamp 1654648307
transform 1 0 31100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_583
timestamp 1654648307
transform 1 0 32600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_584
timestamp 1654648307
transform 1 0 34100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_503
timestamp 1654648307
transform 1 0 32600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_504
timestamp 1654648307
transform 1 0 34100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_585
timestamp 1654648307
transform 1 0 35600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_586
timestamp 1654648307
transform 1 0 37100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_505
timestamp 1654648307
transform 1 0 35600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_506
timestamp 1654648307
transform 1 0 37100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_587
timestamp 1654648307
transform 1 0 38600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_588
timestamp 1654648307
transform 1 0 40100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_507
timestamp 1654648307
transform 1 0 38600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_508
timestamp 1654648307
transform 1 0 40100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_589
timestamp 1654648307
transform 1 0 41600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_590
timestamp 1654648307
transform 1 0 43100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_509
timestamp 1654648307
transform 1 0 41600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_510
timestamp 1654648307
transform 1 0 43100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_591
timestamp 1654648307
transform 1 0 44600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_592
timestamp 1654648307
transform 1 0 46100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_511
timestamp 1654648307
transform 1 0 44600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_512
timestamp 1654648307
transform 1 0 46100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_593
timestamp 1654648307
transform 1 0 47600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_594
timestamp 1654648307
transform 1 0 49100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_513
timestamp 1654648307
transform 1 0 47600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_514
timestamp 1654648307
transform 1 0 49100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_595
timestamp 1654648307
transform 1 0 50600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_596
timestamp 1654648307
transform 1 0 52100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_515
timestamp 1654648307
transform 1 0 50600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_516
timestamp 1654648307
transform 1 0 52100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_597
timestamp 1654648307
transform 1 0 53600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_598
timestamp 1654648307
transform 1 0 55100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_517
timestamp 1654648307
transform 1 0 53600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_518
timestamp 1654648307
transform 1 0 55100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_599
timestamp 1654648307
transform 1 0 56600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_600
timestamp 1654648307
transform 1 0 58100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_519
timestamp 1654648307
transform 1 0 56600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_520
timestamp 1654648307
transform 1 0 58100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_601
timestamp 1654648307
transform 1 0 59600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_602
timestamp 1654648307
transform 1 0 61100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_521
timestamp 1654648307
transform 1 0 59600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_522
timestamp 1654648307
transform 1 0 61100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_603
timestamp 1654648307
transform 1 0 62600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_604
timestamp 1654648307
transform 1 0 64100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_523
timestamp 1654648307
transform 1 0 62600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_524
timestamp 1654648307
transform 1 0 64100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_605
timestamp 1654648307
transform 1 0 65600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_606
timestamp 1654648307
transform 1 0 67100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_525
timestamp 1654648307
transform 1 0 65600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_526
timestamp 1654648307
transform 1 0 67100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_607
timestamp 1654648307
transform 1 0 68600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_608
timestamp 1654648307
transform 1 0 70100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_527
timestamp 1654648307
transform 1 0 68600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_528
timestamp 1654648307
transform 1 0 70100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_609
timestamp 1654648307
transform 1 0 71600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_610
timestamp 1654648307
transform 1 0 73100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_529
timestamp 1654648307
transform 1 0 71600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_530
timestamp 1654648307
transform 1 0 73100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_611
timestamp 1654648307
transform 1 0 74600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_612
timestamp 1654648307
transform 1 0 76100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_531
timestamp 1654648307
transform 1 0 74600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_532
timestamp 1654648307
transform 1 0 76100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_613
timestamp 1654648307
transform 1 0 77600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_614
timestamp 1654648307
transform 1 0 79100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_533
timestamp 1654648307
transform 1 0 77600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_534
timestamp 1654648307
transform 1 0 79100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_615
timestamp 1654648307
transform 1 0 80600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_616
timestamp 1654648307
transform 1 0 82100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_535
timestamp 1654648307
transform 1 0 80600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_536
timestamp 1654648307
transform 1 0 82100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_617
timestamp 1654648307
transform 1 0 83600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_618
timestamp 1654648307
transform 1 0 85100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_537
timestamp 1654648307
transform 1 0 83600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_538
timestamp 1654648307
transform 1 0 85100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_619
timestamp 1654648307
transform 1 0 86600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_620
timestamp 1654648307
transform 1 0 88100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_539
timestamp 1654648307
transform 1 0 86600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_540
timestamp 1654648307
transform 1 0 88100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_621
timestamp 1654648307
transform 1 0 89600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_622
timestamp 1654648307
transform 1 0 91100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_541
timestamp 1654648307
transform 1 0 89600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_542
timestamp 1654648307
transform 1 0 91100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_623
timestamp 1654648307
transform 1 0 92600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_624
timestamp 1654648307
transform 1 0 94100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_543
timestamp 1654648307
transform 1 0 92600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_544
timestamp 1654648307
transform 1 0 94100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_625
timestamp 1654648307
transform 1 0 95600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_626
timestamp 1654648307
transform 1 0 97100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_545
timestamp 1654648307
transform 1 0 95600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_546
timestamp 1654648307
transform 1 0 97100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_627
timestamp 1654648307
transform 1 0 98600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_628
timestamp 1654648307
transform 1 0 100100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_547
timestamp 1654648307
transform 1 0 98600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_548
timestamp 1654648307
transform 1 0 100100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_629
timestamp 1654648307
transform 1 0 101600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_630
timestamp 1654648307
transform 1 0 103100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_549
timestamp 1654648307
transform 1 0 101600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_550
timestamp 1654648307
transform 1 0 103100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_631
timestamp 1654648307
transform 1 0 104600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_632
timestamp 1654648307
transform 1 0 106100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_551
timestamp 1654648307
transform 1 0 104600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_552
timestamp 1654648307
transform 1 0 106100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_633
timestamp 1654648307
transform 1 0 107600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_634
timestamp 1654648307
transform 1 0 109100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_553
timestamp 1654648307
transform 1 0 107600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_554
timestamp 1654648307
transform 1 0 109100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_635
timestamp 1654648307
transform 1 0 110600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_636
timestamp 1654648307
transform 1 0 112100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_555
timestamp 1654648307
transform 1 0 110600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_556
timestamp 1654648307
transform 1 0 112100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_637
timestamp 1654648307
transform 1 0 113600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_638
timestamp 1654648307
transform 1 0 115100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_557
timestamp 1654648307
transform 1 0 113600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_558
timestamp 1654648307
transform 1 0 115100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_639
timestamp 1654648307
transform 1 0 116600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_559
timestamp 1654648307
transform 1 0 116600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_400
timestamp 1654648307
transform 1 0 -1900 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_320
timestamp 1654648307
transform 1 0 -1900 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_401
timestamp 1654648307
transform 1 0 -400 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_402
timestamp 1654648307
transform 1 0 1100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_321
timestamp 1654648307
transform 1 0 -400 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_322
timestamp 1654648307
transform 1 0 1100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_403
timestamp 1654648307
transform 1 0 2600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_404
timestamp 1654648307
transform 1 0 4100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_323
timestamp 1654648307
transform 1 0 2600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_324
timestamp 1654648307
transform 1 0 4100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_405
timestamp 1654648307
transform 1 0 5600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_406
timestamp 1654648307
transform 1 0 7100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_325
timestamp 1654648307
transform 1 0 5600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_326
timestamp 1654648307
transform 1 0 7100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_407
timestamp 1654648307
transform 1 0 8600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_408
timestamp 1654648307
transform 1 0 10100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_327
timestamp 1654648307
transform 1 0 8600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_328
timestamp 1654648307
transform 1 0 10100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_409
timestamp 1654648307
transform 1 0 11600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_410
timestamp 1654648307
transform 1 0 13100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_329
timestamp 1654648307
transform 1 0 11600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_330
timestamp 1654648307
transform 1 0 13100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_411
timestamp 1654648307
transform 1 0 14600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_412
timestamp 1654648307
transform 1 0 16100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_331
timestamp 1654648307
transform 1 0 14600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_332
timestamp 1654648307
transform 1 0 16100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_413
timestamp 1654648307
transform 1 0 17600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_414
timestamp 1654648307
transform 1 0 19100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_333
timestamp 1654648307
transform 1 0 17600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_334
timestamp 1654648307
transform 1 0 19100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_415
timestamp 1654648307
transform 1 0 20600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_416
timestamp 1654648307
transform 1 0 22100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_335
timestamp 1654648307
transform 1 0 20600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_336
timestamp 1654648307
transform 1 0 22100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_417
timestamp 1654648307
transform 1 0 23600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_418
timestamp 1654648307
transform 1 0 25100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_337
timestamp 1654648307
transform 1 0 23600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_338
timestamp 1654648307
transform 1 0 25100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_419
timestamp 1654648307
transform 1 0 26600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_420
timestamp 1654648307
transform 1 0 28100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_339
timestamp 1654648307
transform 1 0 26600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_340
timestamp 1654648307
transform 1 0 28100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_421
timestamp 1654648307
transform 1 0 29600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_422
timestamp 1654648307
transform 1 0 31100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_341
timestamp 1654648307
transform 1 0 29600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_342
timestamp 1654648307
transform 1 0 31100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_423
timestamp 1654648307
transform 1 0 32600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_424
timestamp 1654648307
transform 1 0 34100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_343
timestamp 1654648307
transform 1 0 32600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_344
timestamp 1654648307
transform 1 0 34100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_425
timestamp 1654648307
transform 1 0 35600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_426
timestamp 1654648307
transform 1 0 37100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_345
timestamp 1654648307
transform 1 0 35600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_346
timestamp 1654648307
transform 1 0 37100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_427
timestamp 1654648307
transform 1 0 38600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_428
timestamp 1654648307
transform 1 0 40100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_347
timestamp 1654648307
transform 1 0 38600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_348
timestamp 1654648307
transform 1 0 40100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_429
timestamp 1654648307
transform 1 0 41600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_430
timestamp 1654648307
transform 1 0 43100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_349
timestamp 1654648307
transform 1 0 41600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_350
timestamp 1654648307
transform 1 0 43100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_431
timestamp 1654648307
transform 1 0 44600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_432
timestamp 1654648307
transform 1 0 46100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_351
timestamp 1654648307
transform 1 0 44600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_352
timestamp 1654648307
transform 1 0 46100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_433
timestamp 1654648307
transform 1 0 47600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_434
timestamp 1654648307
transform 1 0 49100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_353
timestamp 1654648307
transform 1 0 47600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_354
timestamp 1654648307
transform 1 0 49100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_435
timestamp 1654648307
transform 1 0 50600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_436
timestamp 1654648307
transform 1 0 52100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_355
timestamp 1654648307
transform 1 0 50600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_356
timestamp 1654648307
transform 1 0 52100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_437
timestamp 1654648307
transform 1 0 53600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_438
timestamp 1654648307
transform 1 0 55100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_357
timestamp 1654648307
transform 1 0 53600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_358
timestamp 1654648307
transform 1 0 55100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_439
timestamp 1654648307
transform 1 0 56600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_440
timestamp 1654648307
transform 1 0 58100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_359
timestamp 1654648307
transform 1 0 56600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_360
timestamp 1654648307
transform 1 0 58100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_441
timestamp 1654648307
transform 1 0 59600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_442
timestamp 1654648307
transform 1 0 61100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_361
timestamp 1654648307
transform 1 0 59600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_362
timestamp 1654648307
transform 1 0 61100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_443
timestamp 1654648307
transform 1 0 62600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_444
timestamp 1654648307
transform 1 0 64100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_363
timestamp 1654648307
transform 1 0 62600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_364
timestamp 1654648307
transform 1 0 64100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_445
timestamp 1654648307
transform 1 0 65600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_446
timestamp 1654648307
transform 1 0 67100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_365
timestamp 1654648307
transform 1 0 65600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_366
timestamp 1654648307
transform 1 0 67100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_447
timestamp 1654648307
transform 1 0 68600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_448
timestamp 1654648307
transform 1 0 70100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_367
timestamp 1654648307
transform 1 0 68600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_368
timestamp 1654648307
transform 1 0 70100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_449
timestamp 1654648307
transform 1 0 71600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_450
timestamp 1654648307
transform 1 0 73100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_369
timestamp 1654648307
transform 1 0 71600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_370
timestamp 1654648307
transform 1 0 73100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_451
timestamp 1654648307
transform 1 0 74600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_452
timestamp 1654648307
transform 1 0 76100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_371
timestamp 1654648307
transform 1 0 74600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_372
timestamp 1654648307
transform 1 0 76100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_453
timestamp 1654648307
transform 1 0 77600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_454
timestamp 1654648307
transform 1 0 79100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_373
timestamp 1654648307
transform 1 0 77600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_374
timestamp 1654648307
transform 1 0 79100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_455
timestamp 1654648307
transform 1 0 80600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_456
timestamp 1654648307
transform 1 0 82100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_375
timestamp 1654648307
transform 1 0 80600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_376
timestamp 1654648307
transform 1 0 82100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_457
timestamp 1654648307
transform 1 0 83600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_458
timestamp 1654648307
transform 1 0 85100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_377
timestamp 1654648307
transform 1 0 83600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_378
timestamp 1654648307
transform 1 0 85100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_459
timestamp 1654648307
transform 1 0 86600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_460
timestamp 1654648307
transform 1 0 88100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_379
timestamp 1654648307
transform 1 0 86600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_380
timestamp 1654648307
transform 1 0 88100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_461
timestamp 1654648307
transform 1 0 89600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_462
timestamp 1654648307
transform 1 0 91100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_381
timestamp 1654648307
transform 1 0 89600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_382
timestamp 1654648307
transform 1 0 91100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_463
timestamp 1654648307
transform 1 0 92600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_464
timestamp 1654648307
transform 1 0 94100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_383
timestamp 1654648307
transform 1 0 92600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_384
timestamp 1654648307
transform 1 0 94100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_465
timestamp 1654648307
transform 1 0 95600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_466
timestamp 1654648307
transform 1 0 97100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_385
timestamp 1654648307
transform 1 0 95600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_386
timestamp 1654648307
transform 1 0 97100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_467
timestamp 1654648307
transform 1 0 98600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_468
timestamp 1654648307
transform 1 0 100100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_387
timestamp 1654648307
transform 1 0 98600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_388
timestamp 1654648307
transform 1 0 100100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_469
timestamp 1654648307
transform 1 0 101600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_470
timestamp 1654648307
transform 1 0 103100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_389
timestamp 1654648307
transform 1 0 101600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_390
timestamp 1654648307
transform 1 0 103100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_471
timestamp 1654648307
transform 1 0 104600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_472
timestamp 1654648307
transform 1 0 106100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_391
timestamp 1654648307
transform 1 0 104600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_392
timestamp 1654648307
transform 1 0 106100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_473
timestamp 1654648307
transform 1 0 107600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_474
timestamp 1654648307
transform 1 0 109100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_393
timestamp 1654648307
transform 1 0 107600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_394
timestamp 1654648307
transform 1 0 109100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_475
timestamp 1654648307
transform 1 0 110600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_476
timestamp 1654648307
transform 1 0 112100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_395
timestamp 1654648307
transform 1 0 110600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_396
timestamp 1654648307
transform 1 0 112100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_477
timestamp 1654648307
transform 1 0 113600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_478
timestamp 1654648307
transform 1 0 115100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_397
timestamp 1654648307
transform 1 0 113600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_398
timestamp 1654648307
transform 1 0 115100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_479
timestamp 1654648307
transform 1 0 116600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_399
timestamp 1654648307
transform 1 0 116600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_240
timestamp 1654648307
transform 1 0 -1900 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_160
timestamp 1654648307
transform 1 0 -1900 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_241
timestamp 1654648307
transform 1 0 -400 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_242
timestamp 1654648307
transform 1 0 1100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_161
timestamp 1654648307
transform 1 0 -400 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_162
timestamp 1654648307
transform 1 0 1100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_243
timestamp 1654648307
transform 1 0 2600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_244
timestamp 1654648307
transform 1 0 4100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_163
timestamp 1654648307
transform 1 0 2600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_164
timestamp 1654648307
transform 1 0 4100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_245
timestamp 1654648307
transform 1 0 5600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_246
timestamp 1654648307
transform 1 0 7100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_165
timestamp 1654648307
transform 1 0 5600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_166
timestamp 1654648307
transform 1 0 7100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_247
timestamp 1654648307
transform 1 0 8600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_248
timestamp 1654648307
transform 1 0 10100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_167
timestamp 1654648307
transform 1 0 8600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_168
timestamp 1654648307
transform 1 0 10100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_249
timestamp 1654648307
transform 1 0 11600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_250
timestamp 1654648307
transform 1 0 13100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_169
timestamp 1654648307
transform 1 0 11600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_170
timestamp 1654648307
transform 1 0 13100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_251
timestamp 1654648307
transform 1 0 14600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_252
timestamp 1654648307
transform 1 0 16100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_171
timestamp 1654648307
transform 1 0 14600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_172
timestamp 1654648307
transform 1 0 16100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_253
timestamp 1654648307
transform 1 0 17600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_254
timestamp 1654648307
transform 1 0 19100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_173
timestamp 1654648307
transform 1 0 17600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_174
timestamp 1654648307
transform 1 0 19100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_255
timestamp 1654648307
transform 1 0 20600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_256
timestamp 1654648307
transform 1 0 22100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_175
timestamp 1654648307
transform 1 0 20600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_176
timestamp 1654648307
transform 1 0 22100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_257
timestamp 1654648307
transform 1 0 23600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_258
timestamp 1654648307
transform 1 0 25100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_177
timestamp 1654648307
transform 1 0 23600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_178
timestamp 1654648307
transform 1 0 25100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_259
timestamp 1654648307
transform 1 0 26600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_260
timestamp 1654648307
transform 1 0 28100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_179
timestamp 1654648307
transform 1 0 26600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_180
timestamp 1654648307
transform 1 0 28100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_261
timestamp 1654648307
transform 1 0 29600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_262
timestamp 1654648307
transform 1 0 31100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_181
timestamp 1654648307
transform 1 0 29600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_182
timestamp 1654648307
transform 1 0 31100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_263
timestamp 1654648307
transform 1 0 32600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_264
timestamp 1654648307
transform 1 0 34100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_183
timestamp 1654648307
transform 1 0 32600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_184
timestamp 1654648307
transform 1 0 34100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_265
timestamp 1654648307
transform 1 0 35600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_266
timestamp 1654648307
transform 1 0 37100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_185
timestamp 1654648307
transform 1 0 35600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_186
timestamp 1654648307
transform 1 0 37100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_267
timestamp 1654648307
transform 1 0 38600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_268
timestamp 1654648307
transform 1 0 40100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_187
timestamp 1654648307
transform 1 0 38600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_188
timestamp 1654648307
transform 1 0 40100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_269
timestamp 1654648307
transform 1 0 41600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_270
timestamp 1654648307
transform 1 0 43100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_189
timestamp 1654648307
transform 1 0 41600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_190
timestamp 1654648307
transform 1 0 43100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_271
timestamp 1654648307
transform 1 0 44600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_272
timestamp 1654648307
transform 1 0 46100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_191
timestamp 1654648307
transform 1 0 44600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_192
timestamp 1654648307
transform 1 0 46100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_273
timestamp 1654648307
transform 1 0 47600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_274
timestamp 1654648307
transform 1 0 49100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_193
timestamp 1654648307
transform 1 0 47600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_194
timestamp 1654648307
transform 1 0 49100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_275
timestamp 1654648307
transform 1 0 50600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_276
timestamp 1654648307
transform 1 0 52100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_195
timestamp 1654648307
transform 1 0 50600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_196
timestamp 1654648307
transform 1 0 52100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_277
timestamp 1654648307
transform 1 0 53600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_278
timestamp 1654648307
transform 1 0 55100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_197
timestamp 1654648307
transform 1 0 53600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_198
timestamp 1654648307
transform 1 0 55100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_279
timestamp 1654648307
transform 1 0 56600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_280
timestamp 1654648307
transform 1 0 58100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_199
timestamp 1654648307
transform 1 0 56600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_200
timestamp 1654648307
transform 1 0 58100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_281
timestamp 1654648307
transform 1 0 59600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_282
timestamp 1654648307
transform 1 0 61100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_201
timestamp 1654648307
transform 1 0 59600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_202
timestamp 1654648307
transform 1 0 61100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_283
timestamp 1654648307
transform 1 0 62600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_284
timestamp 1654648307
transform 1 0 64100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_203
timestamp 1654648307
transform 1 0 62600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_204
timestamp 1654648307
transform 1 0 64100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_285
timestamp 1654648307
transform 1 0 65600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_286
timestamp 1654648307
transform 1 0 67100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_205
timestamp 1654648307
transform 1 0 65600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_206
timestamp 1654648307
transform 1 0 67100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_287
timestamp 1654648307
transform 1 0 68600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_288
timestamp 1654648307
transform 1 0 70100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_207
timestamp 1654648307
transform 1 0 68600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_208
timestamp 1654648307
transform 1 0 70100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_289
timestamp 1654648307
transform 1 0 71600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_290
timestamp 1654648307
transform 1 0 73100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_209
timestamp 1654648307
transform 1 0 71600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_210
timestamp 1654648307
transform 1 0 73100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_291
timestamp 1654648307
transform 1 0 74600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_292
timestamp 1654648307
transform 1 0 76100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_211
timestamp 1654648307
transform 1 0 74600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_212
timestamp 1654648307
transform 1 0 76100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_293
timestamp 1654648307
transform 1 0 77600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_294
timestamp 1654648307
transform 1 0 79100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_213
timestamp 1654648307
transform 1 0 77600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_214
timestamp 1654648307
transform 1 0 79100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_295
timestamp 1654648307
transform 1 0 80600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_296
timestamp 1654648307
transform 1 0 82100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_215
timestamp 1654648307
transform 1 0 80600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_216
timestamp 1654648307
transform 1 0 82100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_297
timestamp 1654648307
transform 1 0 83600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_298
timestamp 1654648307
transform 1 0 85100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_217
timestamp 1654648307
transform 1 0 83600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_218
timestamp 1654648307
transform 1 0 85100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_299
timestamp 1654648307
transform 1 0 86600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_300
timestamp 1654648307
transform 1 0 88100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_219
timestamp 1654648307
transform 1 0 86600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_220
timestamp 1654648307
transform 1 0 88100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_301
timestamp 1654648307
transform 1 0 89600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_302
timestamp 1654648307
transform 1 0 91100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_221
timestamp 1654648307
transform 1 0 89600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_222
timestamp 1654648307
transform 1 0 91100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_303
timestamp 1654648307
transform 1 0 92600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_304
timestamp 1654648307
transform 1 0 94100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_223
timestamp 1654648307
transform 1 0 92600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_224
timestamp 1654648307
transform 1 0 94100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_305
timestamp 1654648307
transform 1 0 95600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_306
timestamp 1654648307
transform 1 0 97100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_225
timestamp 1654648307
transform 1 0 95600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_226
timestamp 1654648307
transform 1 0 97100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_307
timestamp 1654648307
transform 1 0 98600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_308
timestamp 1654648307
transform 1 0 100100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_227
timestamp 1654648307
transform 1 0 98600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_228
timestamp 1654648307
transform 1 0 100100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_309
timestamp 1654648307
transform 1 0 101600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_310
timestamp 1654648307
transform 1 0 103100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_229
timestamp 1654648307
transform 1 0 101600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_230
timestamp 1654648307
transform 1 0 103100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_311
timestamp 1654648307
transform 1 0 104600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_312
timestamp 1654648307
transform 1 0 106100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_231
timestamp 1654648307
transform 1 0 104600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_232
timestamp 1654648307
transform 1 0 106100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_313
timestamp 1654648307
transform 1 0 107600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_314
timestamp 1654648307
transform 1 0 109100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_233
timestamp 1654648307
transform 1 0 107600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_234
timestamp 1654648307
transform 1 0 109100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_315
timestamp 1654648307
transform 1 0 110600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_316
timestamp 1654648307
transform 1 0 112100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_235
timestamp 1654648307
transform 1 0 110600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_236
timestamp 1654648307
transform 1 0 112100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_317
timestamp 1654648307
transform 1 0 113600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_318
timestamp 1654648307
transform 1 0 115100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_237
timestamp 1654648307
transform 1 0 113600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_238
timestamp 1654648307
transform 1 0 115100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_319
timestamp 1654648307
transform 1 0 116600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_239
timestamp 1654648307
transform 1 0 116600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_80
timestamp 1654648307
transform 1 0 -1900 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_0
timestamp 1654648307
transform 1 0 -1900 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_81
timestamp 1654648307
transform 1 0 -400 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_82
timestamp 1654648307
transform 1 0 1100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_1
timestamp 1654648307
transform 1 0 -400 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_2
timestamp 1654648307
transform 1 0 1100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_83
timestamp 1654648307
transform 1 0 2600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_84
timestamp 1654648307
transform 1 0 4100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_3
timestamp 1654648307
transform 1 0 2600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_4
timestamp 1654648307
transform 1 0 4100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_85
timestamp 1654648307
transform 1 0 5600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_86
timestamp 1654648307
transform 1 0 7100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_5
timestamp 1654648307
transform 1 0 5600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_6
timestamp 1654648307
transform 1 0 7100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_87
timestamp 1654648307
transform 1 0 8600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_88
timestamp 1654648307
transform 1 0 10100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_7
timestamp 1654648307
transform 1 0 8600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_8
timestamp 1654648307
transform 1 0 10100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_89
timestamp 1654648307
transform 1 0 11600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_90
timestamp 1654648307
transform 1 0 13100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_9
timestamp 1654648307
transform 1 0 11600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_10
timestamp 1654648307
transform 1 0 13100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_91
timestamp 1654648307
transform 1 0 14600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_92
timestamp 1654648307
transform 1 0 16100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_11
timestamp 1654648307
transform 1 0 14600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_12
timestamp 1654648307
transform 1 0 16100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_93
timestamp 1654648307
transform 1 0 17600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_94
timestamp 1654648307
transform 1 0 19100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_13
timestamp 1654648307
transform 1 0 17600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_14
timestamp 1654648307
transform 1 0 19100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_95
timestamp 1654648307
transform 1 0 20600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_96
timestamp 1654648307
transform 1 0 22100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_15
timestamp 1654648307
transform 1 0 20600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_16
timestamp 1654648307
transform 1 0 22100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_97
timestamp 1654648307
transform 1 0 23600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_98
timestamp 1654648307
transform 1 0 25100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_17
timestamp 1654648307
transform 1 0 23600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_18
timestamp 1654648307
transform 1 0 25100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_99
timestamp 1654648307
transform 1 0 26600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_100
timestamp 1654648307
transform 1 0 28100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_19
timestamp 1654648307
transform 1 0 26600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_20
timestamp 1654648307
transform 1 0 28100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_101
timestamp 1654648307
transform 1 0 29600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_102
timestamp 1654648307
transform 1 0 31100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_21
timestamp 1654648307
transform 1 0 29600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_22
timestamp 1654648307
transform 1 0 31100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_103
timestamp 1654648307
transform 1 0 32600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_104
timestamp 1654648307
transform 1 0 34100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_23
timestamp 1654648307
transform 1 0 32600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_24
timestamp 1654648307
transform 1 0 34100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_105
timestamp 1654648307
transform 1 0 35600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_106
timestamp 1654648307
transform 1 0 37100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_25
timestamp 1654648307
transform 1 0 35600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_26
timestamp 1654648307
transform 1 0 37100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_107
timestamp 1654648307
transform 1 0 38600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_108
timestamp 1654648307
transform 1 0 40100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_27
timestamp 1654648307
transform 1 0 38600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_28
timestamp 1654648307
transform 1 0 40100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_109
timestamp 1654648307
transform 1 0 41600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_110
timestamp 1654648307
transform 1 0 43100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_29
timestamp 1654648307
transform 1 0 41600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_30
timestamp 1654648307
transform 1 0 43100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_111
timestamp 1654648307
transform 1 0 44600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_112
timestamp 1654648307
transform 1 0 46100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_31
timestamp 1654648307
transform 1 0 44600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_32
timestamp 1654648307
transform 1 0 46100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_113
timestamp 1654648307
transform 1 0 47600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_114
timestamp 1654648307
transform 1 0 49100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_33
timestamp 1654648307
transform 1 0 47600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_34
timestamp 1654648307
transform 1 0 49100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_115
timestamp 1654648307
transform 1 0 50600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_116
timestamp 1654648307
transform 1 0 52100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_35
timestamp 1654648307
transform 1 0 50600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_36
timestamp 1654648307
transform 1 0 52100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_117
timestamp 1654648307
transform 1 0 53600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_118
timestamp 1654648307
transform 1 0 55100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_37
timestamp 1654648307
transform 1 0 53600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_38
timestamp 1654648307
transform 1 0 55100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_119
timestamp 1654648307
transform 1 0 56600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_120
timestamp 1654648307
transform 1 0 58100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_39
timestamp 1654648307
transform 1 0 56600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_40
timestamp 1654648307
transform 1 0 58100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_121
timestamp 1654648307
transform 1 0 59600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_122
timestamp 1654648307
transform 1 0 61100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_41
timestamp 1654648307
transform 1 0 59600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_42
timestamp 1654648307
transform 1 0 61100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_123
timestamp 1654648307
transform 1 0 62600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_124
timestamp 1654648307
transform 1 0 64100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_43
timestamp 1654648307
transform 1 0 62600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_44
timestamp 1654648307
transform 1 0 64100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_125
timestamp 1654648307
transform 1 0 65600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_126
timestamp 1654648307
transform 1 0 67100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_45
timestamp 1654648307
transform 1 0 65600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_46
timestamp 1654648307
transform 1 0 67100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_127
timestamp 1654648307
transform 1 0 68600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_128
timestamp 1654648307
transform 1 0 70100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_47
timestamp 1654648307
transform 1 0 68600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_48
timestamp 1654648307
transform 1 0 70100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_129
timestamp 1654648307
transform 1 0 71600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_130
timestamp 1654648307
transform 1 0 73100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_49
timestamp 1654648307
transform 1 0 71600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_50
timestamp 1654648307
transform 1 0 73100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_131
timestamp 1654648307
transform 1 0 74600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_132
timestamp 1654648307
transform 1 0 76100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_51
timestamp 1654648307
transform 1 0 74600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_52
timestamp 1654648307
transform 1 0 76100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_133
timestamp 1654648307
transform 1 0 77600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_134
timestamp 1654648307
transform 1 0 79100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_53
timestamp 1654648307
transform 1 0 77600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_54
timestamp 1654648307
transform 1 0 79100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_135
timestamp 1654648307
transform 1 0 80600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_136
timestamp 1654648307
transform 1 0 82100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_55
timestamp 1654648307
transform 1 0 80600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_56
timestamp 1654648307
transform 1 0 82100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_137
timestamp 1654648307
transform 1 0 83600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_138
timestamp 1654648307
transform 1 0 85100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_57
timestamp 1654648307
transform 1 0 83600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_58
timestamp 1654648307
transform 1 0 85100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_139
timestamp 1654648307
transform 1 0 86600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_140
timestamp 1654648307
transform 1 0 88100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_59
timestamp 1654648307
transform 1 0 86600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_60
timestamp 1654648307
transform 1 0 88100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_141
timestamp 1654648307
transform 1 0 89600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_142
timestamp 1654648307
transform 1 0 91100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_61
timestamp 1654648307
transform 1 0 89600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_62
timestamp 1654648307
transform 1 0 91100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_143
timestamp 1654648307
transform 1 0 92600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_144
timestamp 1654648307
transform 1 0 94100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_63
timestamp 1654648307
transform 1 0 92600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_64
timestamp 1654648307
transform 1 0 94100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_145
timestamp 1654648307
transform 1 0 95600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_146
timestamp 1654648307
transform 1 0 97100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_65
timestamp 1654648307
transform 1 0 95600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_66
timestamp 1654648307
transform 1 0 97100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_147
timestamp 1654648307
transform 1 0 98600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_148
timestamp 1654648307
transform 1 0 100100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_67
timestamp 1654648307
transform 1 0 98600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_68
timestamp 1654648307
transform 1 0 100100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_149
timestamp 1654648307
transform 1 0 101600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_150
timestamp 1654648307
transform 1 0 103100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_69
timestamp 1654648307
transform 1 0 101600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_70
timestamp 1654648307
transform 1 0 103100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_151
timestamp 1654648307
transform 1 0 104600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_152
timestamp 1654648307
transform 1 0 106100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_71
timestamp 1654648307
transform 1 0 104600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_72
timestamp 1654648307
transform 1 0 106100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_153
timestamp 1654648307
transform 1 0 107600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_154
timestamp 1654648307
transform 1 0 109100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_73
timestamp 1654648307
transform 1 0 107600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_74
timestamp 1654648307
transform 1 0 109100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_155
timestamp 1654648307
transform 1 0 110600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_156
timestamp 1654648307
transform 1 0 112100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_75
timestamp 1654648307
transform 1 0 110600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_76
timestamp 1654648307
transform 1 0 112100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_157
timestamp 1654648307
transform 1 0 113600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_158
timestamp 1654648307
transform 1 0 115100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_77
timestamp 1654648307
transform 1 0 113600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_78
timestamp 1654648307
transform 1 0 115100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_159
timestamp 1654648307
transform 1 0 116600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_79
timestamp 1654648307
transform 1 0 116600 0 1 1350
box 1820 -1430 3480 230
<< labels >>
rlabel metal5 520 520 620 620 1 PIX0_IN
port 1 n
rlabel metal4 -1500 1775 -1500 1830 1 VBIAS
port 2 n
rlabel metal2 -1500 1675 -1500 1725 3 VREF
port 3 e
rlabel metal2 0 2020 0 2020 1 NB2
port 4 n
rlabel metal1 -1000 0 -1000 0 1 VDD
port 5 n
rlabel space -580 2875 -580 2875 5 SF_IB
port 6 s
rlabel metal2 -370 1780 -370 1780 1 NB1
port 7 n
rlabel metal2 -1500 740 -1500 785 3 ROW_SEL0
port 8 e
rlabel metal5 -1000 1420 -1000 1420 1 GRING
port 9 n
rlabel metal5 2020 520 2120 620 1 PIX1_IN
port 10 n
rlabel metal5 3520 520 3620 620 1 PIX2_IN
port 11 n
rlabel metal5 5020 520 5120 620 1 PIX3_IN
port 12 n
rlabel metal5 6520 520 6620 620 1 PIX4_IN
port 13 n
rlabel metal5 8020 520 8120 620 1 PIX5_IN
port 14 n
rlabel metal5 9520 520 9620 620 1 PIX6_IN
port 15 n
rlabel metal5 11020 520 11120 620 1 PIX7_IN
port 16 n
rlabel metal5 12520 520 12620 620 1 PIX8_IN
port 17 n
rlabel metal5 14020 520 14120 620 1 PIX9_IN
port 18 n
rlabel metal5 15520 520 15620 620 1 PIX10_IN
port 19 n
rlabel metal5 17020 520 17120 620 1 PIX11_IN
port 20 n
rlabel metal5 18520 520 18620 620 1 PIX12_IN
port 21 n
rlabel metal5 20020 520 20120 620 1 PIX13_IN
port 22 n
rlabel metal5 21520 520 21620 620 1 PIX14_IN
port 23 n
rlabel metal5 23020 520 23120 620 1 PIX15_IN
port 24 n
rlabel metal5 24520 520 24620 620 1 PIX16_IN
port 25 n
rlabel metal5 26020 520 26120 620 1 PIX17_IN
port 26 n
rlabel metal5 27520 520 27620 620 1 PIX18_IN
port 27 n
rlabel metal5 29020 520 29120 620 1 PIX19_IN
port 28 n
rlabel metal5 30520 520 30620 620 1 PIX20_IN
port 29 n
rlabel metal5 32020 520 32120 620 1 PIX21_IN
port 30 n
rlabel metal5 33520 520 33620 620 1 PIX22_IN
port 31 n
rlabel metal5 35020 520 35120 620 1 PIX23_IN
port 32 n
rlabel metal5 36520 520 36620 620 1 PIX24_IN
port 33 n
rlabel metal5 38020 520 38120 620 1 PIX25_IN
port 34 n
rlabel metal5 39520 520 39620 620 1 PIX26_IN
port 35 n
rlabel metal5 41020 520 41120 620 1 PIX27_IN
port 36 n
rlabel metal5 42520 520 42620 620 1 PIX28_IN
port 37 n
rlabel metal5 44020 520 44120 620 1 PIX29_IN
port 38 n
rlabel metal5 45520 520 45620 620 1 PIX30_IN
port 39 n
rlabel metal5 47020 520 47120 620 1 PIX31_IN
port 40 n
rlabel metal5 48520 520 48620 620 1 PIX32_IN
port 41 n
rlabel metal5 50020 520 50120 620 1 PIX33_IN
port 42 n
rlabel metal5 51520 520 51620 620 1 PIX34_IN
port 43 n
rlabel metal5 53020 520 53120 620 1 PIX35_IN
port 44 n
rlabel metal5 54520 520 54620 620 1 PIX36_IN
port 45 n
rlabel metal5 56020 520 56120 620 1 PIX37_IN
port 46 n
rlabel metal5 57520 520 57620 620 1 PIX38_IN
port 47 n
rlabel metal5 59020 520 59120 620 1 PIX39_IN
port 48 n
rlabel metal5 60520 520 60620 620 1 PIX40_IN
port 49 n
rlabel metal5 62020 520 62120 620 1 PIX41_IN
port 50 n
rlabel metal5 63520 520 63620 620 1 PIX42_IN
port 51 n
rlabel metal5 65020 520 65120 620 1 PIX43_IN
port 52 n
rlabel metal5 66520 520 66620 620 1 PIX44_IN
port 53 n
rlabel metal5 68020 520 68120 620 1 PIX45_IN
port 54 n
rlabel metal5 69520 520 69620 620 1 PIX46_IN
port 55 n
rlabel metal5 71020 520 71120 620 1 PIX47_IN
port 56 n
rlabel metal5 72520 520 72620 620 1 PIX48_IN
port 57 n
rlabel metal5 74020 520 74120 620 1 PIX49_IN
port 58 n
rlabel metal5 75520 520 75620 620 1 PIX50_IN
port 59 n
rlabel metal5 77020 520 77120 620 1 PIX51_IN
port 60 n
rlabel metal5 78520 520 78620 620 1 PIX52_IN
port 61 n
rlabel metal5 80020 520 80120 620 1 PIX53_IN
port 62 n
rlabel metal5 81520 520 81620 620 1 PIX54_IN
port 63 n
rlabel metal5 83020 520 83120 620 1 PIX55_IN
port 64 n
rlabel metal5 84520 520 84620 620 1 PIX56_IN
port 65 n
rlabel metal5 86020 520 86120 620 1 PIX57_IN
port 66 n
rlabel metal5 87520 520 87620 620 1 PIX58_IN
port 67 n
rlabel metal5 89020 520 89120 620 1 PIX59_IN
port 68 n
rlabel metal5 90520 520 90620 620 1 PIX60_IN
port 69 n
rlabel metal5 92020 520 92120 620 1 PIX61_IN
port 70 n
rlabel metal5 93520 520 93620 620 1 PIX62_IN
port 71 n
rlabel metal5 95020 520 95120 620 1 PIX63_IN
port 72 n
rlabel metal5 96520 520 96620 620 1 PIX64_IN
port 73 n
rlabel metal5 98020 520 98120 620 1 PIX65_IN
port 74 n
rlabel metal5 99520 520 99620 620 1 PIX66_IN
port 75 n
rlabel metal5 101020 520 101120 620 1 PIX67_IN
port 76 n
rlabel metal5 102520 520 102620 620 1 PIX68_IN
port 77 n
rlabel metal5 104020 520 104120 620 1 PIX69_IN
port 78 n
rlabel metal5 105520 520 105620 620 1 PIX70_IN
port 79 n
rlabel metal5 107020 520 107120 620 1 PIX71_IN
port 80 n
rlabel metal5 108520 520 108620 620 1 PIX72_IN
port 81 n
rlabel metal5 110020 520 110120 620 1 PIX73_IN
port 82 n
rlabel metal5 111520 520 111620 620 1 PIX74_IN
port 83 n
rlabel metal5 113020 520 113120 620 1 PIX75_IN
port 84 n
rlabel metal5 114520 520 114620 620 1 PIX76_IN
port 85 n
rlabel metal5 116020 520 116120 620 1 PIX77_IN
port 86 n
rlabel metal5 117520 520 117620 620 1 PIX78_IN
port 87 n
rlabel metal5 119020 520 119120 620 1 PIX79_IN
port 88 n
rlabel metal1 120200 15 120200 15 1 GND
port 89 n
rlabel metal5 520 -980 620 -880 1 PIX80_IN
port 90 n
rlabel metal2 -1500 -760 -1500 -715 3 ROW_SEL1
port 91 e
rlabel metal5 2020 -980 2120 -880 1 PIX81_IN
port 92 n
rlabel metal5 3520 -980 3620 -880 1 PIX82_IN
port 93 n
rlabel metal5 5020 -980 5120 -880 1 PIX83_IN
port 94 n
rlabel metal5 6520 -980 6620 -880 1 PIX84_IN
port 95 n
rlabel metal5 8020 -980 8120 -880 1 PIX85_IN
port 96 n
rlabel metal5 9520 -980 9620 -880 1 PIX86_IN
port 97 n
rlabel metal5 11020 -980 11120 -880 1 PIX87_IN
port 98 n
rlabel metal5 12520 -980 12620 -880 1 PIX88_IN
port 99 n
rlabel metal5 14020 -980 14120 -880 1 PIX89_IN
port 100 n
rlabel metal5 15520 -980 15620 -880 1 PIX90_IN
port 101 n
rlabel metal5 17020 -980 17120 -880 1 PIX91_IN
port 102 n
rlabel metal5 18520 -980 18620 -880 1 PIX92_IN
port 103 n
rlabel metal5 20020 -980 20120 -880 1 PIX93_IN
port 104 n
rlabel metal5 21520 -980 21620 -880 1 PIX94_IN
port 105 n
rlabel metal5 23020 -980 23120 -880 1 PIX95_IN
port 106 n
rlabel metal5 24520 -980 24620 -880 1 PIX96_IN
port 107 n
rlabel metal5 26020 -980 26120 -880 1 PIX97_IN
port 108 n
rlabel metal5 27520 -980 27620 -880 1 PIX98_IN
port 109 n
rlabel metal5 29020 -980 29120 -880 1 PIX99_IN
port 110 n
rlabel metal5 30520 -980 30620 -880 1 PIX100_IN
port 111 n
rlabel metal5 32020 -980 32120 -880 1 PIX101_IN
port 112 n
rlabel metal5 33520 -980 33620 -880 1 PIX102_IN
port 113 n
rlabel metal5 35020 -980 35120 -880 1 PIX103_IN
port 114 n
rlabel metal5 36520 -980 36620 -880 1 PIX104_IN
port 115 n
rlabel metal5 38020 -980 38120 -880 1 PIX105_IN
port 116 n
rlabel metal5 39520 -980 39620 -880 1 PIX106_IN
port 117 n
rlabel metal5 41020 -980 41120 -880 1 PIX107_IN
port 118 n
rlabel metal5 42520 -980 42620 -880 1 PIX108_IN
port 119 n
rlabel metal5 44020 -980 44120 -880 1 PIX109_IN
port 120 n
rlabel metal5 45520 -980 45620 -880 1 PIX110_IN
port 121 n
rlabel metal5 47020 -980 47120 -880 1 PIX111_IN
port 122 n
rlabel metal5 48520 -980 48620 -880 1 PIX112_IN
port 123 n
rlabel metal5 50020 -980 50120 -880 1 PIX113_IN
port 124 n
rlabel metal5 51520 -980 51620 -880 1 PIX114_IN
port 125 n
rlabel metal5 53020 -980 53120 -880 1 PIX115_IN
port 126 n
rlabel metal5 54520 -980 54620 -880 1 PIX116_IN
port 127 n
rlabel metal5 56020 -980 56120 -880 1 PIX117_IN
port 128 n
rlabel metal5 57520 -980 57620 -880 1 PIX118_IN
port 129 n
rlabel metal5 59020 -980 59120 -880 1 PIX119_IN
port 130 n
rlabel metal5 60520 -980 60620 -880 1 PIX120_IN
port 131 n
rlabel metal5 62020 -980 62120 -880 1 PIX121_IN
port 132 n
rlabel metal5 63520 -980 63620 -880 1 PIX122_IN
port 133 n
rlabel metal5 65020 -980 65120 -880 1 PIX123_IN
port 134 n
rlabel metal5 66520 -980 66620 -880 1 PIX124_IN
port 135 n
rlabel metal5 68020 -980 68120 -880 1 PIX125_IN
port 136 n
rlabel metal5 69520 -980 69620 -880 1 PIX126_IN
port 137 n
rlabel metal5 71020 -980 71120 -880 1 PIX127_IN
port 138 n
rlabel metal5 72520 -980 72620 -880 1 PIX128_IN
port 139 n
rlabel metal5 74020 -980 74120 -880 1 PIX129_IN
port 140 n
rlabel metal5 75520 -980 75620 -880 1 PIX130_IN
port 141 n
rlabel metal5 77020 -980 77120 -880 1 PIX131_IN
port 142 n
rlabel metal5 78520 -980 78620 -880 1 PIX132_IN
port 143 n
rlabel metal5 80020 -980 80120 -880 1 PIX133_IN
port 144 n
rlabel metal5 81520 -980 81620 -880 1 PIX134_IN
port 145 n
rlabel metal5 83020 -980 83120 -880 1 PIX135_IN
port 146 n
rlabel metal5 84520 -980 84620 -880 1 PIX136_IN
port 147 n
rlabel metal5 86020 -980 86120 -880 1 PIX137_IN
port 148 n
rlabel metal5 87520 -980 87620 -880 1 PIX138_IN
port 149 n
rlabel metal5 89020 -980 89120 -880 1 PIX139_IN
port 150 n
rlabel metal5 90520 -980 90620 -880 1 PIX140_IN
port 151 n
rlabel metal5 92020 -980 92120 -880 1 PIX141_IN
port 152 n
rlabel metal5 93520 -980 93620 -880 1 PIX142_IN
port 153 n
rlabel metal5 95020 -980 95120 -880 1 PIX143_IN
port 154 n
rlabel metal5 96520 -980 96620 -880 1 PIX144_IN
port 155 n
rlabel metal5 98020 -980 98120 -880 1 PIX145_IN
port 156 n
rlabel metal5 99520 -980 99620 -880 1 PIX146_IN
port 157 n
rlabel metal5 101020 -980 101120 -880 1 PIX147_IN
port 158 n
rlabel metal5 102520 -980 102620 -880 1 PIX148_IN
port 159 n
rlabel metal5 104020 -980 104120 -880 1 PIX149_IN
port 160 n
rlabel metal5 105520 -980 105620 -880 1 PIX150_IN
port 161 n
rlabel metal5 107020 -980 107120 -880 1 PIX151_IN
port 162 n
rlabel metal5 108520 -980 108620 -880 1 PIX152_IN
port 163 n
rlabel metal5 110020 -980 110120 -880 1 PIX153_IN
port 164 n
rlabel metal5 111520 -980 111620 -880 1 PIX154_IN
port 165 n
rlabel metal5 113020 -980 113120 -880 1 PIX155_IN
port 166 n
rlabel metal5 114520 -980 114620 -880 1 PIX156_IN
port 167 n
rlabel metal5 116020 -980 116120 -880 1 PIX157_IN
port 168 n
rlabel metal5 117520 -980 117620 -880 1 PIX158_IN
port 169 n
rlabel metal5 119020 -980 119120 -880 1 PIX159_IN
port 170 n
rlabel metal5 520 -2480 620 -2380 1 PIX160_IN
port 171 n
rlabel metal2 -1500 -2260 -1500 -2215 3 ROW_SEL2
port 172 e
rlabel metal5 2020 -2480 2120 -2380 1 PIX161_IN
port 173 n
rlabel metal5 3520 -2480 3620 -2380 1 PIX162_IN
port 174 n
rlabel metal5 5020 -2480 5120 -2380 1 PIX163_IN
port 175 n
rlabel metal5 6520 -2480 6620 -2380 1 PIX164_IN
port 176 n
rlabel metal5 8020 -2480 8120 -2380 1 PIX165_IN
port 177 n
rlabel metal5 9520 -2480 9620 -2380 1 PIX166_IN
port 178 n
rlabel metal5 11020 -2480 11120 -2380 1 PIX167_IN
port 179 n
rlabel metal5 12520 -2480 12620 -2380 1 PIX168_IN
port 180 n
rlabel metal5 14020 -2480 14120 -2380 1 PIX169_IN
port 181 n
rlabel metal5 15520 -2480 15620 -2380 1 PIX170_IN
port 182 n
rlabel metal5 17020 -2480 17120 -2380 1 PIX171_IN
port 183 n
rlabel metal5 18520 -2480 18620 -2380 1 PIX172_IN
port 184 n
rlabel metal5 20020 -2480 20120 -2380 1 PIX173_IN
port 185 n
rlabel metal5 21520 -2480 21620 -2380 1 PIX174_IN
port 186 n
rlabel metal5 23020 -2480 23120 -2380 1 PIX175_IN
port 187 n
rlabel metal5 24520 -2480 24620 -2380 1 PIX176_IN
port 188 n
rlabel metal5 26020 -2480 26120 -2380 1 PIX177_IN
port 189 n
rlabel metal5 27520 -2480 27620 -2380 1 PIX178_IN
port 190 n
rlabel metal5 29020 -2480 29120 -2380 1 PIX179_IN
port 191 n
rlabel metal5 30520 -2480 30620 -2380 1 PIX180_IN
port 192 n
rlabel metal5 32020 -2480 32120 -2380 1 PIX181_IN
port 193 n
rlabel metal5 33520 -2480 33620 -2380 1 PIX182_IN
port 194 n
rlabel metal5 35020 -2480 35120 -2380 1 PIX183_IN
port 195 n
rlabel metal5 36520 -2480 36620 -2380 1 PIX184_IN
port 196 n
rlabel metal5 38020 -2480 38120 -2380 1 PIX185_IN
port 197 n
rlabel metal5 39520 -2480 39620 -2380 1 PIX186_IN
port 198 n
rlabel metal5 41020 -2480 41120 -2380 1 PIX187_IN
port 199 n
rlabel metal5 42520 -2480 42620 -2380 1 PIX188_IN
port 200 n
rlabel metal5 44020 -2480 44120 -2380 1 PIX189_IN
port 201 n
rlabel metal5 45520 -2480 45620 -2380 1 PIX190_IN
port 202 n
rlabel metal5 47020 -2480 47120 -2380 1 PIX191_IN
port 203 n
rlabel metal5 48520 -2480 48620 -2380 1 PIX192_IN
port 204 n
rlabel metal5 50020 -2480 50120 -2380 1 PIX193_IN
port 205 n
rlabel metal5 51520 -2480 51620 -2380 1 PIX194_IN
port 206 n
rlabel metal5 53020 -2480 53120 -2380 1 PIX195_IN
port 207 n
rlabel metal5 54520 -2480 54620 -2380 1 PIX196_IN
port 208 n
rlabel metal5 56020 -2480 56120 -2380 1 PIX197_IN
port 209 n
rlabel metal5 57520 -2480 57620 -2380 1 PIX198_IN
port 210 n
rlabel metal5 59020 -2480 59120 -2380 1 PIX199_IN
port 211 n
rlabel metal5 60520 -2480 60620 -2380 1 PIX200_IN
port 212 n
rlabel metal5 62020 -2480 62120 -2380 1 PIX201_IN
port 213 n
rlabel metal5 63520 -2480 63620 -2380 1 PIX202_IN
port 214 n
rlabel metal5 65020 -2480 65120 -2380 1 PIX203_IN
port 215 n
rlabel metal5 66520 -2480 66620 -2380 1 PIX204_IN
port 216 n
rlabel metal5 68020 -2480 68120 -2380 1 PIX205_IN
port 217 n
rlabel metal5 69520 -2480 69620 -2380 1 PIX206_IN
port 218 n
rlabel metal5 71020 -2480 71120 -2380 1 PIX207_IN
port 219 n
rlabel metal5 72520 -2480 72620 -2380 1 PIX208_IN
port 220 n
rlabel metal5 74020 -2480 74120 -2380 1 PIX209_IN
port 221 n
rlabel metal5 75520 -2480 75620 -2380 1 PIX210_IN
port 222 n
rlabel metal5 77020 -2480 77120 -2380 1 PIX211_IN
port 223 n
rlabel metal5 78520 -2480 78620 -2380 1 PIX212_IN
port 224 n
rlabel metal5 80020 -2480 80120 -2380 1 PIX213_IN
port 225 n
rlabel metal5 81520 -2480 81620 -2380 1 PIX214_IN
port 226 n
rlabel metal5 83020 -2480 83120 -2380 1 PIX215_IN
port 227 n
rlabel metal5 84520 -2480 84620 -2380 1 PIX216_IN
port 228 n
rlabel metal5 86020 -2480 86120 -2380 1 PIX217_IN
port 229 n
rlabel metal5 87520 -2480 87620 -2380 1 PIX218_IN
port 230 n
rlabel metal5 89020 -2480 89120 -2380 1 PIX219_IN
port 231 n
rlabel metal5 90520 -2480 90620 -2380 1 PIX220_IN
port 232 n
rlabel metal5 92020 -2480 92120 -2380 1 PIX221_IN
port 233 n
rlabel metal5 93520 -2480 93620 -2380 1 PIX222_IN
port 234 n
rlabel metal5 95020 -2480 95120 -2380 1 PIX223_IN
port 235 n
rlabel metal5 96520 -2480 96620 -2380 1 PIX224_IN
port 236 n
rlabel metal5 98020 -2480 98120 -2380 1 PIX225_IN
port 237 n
rlabel metal5 99520 -2480 99620 -2380 1 PIX226_IN
port 238 n
rlabel metal5 101020 -2480 101120 -2380 1 PIX227_IN
port 239 n
rlabel metal5 102520 -2480 102620 -2380 1 PIX228_IN
port 240 n
rlabel metal5 104020 -2480 104120 -2380 1 PIX229_IN
port 241 n
rlabel metal5 105520 -2480 105620 -2380 1 PIX230_IN
port 242 n
rlabel metal5 107020 -2480 107120 -2380 1 PIX231_IN
port 243 n
rlabel metal5 108520 -2480 108620 -2380 1 PIX232_IN
port 244 n
rlabel metal5 110020 -2480 110120 -2380 1 PIX233_IN
port 245 n
rlabel metal5 111520 -2480 111620 -2380 1 PIX234_IN
port 246 n
rlabel metal5 113020 -2480 113120 -2380 1 PIX235_IN
port 247 n
rlabel metal5 114520 -2480 114620 -2380 1 PIX236_IN
port 248 n
rlabel metal5 116020 -2480 116120 -2380 1 PIX237_IN
port 249 n
rlabel metal5 117520 -2480 117620 -2380 1 PIX238_IN
port 250 n
rlabel metal5 119020 -2480 119120 -2380 1 PIX239_IN
port 251 n
rlabel metal5 520 -3980 620 -3880 1 PIX240_IN
port 252 n
rlabel metal2 -1500 -3760 -1500 -3715 3 ROW_SEL3
port 253 e
rlabel metal5 2020 -3980 2120 -3880 1 PIX241_IN
port 254 n
rlabel metal5 3520 -3980 3620 -3880 1 PIX242_IN
port 255 n
rlabel metal5 5020 -3980 5120 -3880 1 PIX243_IN
port 256 n
rlabel metal5 6520 -3980 6620 -3880 1 PIX244_IN
port 257 n
rlabel metal5 8020 -3980 8120 -3880 1 PIX245_IN
port 258 n
rlabel metal5 9520 -3980 9620 -3880 1 PIX246_IN
port 259 n
rlabel metal5 11020 -3980 11120 -3880 1 PIX247_IN
port 260 n
rlabel metal5 12520 -3980 12620 -3880 1 PIX248_IN
port 261 n
rlabel metal5 14020 -3980 14120 -3880 1 PIX249_IN
port 262 n
rlabel metal5 15520 -3980 15620 -3880 1 PIX250_IN
port 263 n
rlabel metal5 17020 -3980 17120 -3880 1 PIX251_IN
port 264 n
rlabel metal5 18520 -3980 18620 -3880 1 PIX252_IN
port 265 n
rlabel metal5 20020 -3980 20120 -3880 1 PIX253_IN
port 266 n
rlabel metal5 21520 -3980 21620 -3880 1 PIX254_IN
port 267 n
rlabel metal5 23020 -3980 23120 -3880 1 PIX255_IN
port 268 n
rlabel metal5 24520 -3980 24620 -3880 1 PIX256_IN
port 269 n
rlabel metal5 26020 -3980 26120 -3880 1 PIX257_IN
port 270 n
rlabel metal5 27520 -3980 27620 -3880 1 PIX258_IN
port 271 n
rlabel metal5 29020 -3980 29120 -3880 1 PIX259_IN
port 272 n
rlabel metal5 30520 -3980 30620 -3880 1 PIX260_IN
port 273 n
rlabel metal5 32020 -3980 32120 -3880 1 PIX261_IN
port 274 n
rlabel metal5 33520 -3980 33620 -3880 1 PIX262_IN
port 275 n
rlabel metal5 35020 -3980 35120 -3880 1 PIX263_IN
port 276 n
rlabel metal5 36520 -3980 36620 -3880 1 PIX264_IN
port 277 n
rlabel metal5 38020 -3980 38120 -3880 1 PIX265_IN
port 278 n
rlabel metal5 39520 -3980 39620 -3880 1 PIX266_IN
port 279 n
rlabel metal5 41020 -3980 41120 -3880 1 PIX267_IN
port 280 n
rlabel metal5 42520 -3980 42620 -3880 1 PIX268_IN
port 281 n
rlabel metal5 44020 -3980 44120 -3880 1 PIX269_IN
port 282 n
rlabel metal5 45520 -3980 45620 -3880 1 PIX270_IN
port 283 n
rlabel metal5 47020 -3980 47120 -3880 1 PIX271_IN
port 284 n
rlabel metal5 48520 -3980 48620 -3880 1 PIX272_IN
port 285 n
rlabel metal5 50020 -3980 50120 -3880 1 PIX273_IN
port 286 n
rlabel metal5 51520 -3980 51620 -3880 1 PIX274_IN
port 287 n
rlabel metal5 53020 -3980 53120 -3880 1 PIX275_IN
port 288 n
rlabel metal5 54520 -3980 54620 -3880 1 PIX276_IN
port 289 n
rlabel metal5 56020 -3980 56120 -3880 1 PIX277_IN
port 290 n
rlabel metal5 57520 -3980 57620 -3880 1 PIX278_IN
port 291 n
rlabel metal5 59020 -3980 59120 -3880 1 PIX279_IN
port 292 n
rlabel metal5 60520 -3980 60620 -3880 1 PIX280_IN
port 293 n
rlabel metal5 62020 -3980 62120 -3880 1 PIX281_IN
port 294 n
rlabel metal5 63520 -3980 63620 -3880 1 PIX282_IN
port 295 n
rlabel metal5 65020 -3980 65120 -3880 1 PIX283_IN
port 296 n
rlabel metal5 66520 -3980 66620 -3880 1 PIX284_IN
port 297 n
rlabel metal5 68020 -3980 68120 -3880 1 PIX285_IN
port 298 n
rlabel metal5 69520 -3980 69620 -3880 1 PIX286_IN
port 299 n
rlabel metal5 71020 -3980 71120 -3880 1 PIX287_IN
port 300 n
rlabel metal5 72520 -3980 72620 -3880 1 PIX288_IN
port 301 n
rlabel metal5 74020 -3980 74120 -3880 1 PIX289_IN
port 302 n
rlabel metal5 75520 -3980 75620 -3880 1 PIX290_IN
port 303 n
rlabel metal5 77020 -3980 77120 -3880 1 PIX291_IN
port 304 n
rlabel metal5 78520 -3980 78620 -3880 1 PIX292_IN
port 305 n
rlabel metal5 80020 -3980 80120 -3880 1 PIX293_IN
port 306 n
rlabel metal5 81520 -3980 81620 -3880 1 PIX294_IN
port 307 n
rlabel metal5 83020 -3980 83120 -3880 1 PIX295_IN
port 308 n
rlabel metal5 84520 -3980 84620 -3880 1 PIX296_IN
port 309 n
rlabel metal5 86020 -3980 86120 -3880 1 PIX297_IN
port 310 n
rlabel metal5 87520 -3980 87620 -3880 1 PIX298_IN
port 311 n
rlabel metal5 89020 -3980 89120 -3880 1 PIX299_IN
port 312 n
rlabel metal5 90520 -3980 90620 -3880 1 PIX300_IN
port 313 n
rlabel metal5 92020 -3980 92120 -3880 1 PIX301_IN
port 314 n
rlabel metal5 93520 -3980 93620 -3880 1 PIX302_IN
port 315 n
rlabel metal5 95020 -3980 95120 -3880 1 PIX303_IN
port 316 n
rlabel metal5 96520 -3980 96620 -3880 1 PIX304_IN
port 317 n
rlabel metal5 98020 -3980 98120 -3880 1 PIX305_IN
port 318 n
rlabel metal5 99520 -3980 99620 -3880 1 PIX306_IN
port 319 n
rlabel metal5 101020 -3980 101120 -3880 1 PIX307_IN
port 320 n
rlabel metal5 102520 -3980 102620 -3880 1 PIX308_IN
port 321 n
rlabel metal5 104020 -3980 104120 -3880 1 PIX309_IN
port 322 n
rlabel metal5 105520 -3980 105620 -3880 1 PIX310_IN
port 323 n
rlabel metal5 107020 -3980 107120 -3880 1 PIX311_IN
port 324 n
rlabel metal5 108520 -3980 108620 -3880 1 PIX312_IN
port 325 n
rlabel metal5 110020 -3980 110120 -3880 1 PIX313_IN
port 326 n
rlabel metal5 111520 -3980 111620 -3880 1 PIX314_IN
port 327 n
rlabel metal5 113020 -3980 113120 -3880 1 PIX315_IN
port 328 n
rlabel metal5 114520 -3980 114620 -3880 1 PIX316_IN
port 329 n
rlabel metal5 116020 -3980 116120 -3880 1 PIX317_IN
port 330 n
rlabel metal5 117520 -3980 117620 -3880 1 PIX318_IN
port 331 n
rlabel metal5 119020 -3980 119120 -3880 1 PIX319_IN
port 332 n
rlabel metal5 520 -5480 620 -5380 1 PIX320_IN
port 333 n
rlabel metal2 -1500 -5260 -1500 -5215 3 ROW_SEL4
port 334 e
rlabel metal5 2020 -5480 2120 -5380 1 PIX321_IN
port 335 n
rlabel metal5 3520 -5480 3620 -5380 1 PIX322_IN
port 336 n
rlabel metal5 5020 -5480 5120 -5380 1 PIX323_IN
port 337 n
rlabel metal5 6520 -5480 6620 -5380 1 PIX324_IN
port 338 n
rlabel metal5 8020 -5480 8120 -5380 1 PIX325_IN
port 339 n
rlabel metal5 9520 -5480 9620 -5380 1 PIX326_IN
port 340 n
rlabel metal5 11020 -5480 11120 -5380 1 PIX327_IN
port 341 n
rlabel metal5 12520 -5480 12620 -5380 1 PIX328_IN
port 342 n
rlabel metal5 14020 -5480 14120 -5380 1 PIX329_IN
port 343 n
rlabel metal5 15520 -5480 15620 -5380 1 PIX330_IN
port 344 n
rlabel metal5 17020 -5480 17120 -5380 1 PIX331_IN
port 345 n
rlabel metal5 18520 -5480 18620 -5380 1 PIX332_IN
port 346 n
rlabel metal5 20020 -5480 20120 -5380 1 PIX333_IN
port 347 n
rlabel metal5 21520 -5480 21620 -5380 1 PIX334_IN
port 348 n
rlabel metal5 23020 -5480 23120 -5380 1 PIX335_IN
port 349 n
rlabel metal5 24520 -5480 24620 -5380 1 PIX336_IN
port 350 n
rlabel metal5 26020 -5480 26120 -5380 1 PIX337_IN
port 351 n
rlabel metal5 27520 -5480 27620 -5380 1 PIX338_IN
port 352 n
rlabel metal5 29020 -5480 29120 -5380 1 PIX339_IN
port 353 n
rlabel metal5 30520 -5480 30620 -5380 1 PIX340_IN
port 354 n
rlabel metal5 32020 -5480 32120 -5380 1 PIX341_IN
port 355 n
rlabel metal5 33520 -5480 33620 -5380 1 PIX342_IN
port 356 n
rlabel metal5 35020 -5480 35120 -5380 1 PIX343_IN
port 357 n
rlabel metal5 36520 -5480 36620 -5380 1 PIX344_IN
port 358 n
rlabel metal5 38020 -5480 38120 -5380 1 PIX345_IN
port 359 n
rlabel metal5 39520 -5480 39620 -5380 1 PIX346_IN
port 360 n
rlabel metal5 41020 -5480 41120 -5380 1 PIX347_IN
port 361 n
rlabel metal5 42520 -5480 42620 -5380 1 PIX348_IN
port 362 n
rlabel metal5 44020 -5480 44120 -5380 1 PIX349_IN
port 363 n
rlabel metal5 45520 -5480 45620 -5380 1 PIX350_IN
port 364 n
rlabel metal5 47020 -5480 47120 -5380 1 PIX351_IN
port 365 n
rlabel metal5 48520 -5480 48620 -5380 1 PIX352_IN
port 366 n
rlabel metal5 50020 -5480 50120 -5380 1 PIX353_IN
port 367 n
rlabel metal5 51520 -5480 51620 -5380 1 PIX354_IN
port 368 n
rlabel metal5 53020 -5480 53120 -5380 1 PIX355_IN
port 369 n
rlabel metal5 54520 -5480 54620 -5380 1 PIX356_IN
port 370 n
rlabel metal5 56020 -5480 56120 -5380 1 PIX357_IN
port 371 n
rlabel metal5 57520 -5480 57620 -5380 1 PIX358_IN
port 372 n
rlabel metal5 59020 -5480 59120 -5380 1 PIX359_IN
port 373 n
rlabel metal5 60520 -5480 60620 -5380 1 PIX360_IN
port 374 n
rlabel metal5 62020 -5480 62120 -5380 1 PIX361_IN
port 375 n
rlabel metal5 63520 -5480 63620 -5380 1 PIX362_IN
port 376 n
rlabel metal5 65020 -5480 65120 -5380 1 PIX363_IN
port 377 n
rlabel metal5 66520 -5480 66620 -5380 1 PIX364_IN
port 378 n
rlabel metal5 68020 -5480 68120 -5380 1 PIX365_IN
port 379 n
rlabel metal5 69520 -5480 69620 -5380 1 PIX366_IN
port 380 n
rlabel metal5 71020 -5480 71120 -5380 1 PIX367_IN
port 381 n
rlabel metal5 72520 -5480 72620 -5380 1 PIX368_IN
port 382 n
rlabel metal5 74020 -5480 74120 -5380 1 PIX369_IN
port 383 n
rlabel metal5 75520 -5480 75620 -5380 1 PIX370_IN
port 384 n
rlabel metal5 77020 -5480 77120 -5380 1 PIX371_IN
port 385 n
rlabel metal5 78520 -5480 78620 -5380 1 PIX372_IN
port 386 n
rlabel metal5 80020 -5480 80120 -5380 1 PIX373_IN
port 387 n
rlabel metal5 81520 -5480 81620 -5380 1 PIX374_IN
port 388 n
rlabel metal5 83020 -5480 83120 -5380 1 PIX375_IN
port 389 n
rlabel metal5 84520 -5480 84620 -5380 1 PIX376_IN
port 390 n
rlabel metal5 86020 -5480 86120 -5380 1 PIX377_IN
port 391 n
rlabel metal5 87520 -5480 87620 -5380 1 PIX378_IN
port 392 n
rlabel metal5 89020 -5480 89120 -5380 1 PIX379_IN
port 393 n
rlabel metal5 90520 -5480 90620 -5380 1 PIX380_IN
port 394 n
rlabel metal5 92020 -5480 92120 -5380 1 PIX381_IN
port 395 n
rlabel metal5 93520 -5480 93620 -5380 1 PIX382_IN
port 396 n
rlabel metal5 95020 -5480 95120 -5380 1 PIX383_IN
port 397 n
rlabel metal5 96520 -5480 96620 -5380 1 PIX384_IN
port 398 n
rlabel metal5 98020 -5480 98120 -5380 1 PIX385_IN
port 399 n
rlabel metal5 99520 -5480 99620 -5380 1 PIX386_IN
port 400 n
rlabel metal5 101020 -5480 101120 -5380 1 PIX387_IN
port 401 n
rlabel metal5 102520 -5480 102620 -5380 1 PIX388_IN
port 402 n
rlabel metal5 104020 -5480 104120 -5380 1 PIX389_IN
port 403 n
rlabel metal5 105520 -5480 105620 -5380 1 PIX390_IN
port 404 n
rlabel metal5 107020 -5480 107120 -5380 1 PIX391_IN
port 405 n
rlabel metal5 108520 -5480 108620 -5380 1 PIX392_IN
port 406 n
rlabel metal5 110020 -5480 110120 -5380 1 PIX393_IN
port 407 n
rlabel metal5 111520 -5480 111620 -5380 1 PIX394_IN
port 408 n
rlabel metal5 113020 -5480 113120 -5380 1 PIX395_IN
port 409 n
rlabel metal5 114520 -5480 114620 -5380 1 PIX396_IN
port 410 n
rlabel metal5 116020 -5480 116120 -5380 1 PIX397_IN
port 411 n
rlabel metal5 117520 -5480 117620 -5380 1 PIX398_IN
port 412 n
rlabel metal5 119020 -5480 119120 -5380 1 PIX399_IN
port 413 n
rlabel metal5 520 -6980 620 -6880 1 PIX400_IN
port 414 n
rlabel metal2 -1500 -6760 -1500 -6715 3 ROW_SEL5
port 415 e
rlabel metal5 2020 -6980 2120 -6880 1 PIX401_IN
port 416 n
rlabel metal5 3520 -6980 3620 -6880 1 PIX402_IN
port 417 n
rlabel metal5 5020 -6980 5120 -6880 1 PIX403_IN
port 418 n
rlabel metal5 6520 -6980 6620 -6880 1 PIX404_IN
port 419 n
rlabel metal5 8020 -6980 8120 -6880 1 PIX405_IN
port 420 n
rlabel metal5 9520 -6980 9620 -6880 1 PIX406_IN
port 421 n
rlabel metal5 11020 -6980 11120 -6880 1 PIX407_IN
port 422 n
rlabel metal5 12520 -6980 12620 -6880 1 PIX408_IN
port 423 n
rlabel metal5 14020 -6980 14120 -6880 1 PIX409_IN
port 424 n
rlabel metal5 15520 -6980 15620 -6880 1 PIX410_IN
port 425 n
rlabel metal5 17020 -6980 17120 -6880 1 PIX411_IN
port 426 n
rlabel metal5 18520 -6980 18620 -6880 1 PIX412_IN
port 427 n
rlabel metal5 20020 -6980 20120 -6880 1 PIX413_IN
port 428 n
rlabel metal5 21520 -6980 21620 -6880 1 PIX414_IN
port 429 n
rlabel metal5 23020 -6980 23120 -6880 1 PIX415_IN
port 430 n
rlabel metal5 24520 -6980 24620 -6880 1 PIX416_IN
port 431 n
rlabel metal5 26020 -6980 26120 -6880 1 PIX417_IN
port 432 n
rlabel metal5 27520 -6980 27620 -6880 1 PIX418_IN
port 433 n
rlabel metal5 29020 -6980 29120 -6880 1 PIX419_IN
port 434 n
rlabel metal5 30520 -6980 30620 -6880 1 PIX420_IN
port 435 n
rlabel metal5 32020 -6980 32120 -6880 1 PIX421_IN
port 436 n
rlabel metal5 33520 -6980 33620 -6880 1 PIX422_IN
port 437 n
rlabel metal5 35020 -6980 35120 -6880 1 PIX423_IN
port 438 n
rlabel metal5 36520 -6980 36620 -6880 1 PIX424_IN
port 439 n
rlabel metal5 38020 -6980 38120 -6880 1 PIX425_IN
port 440 n
rlabel metal5 39520 -6980 39620 -6880 1 PIX426_IN
port 441 n
rlabel metal5 41020 -6980 41120 -6880 1 PIX427_IN
port 442 n
rlabel metal5 42520 -6980 42620 -6880 1 PIX428_IN
port 443 n
rlabel metal5 44020 -6980 44120 -6880 1 PIX429_IN
port 444 n
rlabel metal5 45520 -6980 45620 -6880 1 PIX430_IN
port 445 n
rlabel metal5 47020 -6980 47120 -6880 1 PIX431_IN
port 446 n
rlabel metal5 48520 -6980 48620 -6880 1 PIX432_IN
port 447 n
rlabel metal5 50020 -6980 50120 -6880 1 PIX433_IN
port 448 n
rlabel metal5 51520 -6980 51620 -6880 1 PIX434_IN
port 449 n
rlabel metal5 53020 -6980 53120 -6880 1 PIX435_IN
port 450 n
rlabel metal5 54520 -6980 54620 -6880 1 PIX436_IN
port 451 n
rlabel metal5 56020 -6980 56120 -6880 1 PIX437_IN
port 452 n
rlabel metal5 57520 -6980 57620 -6880 1 PIX438_IN
port 453 n
rlabel metal5 59020 -6980 59120 -6880 1 PIX439_IN
port 454 n
rlabel metal5 60520 -6980 60620 -6880 1 PIX440_IN
port 455 n
rlabel metal5 62020 -6980 62120 -6880 1 PIX441_IN
port 456 n
rlabel metal5 63520 -6980 63620 -6880 1 PIX442_IN
port 457 n
rlabel metal5 65020 -6980 65120 -6880 1 PIX443_IN
port 458 n
rlabel metal5 66520 -6980 66620 -6880 1 PIX444_IN
port 459 n
rlabel metal5 68020 -6980 68120 -6880 1 PIX445_IN
port 460 n
rlabel metal5 69520 -6980 69620 -6880 1 PIX446_IN
port 461 n
rlabel metal5 71020 -6980 71120 -6880 1 PIX447_IN
port 462 n
rlabel metal5 72520 -6980 72620 -6880 1 PIX448_IN
port 463 n
rlabel metal5 74020 -6980 74120 -6880 1 PIX449_IN
port 464 n
rlabel metal5 75520 -6980 75620 -6880 1 PIX450_IN
port 465 n
rlabel metal5 77020 -6980 77120 -6880 1 PIX451_IN
port 466 n
rlabel metal5 78520 -6980 78620 -6880 1 PIX452_IN
port 467 n
rlabel metal5 80020 -6980 80120 -6880 1 PIX453_IN
port 468 n
rlabel metal5 81520 -6980 81620 -6880 1 PIX454_IN
port 469 n
rlabel metal5 83020 -6980 83120 -6880 1 PIX455_IN
port 470 n
rlabel metal5 84520 -6980 84620 -6880 1 PIX456_IN
port 471 n
rlabel metal5 86020 -6980 86120 -6880 1 PIX457_IN
port 472 n
rlabel metal5 87520 -6980 87620 -6880 1 PIX458_IN
port 473 n
rlabel metal5 89020 -6980 89120 -6880 1 PIX459_IN
port 474 n
rlabel metal5 90520 -6980 90620 -6880 1 PIX460_IN
port 475 n
rlabel metal5 92020 -6980 92120 -6880 1 PIX461_IN
port 476 n
rlabel metal5 93520 -6980 93620 -6880 1 PIX462_IN
port 477 n
rlabel metal5 95020 -6980 95120 -6880 1 PIX463_IN
port 478 n
rlabel metal5 96520 -6980 96620 -6880 1 PIX464_IN
port 479 n
rlabel metal5 98020 -6980 98120 -6880 1 PIX465_IN
port 480 n
rlabel metal5 99520 -6980 99620 -6880 1 PIX466_IN
port 481 n
rlabel metal5 101020 -6980 101120 -6880 1 PIX467_IN
port 482 n
rlabel metal5 102520 -6980 102620 -6880 1 PIX468_IN
port 483 n
rlabel metal5 104020 -6980 104120 -6880 1 PIX469_IN
port 484 n
rlabel metal5 105520 -6980 105620 -6880 1 PIX470_IN
port 485 n
rlabel metal5 107020 -6980 107120 -6880 1 PIX471_IN
port 486 n
rlabel metal5 108520 -6980 108620 -6880 1 PIX472_IN
port 487 n
rlabel metal5 110020 -6980 110120 -6880 1 PIX473_IN
port 488 n
rlabel metal5 111520 -6980 111620 -6880 1 PIX474_IN
port 489 n
rlabel metal5 113020 -6980 113120 -6880 1 PIX475_IN
port 490 n
rlabel metal5 114520 -6980 114620 -6880 1 PIX476_IN
port 491 n
rlabel metal5 116020 -6980 116120 -6880 1 PIX477_IN
port 492 n
rlabel metal5 117520 -6980 117620 -6880 1 PIX478_IN
port 493 n
rlabel metal5 119020 -6980 119120 -6880 1 PIX479_IN
port 494 n
rlabel metal5 520 -8480 620 -8380 1 PIX480_IN
port 495 n
rlabel metal2 -1500 -8260 -1500 -8215 3 ROW_SEL6
port 496 e
rlabel metal5 2020 -8480 2120 -8380 1 PIX481_IN
port 497 n
rlabel metal5 3520 -8480 3620 -8380 1 PIX482_IN
port 498 n
rlabel metal5 5020 -8480 5120 -8380 1 PIX483_IN
port 499 n
rlabel metal5 6520 -8480 6620 -8380 1 PIX484_IN
port 500 n
rlabel metal5 8020 -8480 8120 -8380 1 PIX485_IN
port 501 n
rlabel metal5 9520 -8480 9620 -8380 1 PIX486_IN
port 502 n
rlabel metal5 11020 -8480 11120 -8380 1 PIX487_IN
port 503 n
rlabel metal5 12520 -8480 12620 -8380 1 PIX488_IN
port 504 n
rlabel metal5 14020 -8480 14120 -8380 1 PIX489_IN
port 505 n
rlabel metal5 15520 -8480 15620 -8380 1 PIX490_IN
port 506 n
rlabel metal5 17020 -8480 17120 -8380 1 PIX491_IN
port 507 n
rlabel metal5 18520 -8480 18620 -8380 1 PIX492_IN
port 508 n
rlabel metal5 20020 -8480 20120 -8380 1 PIX493_IN
port 509 n
rlabel metal5 21520 -8480 21620 -8380 1 PIX494_IN
port 510 n
rlabel metal5 23020 -8480 23120 -8380 1 PIX495_IN
port 511 n
rlabel metal5 24520 -8480 24620 -8380 1 PIX496_IN
port 512 n
rlabel metal5 26020 -8480 26120 -8380 1 PIX497_IN
port 513 n
rlabel metal5 27520 -8480 27620 -8380 1 PIX498_IN
port 514 n
rlabel metal5 29020 -8480 29120 -8380 1 PIX499_IN
port 515 n
rlabel metal5 30520 -8480 30620 -8380 1 PIX500_IN
port 516 n
rlabel metal5 32020 -8480 32120 -8380 1 PIX501_IN
port 517 n
rlabel metal5 33520 -8480 33620 -8380 1 PIX502_IN
port 518 n
rlabel metal5 35020 -8480 35120 -8380 1 PIX503_IN
port 519 n
rlabel metal5 36520 -8480 36620 -8380 1 PIX504_IN
port 520 n
rlabel metal5 38020 -8480 38120 -8380 1 PIX505_IN
port 521 n
rlabel metal5 39520 -8480 39620 -8380 1 PIX506_IN
port 522 n
rlabel metal5 41020 -8480 41120 -8380 1 PIX507_IN
port 523 n
rlabel metal5 42520 -8480 42620 -8380 1 PIX508_IN
port 524 n
rlabel metal5 44020 -8480 44120 -8380 1 PIX509_IN
port 525 n
rlabel metal5 45520 -8480 45620 -8380 1 PIX510_IN
port 526 n
rlabel metal5 47020 -8480 47120 -8380 1 PIX511_IN
port 527 n
rlabel metal5 48520 -8480 48620 -8380 1 PIX512_IN
port 528 n
rlabel metal5 50020 -8480 50120 -8380 1 PIX513_IN
port 529 n
rlabel metal5 51520 -8480 51620 -8380 1 PIX514_IN
port 530 n
rlabel metal5 53020 -8480 53120 -8380 1 PIX515_IN
port 531 n
rlabel metal5 54520 -8480 54620 -8380 1 PIX516_IN
port 532 n
rlabel metal5 56020 -8480 56120 -8380 1 PIX517_IN
port 533 n
rlabel metal5 57520 -8480 57620 -8380 1 PIX518_IN
port 534 n
rlabel metal5 59020 -8480 59120 -8380 1 PIX519_IN
port 535 n
rlabel metal5 60520 -8480 60620 -8380 1 PIX520_IN
port 536 n
rlabel metal5 62020 -8480 62120 -8380 1 PIX521_IN
port 537 n
rlabel metal5 63520 -8480 63620 -8380 1 PIX522_IN
port 538 n
rlabel metal5 65020 -8480 65120 -8380 1 PIX523_IN
port 539 n
rlabel metal5 66520 -8480 66620 -8380 1 PIX524_IN
port 540 n
rlabel metal5 68020 -8480 68120 -8380 1 PIX525_IN
port 541 n
rlabel metal5 69520 -8480 69620 -8380 1 PIX526_IN
port 542 n
rlabel metal5 71020 -8480 71120 -8380 1 PIX527_IN
port 543 n
rlabel metal5 72520 -8480 72620 -8380 1 PIX528_IN
port 544 n
rlabel metal5 74020 -8480 74120 -8380 1 PIX529_IN
port 545 n
rlabel metal5 75520 -8480 75620 -8380 1 PIX530_IN
port 546 n
rlabel metal5 77020 -8480 77120 -8380 1 PIX531_IN
port 547 n
rlabel metal5 78520 -8480 78620 -8380 1 PIX532_IN
port 548 n
rlabel metal5 80020 -8480 80120 -8380 1 PIX533_IN
port 549 n
rlabel metal5 81520 -8480 81620 -8380 1 PIX534_IN
port 550 n
rlabel metal5 83020 -8480 83120 -8380 1 PIX535_IN
port 551 n
rlabel metal5 84520 -8480 84620 -8380 1 PIX536_IN
port 552 n
rlabel metal5 86020 -8480 86120 -8380 1 PIX537_IN
port 553 n
rlabel metal5 87520 -8480 87620 -8380 1 PIX538_IN
port 554 n
rlabel metal5 89020 -8480 89120 -8380 1 PIX539_IN
port 555 n
rlabel metal5 90520 -8480 90620 -8380 1 PIX540_IN
port 556 n
rlabel metal5 92020 -8480 92120 -8380 1 PIX541_IN
port 557 n
rlabel metal5 93520 -8480 93620 -8380 1 PIX542_IN
port 558 n
rlabel metal5 95020 -8480 95120 -8380 1 PIX543_IN
port 559 n
rlabel metal5 96520 -8480 96620 -8380 1 PIX544_IN
port 560 n
rlabel metal5 98020 -8480 98120 -8380 1 PIX545_IN
port 561 n
rlabel metal5 99520 -8480 99620 -8380 1 PIX546_IN
port 562 n
rlabel metal5 101020 -8480 101120 -8380 1 PIX547_IN
port 563 n
rlabel metal5 102520 -8480 102620 -8380 1 PIX548_IN
port 564 n
rlabel metal5 104020 -8480 104120 -8380 1 PIX549_IN
port 565 n
rlabel metal5 105520 -8480 105620 -8380 1 PIX550_IN
port 566 n
rlabel metal5 107020 -8480 107120 -8380 1 PIX551_IN
port 567 n
rlabel metal5 108520 -8480 108620 -8380 1 PIX552_IN
port 568 n
rlabel metal5 110020 -8480 110120 -8380 1 PIX553_IN
port 569 n
rlabel metal5 111520 -8480 111620 -8380 1 PIX554_IN
port 570 n
rlabel metal5 113020 -8480 113120 -8380 1 PIX555_IN
port 571 n
rlabel metal5 114520 -8480 114620 -8380 1 PIX556_IN
port 572 n
rlabel metal5 116020 -8480 116120 -8380 1 PIX557_IN
port 573 n
rlabel metal5 117520 -8480 117620 -8380 1 PIX558_IN
port 574 n
rlabel metal5 119020 -8480 119120 -8380 1 PIX559_IN
port 575 n
rlabel metal5 520 -9980 620 -9880 1 PIX560_IN
port 576 n
rlabel metal2 -1500 -9760 -1500 -9715 3 ROW_SEL7
port 577 e
rlabel metal5 2020 -9980 2120 -9880 1 PIX561_IN
port 578 n
rlabel metal5 3520 -9980 3620 -9880 1 PIX562_IN
port 579 n
rlabel metal5 5020 -9980 5120 -9880 1 PIX563_IN
port 580 n
rlabel metal5 6520 -9980 6620 -9880 1 PIX564_IN
port 581 n
rlabel metal5 8020 -9980 8120 -9880 1 PIX565_IN
port 582 n
rlabel metal5 9520 -9980 9620 -9880 1 PIX566_IN
port 583 n
rlabel metal5 11020 -9980 11120 -9880 1 PIX567_IN
port 584 n
rlabel metal5 12520 -9980 12620 -9880 1 PIX568_IN
port 585 n
rlabel metal5 14020 -9980 14120 -9880 1 PIX569_IN
port 586 n
rlabel metal5 15520 -9980 15620 -9880 1 PIX570_IN
port 587 n
rlabel metal5 17020 -9980 17120 -9880 1 PIX571_IN
port 588 n
rlabel metal5 18520 -9980 18620 -9880 1 PIX572_IN
port 589 n
rlabel metal5 20020 -9980 20120 -9880 1 PIX573_IN
port 590 n
rlabel metal5 21520 -9980 21620 -9880 1 PIX574_IN
port 591 n
rlabel metal5 23020 -9980 23120 -9880 1 PIX575_IN
port 592 n
rlabel metal5 24520 -9980 24620 -9880 1 PIX576_IN
port 593 n
rlabel metal5 26020 -9980 26120 -9880 1 PIX577_IN
port 594 n
rlabel metal5 27520 -9980 27620 -9880 1 PIX578_IN
port 595 n
rlabel metal5 29020 -9980 29120 -9880 1 PIX579_IN
port 596 n
rlabel metal5 30520 -9980 30620 -9880 1 PIX580_IN
port 597 n
rlabel metal5 32020 -9980 32120 -9880 1 PIX581_IN
port 598 n
rlabel metal5 33520 -9980 33620 -9880 1 PIX582_IN
port 599 n
rlabel metal5 35020 -9980 35120 -9880 1 PIX583_IN
port 600 n
rlabel metal5 36520 -9980 36620 -9880 1 PIX584_IN
port 601 n
rlabel metal5 38020 -9980 38120 -9880 1 PIX585_IN
port 602 n
rlabel metal5 39520 -9980 39620 -9880 1 PIX586_IN
port 603 n
rlabel metal5 41020 -9980 41120 -9880 1 PIX587_IN
port 604 n
rlabel metal5 42520 -9980 42620 -9880 1 PIX588_IN
port 605 n
rlabel metal5 44020 -9980 44120 -9880 1 PIX589_IN
port 606 n
rlabel metal5 45520 -9980 45620 -9880 1 PIX590_IN
port 607 n
rlabel metal5 47020 -9980 47120 -9880 1 PIX591_IN
port 608 n
rlabel metal5 48520 -9980 48620 -9880 1 PIX592_IN
port 609 n
rlabel metal5 50020 -9980 50120 -9880 1 PIX593_IN
port 610 n
rlabel metal5 51520 -9980 51620 -9880 1 PIX594_IN
port 611 n
rlabel metal5 53020 -9980 53120 -9880 1 PIX595_IN
port 612 n
rlabel metal5 54520 -9980 54620 -9880 1 PIX596_IN
port 613 n
rlabel metal5 56020 -9980 56120 -9880 1 PIX597_IN
port 614 n
rlabel metal5 57520 -9980 57620 -9880 1 PIX598_IN
port 615 n
rlabel metal5 59020 -9980 59120 -9880 1 PIX599_IN
port 616 n
rlabel metal5 60520 -9980 60620 -9880 1 PIX600_IN
port 617 n
rlabel metal5 62020 -9980 62120 -9880 1 PIX601_IN
port 618 n
rlabel metal5 63520 -9980 63620 -9880 1 PIX602_IN
port 619 n
rlabel metal5 65020 -9980 65120 -9880 1 PIX603_IN
port 620 n
rlabel metal5 66520 -9980 66620 -9880 1 PIX604_IN
port 621 n
rlabel metal5 68020 -9980 68120 -9880 1 PIX605_IN
port 622 n
rlabel metal5 69520 -9980 69620 -9880 1 PIX606_IN
port 623 n
rlabel metal5 71020 -9980 71120 -9880 1 PIX607_IN
port 624 n
rlabel metal5 72520 -9980 72620 -9880 1 PIX608_IN
port 625 n
rlabel metal5 74020 -9980 74120 -9880 1 PIX609_IN
port 626 n
rlabel metal5 75520 -9980 75620 -9880 1 PIX610_IN
port 627 n
rlabel metal5 77020 -9980 77120 -9880 1 PIX611_IN
port 628 n
rlabel metal5 78520 -9980 78620 -9880 1 PIX612_IN
port 629 n
rlabel metal5 80020 -9980 80120 -9880 1 PIX613_IN
port 630 n
rlabel metal5 81520 -9980 81620 -9880 1 PIX614_IN
port 631 n
rlabel metal5 83020 -9980 83120 -9880 1 PIX615_IN
port 632 n
rlabel metal5 84520 -9980 84620 -9880 1 PIX616_IN
port 633 n
rlabel metal5 86020 -9980 86120 -9880 1 PIX617_IN
port 634 n
rlabel metal5 87520 -9980 87620 -9880 1 PIX618_IN
port 635 n
rlabel metal5 89020 -9980 89120 -9880 1 PIX619_IN
port 636 n
rlabel metal5 90520 -9980 90620 -9880 1 PIX620_IN
port 637 n
rlabel metal5 92020 -9980 92120 -9880 1 PIX621_IN
port 638 n
rlabel metal5 93520 -9980 93620 -9880 1 PIX622_IN
port 639 n
rlabel metal5 95020 -9980 95120 -9880 1 PIX623_IN
port 640 n
rlabel metal5 96520 -9980 96620 -9880 1 PIX624_IN
port 641 n
rlabel metal5 98020 -9980 98120 -9880 1 PIX625_IN
port 642 n
rlabel metal5 99520 -9980 99620 -9880 1 PIX626_IN
port 643 n
rlabel metal5 101020 -9980 101120 -9880 1 PIX627_IN
port 644 n
rlabel metal5 102520 -9980 102620 -9880 1 PIX628_IN
port 645 n
rlabel metal5 104020 -9980 104120 -9880 1 PIX629_IN
port 646 n
rlabel metal5 105520 -9980 105620 -9880 1 PIX630_IN
port 647 n
rlabel metal5 107020 -9980 107120 -9880 1 PIX631_IN
port 648 n
rlabel metal5 108520 -9980 108620 -9880 1 PIX632_IN
port 649 n
rlabel metal5 110020 -9980 110120 -9880 1 PIX633_IN
port 650 n
rlabel metal5 111520 -9980 111620 -9880 1 PIX634_IN
port 651 n
rlabel metal5 113020 -9980 113120 -9880 1 PIX635_IN
port 652 n
rlabel metal5 114520 -9980 114620 -9880 1 PIX636_IN
port 653 n
rlabel metal5 116020 -9980 116120 -9880 1 PIX637_IN
port 654 n
rlabel metal5 117520 -9980 117620 -9880 1 PIX638_IN
port 655 n
rlabel metal5 119020 -9980 119120 -9880 1 PIX639_IN
port 656 n
rlabel metal5 520 -11480 620 -11380 1 PIX640_IN
port 657 n
rlabel metal2 -1500 -11260 -1500 -11215 3 ROW_SEL8
port 658 e
rlabel metal5 2020 -11480 2120 -11380 1 PIX641_IN
port 659 n
rlabel metal5 3520 -11480 3620 -11380 1 PIX642_IN
port 660 n
rlabel metal5 5020 -11480 5120 -11380 1 PIX643_IN
port 661 n
rlabel metal5 6520 -11480 6620 -11380 1 PIX644_IN
port 662 n
rlabel metal5 8020 -11480 8120 -11380 1 PIX645_IN
port 663 n
rlabel metal5 9520 -11480 9620 -11380 1 PIX646_IN
port 664 n
rlabel metal5 11020 -11480 11120 -11380 1 PIX647_IN
port 665 n
rlabel metal5 12520 -11480 12620 -11380 1 PIX648_IN
port 666 n
rlabel metal5 14020 -11480 14120 -11380 1 PIX649_IN
port 667 n
rlabel metal5 15520 -11480 15620 -11380 1 PIX650_IN
port 668 n
rlabel metal5 17020 -11480 17120 -11380 1 PIX651_IN
port 669 n
rlabel metal5 18520 -11480 18620 -11380 1 PIX652_IN
port 670 n
rlabel metal5 20020 -11480 20120 -11380 1 PIX653_IN
port 671 n
rlabel metal5 21520 -11480 21620 -11380 1 PIX654_IN
port 672 n
rlabel metal5 23020 -11480 23120 -11380 1 PIX655_IN
port 673 n
rlabel metal5 24520 -11480 24620 -11380 1 PIX656_IN
port 674 n
rlabel metal5 26020 -11480 26120 -11380 1 PIX657_IN
port 675 n
rlabel metal5 27520 -11480 27620 -11380 1 PIX658_IN
port 676 n
rlabel metal5 29020 -11480 29120 -11380 1 PIX659_IN
port 677 n
rlabel metal5 30520 -11480 30620 -11380 1 PIX660_IN
port 678 n
rlabel metal5 32020 -11480 32120 -11380 1 PIX661_IN
port 679 n
rlabel metal5 33520 -11480 33620 -11380 1 PIX662_IN
port 680 n
rlabel metal5 35020 -11480 35120 -11380 1 PIX663_IN
port 681 n
rlabel metal5 36520 -11480 36620 -11380 1 PIX664_IN
port 682 n
rlabel metal5 38020 -11480 38120 -11380 1 PIX665_IN
port 683 n
rlabel metal5 39520 -11480 39620 -11380 1 PIX666_IN
port 684 n
rlabel metal5 41020 -11480 41120 -11380 1 PIX667_IN
port 685 n
rlabel metal5 42520 -11480 42620 -11380 1 PIX668_IN
port 686 n
rlabel metal5 44020 -11480 44120 -11380 1 PIX669_IN
port 687 n
rlabel metal5 45520 -11480 45620 -11380 1 PIX670_IN
port 688 n
rlabel metal5 47020 -11480 47120 -11380 1 PIX671_IN
port 689 n
rlabel metal5 48520 -11480 48620 -11380 1 PIX672_IN
port 690 n
rlabel metal5 50020 -11480 50120 -11380 1 PIX673_IN
port 691 n
rlabel metal5 51520 -11480 51620 -11380 1 PIX674_IN
port 692 n
rlabel metal5 53020 -11480 53120 -11380 1 PIX675_IN
port 693 n
rlabel metal5 54520 -11480 54620 -11380 1 PIX676_IN
port 694 n
rlabel metal5 56020 -11480 56120 -11380 1 PIX677_IN
port 695 n
rlabel metal5 57520 -11480 57620 -11380 1 PIX678_IN
port 696 n
rlabel metal5 59020 -11480 59120 -11380 1 PIX679_IN
port 697 n
rlabel metal5 60520 -11480 60620 -11380 1 PIX680_IN
port 698 n
rlabel metal5 62020 -11480 62120 -11380 1 PIX681_IN
port 699 n
rlabel metal5 63520 -11480 63620 -11380 1 PIX682_IN
port 700 n
rlabel metal5 65020 -11480 65120 -11380 1 PIX683_IN
port 701 n
rlabel metal5 66520 -11480 66620 -11380 1 PIX684_IN
port 702 n
rlabel metal5 68020 -11480 68120 -11380 1 PIX685_IN
port 703 n
rlabel metal5 69520 -11480 69620 -11380 1 PIX686_IN
port 704 n
rlabel metal5 71020 -11480 71120 -11380 1 PIX687_IN
port 705 n
rlabel metal5 72520 -11480 72620 -11380 1 PIX688_IN
port 706 n
rlabel metal5 74020 -11480 74120 -11380 1 PIX689_IN
port 707 n
rlabel metal5 75520 -11480 75620 -11380 1 PIX690_IN
port 708 n
rlabel metal5 77020 -11480 77120 -11380 1 PIX691_IN
port 709 n
rlabel metal5 78520 -11480 78620 -11380 1 PIX692_IN
port 710 n
rlabel metal5 80020 -11480 80120 -11380 1 PIX693_IN
port 711 n
rlabel metal5 81520 -11480 81620 -11380 1 PIX694_IN
port 712 n
rlabel metal5 83020 -11480 83120 -11380 1 PIX695_IN
port 713 n
rlabel metal5 84520 -11480 84620 -11380 1 PIX696_IN
port 714 n
rlabel metal5 86020 -11480 86120 -11380 1 PIX697_IN
port 715 n
rlabel metal5 87520 -11480 87620 -11380 1 PIX698_IN
port 716 n
rlabel metal5 89020 -11480 89120 -11380 1 PIX699_IN
port 717 n
rlabel metal5 90520 -11480 90620 -11380 1 PIX700_IN
port 718 n
rlabel metal5 92020 -11480 92120 -11380 1 PIX701_IN
port 719 n
rlabel metal5 93520 -11480 93620 -11380 1 PIX702_IN
port 720 n
rlabel metal5 95020 -11480 95120 -11380 1 PIX703_IN
port 721 n
rlabel metal5 96520 -11480 96620 -11380 1 PIX704_IN
port 722 n
rlabel metal5 98020 -11480 98120 -11380 1 PIX705_IN
port 723 n
rlabel metal5 99520 -11480 99620 -11380 1 PIX706_IN
port 724 n
rlabel metal5 101020 -11480 101120 -11380 1 PIX707_IN
port 725 n
rlabel metal5 102520 -11480 102620 -11380 1 PIX708_IN
port 726 n
rlabel metal5 104020 -11480 104120 -11380 1 PIX709_IN
port 727 n
rlabel metal5 105520 -11480 105620 -11380 1 PIX710_IN
port 728 n
rlabel metal5 107020 -11480 107120 -11380 1 PIX711_IN
port 729 n
rlabel metal5 108520 -11480 108620 -11380 1 PIX712_IN
port 730 n
rlabel metal5 110020 -11480 110120 -11380 1 PIX713_IN
port 731 n
rlabel metal5 111520 -11480 111620 -11380 1 PIX714_IN
port 732 n
rlabel metal5 113020 -11480 113120 -11380 1 PIX715_IN
port 733 n
rlabel metal5 114520 -11480 114620 -11380 1 PIX716_IN
port 734 n
rlabel metal5 116020 -11480 116120 -11380 1 PIX717_IN
port 735 n
rlabel metal5 117520 -11480 117620 -11380 1 PIX718_IN
port 736 n
rlabel metal5 119020 -11480 119120 -11380 1 PIX719_IN
port 737 n
rlabel metal5 520 -12980 620 -12880 1 PIX720_IN
port 738 n
rlabel metal2 -1500 -12760 -1500 -12715 3 ROW_SEL9
port 739 e
rlabel metal5 2020 -12980 2120 -12880 1 PIX721_IN
port 740 n
rlabel metal5 3520 -12980 3620 -12880 1 PIX722_IN
port 741 n
rlabel metal5 5020 -12980 5120 -12880 1 PIX723_IN
port 742 n
rlabel metal5 6520 -12980 6620 -12880 1 PIX724_IN
port 743 n
rlabel metal5 8020 -12980 8120 -12880 1 PIX725_IN
port 744 n
rlabel metal5 9520 -12980 9620 -12880 1 PIX726_IN
port 745 n
rlabel metal5 11020 -12980 11120 -12880 1 PIX727_IN
port 746 n
rlabel metal5 12520 -12980 12620 -12880 1 PIX728_IN
port 747 n
rlabel metal5 14020 -12980 14120 -12880 1 PIX729_IN
port 748 n
rlabel metal5 15520 -12980 15620 -12880 1 PIX730_IN
port 749 n
rlabel metal5 17020 -12980 17120 -12880 1 PIX731_IN
port 750 n
rlabel metal5 18520 -12980 18620 -12880 1 PIX732_IN
port 751 n
rlabel metal5 20020 -12980 20120 -12880 1 PIX733_IN
port 752 n
rlabel metal5 21520 -12980 21620 -12880 1 PIX734_IN
port 753 n
rlabel metal5 23020 -12980 23120 -12880 1 PIX735_IN
port 754 n
rlabel metal5 24520 -12980 24620 -12880 1 PIX736_IN
port 755 n
rlabel metal5 26020 -12980 26120 -12880 1 PIX737_IN
port 756 n
rlabel metal5 27520 -12980 27620 -12880 1 PIX738_IN
port 757 n
rlabel metal5 29020 -12980 29120 -12880 1 PIX739_IN
port 758 n
rlabel metal5 30520 -12980 30620 -12880 1 PIX740_IN
port 759 n
rlabel metal5 32020 -12980 32120 -12880 1 PIX741_IN
port 760 n
rlabel metal5 33520 -12980 33620 -12880 1 PIX742_IN
port 761 n
rlabel metal5 35020 -12980 35120 -12880 1 PIX743_IN
port 762 n
rlabel metal5 36520 -12980 36620 -12880 1 PIX744_IN
port 763 n
rlabel metal5 38020 -12980 38120 -12880 1 PIX745_IN
port 764 n
rlabel metal5 39520 -12980 39620 -12880 1 PIX746_IN
port 765 n
rlabel metal5 41020 -12980 41120 -12880 1 PIX747_IN
port 766 n
rlabel metal5 42520 -12980 42620 -12880 1 PIX748_IN
port 767 n
rlabel metal5 44020 -12980 44120 -12880 1 PIX749_IN
port 768 n
rlabel metal5 45520 -12980 45620 -12880 1 PIX750_IN
port 769 n
rlabel metal5 47020 -12980 47120 -12880 1 PIX751_IN
port 770 n
rlabel metal5 48520 -12980 48620 -12880 1 PIX752_IN
port 771 n
rlabel metal5 50020 -12980 50120 -12880 1 PIX753_IN
port 772 n
rlabel metal5 51520 -12980 51620 -12880 1 PIX754_IN
port 773 n
rlabel metal5 53020 -12980 53120 -12880 1 PIX755_IN
port 774 n
rlabel metal5 54520 -12980 54620 -12880 1 PIX756_IN
port 775 n
rlabel metal5 56020 -12980 56120 -12880 1 PIX757_IN
port 776 n
rlabel metal5 57520 -12980 57620 -12880 1 PIX758_IN
port 777 n
rlabel metal5 59020 -12980 59120 -12880 1 PIX759_IN
port 778 n
rlabel metal5 60520 -12980 60620 -12880 1 PIX760_IN
port 779 n
rlabel metal5 62020 -12980 62120 -12880 1 PIX761_IN
port 780 n
rlabel metal5 63520 -12980 63620 -12880 1 PIX762_IN
port 781 n
rlabel metal5 65020 -12980 65120 -12880 1 PIX763_IN
port 782 n
rlabel metal5 66520 -12980 66620 -12880 1 PIX764_IN
port 783 n
rlabel metal5 68020 -12980 68120 -12880 1 PIX765_IN
port 784 n
rlabel metal5 69520 -12980 69620 -12880 1 PIX766_IN
port 785 n
rlabel metal5 71020 -12980 71120 -12880 1 PIX767_IN
port 786 n
rlabel metal5 72520 -12980 72620 -12880 1 PIX768_IN
port 787 n
rlabel metal5 74020 -12980 74120 -12880 1 PIX769_IN
port 788 n
rlabel metal5 75520 -12980 75620 -12880 1 PIX770_IN
port 789 n
rlabel metal5 77020 -12980 77120 -12880 1 PIX771_IN
port 790 n
rlabel metal5 78520 -12980 78620 -12880 1 PIX772_IN
port 791 n
rlabel metal5 80020 -12980 80120 -12880 1 PIX773_IN
port 792 n
rlabel metal5 81520 -12980 81620 -12880 1 PIX774_IN
port 793 n
rlabel metal5 83020 -12980 83120 -12880 1 PIX775_IN
port 794 n
rlabel metal5 84520 -12980 84620 -12880 1 PIX776_IN
port 795 n
rlabel metal5 86020 -12980 86120 -12880 1 PIX777_IN
port 796 n
rlabel metal5 87520 -12980 87620 -12880 1 PIX778_IN
port 797 n
rlabel metal5 89020 -12980 89120 -12880 1 PIX779_IN
port 798 n
rlabel metal5 90520 -12980 90620 -12880 1 PIX780_IN
port 799 n
rlabel metal5 92020 -12980 92120 -12880 1 PIX781_IN
port 800 n
rlabel metal5 93520 -12980 93620 -12880 1 PIX782_IN
port 801 n
rlabel metal5 95020 -12980 95120 -12880 1 PIX783_IN
port 802 n
rlabel metal5 96520 -12980 96620 -12880 1 PIX784_IN
port 803 n
rlabel metal5 98020 -12980 98120 -12880 1 PIX785_IN
port 804 n
rlabel metal5 99520 -12980 99620 -12880 1 PIX786_IN
port 805 n
rlabel metal5 101020 -12980 101120 -12880 1 PIX787_IN
port 806 n
rlabel metal5 102520 -12980 102620 -12880 1 PIX788_IN
port 807 n
rlabel metal5 104020 -12980 104120 -12880 1 PIX789_IN
port 808 n
rlabel metal5 105520 -12980 105620 -12880 1 PIX790_IN
port 809 n
rlabel metal5 107020 -12980 107120 -12880 1 PIX791_IN
port 810 n
rlabel metal5 108520 -12980 108620 -12880 1 PIX792_IN
port 811 n
rlabel metal5 110020 -12980 110120 -12880 1 PIX793_IN
port 812 n
rlabel metal5 111520 -12980 111620 -12880 1 PIX794_IN
port 813 n
rlabel metal5 113020 -12980 113120 -12880 1 PIX795_IN
port 814 n
rlabel metal5 114520 -12980 114620 -12880 1 PIX796_IN
port 815 n
rlabel metal5 116020 -12980 116120 -12880 1 PIX797_IN
port 816 n
rlabel metal5 117520 -12980 117620 -12880 1 PIX798_IN
port 817 n
rlabel metal5 119020 -12980 119120 -12880 1 PIX799_IN
port 818 n
rlabel metal5 520 -14480 620 -14380 1 PIX800_IN
port 819 n
rlabel metal2 -1500 -14260 -1500 -14215 3 ROW_SEL10
port 820 e
rlabel metal5 2020 -14480 2120 -14380 1 PIX801_IN
port 821 n
rlabel metal5 3520 -14480 3620 -14380 1 PIX802_IN
port 822 n
rlabel metal5 5020 -14480 5120 -14380 1 PIX803_IN
port 823 n
rlabel metal5 6520 -14480 6620 -14380 1 PIX804_IN
port 824 n
rlabel metal5 8020 -14480 8120 -14380 1 PIX805_IN
port 825 n
rlabel metal5 9520 -14480 9620 -14380 1 PIX806_IN
port 826 n
rlabel metal5 11020 -14480 11120 -14380 1 PIX807_IN
port 827 n
rlabel metal5 12520 -14480 12620 -14380 1 PIX808_IN
port 828 n
rlabel metal5 14020 -14480 14120 -14380 1 PIX809_IN
port 829 n
rlabel metal5 15520 -14480 15620 -14380 1 PIX810_IN
port 830 n
rlabel metal5 17020 -14480 17120 -14380 1 PIX811_IN
port 831 n
rlabel metal5 18520 -14480 18620 -14380 1 PIX812_IN
port 832 n
rlabel metal5 20020 -14480 20120 -14380 1 PIX813_IN
port 833 n
rlabel metal5 21520 -14480 21620 -14380 1 PIX814_IN
port 834 n
rlabel metal5 23020 -14480 23120 -14380 1 PIX815_IN
port 835 n
rlabel metal5 24520 -14480 24620 -14380 1 PIX816_IN
port 836 n
rlabel metal5 26020 -14480 26120 -14380 1 PIX817_IN
port 837 n
rlabel metal5 27520 -14480 27620 -14380 1 PIX818_IN
port 838 n
rlabel metal5 29020 -14480 29120 -14380 1 PIX819_IN
port 839 n
rlabel metal5 30520 -14480 30620 -14380 1 PIX820_IN
port 840 n
rlabel metal5 32020 -14480 32120 -14380 1 PIX821_IN
port 841 n
rlabel metal5 33520 -14480 33620 -14380 1 PIX822_IN
port 842 n
rlabel metal5 35020 -14480 35120 -14380 1 PIX823_IN
port 843 n
rlabel metal5 36520 -14480 36620 -14380 1 PIX824_IN
port 844 n
rlabel metal5 38020 -14480 38120 -14380 1 PIX825_IN
port 845 n
rlabel metal5 39520 -14480 39620 -14380 1 PIX826_IN
port 846 n
rlabel metal5 41020 -14480 41120 -14380 1 PIX827_IN
port 847 n
rlabel metal5 42520 -14480 42620 -14380 1 PIX828_IN
port 848 n
rlabel metal5 44020 -14480 44120 -14380 1 PIX829_IN
port 849 n
rlabel metal5 45520 -14480 45620 -14380 1 PIX830_IN
port 850 n
rlabel metal5 47020 -14480 47120 -14380 1 PIX831_IN
port 851 n
rlabel metal5 48520 -14480 48620 -14380 1 PIX832_IN
port 852 n
rlabel metal5 50020 -14480 50120 -14380 1 PIX833_IN
port 853 n
rlabel metal5 51520 -14480 51620 -14380 1 PIX834_IN
port 854 n
rlabel metal5 53020 -14480 53120 -14380 1 PIX835_IN
port 855 n
rlabel metal5 54520 -14480 54620 -14380 1 PIX836_IN
port 856 n
rlabel metal5 56020 -14480 56120 -14380 1 PIX837_IN
port 857 n
rlabel metal5 57520 -14480 57620 -14380 1 PIX838_IN
port 858 n
rlabel metal5 59020 -14480 59120 -14380 1 PIX839_IN
port 859 n
rlabel metal5 60520 -14480 60620 -14380 1 PIX840_IN
port 860 n
rlabel metal5 62020 -14480 62120 -14380 1 PIX841_IN
port 861 n
rlabel metal5 63520 -14480 63620 -14380 1 PIX842_IN
port 862 n
rlabel metal5 65020 -14480 65120 -14380 1 PIX843_IN
port 863 n
rlabel metal5 66520 -14480 66620 -14380 1 PIX844_IN
port 864 n
rlabel metal5 68020 -14480 68120 -14380 1 PIX845_IN
port 865 n
rlabel metal5 69520 -14480 69620 -14380 1 PIX846_IN
port 866 n
rlabel metal5 71020 -14480 71120 -14380 1 PIX847_IN
port 867 n
rlabel metal5 72520 -14480 72620 -14380 1 PIX848_IN
port 868 n
rlabel metal5 74020 -14480 74120 -14380 1 PIX849_IN
port 869 n
rlabel metal5 75520 -14480 75620 -14380 1 PIX850_IN
port 870 n
rlabel metal5 77020 -14480 77120 -14380 1 PIX851_IN
port 871 n
rlabel metal5 78520 -14480 78620 -14380 1 PIX852_IN
port 872 n
rlabel metal5 80020 -14480 80120 -14380 1 PIX853_IN
port 873 n
rlabel metal5 81520 -14480 81620 -14380 1 PIX854_IN
port 874 n
rlabel metal5 83020 -14480 83120 -14380 1 PIX855_IN
port 875 n
rlabel metal5 84520 -14480 84620 -14380 1 PIX856_IN
port 876 n
rlabel metal5 86020 -14480 86120 -14380 1 PIX857_IN
port 877 n
rlabel metal5 87520 -14480 87620 -14380 1 PIX858_IN
port 878 n
rlabel metal5 89020 -14480 89120 -14380 1 PIX859_IN
port 879 n
rlabel metal5 90520 -14480 90620 -14380 1 PIX860_IN
port 880 n
rlabel metal5 92020 -14480 92120 -14380 1 PIX861_IN
port 881 n
rlabel metal5 93520 -14480 93620 -14380 1 PIX862_IN
port 882 n
rlabel metal5 95020 -14480 95120 -14380 1 PIX863_IN
port 883 n
rlabel metal5 96520 -14480 96620 -14380 1 PIX864_IN
port 884 n
rlabel metal5 98020 -14480 98120 -14380 1 PIX865_IN
port 885 n
rlabel metal5 99520 -14480 99620 -14380 1 PIX866_IN
port 886 n
rlabel metal5 101020 -14480 101120 -14380 1 PIX867_IN
port 887 n
rlabel metal5 102520 -14480 102620 -14380 1 PIX868_IN
port 888 n
rlabel metal5 104020 -14480 104120 -14380 1 PIX869_IN
port 889 n
rlabel metal5 105520 -14480 105620 -14380 1 PIX870_IN
port 890 n
rlabel metal5 107020 -14480 107120 -14380 1 PIX871_IN
port 891 n
rlabel metal5 108520 -14480 108620 -14380 1 PIX872_IN
port 892 n
rlabel metal5 110020 -14480 110120 -14380 1 PIX873_IN
port 893 n
rlabel metal5 111520 -14480 111620 -14380 1 PIX874_IN
port 894 n
rlabel metal5 113020 -14480 113120 -14380 1 PIX875_IN
port 895 n
rlabel metal5 114520 -14480 114620 -14380 1 PIX876_IN
port 896 n
rlabel metal5 116020 -14480 116120 -14380 1 PIX877_IN
port 897 n
rlabel metal5 117520 -14480 117620 -14380 1 PIX878_IN
port 898 n
rlabel metal5 119020 -14480 119120 -14380 1 PIX879_IN
port 899 n
rlabel metal5 520 -15980 620 -15880 1 PIX880_IN
port 900 n
rlabel metal2 -1500 -15760 -1500 -15715 3 ROW_SEL11
port 901 e
rlabel metal5 2020 -15980 2120 -15880 1 PIX881_IN
port 902 n
rlabel metal5 3520 -15980 3620 -15880 1 PIX882_IN
port 903 n
rlabel metal5 5020 -15980 5120 -15880 1 PIX883_IN
port 904 n
rlabel metal5 6520 -15980 6620 -15880 1 PIX884_IN
port 905 n
rlabel metal5 8020 -15980 8120 -15880 1 PIX885_IN
port 906 n
rlabel metal5 9520 -15980 9620 -15880 1 PIX886_IN
port 907 n
rlabel metal5 11020 -15980 11120 -15880 1 PIX887_IN
port 908 n
rlabel metal5 12520 -15980 12620 -15880 1 PIX888_IN
port 909 n
rlabel metal5 14020 -15980 14120 -15880 1 PIX889_IN
port 910 n
rlabel metal5 15520 -15980 15620 -15880 1 PIX890_IN
port 911 n
rlabel metal5 17020 -15980 17120 -15880 1 PIX891_IN
port 912 n
rlabel metal5 18520 -15980 18620 -15880 1 PIX892_IN
port 913 n
rlabel metal5 20020 -15980 20120 -15880 1 PIX893_IN
port 914 n
rlabel metal5 21520 -15980 21620 -15880 1 PIX894_IN
port 915 n
rlabel metal5 23020 -15980 23120 -15880 1 PIX895_IN
port 916 n
rlabel metal5 24520 -15980 24620 -15880 1 PIX896_IN
port 917 n
rlabel metal5 26020 -15980 26120 -15880 1 PIX897_IN
port 918 n
rlabel metal5 27520 -15980 27620 -15880 1 PIX898_IN
port 919 n
rlabel metal5 29020 -15980 29120 -15880 1 PIX899_IN
port 920 n
rlabel metal5 30520 -15980 30620 -15880 1 PIX900_IN
port 921 n
rlabel metal5 32020 -15980 32120 -15880 1 PIX901_IN
port 922 n
rlabel metal5 33520 -15980 33620 -15880 1 PIX902_IN
port 923 n
rlabel metal5 35020 -15980 35120 -15880 1 PIX903_IN
port 924 n
rlabel metal5 36520 -15980 36620 -15880 1 PIX904_IN
port 925 n
rlabel metal5 38020 -15980 38120 -15880 1 PIX905_IN
port 926 n
rlabel metal5 39520 -15980 39620 -15880 1 PIX906_IN
port 927 n
rlabel metal5 41020 -15980 41120 -15880 1 PIX907_IN
port 928 n
rlabel metal5 42520 -15980 42620 -15880 1 PIX908_IN
port 929 n
rlabel metal5 44020 -15980 44120 -15880 1 PIX909_IN
port 930 n
rlabel metal5 45520 -15980 45620 -15880 1 PIX910_IN
port 931 n
rlabel metal5 47020 -15980 47120 -15880 1 PIX911_IN
port 932 n
rlabel metal5 48520 -15980 48620 -15880 1 PIX912_IN
port 933 n
rlabel metal5 50020 -15980 50120 -15880 1 PIX913_IN
port 934 n
rlabel metal5 51520 -15980 51620 -15880 1 PIX914_IN
port 935 n
rlabel metal5 53020 -15980 53120 -15880 1 PIX915_IN
port 936 n
rlabel metal5 54520 -15980 54620 -15880 1 PIX916_IN
port 937 n
rlabel metal5 56020 -15980 56120 -15880 1 PIX917_IN
port 938 n
rlabel metal5 57520 -15980 57620 -15880 1 PIX918_IN
port 939 n
rlabel metal5 59020 -15980 59120 -15880 1 PIX919_IN
port 940 n
rlabel metal5 60520 -15980 60620 -15880 1 PIX920_IN
port 941 n
rlabel metal5 62020 -15980 62120 -15880 1 PIX921_IN
port 942 n
rlabel metal5 63520 -15980 63620 -15880 1 PIX922_IN
port 943 n
rlabel metal5 65020 -15980 65120 -15880 1 PIX923_IN
port 944 n
rlabel metal5 66520 -15980 66620 -15880 1 PIX924_IN
port 945 n
rlabel metal5 68020 -15980 68120 -15880 1 PIX925_IN
port 946 n
rlabel metal5 69520 -15980 69620 -15880 1 PIX926_IN
port 947 n
rlabel metal5 71020 -15980 71120 -15880 1 PIX927_IN
port 948 n
rlabel metal5 72520 -15980 72620 -15880 1 PIX928_IN
port 949 n
rlabel metal5 74020 -15980 74120 -15880 1 PIX929_IN
port 950 n
rlabel metal5 75520 -15980 75620 -15880 1 PIX930_IN
port 951 n
rlabel metal5 77020 -15980 77120 -15880 1 PIX931_IN
port 952 n
rlabel metal5 78520 -15980 78620 -15880 1 PIX932_IN
port 953 n
rlabel metal5 80020 -15980 80120 -15880 1 PIX933_IN
port 954 n
rlabel metal5 81520 -15980 81620 -15880 1 PIX934_IN
port 955 n
rlabel metal5 83020 -15980 83120 -15880 1 PIX935_IN
port 956 n
rlabel metal5 84520 -15980 84620 -15880 1 PIX936_IN
port 957 n
rlabel metal5 86020 -15980 86120 -15880 1 PIX937_IN
port 958 n
rlabel metal5 87520 -15980 87620 -15880 1 PIX938_IN
port 959 n
rlabel metal5 89020 -15980 89120 -15880 1 PIX939_IN
port 960 n
rlabel metal5 90520 -15980 90620 -15880 1 PIX940_IN
port 961 n
rlabel metal5 92020 -15980 92120 -15880 1 PIX941_IN
port 962 n
rlabel metal5 93520 -15980 93620 -15880 1 PIX942_IN
port 963 n
rlabel metal5 95020 -15980 95120 -15880 1 PIX943_IN
port 964 n
rlabel metal5 96520 -15980 96620 -15880 1 PIX944_IN
port 965 n
rlabel metal5 98020 -15980 98120 -15880 1 PIX945_IN
port 966 n
rlabel metal5 99520 -15980 99620 -15880 1 PIX946_IN
port 967 n
rlabel metal5 101020 -15980 101120 -15880 1 PIX947_IN
port 968 n
rlabel metal5 102520 -15980 102620 -15880 1 PIX948_IN
port 969 n
rlabel metal5 104020 -15980 104120 -15880 1 PIX949_IN
port 970 n
rlabel metal5 105520 -15980 105620 -15880 1 PIX950_IN
port 971 n
rlabel metal5 107020 -15980 107120 -15880 1 PIX951_IN
port 972 n
rlabel metal5 108520 -15980 108620 -15880 1 PIX952_IN
port 973 n
rlabel metal5 110020 -15980 110120 -15880 1 PIX953_IN
port 974 n
rlabel metal5 111520 -15980 111620 -15880 1 PIX954_IN
port 975 n
rlabel metal5 113020 -15980 113120 -15880 1 PIX955_IN
port 976 n
rlabel metal5 114520 -15980 114620 -15880 1 PIX956_IN
port 977 n
rlabel metal5 116020 -15980 116120 -15880 1 PIX957_IN
port 978 n
rlabel metal5 117520 -15980 117620 -15880 1 PIX958_IN
port 979 n
rlabel metal5 119020 -15980 119120 -15880 1 PIX959_IN
port 980 n
rlabel metal5 520 -17480 620 -17380 1 PIX960_IN
port 981 n
rlabel metal2 -1500 -17260 -1500 -17215 3 ROW_SEL12
port 982 e
rlabel metal5 2020 -17480 2120 -17380 1 PIX961_IN
port 983 n
rlabel metal5 3520 -17480 3620 -17380 1 PIX962_IN
port 984 n
rlabel metal5 5020 -17480 5120 -17380 1 PIX963_IN
port 985 n
rlabel metal5 6520 -17480 6620 -17380 1 PIX964_IN
port 986 n
rlabel metal5 8020 -17480 8120 -17380 1 PIX965_IN
port 987 n
rlabel metal5 9520 -17480 9620 -17380 1 PIX966_IN
port 988 n
rlabel metal5 11020 -17480 11120 -17380 1 PIX967_IN
port 989 n
rlabel metal5 12520 -17480 12620 -17380 1 PIX968_IN
port 990 n
rlabel metal5 14020 -17480 14120 -17380 1 PIX969_IN
port 991 n
rlabel metal5 15520 -17480 15620 -17380 1 PIX970_IN
port 992 n
rlabel metal5 17020 -17480 17120 -17380 1 PIX971_IN
port 993 n
rlabel metal5 18520 -17480 18620 -17380 1 PIX972_IN
port 994 n
rlabel metal5 20020 -17480 20120 -17380 1 PIX973_IN
port 995 n
rlabel metal5 21520 -17480 21620 -17380 1 PIX974_IN
port 996 n
rlabel metal5 23020 -17480 23120 -17380 1 PIX975_IN
port 997 n
rlabel metal5 24520 -17480 24620 -17380 1 PIX976_IN
port 998 n
rlabel metal5 26020 -17480 26120 -17380 1 PIX977_IN
port 999 n
rlabel metal5 27520 -17480 27620 -17380 1 PIX978_IN
port 1000 n
rlabel metal5 29020 -17480 29120 -17380 1 PIX979_IN
port 1001 n
rlabel metal5 30520 -17480 30620 -17380 1 PIX980_IN
port 1002 n
rlabel metal5 32020 -17480 32120 -17380 1 PIX981_IN
port 1003 n
rlabel metal5 33520 -17480 33620 -17380 1 PIX982_IN
port 1004 n
rlabel metal5 35020 -17480 35120 -17380 1 PIX983_IN
port 1005 n
rlabel metal5 36520 -17480 36620 -17380 1 PIX984_IN
port 1006 n
rlabel metal5 38020 -17480 38120 -17380 1 PIX985_IN
port 1007 n
rlabel metal5 39520 -17480 39620 -17380 1 PIX986_IN
port 1008 n
rlabel metal5 41020 -17480 41120 -17380 1 PIX987_IN
port 1009 n
rlabel metal5 42520 -17480 42620 -17380 1 PIX988_IN
port 1010 n
rlabel metal5 44020 -17480 44120 -17380 1 PIX989_IN
port 1011 n
rlabel metal5 45520 -17480 45620 -17380 1 PIX990_IN
port 1012 n
rlabel metal5 47020 -17480 47120 -17380 1 PIX991_IN
port 1013 n
rlabel metal5 48520 -17480 48620 -17380 1 PIX992_IN
port 1014 n
rlabel metal5 50020 -17480 50120 -17380 1 PIX993_IN
port 1015 n
rlabel metal5 51520 -17480 51620 -17380 1 PIX994_IN
port 1016 n
rlabel metal5 53020 -17480 53120 -17380 1 PIX995_IN
port 1017 n
rlabel metal5 54520 -17480 54620 -17380 1 PIX996_IN
port 1018 n
rlabel metal5 56020 -17480 56120 -17380 1 PIX997_IN
port 1019 n
rlabel metal5 57520 -17480 57620 -17380 1 PIX998_IN
port 1020 n
rlabel metal5 59020 -17480 59120 -17380 1 PIX999_IN
port 1021 n
rlabel metal5 60520 -17480 60620 -17380 1 PIX1000_IN
port 1022 n
rlabel metal5 62020 -17480 62120 -17380 1 PIX1001_IN
port 1023 n
rlabel metal5 63520 -17480 63620 -17380 1 PIX1002_IN
port 1024 n
rlabel metal5 65020 -17480 65120 -17380 1 PIX1003_IN
port 1025 n
rlabel metal5 66520 -17480 66620 -17380 1 PIX1004_IN
port 1026 n
rlabel metal5 68020 -17480 68120 -17380 1 PIX1005_IN
port 1027 n
rlabel metal5 69520 -17480 69620 -17380 1 PIX1006_IN
port 1028 n
rlabel metal5 71020 -17480 71120 -17380 1 PIX1007_IN
port 1029 n
rlabel metal5 72520 -17480 72620 -17380 1 PIX1008_IN
port 1030 n
rlabel metal5 74020 -17480 74120 -17380 1 PIX1009_IN
port 1031 n
rlabel metal5 75520 -17480 75620 -17380 1 PIX1010_IN
port 1032 n
rlabel metal5 77020 -17480 77120 -17380 1 PIX1011_IN
port 1033 n
rlabel metal5 78520 -17480 78620 -17380 1 PIX1012_IN
port 1034 n
rlabel metal5 80020 -17480 80120 -17380 1 PIX1013_IN
port 1035 n
rlabel metal5 81520 -17480 81620 -17380 1 PIX1014_IN
port 1036 n
rlabel metal5 83020 -17480 83120 -17380 1 PIX1015_IN
port 1037 n
rlabel metal5 84520 -17480 84620 -17380 1 PIX1016_IN
port 1038 n
rlabel metal5 86020 -17480 86120 -17380 1 PIX1017_IN
port 1039 n
rlabel metal5 87520 -17480 87620 -17380 1 PIX1018_IN
port 1040 n
rlabel metal5 89020 -17480 89120 -17380 1 PIX1019_IN
port 1041 n
rlabel metal5 90520 -17480 90620 -17380 1 PIX1020_IN
port 1042 n
rlabel metal5 92020 -17480 92120 -17380 1 PIX1021_IN
port 1043 n
rlabel metal5 93520 -17480 93620 -17380 1 PIX1022_IN
port 1044 n
rlabel metal5 95020 -17480 95120 -17380 1 PIX1023_IN
port 1045 n
rlabel metal5 96520 -17480 96620 -17380 1 PIX1024_IN
port 1046 n
rlabel metal5 98020 -17480 98120 -17380 1 PIX1025_IN
port 1047 n
rlabel metal5 99520 -17480 99620 -17380 1 PIX1026_IN
port 1048 n
rlabel metal5 101020 -17480 101120 -17380 1 PIX1027_IN
port 1049 n
rlabel metal5 102520 -17480 102620 -17380 1 PIX1028_IN
port 1050 n
rlabel metal5 104020 -17480 104120 -17380 1 PIX1029_IN
port 1051 n
rlabel metal5 105520 -17480 105620 -17380 1 PIX1030_IN
port 1052 n
rlabel metal5 107020 -17480 107120 -17380 1 PIX1031_IN
port 1053 n
rlabel metal5 108520 -17480 108620 -17380 1 PIX1032_IN
port 1054 n
rlabel metal5 110020 -17480 110120 -17380 1 PIX1033_IN
port 1055 n
rlabel metal5 111520 -17480 111620 -17380 1 PIX1034_IN
port 1056 n
rlabel metal5 113020 -17480 113120 -17380 1 PIX1035_IN
port 1057 n
rlabel metal5 114520 -17480 114620 -17380 1 PIX1036_IN
port 1058 n
rlabel metal5 116020 -17480 116120 -17380 1 PIX1037_IN
port 1059 n
rlabel metal5 117520 -17480 117620 -17380 1 PIX1038_IN
port 1060 n
rlabel metal5 119020 -17480 119120 -17380 1 PIX1039_IN
port 1061 n
rlabel metal5 520 -18980 620 -18880 1 PIX1040_IN
port 1062 n
rlabel metal2 -1500 -18760 -1500 -18715 3 ROW_SEL13
port 1063 e
rlabel metal5 2020 -18980 2120 -18880 1 PIX1041_IN
port 1064 n
rlabel metal5 3520 -18980 3620 -18880 1 PIX1042_IN
port 1065 n
rlabel metal5 5020 -18980 5120 -18880 1 PIX1043_IN
port 1066 n
rlabel metal5 6520 -18980 6620 -18880 1 PIX1044_IN
port 1067 n
rlabel metal5 8020 -18980 8120 -18880 1 PIX1045_IN
port 1068 n
rlabel metal5 9520 -18980 9620 -18880 1 PIX1046_IN
port 1069 n
rlabel metal5 11020 -18980 11120 -18880 1 PIX1047_IN
port 1070 n
rlabel metal5 12520 -18980 12620 -18880 1 PIX1048_IN
port 1071 n
rlabel metal5 14020 -18980 14120 -18880 1 PIX1049_IN
port 1072 n
rlabel metal5 15520 -18980 15620 -18880 1 PIX1050_IN
port 1073 n
rlabel metal5 17020 -18980 17120 -18880 1 PIX1051_IN
port 1074 n
rlabel metal5 18520 -18980 18620 -18880 1 PIX1052_IN
port 1075 n
rlabel metal5 20020 -18980 20120 -18880 1 PIX1053_IN
port 1076 n
rlabel metal5 21520 -18980 21620 -18880 1 PIX1054_IN
port 1077 n
rlabel metal5 23020 -18980 23120 -18880 1 PIX1055_IN
port 1078 n
rlabel metal5 24520 -18980 24620 -18880 1 PIX1056_IN
port 1079 n
rlabel metal5 26020 -18980 26120 -18880 1 PIX1057_IN
port 1080 n
rlabel metal5 27520 -18980 27620 -18880 1 PIX1058_IN
port 1081 n
rlabel metal5 29020 -18980 29120 -18880 1 PIX1059_IN
port 1082 n
rlabel metal5 30520 -18980 30620 -18880 1 PIX1060_IN
port 1083 n
rlabel metal5 32020 -18980 32120 -18880 1 PIX1061_IN
port 1084 n
rlabel metal5 33520 -18980 33620 -18880 1 PIX1062_IN
port 1085 n
rlabel metal5 35020 -18980 35120 -18880 1 PIX1063_IN
port 1086 n
rlabel metal5 36520 -18980 36620 -18880 1 PIX1064_IN
port 1087 n
rlabel metal5 38020 -18980 38120 -18880 1 PIX1065_IN
port 1088 n
rlabel metal5 39520 -18980 39620 -18880 1 PIX1066_IN
port 1089 n
rlabel metal5 41020 -18980 41120 -18880 1 PIX1067_IN
port 1090 n
rlabel metal5 42520 -18980 42620 -18880 1 PIX1068_IN
port 1091 n
rlabel metal5 44020 -18980 44120 -18880 1 PIX1069_IN
port 1092 n
rlabel metal5 45520 -18980 45620 -18880 1 PIX1070_IN
port 1093 n
rlabel metal5 47020 -18980 47120 -18880 1 PIX1071_IN
port 1094 n
rlabel metal5 48520 -18980 48620 -18880 1 PIX1072_IN
port 1095 n
rlabel metal5 50020 -18980 50120 -18880 1 PIX1073_IN
port 1096 n
rlabel metal5 51520 -18980 51620 -18880 1 PIX1074_IN
port 1097 n
rlabel metal5 53020 -18980 53120 -18880 1 PIX1075_IN
port 1098 n
rlabel metal5 54520 -18980 54620 -18880 1 PIX1076_IN
port 1099 n
rlabel metal5 56020 -18980 56120 -18880 1 PIX1077_IN
port 1100 n
rlabel metal5 57520 -18980 57620 -18880 1 PIX1078_IN
port 1101 n
rlabel metal5 59020 -18980 59120 -18880 1 PIX1079_IN
port 1102 n
rlabel metal5 60520 -18980 60620 -18880 1 PIX1080_IN
port 1103 n
rlabel metal5 62020 -18980 62120 -18880 1 PIX1081_IN
port 1104 n
rlabel metal5 63520 -18980 63620 -18880 1 PIX1082_IN
port 1105 n
rlabel metal5 65020 -18980 65120 -18880 1 PIX1083_IN
port 1106 n
rlabel metal5 66520 -18980 66620 -18880 1 PIX1084_IN
port 1107 n
rlabel metal5 68020 -18980 68120 -18880 1 PIX1085_IN
port 1108 n
rlabel metal5 69520 -18980 69620 -18880 1 PIX1086_IN
port 1109 n
rlabel metal5 71020 -18980 71120 -18880 1 PIX1087_IN
port 1110 n
rlabel metal5 72520 -18980 72620 -18880 1 PIX1088_IN
port 1111 n
rlabel metal5 74020 -18980 74120 -18880 1 PIX1089_IN
port 1112 n
rlabel metal5 75520 -18980 75620 -18880 1 PIX1090_IN
port 1113 n
rlabel metal5 77020 -18980 77120 -18880 1 PIX1091_IN
port 1114 n
rlabel metal5 78520 -18980 78620 -18880 1 PIX1092_IN
port 1115 n
rlabel metal5 80020 -18980 80120 -18880 1 PIX1093_IN
port 1116 n
rlabel metal5 81520 -18980 81620 -18880 1 PIX1094_IN
port 1117 n
rlabel metal5 83020 -18980 83120 -18880 1 PIX1095_IN
port 1118 n
rlabel metal5 84520 -18980 84620 -18880 1 PIX1096_IN
port 1119 n
rlabel metal5 86020 -18980 86120 -18880 1 PIX1097_IN
port 1120 n
rlabel metal5 87520 -18980 87620 -18880 1 PIX1098_IN
port 1121 n
rlabel metal5 89020 -18980 89120 -18880 1 PIX1099_IN
port 1122 n
rlabel metal5 90520 -18980 90620 -18880 1 PIX1100_IN
port 1123 n
rlabel metal5 92020 -18980 92120 -18880 1 PIX1101_IN
port 1124 n
rlabel metal5 93520 -18980 93620 -18880 1 PIX1102_IN
port 1125 n
rlabel metal5 95020 -18980 95120 -18880 1 PIX1103_IN
port 1126 n
rlabel metal5 96520 -18980 96620 -18880 1 PIX1104_IN
port 1127 n
rlabel metal5 98020 -18980 98120 -18880 1 PIX1105_IN
port 1128 n
rlabel metal5 99520 -18980 99620 -18880 1 PIX1106_IN
port 1129 n
rlabel metal5 101020 -18980 101120 -18880 1 PIX1107_IN
port 1130 n
rlabel metal5 102520 -18980 102620 -18880 1 PIX1108_IN
port 1131 n
rlabel metal5 104020 -18980 104120 -18880 1 PIX1109_IN
port 1132 n
rlabel metal5 105520 -18980 105620 -18880 1 PIX1110_IN
port 1133 n
rlabel metal5 107020 -18980 107120 -18880 1 PIX1111_IN
port 1134 n
rlabel metal5 108520 -18980 108620 -18880 1 PIX1112_IN
port 1135 n
rlabel metal5 110020 -18980 110120 -18880 1 PIX1113_IN
port 1136 n
rlabel metal5 111520 -18980 111620 -18880 1 PIX1114_IN
port 1137 n
rlabel metal5 113020 -18980 113120 -18880 1 PIX1115_IN
port 1138 n
rlabel metal5 114520 -18980 114620 -18880 1 PIX1116_IN
port 1139 n
rlabel metal5 116020 -18980 116120 -18880 1 PIX1117_IN
port 1140 n
rlabel metal5 117520 -18980 117620 -18880 1 PIX1118_IN
port 1141 n
rlabel metal5 119020 -18980 119120 -18880 1 PIX1119_IN
port 1142 n
rlabel metal5 520 -20480 620 -20380 1 PIX1120_IN
port 1143 n
rlabel metal2 -1500 -20260 -1500 -20215 3 ROW_SEL14
port 1144 e
rlabel metal5 2020 -20480 2120 -20380 1 PIX1121_IN
port 1145 n
rlabel metal5 3520 -20480 3620 -20380 1 PIX1122_IN
port 1146 n
rlabel metal5 5020 -20480 5120 -20380 1 PIX1123_IN
port 1147 n
rlabel metal5 6520 -20480 6620 -20380 1 PIX1124_IN
port 1148 n
rlabel metal5 8020 -20480 8120 -20380 1 PIX1125_IN
port 1149 n
rlabel metal5 9520 -20480 9620 -20380 1 PIX1126_IN
port 1150 n
rlabel metal5 11020 -20480 11120 -20380 1 PIX1127_IN
port 1151 n
rlabel metal5 12520 -20480 12620 -20380 1 PIX1128_IN
port 1152 n
rlabel metal5 14020 -20480 14120 -20380 1 PIX1129_IN
port 1153 n
rlabel metal5 15520 -20480 15620 -20380 1 PIX1130_IN
port 1154 n
rlabel metal5 17020 -20480 17120 -20380 1 PIX1131_IN
port 1155 n
rlabel metal5 18520 -20480 18620 -20380 1 PIX1132_IN
port 1156 n
rlabel metal5 20020 -20480 20120 -20380 1 PIX1133_IN
port 1157 n
rlabel metal5 21520 -20480 21620 -20380 1 PIX1134_IN
port 1158 n
rlabel metal5 23020 -20480 23120 -20380 1 PIX1135_IN
port 1159 n
rlabel metal5 24520 -20480 24620 -20380 1 PIX1136_IN
port 1160 n
rlabel metal5 26020 -20480 26120 -20380 1 PIX1137_IN
port 1161 n
rlabel metal5 27520 -20480 27620 -20380 1 PIX1138_IN
port 1162 n
rlabel metal5 29020 -20480 29120 -20380 1 PIX1139_IN
port 1163 n
rlabel metal5 30520 -20480 30620 -20380 1 PIX1140_IN
port 1164 n
rlabel metal5 32020 -20480 32120 -20380 1 PIX1141_IN
port 1165 n
rlabel metal5 33520 -20480 33620 -20380 1 PIX1142_IN
port 1166 n
rlabel metal5 35020 -20480 35120 -20380 1 PIX1143_IN
port 1167 n
rlabel metal5 36520 -20480 36620 -20380 1 PIX1144_IN
port 1168 n
rlabel metal5 38020 -20480 38120 -20380 1 PIX1145_IN
port 1169 n
rlabel metal5 39520 -20480 39620 -20380 1 PIX1146_IN
port 1170 n
rlabel metal5 41020 -20480 41120 -20380 1 PIX1147_IN
port 1171 n
rlabel metal5 42520 -20480 42620 -20380 1 PIX1148_IN
port 1172 n
rlabel metal5 44020 -20480 44120 -20380 1 PIX1149_IN
port 1173 n
rlabel metal5 45520 -20480 45620 -20380 1 PIX1150_IN
port 1174 n
rlabel metal5 47020 -20480 47120 -20380 1 PIX1151_IN
port 1175 n
rlabel metal5 48520 -20480 48620 -20380 1 PIX1152_IN
port 1176 n
rlabel metal5 50020 -20480 50120 -20380 1 PIX1153_IN
port 1177 n
rlabel metal5 51520 -20480 51620 -20380 1 PIX1154_IN
port 1178 n
rlabel metal5 53020 -20480 53120 -20380 1 PIX1155_IN
port 1179 n
rlabel metal5 54520 -20480 54620 -20380 1 PIX1156_IN
port 1180 n
rlabel metal5 56020 -20480 56120 -20380 1 PIX1157_IN
port 1181 n
rlabel metal5 57520 -20480 57620 -20380 1 PIX1158_IN
port 1182 n
rlabel metal5 59020 -20480 59120 -20380 1 PIX1159_IN
port 1183 n
rlabel metal5 60520 -20480 60620 -20380 1 PIX1160_IN
port 1184 n
rlabel metal5 62020 -20480 62120 -20380 1 PIX1161_IN
port 1185 n
rlabel metal5 63520 -20480 63620 -20380 1 PIX1162_IN
port 1186 n
rlabel metal5 65020 -20480 65120 -20380 1 PIX1163_IN
port 1187 n
rlabel metal5 66520 -20480 66620 -20380 1 PIX1164_IN
port 1188 n
rlabel metal5 68020 -20480 68120 -20380 1 PIX1165_IN
port 1189 n
rlabel metal5 69520 -20480 69620 -20380 1 PIX1166_IN
port 1190 n
rlabel metal5 71020 -20480 71120 -20380 1 PIX1167_IN
port 1191 n
rlabel metal5 72520 -20480 72620 -20380 1 PIX1168_IN
port 1192 n
rlabel metal5 74020 -20480 74120 -20380 1 PIX1169_IN
port 1193 n
rlabel metal5 75520 -20480 75620 -20380 1 PIX1170_IN
port 1194 n
rlabel metal5 77020 -20480 77120 -20380 1 PIX1171_IN
port 1195 n
rlabel metal5 78520 -20480 78620 -20380 1 PIX1172_IN
port 1196 n
rlabel metal5 80020 -20480 80120 -20380 1 PIX1173_IN
port 1197 n
rlabel metal5 81520 -20480 81620 -20380 1 PIX1174_IN
port 1198 n
rlabel metal5 83020 -20480 83120 -20380 1 PIX1175_IN
port 1199 n
rlabel metal5 84520 -20480 84620 -20380 1 PIX1176_IN
port 1200 n
rlabel metal5 86020 -20480 86120 -20380 1 PIX1177_IN
port 1201 n
rlabel metal5 87520 -20480 87620 -20380 1 PIX1178_IN
port 1202 n
rlabel metal5 89020 -20480 89120 -20380 1 PIX1179_IN
port 1203 n
rlabel metal5 90520 -20480 90620 -20380 1 PIX1180_IN
port 1204 n
rlabel metal5 92020 -20480 92120 -20380 1 PIX1181_IN
port 1205 n
rlabel metal5 93520 -20480 93620 -20380 1 PIX1182_IN
port 1206 n
rlabel metal5 95020 -20480 95120 -20380 1 PIX1183_IN
port 1207 n
rlabel metal5 96520 -20480 96620 -20380 1 PIX1184_IN
port 1208 n
rlabel metal5 98020 -20480 98120 -20380 1 PIX1185_IN
port 1209 n
rlabel metal5 99520 -20480 99620 -20380 1 PIX1186_IN
port 1210 n
rlabel metal5 101020 -20480 101120 -20380 1 PIX1187_IN
port 1211 n
rlabel metal5 102520 -20480 102620 -20380 1 PIX1188_IN
port 1212 n
rlabel metal5 104020 -20480 104120 -20380 1 PIX1189_IN
port 1213 n
rlabel metal5 105520 -20480 105620 -20380 1 PIX1190_IN
port 1214 n
rlabel metal5 107020 -20480 107120 -20380 1 PIX1191_IN
port 1215 n
rlabel metal5 108520 -20480 108620 -20380 1 PIX1192_IN
port 1216 n
rlabel metal5 110020 -20480 110120 -20380 1 PIX1193_IN
port 1217 n
rlabel metal5 111520 -20480 111620 -20380 1 PIX1194_IN
port 1218 n
rlabel metal5 113020 -20480 113120 -20380 1 PIX1195_IN
port 1219 n
rlabel metal5 114520 -20480 114620 -20380 1 PIX1196_IN
port 1220 n
rlabel metal5 116020 -20480 116120 -20380 1 PIX1197_IN
port 1221 n
rlabel metal5 117520 -20480 117620 -20380 1 PIX1198_IN
port 1222 n
rlabel metal5 119020 -20480 119120 -20380 1 PIX1199_IN
port 1223 n
rlabel metal5 520 -21980 620 -21880 1 PIX1200_IN
port 1224 n
rlabel metal2 -1500 -21760 -1500 -21715 3 ROW_SEL15
port 1225 e
rlabel metal5 2020 -21980 2120 -21880 1 PIX1201_IN
port 1226 n
rlabel metal5 3520 -21980 3620 -21880 1 PIX1202_IN
port 1227 n
rlabel metal5 5020 -21980 5120 -21880 1 PIX1203_IN
port 1228 n
rlabel metal5 6520 -21980 6620 -21880 1 PIX1204_IN
port 1229 n
rlabel metal5 8020 -21980 8120 -21880 1 PIX1205_IN
port 1230 n
rlabel metal5 9520 -21980 9620 -21880 1 PIX1206_IN
port 1231 n
rlabel metal5 11020 -21980 11120 -21880 1 PIX1207_IN
port 1232 n
rlabel metal5 12520 -21980 12620 -21880 1 PIX1208_IN
port 1233 n
rlabel metal5 14020 -21980 14120 -21880 1 PIX1209_IN
port 1234 n
rlabel metal5 15520 -21980 15620 -21880 1 PIX1210_IN
port 1235 n
rlabel metal5 17020 -21980 17120 -21880 1 PIX1211_IN
port 1236 n
rlabel metal5 18520 -21980 18620 -21880 1 PIX1212_IN
port 1237 n
rlabel metal5 20020 -21980 20120 -21880 1 PIX1213_IN
port 1238 n
rlabel metal5 21520 -21980 21620 -21880 1 PIX1214_IN
port 1239 n
rlabel metal5 23020 -21980 23120 -21880 1 PIX1215_IN
port 1240 n
rlabel metal5 24520 -21980 24620 -21880 1 PIX1216_IN
port 1241 n
rlabel metal5 26020 -21980 26120 -21880 1 PIX1217_IN
port 1242 n
rlabel metal5 27520 -21980 27620 -21880 1 PIX1218_IN
port 1243 n
rlabel metal5 29020 -21980 29120 -21880 1 PIX1219_IN
port 1244 n
rlabel metal5 30520 -21980 30620 -21880 1 PIX1220_IN
port 1245 n
rlabel metal5 32020 -21980 32120 -21880 1 PIX1221_IN
port 1246 n
rlabel metal5 33520 -21980 33620 -21880 1 PIX1222_IN
port 1247 n
rlabel metal5 35020 -21980 35120 -21880 1 PIX1223_IN
port 1248 n
rlabel metal5 36520 -21980 36620 -21880 1 PIX1224_IN
port 1249 n
rlabel metal5 38020 -21980 38120 -21880 1 PIX1225_IN
port 1250 n
rlabel metal5 39520 -21980 39620 -21880 1 PIX1226_IN
port 1251 n
rlabel metal5 41020 -21980 41120 -21880 1 PIX1227_IN
port 1252 n
rlabel metal5 42520 -21980 42620 -21880 1 PIX1228_IN
port 1253 n
rlabel metal5 44020 -21980 44120 -21880 1 PIX1229_IN
port 1254 n
rlabel metal5 45520 -21980 45620 -21880 1 PIX1230_IN
port 1255 n
rlabel metal5 47020 -21980 47120 -21880 1 PIX1231_IN
port 1256 n
rlabel metal5 48520 -21980 48620 -21880 1 PIX1232_IN
port 1257 n
rlabel metal5 50020 -21980 50120 -21880 1 PIX1233_IN
port 1258 n
rlabel metal5 51520 -21980 51620 -21880 1 PIX1234_IN
port 1259 n
rlabel metal5 53020 -21980 53120 -21880 1 PIX1235_IN
port 1260 n
rlabel metal5 54520 -21980 54620 -21880 1 PIX1236_IN
port 1261 n
rlabel metal5 56020 -21980 56120 -21880 1 PIX1237_IN
port 1262 n
rlabel metal5 57520 -21980 57620 -21880 1 PIX1238_IN
port 1263 n
rlabel metal5 59020 -21980 59120 -21880 1 PIX1239_IN
port 1264 n
rlabel metal5 60520 -21980 60620 -21880 1 PIX1240_IN
port 1265 n
rlabel metal5 62020 -21980 62120 -21880 1 PIX1241_IN
port 1266 n
rlabel metal5 63520 -21980 63620 -21880 1 PIX1242_IN
port 1267 n
rlabel metal5 65020 -21980 65120 -21880 1 PIX1243_IN
port 1268 n
rlabel metal5 66520 -21980 66620 -21880 1 PIX1244_IN
port 1269 n
rlabel metal5 68020 -21980 68120 -21880 1 PIX1245_IN
port 1270 n
rlabel metal5 69520 -21980 69620 -21880 1 PIX1246_IN
port 1271 n
rlabel metal5 71020 -21980 71120 -21880 1 PIX1247_IN
port 1272 n
rlabel metal5 72520 -21980 72620 -21880 1 PIX1248_IN
port 1273 n
rlabel metal5 74020 -21980 74120 -21880 1 PIX1249_IN
port 1274 n
rlabel metal5 75520 -21980 75620 -21880 1 PIX1250_IN
port 1275 n
rlabel metal5 77020 -21980 77120 -21880 1 PIX1251_IN
port 1276 n
rlabel metal5 78520 -21980 78620 -21880 1 PIX1252_IN
port 1277 n
rlabel metal5 80020 -21980 80120 -21880 1 PIX1253_IN
port 1278 n
rlabel metal5 81520 -21980 81620 -21880 1 PIX1254_IN
port 1279 n
rlabel metal5 83020 -21980 83120 -21880 1 PIX1255_IN
port 1280 n
rlabel metal5 84520 -21980 84620 -21880 1 PIX1256_IN
port 1281 n
rlabel metal5 86020 -21980 86120 -21880 1 PIX1257_IN
port 1282 n
rlabel metal5 87520 -21980 87620 -21880 1 PIX1258_IN
port 1283 n
rlabel metal5 89020 -21980 89120 -21880 1 PIX1259_IN
port 1284 n
rlabel metal5 90520 -21980 90620 -21880 1 PIX1260_IN
port 1285 n
rlabel metal5 92020 -21980 92120 -21880 1 PIX1261_IN
port 1286 n
rlabel metal5 93520 -21980 93620 -21880 1 PIX1262_IN
port 1287 n
rlabel metal5 95020 -21980 95120 -21880 1 PIX1263_IN
port 1288 n
rlabel metal5 96520 -21980 96620 -21880 1 PIX1264_IN
port 1289 n
rlabel metal5 98020 -21980 98120 -21880 1 PIX1265_IN
port 1290 n
rlabel metal5 99520 -21980 99620 -21880 1 PIX1266_IN
port 1291 n
rlabel metal5 101020 -21980 101120 -21880 1 PIX1267_IN
port 1292 n
rlabel metal5 102520 -21980 102620 -21880 1 PIX1268_IN
port 1293 n
rlabel metal5 104020 -21980 104120 -21880 1 PIX1269_IN
port 1294 n
rlabel metal5 105520 -21980 105620 -21880 1 PIX1270_IN
port 1295 n
rlabel metal5 107020 -21980 107120 -21880 1 PIX1271_IN
port 1296 n
rlabel metal5 108520 -21980 108620 -21880 1 PIX1272_IN
port 1297 n
rlabel metal5 110020 -21980 110120 -21880 1 PIX1273_IN
port 1298 n
rlabel metal5 111520 -21980 111620 -21880 1 PIX1274_IN
port 1299 n
rlabel metal5 113020 -21980 113120 -21880 1 PIX1275_IN
port 1300 n
rlabel metal5 114520 -21980 114620 -21880 1 PIX1276_IN
port 1301 n
rlabel metal5 116020 -21980 116120 -21880 1 PIX1277_IN
port 1302 n
rlabel metal5 117520 -21980 117620 -21880 1 PIX1278_IN
port 1303 n
rlabel metal5 119020 -21980 119120 -21880 1 PIX1279_IN
port 1304 n
rlabel metal5 520 -23480 620 -23380 1 PIX1280_IN
port 1305 n
rlabel metal2 -1500 -23260 -1500 -23215 3 ROW_SEL16
port 1306 e
rlabel metal5 2020 -23480 2120 -23380 1 PIX1281_IN
port 1307 n
rlabel metal5 3520 -23480 3620 -23380 1 PIX1282_IN
port 1308 n
rlabel metal5 5020 -23480 5120 -23380 1 PIX1283_IN
port 1309 n
rlabel metal5 6520 -23480 6620 -23380 1 PIX1284_IN
port 1310 n
rlabel metal5 8020 -23480 8120 -23380 1 PIX1285_IN
port 1311 n
rlabel metal5 9520 -23480 9620 -23380 1 PIX1286_IN
port 1312 n
rlabel metal5 11020 -23480 11120 -23380 1 PIX1287_IN
port 1313 n
rlabel metal5 12520 -23480 12620 -23380 1 PIX1288_IN
port 1314 n
rlabel metal5 14020 -23480 14120 -23380 1 PIX1289_IN
port 1315 n
rlabel metal5 15520 -23480 15620 -23380 1 PIX1290_IN
port 1316 n
rlabel metal5 17020 -23480 17120 -23380 1 PIX1291_IN
port 1317 n
rlabel metal5 18520 -23480 18620 -23380 1 PIX1292_IN
port 1318 n
rlabel metal5 20020 -23480 20120 -23380 1 PIX1293_IN
port 1319 n
rlabel metal5 21520 -23480 21620 -23380 1 PIX1294_IN
port 1320 n
rlabel metal5 23020 -23480 23120 -23380 1 PIX1295_IN
port 1321 n
rlabel metal5 24520 -23480 24620 -23380 1 PIX1296_IN
port 1322 n
rlabel metal5 26020 -23480 26120 -23380 1 PIX1297_IN
port 1323 n
rlabel metal5 27520 -23480 27620 -23380 1 PIX1298_IN
port 1324 n
rlabel metal5 29020 -23480 29120 -23380 1 PIX1299_IN
port 1325 n
rlabel metal5 30520 -23480 30620 -23380 1 PIX1300_IN
port 1326 n
rlabel metal5 32020 -23480 32120 -23380 1 PIX1301_IN
port 1327 n
rlabel metal5 33520 -23480 33620 -23380 1 PIX1302_IN
port 1328 n
rlabel metal5 35020 -23480 35120 -23380 1 PIX1303_IN
port 1329 n
rlabel metal5 36520 -23480 36620 -23380 1 PIX1304_IN
port 1330 n
rlabel metal5 38020 -23480 38120 -23380 1 PIX1305_IN
port 1331 n
rlabel metal5 39520 -23480 39620 -23380 1 PIX1306_IN
port 1332 n
rlabel metal5 41020 -23480 41120 -23380 1 PIX1307_IN
port 1333 n
rlabel metal5 42520 -23480 42620 -23380 1 PIX1308_IN
port 1334 n
rlabel metal5 44020 -23480 44120 -23380 1 PIX1309_IN
port 1335 n
rlabel metal5 45520 -23480 45620 -23380 1 PIX1310_IN
port 1336 n
rlabel metal5 47020 -23480 47120 -23380 1 PIX1311_IN
port 1337 n
rlabel metal5 48520 -23480 48620 -23380 1 PIX1312_IN
port 1338 n
rlabel metal5 50020 -23480 50120 -23380 1 PIX1313_IN
port 1339 n
rlabel metal5 51520 -23480 51620 -23380 1 PIX1314_IN
port 1340 n
rlabel metal5 53020 -23480 53120 -23380 1 PIX1315_IN
port 1341 n
rlabel metal5 54520 -23480 54620 -23380 1 PIX1316_IN
port 1342 n
rlabel metal5 56020 -23480 56120 -23380 1 PIX1317_IN
port 1343 n
rlabel metal5 57520 -23480 57620 -23380 1 PIX1318_IN
port 1344 n
rlabel metal5 59020 -23480 59120 -23380 1 PIX1319_IN
port 1345 n
rlabel metal5 60520 -23480 60620 -23380 1 PIX1320_IN
port 1346 n
rlabel metal5 62020 -23480 62120 -23380 1 PIX1321_IN
port 1347 n
rlabel metal5 63520 -23480 63620 -23380 1 PIX1322_IN
port 1348 n
rlabel metal5 65020 -23480 65120 -23380 1 PIX1323_IN
port 1349 n
rlabel metal5 66520 -23480 66620 -23380 1 PIX1324_IN
port 1350 n
rlabel metal5 68020 -23480 68120 -23380 1 PIX1325_IN
port 1351 n
rlabel metal5 69520 -23480 69620 -23380 1 PIX1326_IN
port 1352 n
rlabel metal5 71020 -23480 71120 -23380 1 PIX1327_IN
port 1353 n
rlabel metal5 72520 -23480 72620 -23380 1 PIX1328_IN
port 1354 n
rlabel metal5 74020 -23480 74120 -23380 1 PIX1329_IN
port 1355 n
rlabel metal5 75520 -23480 75620 -23380 1 PIX1330_IN
port 1356 n
rlabel metal5 77020 -23480 77120 -23380 1 PIX1331_IN
port 1357 n
rlabel metal5 78520 -23480 78620 -23380 1 PIX1332_IN
port 1358 n
rlabel metal5 80020 -23480 80120 -23380 1 PIX1333_IN
port 1359 n
rlabel metal5 81520 -23480 81620 -23380 1 PIX1334_IN
port 1360 n
rlabel metal5 83020 -23480 83120 -23380 1 PIX1335_IN
port 1361 n
rlabel metal5 84520 -23480 84620 -23380 1 PIX1336_IN
port 1362 n
rlabel metal5 86020 -23480 86120 -23380 1 PIX1337_IN
port 1363 n
rlabel metal5 87520 -23480 87620 -23380 1 PIX1338_IN
port 1364 n
rlabel metal5 89020 -23480 89120 -23380 1 PIX1339_IN
port 1365 n
rlabel metal5 90520 -23480 90620 -23380 1 PIX1340_IN
port 1366 n
rlabel metal5 92020 -23480 92120 -23380 1 PIX1341_IN
port 1367 n
rlabel metal5 93520 -23480 93620 -23380 1 PIX1342_IN
port 1368 n
rlabel metal5 95020 -23480 95120 -23380 1 PIX1343_IN
port 1369 n
rlabel metal5 96520 -23480 96620 -23380 1 PIX1344_IN
port 1370 n
rlabel metal5 98020 -23480 98120 -23380 1 PIX1345_IN
port 1371 n
rlabel metal5 99520 -23480 99620 -23380 1 PIX1346_IN
port 1372 n
rlabel metal5 101020 -23480 101120 -23380 1 PIX1347_IN
port 1373 n
rlabel metal5 102520 -23480 102620 -23380 1 PIX1348_IN
port 1374 n
rlabel metal5 104020 -23480 104120 -23380 1 PIX1349_IN
port 1375 n
rlabel metal5 105520 -23480 105620 -23380 1 PIX1350_IN
port 1376 n
rlabel metal5 107020 -23480 107120 -23380 1 PIX1351_IN
port 1377 n
rlabel metal5 108520 -23480 108620 -23380 1 PIX1352_IN
port 1378 n
rlabel metal5 110020 -23480 110120 -23380 1 PIX1353_IN
port 1379 n
rlabel metal5 111520 -23480 111620 -23380 1 PIX1354_IN
port 1380 n
rlabel metal5 113020 -23480 113120 -23380 1 PIX1355_IN
port 1381 n
rlabel metal5 114520 -23480 114620 -23380 1 PIX1356_IN
port 1382 n
rlabel metal5 116020 -23480 116120 -23380 1 PIX1357_IN
port 1383 n
rlabel metal5 117520 -23480 117620 -23380 1 PIX1358_IN
port 1384 n
rlabel metal5 119020 -23480 119120 -23380 1 PIX1359_IN
port 1385 n
rlabel metal5 520 -24980 620 -24880 1 PIX1360_IN
port 1386 n
rlabel metal2 -1500 -24760 -1500 -24715 3 ROW_SEL17
port 1387 e
rlabel metal5 2020 -24980 2120 -24880 1 PIX1361_IN
port 1388 n
rlabel metal5 3520 -24980 3620 -24880 1 PIX1362_IN
port 1389 n
rlabel metal5 5020 -24980 5120 -24880 1 PIX1363_IN
port 1390 n
rlabel metal5 6520 -24980 6620 -24880 1 PIX1364_IN
port 1391 n
rlabel metal5 8020 -24980 8120 -24880 1 PIX1365_IN
port 1392 n
rlabel metal5 9520 -24980 9620 -24880 1 PIX1366_IN
port 1393 n
rlabel metal5 11020 -24980 11120 -24880 1 PIX1367_IN
port 1394 n
rlabel metal5 12520 -24980 12620 -24880 1 PIX1368_IN
port 1395 n
rlabel metal5 14020 -24980 14120 -24880 1 PIX1369_IN
port 1396 n
rlabel metal5 15520 -24980 15620 -24880 1 PIX1370_IN
port 1397 n
rlabel metal5 17020 -24980 17120 -24880 1 PIX1371_IN
port 1398 n
rlabel metal5 18520 -24980 18620 -24880 1 PIX1372_IN
port 1399 n
rlabel metal5 20020 -24980 20120 -24880 1 PIX1373_IN
port 1400 n
rlabel metal5 21520 -24980 21620 -24880 1 PIX1374_IN
port 1401 n
rlabel metal5 23020 -24980 23120 -24880 1 PIX1375_IN
port 1402 n
rlabel metal5 24520 -24980 24620 -24880 1 PIX1376_IN
port 1403 n
rlabel metal5 26020 -24980 26120 -24880 1 PIX1377_IN
port 1404 n
rlabel metal5 27520 -24980 27620 -24880 1 PIX1378_IN
port 1405 n
rlabel metal5 29020 -24980 29120 -24880 1 PIX1379_IN
port 1406 n
rlabel metal5 30520 -24980 30620 -24880 1 PIX1380_IN
port 1407 n
rlabel metal5 32020 -24980 32120 -24880 1 PIX1381_IN
port 1408 n
rlabel metal5 33520 -24980 33620 -24880 1 PIX1382_IN
port 1409 n
rlabel metal5 35020 -24980 35120 -24880 1 PIX1383_IN
port 1410 n
rlabel metal5 36520 -24980 36620 -24880 1 PIX1384_IN
port 1411 n
rlabel metal5 38020 -24980 38120 -24880 1 PIX1385_IN
port 1412 n
rlabel metal5 39520 -24980 39620 -24880 1 PIX1386_IN
port 1413 n
rlabel metal5 41020 -24980 41120 -24880 1 PIX1387_IN
port 1414 n
rlabel metal5 42520 -24980 42620 -24880 1 PIX1388_IN
port 1415 n
rlabel metal5 44020 -24980 44120 -24880 1 PIX1389_IN
port 1416 n
rlabel metal5 45520 -24980 45620 -24880 1 PIX1390_IN
port 1417 n
rlabel metal5 47020 -24980 47120 -24880 1 PIX1391_IN
port 1418 n
rlabel metal5 48520 -24980 48620 -24880 1 PIX1392_IN
port 1419 n
rlabel metal5 50020 -24980 50120 -24880 1 PIX1393_IN
port 1420 n
rlabel metal5 51520 -24980 51620 -24880 1 PIX1394_IN
port 1421 n
rlabel metal5 53020 -24980 53120 -24880 1 PIX1395_IN
port 1422 n
rlabel metal5 54520 -24980 54620 -24880 1 PIX1396_IN
port 1423 n
rlabel metal5 56020 -24980 56120 -24880 1 PIX1397_IN
port 1424 n
rlabel metal5 57520 -24980 57620 -24880 1 PIX1398_IN
port 1425 n
rlabel metal5 59020 -24980 59120 -24880 1 PIX1399_IN
port 1426 n
rlabel metal5 60520 -24980 60620 -24880 1 PIX1400_IN
port 1427 n
rlabel metal5 62020 -24980 62120 -24880 1 PIX1401_IN
port 1428 n
rlabel metal5 63520 -24980 63620 -24880 1 PIX1402_IN
port 1429 n
rlabel metal5 65020 -24980 65120 -24880 1 PIX1403_IN
port 1430 n
rlabel metal5 66520 -24980 66620 -24880 1 PIX1404_IN
port 1431 n
rlabel metal5 68020 -24980 68120 -24880 1 PIX1405_IN
port 1432 n
rlabel metal5 69520 -24980 69620 -24880 1 PIX1406_IN
port 1433 n
rlabel metal5 71020 -24980 71120 -24880 1 PIX1407_IN
port 1434 n
rlabel metal5 72520 -24980 72620 -24880 1 PIX1408_IN
port 1435 n
rlabel metal5 74020 -24980 74120 -24880 1 PIX1409_IN
port 1436 n
rlabel metal5 75520 -24980 75620 -24880 1 PIX1410_IN
port 1437 n
rlabel metal5 77020 -24980 77120 -24880 1 PIX1411_IN
port 1438 n
rlabel metal5 78520 -24980 78620 -24880 1 PIX1412_IN
port 1439 n
rlabel metal5 80020 -24980 80120 -24880 1 PIX1413_IN
port 1440 n
rlabel metal5 81520 -24980 81620 -24880 1 PIX1414_IN
port 1441 n
rlabel metal5 83020 -24980 83120 -24880 1 PIX1415_IN
port 1442 n
rlabel metal5 84520 -24980 84620 -24880 1 PIX1416_IN
port 1443 n
rlabel metal5 86020 -24980 86120 -24880 1 PIX1417_IN
port 1444 n
rlabel metal5 87520 -24980 87620 -24880 1 PIX1418_IN
port 1445 n
rlabel metal5 89020 -24980 89120 -24880 1 PIX1419_IN
port 1446 n
rlabel metal5 90520 -24980 90620 -24880 1 PIX1420_IN
port 1447 n
rlabel metal5 92020 -24980 92120 -24880 1 PIX1421_IN
port 1448 n
rlabel metal5 93520 -24980 93620 -24880 1 PIX1422_IN
port 1449 n
rlabel metal5 95020 -24980 95120 -24880 1 PIX1423_IN
port 1450 n
rlabel metal5 96520 -24980 96620 -24880 1 PIX1424_IN
port 1451 n
rlabel metal5 98020 -24980 98120 -24880 1 PIX1425_IN
port 1452 n
rlabel metal5 99520 -24980 99620 -24880 1 PIX1426_IN
port 1453 n
rlabel metal5 101020 -24980 101120 -24880 1 PIX1427_IN
port 1454 n
rlabel metal5 102520 -24980 102620 -24880 1 PIX1428_IN
port 1455 n
rlabel metal5 104020 -24980 104120 -24880 1 PIX1429_IN
port 1456 n
rlabel metal5 105520 -24980 105620 -24880 1 PIX1430_IN
port 1457 n
rlabel metal5 107020 -24980 107120 -24880 1 PIX1431_IN
port 1458 n
rlabel metal5 108520 -24980 108620 -24880 1 PIX1432_IN
port 1459 n
rlabel metal5 110020 -24980 110120 -24880 1 PIX1433_IN
port 1460 n
rlabel metal5 111520 -24980 111620 -24880 1 PIX1434_IN
port 1461 n
rlabel metal5 113020 -24980 113120 -24880 1 PIX1435_IN
port 1462 n
rlabel metal5 114520 -24980 114620 -24880 1 PIX1436_IN
port 1463 n
rlabel metal5 116020 -24980 116120 -24880 1 PIX1437_IN
port 1464 n
rlabel metal5 117520 -24980 117620 -24880 1 PIX1438_IN
port 1465 n
rlabel metal5 119020 -24980 119120 -24880 1 PIX1439_IN
port 1466 n
rlabel metal5 520 -26480 620 -26380 1 PIX1440_IN
port 1467 n
rlabel metal2 -1500 -26260 -1500 -26215 3 ROW_SEL18
port 1468 e
rlabel metal5 2020 -26480 2120 -26380 1 PIX1441_IN
port 1469 n
rlabel metal5 3520 -26480 3620 -26380 1 PIX1442_IN
port 1470 n
rlabel metal5 5020 -26480 5120 -26380 1 PIX1443_IN
port 1471 n
rlabel metal5 6520 -26480 6620 -26380 1 PIX1444_IN
port 1472 n
rlabel metal5 8020 -26480 8120 -26380 1 PIX1445_IN
port 1473 n
rlabel metal5 9520 -26480 9620 -26380 1 PIX1446_IN
port 1474 n
rlabel metal5 11020 -26480 11120 -26380 1 PIX1447_IN
port 1475 n
rlabel metal5 12520 -26480 12620 -26380 1 PIX1448_IN
port 1476 n
rlabel metal5 14020 -26480 14120 -26380 1 PIX1449_IN
port 1477 n
rlabel metal5 15520 -26480 15620 -26380 1 PIX1450_IN
port 1478 n
rlabel metal5 17020 -26480 17120 -26380 1 PIX1451_IN
port 1479 n
rlabel metal5 18520 -26480 18620 -26380 1 PIX1452_IN
port 1480 n
rlabel metal5 20020 -26480 20120 -26380 1 PIX1453_IN
port 1481 n
rlabel metal5 21520 -26480 21620 -26380 1 PIX1454_IN
port 1482 n
rlabel metal5 23020 -26480 23120 -26380 1 PIX1455_IN
port 1483 n
rlabel metal5 24520 -26480 24620 -26380 1 PIX1456_IN
port 1484 n
rlabel metal5 26020 -26480 26120 -26380 1 PIX1457_IN
port 1485 n
rlabel metal5 27520 -26480 27620 -26380 1 PIX1458_IN
port 1486 n
rlabel metal5 29020 -26480 29120 -26380 1 PIX1459_IN
port 1487 n
rlabel metal5 30520 -26480 30620 -26380 1 PIX1460_IN
port 1488 n
rlabel metal5 32020 -26480 32120 -26380 1 PIX1461_IN
port 1489 n
rlabel metal5 33520 -26480 33620 -26380 1 PIX1462_IN
port 1490 n
rlabel metal5 35020 -26480 35120 -26380 1 PIX1463_IN
port 1491 n
rlabel metal5 36520 -26480 36620 -26380 1 PIX1464_IN
port 1492 n
rlabel metal5 38020 -26480 38120 -26380 1 PIX1465_IN
port 1493 n
rlabel metal5 39520 -26480 39620 -26380 1 PIX1466_IN
port 1494 n
rlabel metal5 41020 -26480 41120 -26380 1 PIX1467_IN
port 1495 n
rlabel metal5 42520 -26480 42620 -26380 1 PIX1468_IN
port 1496 n
rlabel metal5 44020 -26480 44120 -26380 1 PIX1469_IN
port 1497 n
rlabel metal5 45520 -26480 45620 -26380 1 PIX1470_IN
port 1498 n
rlabel metal5 47020 -26480 47120 -26380 1 PIX1471_IN
port 1499 n
rlabel metal5 48520 -26480 48620 -26380 1 PIX1472_IN
port 1500 n
rlabel metal5 50020 -26480 50120 -26380 1 PIX1473_IN
port 1501 n
rlabel metal5 51520 -26480 51620 -26380 1 PIX1474_IN
port 1502 n
rlabel metal5 53020 -26480 53120 -26380 1 PIX1475_IN
port 1503 n
rlabel metal5 54520 -26480 54620 -26380 1 PIX1476_IN
port 1504 n
rlabel metal5 56020 -26480 56120 -26380 1 PIX1477_IN
port 1505 n
rlabel metal5 57520 -26480 57620 -26380 1 PIX1478_IN
port 1506 n
rlabel metal5 59020 -26480 59120 -26380 1 PIX1479_IN
port 1507 n
rlabel metal5 60520 -26480 60620 -26380 1 PIX1480_IN
port 1508 n
rlabel metal5 62020 -26480 62120 -26380 1 PIX1481_IN
port 1509 n
rlabel metal5 63520 -26480 63620 -26380 1 PIX1482_IN
port 1510 n
rlabel metal5 65020 -26480 65120 -26380 1 PIX1483_IN
port 1511 n
rlabel metal5 66520 -26480 66620 -26380 1 PIX1484_IN
port 1512 n
rlabel metal5 68020 -26480 68120 -26380 1 PIX1485_IN
port 1513 n
rlabel metal5 69520 -26480 69620 -26380 1 PIX1486_IN
port 1514 n
rlabel metal5 71020 -26480 71120 -26380 1 PIX1487_IN
port 1515 n
rlabel metal5 72520 -26480 72620 -26380 1 PIX1488_IN
port 1516 n
rlabel metal5 74020 -26480 74120 -26380 1 PIX1489_IN
port 1517 n
rlabel metal5 75520 -26480 75620 -26380 1 PIX1490_IN
port 1518 n
rlabel metal5 77020 -26480 77120 -26380 1 PIX1491_IN
port 1519 n
rlabel metal5 78520 -26480 78620 -26380 1 PIX1492_IN
port 1520 n
rlabel metal5 80020 -26480 80120 -26380 1 PIX1493_IN
port 1521 n
rlabel metal5 81520 -26480 81620 -26380 1 PIX1494_IN
port 1522 n
rlabel metal5 83020 -26480 83120 -26380 1 PIX1495_IN
port 1523 n
rlabel metal5 84520 -26480 84620 -26380 1 PIX1496_IN
port 1524 n
rlabel metal5 86020 -26480 86120 -26380 1 PIX1497_IN
port 1525 n
rlabel metal5 87520 -26480 87620 -26380 1 PIX1498_IN
port 1526 n
rlabel metal5 89020 -26480 89120 -26380 1 PIX1499_IN
port 1527 n
rlabel metal5 90520 -26480 90620 -26380 1 PIX1500_IN
port 1528 n
rlabel metal5 92020 -26480 92120 -26380 1 PIX1501_IN
port 1529 n
rlabel metal5 93520 -26480 93620 -26380 1 PIX1502_IN
port 1530 n
rlabel metal5 95020 -26480 95120 -26380 1 PIX1503_IN
port 1531 n
rlabel metal5 96520 -26480 96620 -26380 1 PIX1504_IN
port 1532 n
rlabel metal5 98020 -26480 98120 -26380 1 PIX1505_IN
port 1533 n
rlabel metal5 99520 -26480 99620 -26380 1 PIX1506_IN
port 1534 n
rlabel metal5 101020 -26480 101120 -26380 1 PIX1507_IN
port 1535 n
rlabel metal5 102520 -26480 102620 -26380 1 PIX1508_IN
port 1536 n
rlabel metal5 104020 -26480 104120 -26380 1 PIX1509_IN
port 1537 n
rlabel metal5 105520 -26480 105620 -26380 1 PIX1510_IN
port 1538 n
rlabel metal5 107020 -26480 107120 -26380 1 PIX1511_IN
port 1539 n
rlabel metal5 108520 -26480 108620 -26380 1 PIX1512_IN
port 1540 n
rlabel metal5 110020 -26480 110120 -26380 1 PIX1513_IN
port 1541 n
rlabel metal5 111520 -26480 111620 -26380 1 PIX1514_IN
port 1542 n
rlabel metal5 113020 -26480 113120 -26380 1 PIX1515_IN
port 1543 n
rlabel metal5 114520 -26480 114620 -26380 1 PIX1516_IN
port 1544 n
rlabel metal5 116020 -26480 116120 -26380 1 PIX1517_IN
port 1545 n
rlabel metal5 117520 -26480 117620 -26380 1 PIX1518_IN
port 1546 n
rlabel metal5 119020 -26480 119120 -26380 1 PIX1519_IN
port 1547 n
rlabel metal5 520 -27980 620 -27880 1 PIX1520_IN
port 1548 n
rlabel metal2 -1500 -27760 -1500 -27715 3 ROW_SEL19
port 1549 e
rlabel metal5 2020 -27980 2120 -27880 1 PIX1521_IN
port 1550 n
rlabel metal5 3520 -27980 3620 -27880 1 PIX1522_IN
port 1551 n
rlabel metal5 5020 -27980 5120 -27880 1 PIX1523_IN
port 1552 n
rlabel metal5 6520 -27980 6620 -27880 1 PIX1524_IN
port 1553 n
rlabel metal5 8020 -27980 8120 -27880 1 PIX1525_IN
port 1554 n
rlabel metal5 9520 -27980 9620 -27880 1 PIX1526_IN
port 1555 n
rlabel metal5 11020 -27980 11120 -27880 1 PIX1527_IN
port 1556 n
rlabel metal5 12520 -27980 12620 -27880 1 PIX1528_IN
port 1557 n
rlabel metal5 14020 -27980 14120 -27880 1 PIX1529_IN
port 1558 n
rlabel metal5 15520 -27980 15620 -27880 1 PIX1530_IN
port 1559 n
rlabel metal5 17020 -27980 17120 -27880 1 PIX1531_IN
port 1560 n
rlabel metal5 18520 -27980 18620 -27880 1 PIX1532_IN
port 1561 n
rlabel metal5 20020 -27980 20120 -27880 1 PIX1533_IN
port 1562 n
rlabel metal5 21520 -27980 21620 -27880 1 PIX1534_IN
port 1563 n
rlabel metal5 23020 -27980 23120 -27880 1 PIX1535_IN
port 1564 n
rlabel metal5 24520 -27980 24620 -27880 1 PIX1536_IN
port 1565 n
rlabel metal5 26020 -27980 26120 -27880 1 PIX1537_IN
port 1566 n
rlabel metal5 27520 -27980 27620 -27880 1 PIX1538_IN
port 1567 n
rlabel metal5 29020 -27980 29120 -27880 1 PIX1539_IN
port 1568 n
rlabel metal5 30520 -27980 30620 -27880 1 PIX1540_IN
port 1569 n
rlabel metal5 32020 -27980 32120 -27880 1 PIX1541_IN
port 1570 n
rlabel metal5 33520 -27980 33620 -27880 1 PIX1542_IN
port 1571 n
rlabel metal5 35020 -27980 35120 -27880 1 PIX1543_IN
port 1572 n
rlabel metal5 36520 -27980 36620 -27880 1 PIX1544_IN
port 1573 n
rlabel metal5 38020 -27980 38120 -27880 1 PIX1545_IN
port 1574 n
rlabel metal5 39520 -27980 39620 -27880 1 PIX1546_IN
port 1575 n
rlabel metal5 41020 -27980 41120 -27880 1 PIX1547_IN
port 1576 n
rlabel metal5 42520 -27980 42620 -27880 1 PIX1548_IN
port 1577 n
rlabel metal5 44020 -27980 44120 -27880 1 PIX1549_IN
port 1578 n
rlabel metal5 45520 -27980 45620 -27880 1 PIX1550_IN
port 1579 n
rlabel metal5 47020 -27980 47120 -27880 1 PIX1551_IN
port 1580 n
rlabel metal5 48520 -27980 48620 -27880 1 PIX1552_IN
port 1581 n
rlabel metal5 50020 -27980 50120 -27880 1 PIX1553_IN
port 1582 n
rlabel metal5 51520 -27980 51620 -27880 1 PIX1554_IN
port 1583 n
rlabel metal5 53020 -27980 53120 -27880 1 PIX1555_IN
port 1584 n
rlabel metal5 54520 -27980 54620 -27880 1 PIX1556_IN
port 1585 n
rlabel metal5 56020 -27980 56120 -27880 1 PIX1557_IN
port 1586 n
rlabel metal5 57520 -27980 57620 -27880 1 PIX1558_IN
port 1587 n
rlabel metal5 59020 -27980 59120 -27880 1 PIX1559_IN
port 1588 n
rlabel metal5 60520 -27980 60620 -27880 1 PIX1560_IN
port 1589 n
rlabel metal5 62020 -27980 62120 -27880 1 PIX1561_IN
port 1590 n
rlabel metal5 63520 -27980 63620 -27880 1 PIX1562_IN
port 1591 n
rlabel metal5 65020 -27980 65120 -27880 1 PIX1563_IN
port 1592 n
rlabel metal5 66520 -27980 66620 -27880 1 PIX1564_IN
port 1593 n
rlabel metal5 68020 -27980 68120 -27880 1 PIX1565_IN
port 1594 n
rlabel metal5 69520 -27980 69620 -27880 1 PIX1566_IN
port 1595 n
rlabel metal5 71020 -27980 71120 -27880 1 PIX1567_IN
port 1596 n
rlabel metal5 72520 -27980 72620 -27880 1 PIX1568_IN
port 1597 n
rlabel metal5 74020 -27980 74120 -27880 1 PIX1569_IN
port 1598 n
rlabel metal5 75520 -27980 75620 -27880 1 PIX1570_IN
port 1599 n
rlabel metal5 77020 -27980 77120 -27880 1 PIX1571_IN
port 1600 n
rlabel metal5 78520 -27980 78620 -27880 1 PIX1572_IN
port 1601 n
rlabel metal5 80020 -27980 80120 -27880 1 PIX1573_IN
port 1602 n
rlabel metal5 81520 -27980 81620 -27880 1 PIX1574_IN
port 1603 n
rlabel metal5 83020 -27980 83120 -27880 1 PIX1575_IN
port 1604 n
rlabel metal5 84520 -27980 84620 -27880 1 PIX1576_IN
port 1605 n
rlabel metal5 86020 -27980 86120 -27880 1 PIX1577_IN
port 1606 n
rlabel metal5 87520 -27980 87620 -27880 1 PIX1578_IN
port 1607 n
rlabel metal5 89020 -27980 89120 -27880 1 PIX1579_IN
port 1608 n
rlabel metal5 90520 -27980 90620 -27880 1 PIX1580_IN
port 1609 n
rlabel metal5 92020 -27980 92120 -27880 1 PIX1581_IN
port 1610 n
rlabel metal5 93520 -27980 93620 -27880 1 PIX1582_IN
port 1611 n
rlabel metal5 95020 -27980 95120 -27880 1 PIX1583_IN
port 1612 n
rlabel metal5 96520 -27980 96620 -27880 1 PIX1584_IN
port 1613 n
rlabel metal5 98020 -27980 98120 -27880 1 PIX1585_IN
port 1614 n
rlabel metal5 99520 -27980 99620 -27880 1 PIX1586_IN
port 1615 n
rlabel metal5 101020 -27980 101120 -27880 1 PIX1587_IN
port 1616 n
rlabel metal5 102520 -27980 102620 -27880 1 PIX1588_IN
port 1617 n
rlabel metal5 104020 -27980 104120 -27880 1 PIX1589_IN
port 1618 n
rlabel metal5 105520 -27980 105620 -27880 1 PIX1590_IN
port 1619 n
rlabel metal5 107020 -27980 107120 -27880 1 PIX1591_IN
port 1620 n
rlabel metal5 108520 -27980 108620 -27880 1 PIX1592_IN
port 1621 n
rlabel metal5 110020 -27980 110120 -27880 1 PIX1593_IN
port 1622 n
rlabel metal5 111520 -27980 111620 -27880 1 PIX1594_IN
port 1623 n
rlabel metal5 113020 -27980 113120 -27880 1 PIX1595_IN
port 1624 n
rlabel metal5 114520 -27980 114620 -27880 1 PIX1596_IN
port 1625 n
rlabel metal5 116020 -27980 116120 -27880 1 PIX1597_IN
port 1626 n
rlabel metal5 117520 -27980 117620 -27880 1 PIX1598_IN
port 1627 n
rlabel metal5 119020 -27980 119120 -27880 1 PIX1599_IN
port 1628 n
rlabel metal5 520 -29480 620 -29380 1 PIX1600_IN
port 1629 n
rlabel metal2 -1500 -29260 -1500 -29215 3 ROW_SEL20
port 1630 e
rlabel metal5 2020 -29480 2120 -29380 1 PIX1601_IN
port 1631 n
rlabel metal5 3520 -29480 3620 -29380 1 PIX1602_IN
port 1632 n
rlabel metal5 5020 -29480 5120 -29380 1 PIX1603_IN
port 1633 n
rlabel metal5 6520 -29480 6620 -29380 1 PIX1604_IN
port 1634 n
rlabel metal5 8020 -29480 8120 -29380 1 PIX1605_IN
port 1635 n
rlabel metal5 9520 -29480 9620 -29380 1 PIX1606_IN
port 1636 n
rlabel metal5 11020 -29480 11120 -29380 1 PIX1607_IN
port 1637 n
rlabel metal5 12520 -29480 12620 -29380 1 PIX1608_IN
port 1638 n
rlabel metal5 14020 -29480 14120 -29380 1 PIX1609_IN
port 1639 n
rlabel metal5 15520 -29480 15620 -29380 1 PIX1610_IN
port 1640 n
rlabel metal5 17020 -29480 17120 -29380 1 PIX1611_IN
port 1641 n
rlabel metal5 18520 -29480 18620 -29380 1 PIX1612_IN
port 1642 n
rlabel metal5 20020 -29480 20120 -29380 1 PIX1613_IN
port 1643 n
rlabel metal5 21520 -29480 21620 -29380 1 PIX1614_IN
port 1644 n
rlabel metal5 23020 -29480 23120 -29380 1 PIX1615_IN
port 1645 n
rlabel metal5 24520 -29480 24620 -29380 1 PIX1616_IN
port 1646 n
rlabel metal5 26020 -29480 26120 -29380 1 PIX1617_IN
port 1647 n
rlabel metal5 27520 -29480 27620 -29380 1 PIX1618_IN
port 1648 n
rlabel metal5 29020 -29480 29120 -29380 1 PIX1619_IN
port 1649 n
rlabel metal5 30520 -29480 30620 -29380 1 PIX1620_IN
port 1650 n
rlabel metal5 32020 -29480 32120 -29380 1 PIX1621_IN
port 1651 n
rlabel metal5 33520 -29480 33620 -29380 1 PIX1622_IN
port 1652 n
rlabel metal5 35020 -29480 35120 -29380 1 PIX1623_IN
port 1653 n
rlabel metal5 36520 -29480 36620 -29380 1 PIX1624_IN
port 1654 n
rlabel metal5 38020 -29480 38120 -29380 1 PIX1625_IN
port 1655 n
rlabel metal5 39520 -29480 39620 -29380 1 PIX1626_IN
port 1656 n
rlabel metal5 41020 -29480 41120 -29380 1 PIX1627_IN
port 1657 n
rlabel metal5 42520 -29480 42620 -29380 1 PIX1628_IN
port 1658 n
rlabel metal5 44020 -29480 44120 -29380 1 PIX1629_IN
port 1659 n
rlabel metal5 45520 -29480 45620 -29380 1 PIX1630_IN
port 1660 n
rlabel metal5 47020 -29480 47120 -29380 1 PIX1631_IN
port 1661 n
rlabel metal5 48520 -29480 48620 -29380 1 PIX1632_IN
port 1662 n
rlabel metal5 50020 -29480 50120 -29380 1 PIX1633_IN
port 1663 n
rlabel metal5 51520 -29480 51620 -29380 1 PIX1634_IN
port 1664 n
rlabel metal5 53020 -29480 53120 -29380 1 PIX1635_IN
port 1665 n
rlabel metal5 54520 -29480 54620 -29380 1 PIX1636_IN
port 1666 n
rlabel metal5 56020 -29480 56120 -29380 1 PIX1637_IN
port 1667 n
rlabel metal5 57520 -29480 57620 -29380 1 PIX1638_IN
port 1668 n
rlabel metal5 59020 -29480 59120 -29380 1 PIX1639_IN
port 1669 n
rlabel metal5 60520 -29480 60620 -29380 1 PIX1640_IN
port 1670 n
rlabel metal5 62020 -29480 62120 -29380 1 PIX1641_IN
port 1671 n
rlabel metal5 63520 -29480 63620 -29380 1 PIX1642_IN
port 1672 n
rlabel metal5 65020 -29480 65120 -29380 1 PIX1643_IN
port 1673 n
rlabel metal5 66520 -29480 66620 -29380 1 PIX1644_IN
port 1674 n
rlabel metal5 68020 -29480 68120 -29380 1 PIX1645_IN
port 1675 n
rlabel metal5 69520 -29480 69620 -29380 1 PIX1646_IN
port 1676 n
rlabel metal5 71020 -29480 71120 -29380 1 PIX1647_IN
port 1677 n
rlabel metal5 72520 -29480 72620 -29380 1 PIX1648_IN
port 1678 n
rlabel metal5 74020 -29480 74120 -29380 1 PIX1649_IN
port 1679 n
rlabel metal5 75520 -29480 75620 -29380 1 PIX1650_IN
port 1680 n
rlabel metal5 77020 -29480 77120 -29380 1 PIX1651_IN
port 1681 n
rlabel metal5 78520 -29480 78620 -29380 1 PIX1652_IN
port 1682 n
rlabel metal5 80020 -29480 80120 -29380 1 PIX1653_IN
port 1683 n
rlabel metal5 81520 -29480 81620 -29380 1 PIX1654_IN
port 1684 n
rlabel metal5 83020 -29480 83120 -29380 1 PIX1655_IN
port 1685 n
rlabel metal5 84520 -29480 84620 -29380 1 PIX1656_IN
port 1686 n
rlabel metal5 86020 -29480 86120 -29380 1 PIX1657_IN
port 1687 n
rlabel metal5 87520 -29480 87620 -29380 1 PIX1658_IN
port 1688 n
rlabel metal5 89020 -29480 89120 -29380 1 PIX1659_IN
port 1689 n
rlabel metal5 90520 -29480 90620 -29380 1 PIX1660_IN
port 1690 n
rlabel metal5 92020 -29480 92120 -29380 1 PIX1661_IN
port 1691 n
rlabel metal5 93520 -29480 93620 -29380 1 PIX1662_IN
port 1692 n
rlabel metal5 95020 -29480 95120 -29380 1 PIX1663_IN
port 1693 n
rlabel metal5 96520 -29480 96620 -29380 1 PIX1664_IN
port 1694 n
rlabel metal5 98020 -29480 98120 -29380 1 PIX1665_IN
port 1695 n
rlabel metal5 99520 -29480 99620 -29380 1 PIX1666_IN
port 1696 n
rlabel metal5 101020 -29480 101120 -29380 1 PIX1667_IN
port 1697 n
rlabel metal5 102520 -29480 102620 -29380 1 PIX1668_IN
port 1698 n
rlabel metal5 104020 -29480 104120 -29380 1 PIX1669_IN
port 1699 n
rlabel metal5 105520 -29480 105620 -29380 1 PIX1670_IN
port 1700 n
rlabel metal5 107020 -29480 107120 -29380 1 PIX1671_IN
port 1701 n
rlabel metal5 108520 -29480 108620 -29380 1 PIX1672_IN
port 1702 n
rlabel metal5 110020 -29480 110120 -29380 1 PIX1673_IN
port 1703 n
rlabel metal5 111520 -29480 111620 -29380 1 PIX1674_IN
port 1704 n
rlabel metal5 113020 -29480 113120 -29380 1 PIX1675_IN
port 1705 n
rlabel metal5 114520 -29480 114620 -29380 1 PIX1676_IN
port 1706 n
rlabel metal5 116020 -29480 116120 -29380 1 PIX1677_IN
port 1707 n
rlabel metal5 117520 -29480 117620 -29380 1 PIX1678_IN
port 1708 n
rlabel metal5 119020 -29480 119120 -29380 1 PIX1679_IN
port 1709 n
rlabel metal5 520 -30980 620 -30880 1 PIX1680_IN
port 1710 n
rlabel metal2 -1500 -30760 -1500 -30715 3 ROW_SEL21
port 1711 e
rlabel metal5 2020 -30980 2120 -30880 1 PIX1681_IN
port 1712 n
rlabel metal5 3520 -30980 3620 -30880 1 PIX1682_IN
port 1713 n
rlabel metal5 5020 -30980 5120 -30880 1 PIX1683_IN
port 1714 n
rlabel metal5 6520 -30980 6620 -30880 1 PIX1684_IN
port 1715 n
rlabel metal5 8020 -30980 8120 -30880 1 PIX1685_IN
port 1716 n
rlabel metal5 9520 -30980 9620 -30880 1 PIX1686_IN
port 1717 n
rlabel metal5 11020 -30980 11120 -30880 1 PIX1687_IN
port 1718 n
rlabel metal5 12520 -30980 12620 -30880 1 PIX1688_IN
port 1719 n
rlabel metal5 14020 -30980 14120 -30880 1 PIX1689_IN
port 1720 n
rlabel metal5 15520 -30980 15620 -30880 1 PIX1690_IN
port 1721 n
rlabel metal5 17020 -30980 17120 -30880 1 PIX1691_IN
port 1722 n
rlabel metal5 18520 -30980 18620 -30880 1 PIX1692_IN
port 1723 n
rlabel metal5 20020 -30980 20120 -30880 1 PIX1693_IN
port 1724 n
rlabel metal5 21520 -30980 21620 -30880 1 PIX1694_IN
port 1725 n
rlabel metal5 23020 -30980 23120 -30880 1 PIX1695_IN
port 1726 n
rlabel metal5 24520 -30980 24620 -30880 1 PIX1696_IN
port 1727 n
rlabel metal5 26020 -30980 26120 -30880 1 PIX1697_IN
port 1728 n
rlabel metal5 27520 -30980 27620 -30880 1 PIX1698_IN
port 1729 n
rlabel metal5 29020 -30980 29120 -30880 1 PIX1699_IN
port 1730 n
rlabel metal5 30520 -30980 30620 -30880 1 PIX1700_IN
port 1731 n
rlabel metal5 32020 -30980 32120 -30880 1 PIX1701_IN
port 1732 n
rlabel metal5 33520 -30980 33620 -30880 1 PIX1702_IN
port 1733 n
rlabel metal5 35020 -30980 35120 -30880 1 PIX1703_IN
port 1734 n
rlabel metal5 36520 -30980 36620 -30880 1 PIX1704_IN
port 1735 n
rlabel metal5 38020 -30980 38120 -30880 1 PIX1705_IN
port 1736 n
rlabel metal5 39520 -30980 39620 -30880 1 PIX1706_IN
port 1737 n
rlabel metal5 41020 -30980 41120 -30880 1 PIX1707_IN
port 1738 n
rlabel metal5 42520 -30980 42620 -30880 1 PIX1708_IN
port 1739 n
rlabel metal5 44020 -30980 44120 -30880 1 PIX1709_IN
port 1740 n
rlabel metal5 45520 -30980 45620 -30880 1 PIX1710_IN
port 1741 n
rlabel metal5 47020 -30980 47120 -30880 1 PIX1711_IN
port 1742 n
rlabel metal5 48520 -30980 48620 -30880 1 PIX1712_IN
port 1743 n
rlabel metal5 50020 -30980 50120 -30880 1 PIX1713_IN
port 1744 n
rlabel metal5 51520 -30980 51620 -30880 1 PIX1714_IN
port 1745 n
rlabel metal5 53020 -30980 53120 -30880 1 PIX1715_IN
port 1746 n
rlabel metal5 54520 -30980 54620 -30880 1 PIX1716_IN
port 1747 n
rlabel metal5 56020 -30980 56120 -30880 1 PIX1717_IN
port 1748 n
rlabel metal5 57520 -30980 57620 -30880 1 PIX1718_IN
port 1749 n
rlabel metal5 59020 -30980 59120 -30880 1 PIX1719_IN
port 1750 n
rlabel metal5 60520 -30980 60620 -30880 1 PIX1720_IN
port 1751 n
rlabel metal5 62020 -30980 62120 -30880 1 PIX1721_IN
port 1752 n
rlabel metal5 63520 -30980 63620 -30880 1 PIX1722_IN
port 1753 n
rlabel metal5 65020 -30980 65120 -30880 1 PIX1723_IN
port 1754 n
rlabel metal5 66520 -30980 66620 -30880 1 PIX1724_IN
port 1755 n
rlabel metal5 68020 -30980 68120 -30880 1 PIX1725_IN
port 1756 n
rlabel metal5 69520 -30980 69620 -30880 1 PIX1726_IN
port 1757 n
rlabel metal5 71020 -30980 71120 -30880 1 PIX1727_IN
port 1758 n
rlabel metal5 72520 -30980 72620 -30880 1 PIX1728_IN
port 1759 n
rlabel metal5 74020 -30980 74120 -30880 1 PIX1729_IN
port 1760 n
rlabel metal5 75520 -30980 75620 -30880 1 PIX1730_IN
port 1761 n
rlabel metal5 77020 -30980 77120 -30880 1 PIX1731_IN
port 1762 n
rlabel metal5 78520 -30980 78620 -30880 1 PIX1732_IN
port 1763 n
rlabel metal5 80020 -30980 80120 -30880 1 PIX1733_IN
port 1764 n
rlabel metal5 81520 -30980 81620 -30880 1 PIX1734_IN
port 1765 n
rlabel metal5 83020 -30980 83120 -30880 1 PIX1735_IN
port 1766 n
rlabel metal5 84520 -30980 84620 -30880 1 PIX1736_IN
port 1767 n
rlabel metal5 86020 -30980 86120 -30880 1 PIX1737_IN
port 1768 n
rlabel metal5 87520 -30980 87620 -30880 1 PIX1738_IN
port 1769 n
rlabel metal5 89020 -30980 89120 -30880 1 PIX1739_IN
port 1770 n
rlabel metal5 90520 -30980 90620 -30880 1 PIX1740_IN
port 1771 n
rlabel metal5 92020 -30980 92120 -30880 1 PIX1741_IN
port 1772 n
rlabel metal5 93520 -30980 93620 -30880 1 PIX1742_IN
port 1773 n
rlabel metal5 95020 -30980 95120 -30880 1 PIX1743_IN
port 1774 n
rlabel metal5 96520 -30980 96620 -30880 1 PIX1744_IN
port 1775 n
rlabel metal5 98020 -30980 98120 -30880 1 PIX1745_IN
port 1776 n
rlabel metal5 99520 -30980 99620 -30880 1 PIX1746_IN
port 1777 n
rlabel metal5 101020 -30980 101120 -30880 1 PIX1747_IN
port 1778 n
rlabel metal5 102520 -30980 102620 -30880 1 PIX1748_IN
port 1779 n
rlabel metal5 104020 -30980 104120 -30880 1 PIX1749_IN
port 1780 n
rlabel metal5 105520 -30980 105620 -30880 1 PIX1750_IN
port 1781 n
rlabel metal5 107020 -30980 107120 -30880 1 PIX1751_IN
port 1782 n
rlabel metal5 108520 -30980 108620 -30880 1 PIX1752_IN
port 1783 n
rlabel metal5 110020 -30980 110120 -30880 1 PIX1753_IN
port 1784 n
rlabel metal5 111520 -30980 111620 -30880 1 PIX1754_IN
port 1785 n
rlabel metal5 113020 -30980 113120 -30880 1 PIX1755_IN
port 1786 n
rlabel metal5 114520 -30980 114620 -30880 1 PIX1756_IN
port 1787 n
rlabel metal5 116020 -30980 116120 -30880 1 PIX1757_IN
port 1788 n
rlabel metal5 117520 -30980 117620 -30880 1 PIX1758_IN
port 1789 n
rlabel metal5 119020 -30980 119120 -30880 1 PIX1759_IN
port 1790 n
rlabel metal5 520 -32480 620 -32380 1 PIX1760_IN
port 1791 n
rlabel metal2 -1500 -32260 -1500 -32215 3 ROW_SEL22
port 1792 e
rlabel metal5 2020 -32480 2120 -32380 1 PIX1761_IN
port 1793 n
rlabel metal5 3520 -32480 3620 -32380 1 PIX1762_IN
port 1794 n
rlabel metal5 5020 -32480 5120 -32380 1 PIX1763_IN
port 1795 n
rlabel metal5 6520 -32480 6620 -32380 1 PIX1764_IN
port 1796 n
rlabel metal5 8020 -32480 8120 -32380 1 PIX1765_IN
port 1797 n
rlabel metal5 9520 -32480 9620 -32380 1 PIX1766_IN
port 1798 n
rlabel metal5 11020 -32480 11120 -32380 1 PIX1767_IN
port 1799 n
rlabel metal5 12520 -32480 12620 -32380 1 PIX1768_IN
port 1800 n
rlabel metal5 14020 -32480 14120 -32380 1 PIX1769_IN
port 1801 n
rlabel metal5 15520 -32480 15620 -32380 1 PIX1770_IN
port 1802 n
rlabel metal5 17020 -32480 17120 -32380 1 PIX1771_IN
port 1803 n
rlabel metal5 18520 -32480 18620 -32380 1 PIX1772_IN
port 1804 n
rlabel metal5 20020 -32480 20120 -32380 1 PIX1773_IN
port 1805 n
rlabel metal5 21520 -32480 21620 -32380 1 PIX1774_IN
port 1806 n
rlabel metal5 23020 -32480 23120 -32380 1 PIX1775_IN
port 1807 n
rlabel metal5 24520 -32480 24620 -32380 1 PIX1776_IN
port 1808 n
rlabel metal5 26020 -32480 26120 -32380 1 PIX1777_IN
port 1809 n
rlabel metal5 27520 -32480 27620 -32380 1 PIX1778_IN
port 1810 n
rlabel metal5 29020 -32480 29120 -32380 1 PIX1779_IN
port 1811 n
rlabel metal5 30520 -32480 30620 -32380 1 PIX1780_IN
port 1812 n
rlabel metal5 32020 -32480 32120 -32380 1 PIX1781_IN
port 1813 n
rlabel metal5 33520 -32480 33620 -32380 1 PIX1782_IN
port 1814 n
rlabel metal5 35020 -32480 35120 -32380 1 PIX1783_IN
port 1815 n
rlabel metal5 36520 -32480 36620 -32380 1 PIX1784_IN
port 1816 n
rlabel metal5 38020 -32480 38120 -32380 1 PIX1785_IN
port 1817 n
rlabel metal5 39520 -32480 39620 -32380 1 PIX1786_IN
port 1818 n
rlabel metal5 41020 -32480 41120 -32380 1 PIX1787_IN
port 1819 n
rlabel metal5 42520 -32480 42620 -32380 1 PIX1788_IN
port 1820 n
rlabel metal5 44020 -32480 44120 -32380 1 PIX1789_IN
port 1821 n
rlabel metal5 45520 -32480 45620 -32380 1 PIX1790_IN
port 1822 n
rlabel metal5 47020 -32480 47120 -32380 1 PIX1791_IN
port 1823 n
rlabel metal5 48520 -32480 48620 -32380 1 PIX1792_IN
port 1824 n
rlabel metal5 50020 -32480 50120 -32380 1 PIX1793_IN
port 1825 n
rlabel metal5 51520 -32480 51620 -32380 1 PIX1794_IN
port 1826 n
rlabel metal5 53020 -32480 53120 -32380 1 PIX1795_IN
port 1827 n
rlabel metal5 54520 -32480 54620 -32380 1 PIX1796_IN
port 1828 n
rlabel metal5 56020 -32480 56120 -32380 1 PIX1797_IN
port 1829 n
rlabel metal5 57520 -32480 57620 -32380 1 PIX1798_IN
port 1830 n
rlabel metal5 59020 -32480 59120 -32380 1 PIX1799_IN
port 1831 n
rlabel metal5 60520 -32480 60620 -32380 1 PIX1800_IN
port 1832 n
rlabel metal5 62020 -32480 62120 -32380 1 PIX1801_IN
port 1833 n
rlabel metal5 63520 -32480 63620 -32380 1 PIX1802_IN
port 1834 n
rlabel metal5 65020 -32480 65120 -32380 1 PIX1803_IN
port 1835 n
rlabel metal5 66520 -32480 66620 -32380 1 PIX1804_IN
port 1836 n
rlabel metal5 68020 -32480 68120 -32380 1 PIX1805_IN
port 1837 n
rlabel metal5 69520 -32480 69620 -32380 1 PIX1806_IN
port 1838 n
rlabel metal5 71020 -32480 71120 -32380 1 PIX1807_IN
port 1839 n
rlabel metal5 72520 -32480 72620 -32380 1 PIX1808_IN
port 1840 n
rlabel metal5 74020 -32480 74120 -32380 1 PIX1809_IN
port 1841 n
rlabel metal5 75520 -32480 75620 -32380 1 PIX1810_IN
port 1842 n
rlabel metal5 77020 -32480 77120 -32380 1 PIX1811_IN
port 1843 n
rlabel metal5 78520 -32480 78620 -32380 1 PIX1812_IN
port 1844 n
rlabel metal5 80020 -32480 80120 -32380 1 PIX1813_IN
port 1845 n
rlabel metal5 81520 -32480 81620 -32380 1 PIX1814_IN
port 1846 n
rlabel metal5 83020 -32480 83120 -32380 1 PIX1815_IN
port 1847 n
rlabel metal5 84520 -32480 84620 -32380 1 PIX1816_IN
port 1848 n
rlabel metal5 86020 -32480 86120 -32380 1 PIX1817_IN
port 1849 n
rlabel metal5 87520 -32480 87620 -32380 1 PIX1818_IN
port 1850 n
rlabel metal5 89020 -32480 89120 -32380 1 PIX1819_IN
port 1851 n
rlabel metal5 90520 -32480 90620 -32380 1 PIX1820_IN
port 1852 n
rlabel metal5 92020 -32480 92120 -32380 1 PIX1821_IN
port 1853 n
rlabel metal5 93520 -32480 93620 -32380 1 PIX1822_IN
port 1854 n
rlabel metal5 95020 -32480 95120 -32380 1 PIX1823_IN
port 1855 n
rlabel metal5 96520 -32480 96620 -32380 1 PIX1824_IN
port 1856 n
rlabel metal5 98020 -32480 98120 -32380 1 PIX1825_IN
port 1857 n
rlabel metal5 99520 -32480 99620 -32380 1 PIX1826_IN
port 1858 n
rlabel metal5 101020 -32480 101120 -32380 1 PIX1827_IN
port 1859 n
rlabel metal5 102520 -32480 102620 -32380 1 PIX1828_IN
port 1860 n
rlabel metal5 104020 -32480 104120 -32380 1 PIX1829_IN
port 1861 n
rlabel metal5 105520 -32480 105620 -32380 1 PIX1830_IN
port 1862 n
rlabel metal5 107020 -32480 107120 -32380 1 PIX1831_IN
port 1863 n
rlabel metal5 108520 -32480 108620 -32380 1 PIX1832_IN
port 1864 n
rlabel metal5 110020 -32480 110120 -32380 1 PIX1833_IN
port 1865 n
rlabel metal5 111520 -32480 111620 -32380 1 PIX1834_IN
port 1866 n
rlabel metal5 113020 -32480 113120 -32380 1 PIX1835_IN
port 1867 n
rlabel metal5 114520 -32480 114620 -32380 1 PIX1836_IN
port 1868 n
rlabel metal5 116020 -32480 116120 -32380 1 PIX1837_IN
port 1869 n
rlabel metal5 117520 -32480 117620 -32380 1 PIX1838_IN
port 1870 n
rlabel metal5 119020 -32480 119120 -32380 1 PIX1839_IN
port 1871 n
rlabel metal5 520 -33980 620 -33880 1 PIX1840_IN
port 1872 n
rlabel metal2 -1500 -33760 -1500 -33715 3 ROW_SEL23
port 1873 e
rlabel metal5 2020 -33980 2120 -33880 1 PIX1841_IN
port 1874 n
rlabel metal5 3520 -33980 3620 -33880 1 PIX1842_IN
port 1875 n
rlabel metal5 5020 -33980 5120 -33880 1 PIX1843_IN
port 1876 n
rlabel metal5 6520 -33980 6620 -33880 1 PIX1844_IN
port 1877 n
rlabel metal5 8020 -33980 8120 -33880 1 PIX1845_IN
port 1878 n
rlabel metal5 9520 -33980 9620 -33880 1 PIX1846_IN
port 1879 n
rlabel metal5 11020 -33980 11120 -33880 1 PIX1847_IN
port 1880 n
rlabel metal5 12520 -33980 12620 -33880 1 PIX1848_IN
port 1881 n
rlabel metal5 14020 -33980 14120 -33880 1 PIX1849_IN
port 1882 n
rlabel metal5 15520 -33980 15620 -33880 1 PIX1850_IN
port 1883 n
rlabel metal5 17020 -33980 17120 -33880 1 PIX1851_IN
port 1884 n
rlabel metal5 18520 -33980 18620 -33880 1 PIX1852_IN
port 1885 n
rlabel metal5 20020 -33980 20120 -33880 1 PIX1853_IN
port 1886 n
rlabel metal5 21520 -33980 21620 -33880 1 PIX1854_IN
port 1887 n
rlabel metal5 23020 -33980 23120 -33880 1 PIX1855_IN
port 1888 n
rlabel metal5 24520 -33980 24620 -33880 1 PIX1856_IN
port 1889 n
rlabel metal5 26020 -33980 26120 -33880 1 PIX1857_IN
port 1890 n
rlabel metal5 27520 -33980 27620 -33880 1 PIX1858_IN
port 1891 n
rlabel metal5 29020 -33980 29120 -33880 1 PIX1859_IN
port 1892 n
rlabel metal5 30520 -33980 30620 -33880 1 PIX1860_IN
port 1893 n
rlabel metal5 32020 -33980 32120 -33880 1 PIX1861_IN
port 1894 n
rlabel metal5 33520 -33980 33620 -33880 1 PIX1862_IN
port 1895 n
rlabel metal5 35020 -33980 35120 -33880 1 PIX1863_IN
port 1896 n
rlabel metal5 36520 -33980 36620 -33880 1 PIX1864_IN
port 1897 n
rlabel metal5 38020 -33980 38120 -33880 1 PIX1865_IN
port 1898 n
rlabel metal5 39520 -33980 39620 -33880 1 PIX1866_IN
port 1899 n
rlabel metal5 41020 -33980 41120 -33880 1 PIX1867_IN
port 1900 n
rlabel metal5 42520 -33980 42620 -33880 1 PIX1868_IN
port 1901 n
rlabel metal5 44020 -33980 44120 -33880 1 PIX1869_IN
port 1902 n
rlabel metal5 45520 -33980 45620 -33880 1 PIX1870_IN
port 1903 n
rlabel metal5 47020 -33980 47120 -33880 1 PIX1871_IN
port 1904 n
rlabel metal5 48520 -33980 48620 -33880 1 PIX1872_IN
port 1905 n
rlabel metal5 50020 -33980 50120 -33880 1 PIX1873_IN
port 1906 n
rlabel metal5 51520 -33980 51620 -33880 1 PIX1874_IN
port 1907 n
rlabel metal5 53020 -33980 53120 -33880 1 PIX1875_IN
port 1908 n
rlabel metal5 54520 -33980 54620 -33880 1 PIX1876_IN
port 1909 n
rlabel metal5 56020 -33980 56120 -33880 1 PIX1877_IN
port 1910 n
rlabel metal5 57520 -33980 57620 -33880 1 PIX1878_IN
port 1911 n
rlabel metal5 59020 -33980 59120 -33880 1 PIX1879_IN
port 1912 n
rlabel metal5 60520 -33980 60620 -33880 1 PIX1880_IN
port 1913 n
rlabel metal5 62020 -33980 62120 -33880 1 PIX1881_IN
port 1914 n
rlabel metal5 63520 -33980 63620 -33880 1 PIX1882_IN
port 1915 n
rlabel metal5 65020 -33980 65120 -33880 1 PIX1883_IN
port 1916 n
rlabel metal5 66520 -33980 66620 -33880 1 PIX1884_IN
port 1917 n
rlabel metal5 68020 -33980 68120 -33880 1 PIX1885_IN
port 1918 n
rlabel metal5 69520 -33980 69620 -33880 1 PIX1886_IN
port 1919 n
rlabel metal5 71020 -33980 71120 -33880 1 PIX1887_IN
port 1920 n
rlabel metal5 72520 -33980 72620 -33880 1 PIX1888_IN
port 1921 n
rlabel metal5 74020 -33980 74120 -33880 1 PIX1889_IN
port 1922 n
rlabel metal5 75520 -33980 75620 -33880 1 PIX1890_IN
port 1923 n
rlabel metal5 77020 -33980 77120 -33880 1 PIX1891_IN
port 1924 n
rlabel metal5 78520 -33980 78620 -33880 1 PIX1892_IN
port 1925 n
rlabel metal5 80020 -33980 80120 -33880 1 PIX1893_IN
port 1926 n
rlabel metal5 81520 -33980 81620 -33880 1 PIX1894_IN
port 1927 n
rlabel metal5 83020 -33980 83120 -33880 1 PIX1895_IN
port 1928 n
rlabel metal5 84520 -33980 84620 -33880 1 PIX1896_IN
port 1929 n
rlabel metal5 86020 -33980 86120 -33880 1 PIX1897_IN
port 1930 n
rlabel metal5 87520 -33980 87620 -33880 1 PIX1898_IN
port 1931 n
rlabel metal5 89020 -33980 89120 -33880 1 PIX1899_IN
port 1932 n
rlabel metal5 90520 -33980 90620 -33880 1 PIX1900_IN
port 1933 n
rlabel metal5 92020 -33980 92120 -33880 1 PIX1901_IN
port 1934 n
rlabel metal5 93520 -33980 93620 -33880 1 PIX1902_IN
port 1935 n
rlabel metal5 95020 -33980 95120 -33880 1 PIX1903_IN
port 1936 n
rlabel metal5 96520 -33980 96620 -33880 1 PIX1904_IN
port 1937 n
rlabel metal5 98020 -33980 98120 -33880 1 PIX1905_IN
port 1938 n
rlabel metal5 99520 -33980 99620 -33880 1 PIX1906_IN
port 1939 n
rlabel metal5 101020 -33980 101120 -33880 1 PIX1907_IN
port 1940 n
rlabel metal5 102520 -33980 102620 -33880 1 PIX1908_IN
port 1941 n
rlabel metal5 104020 -33980 104120 -33880 1 PIX1909_IN
port 1942 n
rlabel metal5 105520 -33980 105620 -33880 1 PIX1910_IN
port 1943 n
rlabel metal5 107020 -33980 107120 -33880 1 PIX1911_IN
port 1944 n
rlabel metal5 108520 -33980 108620 -33880 1 PIX1912_IN
port 1945 n
rlabel metal5 110020 -33980 110120 -33880 1 PIX1913_IN
port 1946 n
rlabel metal5 111520 -33980 111620 -33880 1 PIX1914_IN
port 1947 n
rlabel metal5 113020 -33980 113120 -33880 1 PIX1915_IN
port 1948 n
rlabel metal5 114520 -33980 114620 -33880 1 PIX1916_IN
port 1949 n
rlabel metal5 116020 -33980 116120 -33880 1 PIX1917_IN
port 1950 n
rlabel metal5 117520 -33980 117620 -33880 1 PIX1918_IN
port 1951 n
rlabel metal5 119020 -33980 119120 -33880 1 PIX1919_IN
port 1952 n
rlabel metal5 520 -35480 620 -35380 1 PIX1920_IN
port 1953 n
rlabel metal2 -1500 -35260 -1500 -35215 3 ROW_SEL24
port 1954 e
rlabel metal5 2020 -35480 2120 -35380 1 PIX1921_IN
port 1955 n
rlabel metal5 3520 -35480 3620 -35380 1 PIX1922_IN
port 1956 n
rlabel metal5 5020 -35480 5120 -35380 1 PIX1923_IN
port 1957 n
rlabel metal5 6520 -35480 6620 -35380 1 PIX1924_IN
port 1958 n
rlabel metal5 8020 -35480 8120 -35380 1 PIX1925_IN
port 1959 n
rlabel metal5 9520 -35480 9620 -35380 1 PIX1926_IN
port 1960 n
rlabel metal5 11020 -35480 11120 -35380 1 PIX1927_IN
port 1961 n
rlabel metal5 12520 -35480 12620 -35380 1 PIX1928_IN
port 1962 n
rlabel metal5 14020 -35480 14120 -35380 1 PIX1929_IN
port 1963 n
rlabel metal5 15520 -35480 15620 -35380 1 PIX1930_IN
port 1964 n
rlabel metal5 17020 -35480 17120 -35380 1 PIX1931_IN
port 1965 n
rlabel metal5 18520 -35480 18620 -35380 1 PIX1932_IN
port 1966 n
rlabel metal5 20020 -35480 20120 -35380 1 PIX1933_IN
port 1967 n
rlabel metal5 21520 -35480 21620 -35380 1 PIX1934_IN
port 1968 n
rlabel metal5 23020 -35480 23120 -35380 1 PIX1935_IN
port 1969 n
rlabel metal5 24520 -35480 24620 -35380 1 PIX1936_IN
port 1970 n
rlabel metal5 26020 -35480 26120 -35380 1 PIX1937_IN
port 1971 n
rlabel metal5 27520 -35480 27620 -35380 1 PIX1938_IN
port 1972 n
rlabel metal5 29020 -35480 29120 -35380 1 PIX1939_IN
port 1973 n
rlabel metal5 30520 -35480 30620 -35380 1 PIX1940_IN
port 1974 n
rlabel metal5 32020 -35480 32120 -35380 1 PIX1941_IN
port 1975 n
rlabel metal5 33520 -35480 33620 -35380 1 PIX1942_IN
port 1976 n
rlabel metal5 35020 -35480 35120 -35380 1 PIX1943_IN
port 1977 n
rlabel metal5 36520 -35480 36620 -35380 1 PIX1944_IN
port 1978 n
rlabel metal5 38020 -35480 38120 -35380 1 PIX1945_IN
port 1979 n
rlabel metal5 39520 -35480 39620 -35380 1 PIX1946_IN
port 1980 n
rlabel metal5 41020 -35480 41120 -35380 1 PIX1947_IN
port 1981 n
rlabel metal5 42520 -35480 42620 -35380 1 PIX1948_IN
port 1982 n
rlabel metal5 44020 -35480 44120 -35380 1 PIX1949_IN
port 1983 n
rlabel metal5 45520 -35480 45620 -35380 1 PIX1950_IN
port 1984 n
rlabel metal5 47020 -35480 47120 -35380 1 PIX1951_IN
port 1985 n
rlabel metal5 48520 -35480 48620 -35380 1 PIX1952_IN
port 1986 n
rlabel metal5 50020 -35480 50120 -35380 1 PIX1953_IN
port 1987 n
rlabel metal5 51520 -35480 51620 -35380 1 PIX1954_IN
port 1988 n
rlabel metal5 53020 -35480 53120 -35380 1 PIX1955_IN
port 1989 n
rlabel metal5 54520 -35480 54620 -35380 1 PIX1956_IN
port 1990 n
rlabel metal5 56020 -35480 56120 -35380 1 PIX1957_IN
port 1991 n
rlabel metal5 57520 -35480 57620 -35380 1 PIX1958_IN
port 1992 n
rlabel metal5 59020 -35480 59120 -35380 1 PIX1959_IN
port 1993 n
rlabel metal5 60520 -35480 60620 -35380 1 PIX1960_IN
port 1994 n
rlabel metal5 62020 -35480 62120 -35380 1 PIX1961_IN
port 1995 n
rlabel metal5 63520 -35480 63620 -35380 1 PIX1962_IN
port 1996 n
rlabel metal5 65020 -35480 65120 -35380 1 PIX1963_IN
port 1997 n
rlabel metal5 66520 -35480 66620 -35380 1 PIX1964_IN
port 1998 n
rlabel metal5 68020 -35480 68120 -35380 1 PIX1965_IN
port 1999 n
rlabel metal5 69520 -35480 69620 -35380 1 PIX1966_IN
port 2000 n
rlabel metal5 71020 -35480 71120 -35380 1 PIX1967_IN
port 2001 n
rlabel metal5 72520 -35480 72620 -35380 1 PIX1968_IN
port 2002 n
rlabel metal5 74020 -35480 74120 -35380 1 PIX1969_IN
port 2003 n
rlabel metal5 75520 -35480 75620 -35380 1 PIX1970_IN
port 2004 n
rlabel metal5 77020 -35480 77120 -35380 1 PIX1971_IN
port 2005 n
rlabel metal5 78520 -35480 78620 -35380 1 PIX1972_IN
port 2006 n
rlabel metal5 80020 -35480 80120 -35380 1 PIX1973_IN
port 2007 n
rlabel metal5 81520 -35480 81620 -35380 1 PIX1974_IN
port 2008 n
rlabel metal5 83020 -35480 83120 -35380 1 PIX1975_IN
port 2009 n
rlabel metal5 84520 -35480 84620 -35380 1 PIX1976_IN
port 2010 n
rlabel metal5 86020 -35480 86120 -35380 1 PIX1977_IN
port 2011 n
rlabel metal5 87520 -35480 87620 -35380 1 PIX1978_IN
port 2012 n
rlabel metal5 89020 -35480 89120 -35380 1 PIX1979_IN
port 2013 n
rlabel metal5 90520 -35480 90620 -35380 1 PIX1980_IN
port 2014 n
rlabel metal5 92020 -35480 92120 -35380 1 PIX1981_IN
port 2015 n
rlabel metal5 93520 -35480 93620 -35380 1 PIX1982_IN
port 2016 n
rlabel metal5 95020 -35480 95120 -35380 1 PIX1983_IN
port 2017 n
rlabel metal5 96520 -35480 96620 -35380 1 PIX1984_IN
port 2018 n
rlabel metal5 98020 -35480 98120 -35380 1 PIX1985_IN
port 2019 n
rlabel metal5 99520 -35480 99620 -35380 1 PIX1986_IN
port 2020 n
rlabel metal5 101020 -35480 101120 -35380 1 PIX1987_IN
port 2021 n
rlabel metal5 102520 -35480 102620 -35380 1 PIX1988_IN
port 2022 n
rlabel metal5 104020 -35480 104120 -35380 1 PIX1989_IN
port 2023 n
rlabel metal5 105520 -35480 105620 -35380 1 PIX1990_IN
port 2024 n
rlabel metal5 107020 -35480 107120 -35380 1 PIX1991_IN
port 2025 n
rlabel metal5 108520 -35480 108620 -35380 1 PIX1992_IN
port 2026 n
rlabel metal5 110020 -35480 110120 -35380 1 PIX1993_IN
port 2027 n
rlabel metal5 111520 -35480 111620 -35380 1 PIX1994_IN
port 2028 n
rlabel metal5 113020 -35480 113120 -35380 1 PIX1995_IN
port 2029 n
rlabel metal5 114520 -35480 114620 -35380 1 PIX1996_IN
port 2030 n
rlabel metal5 116020 -35480 116120 -35380 1 PIX1997_IN
port 2031 n
rlabel metal5 117520 -35480 117620 -35380 1 PIX1998_IN
port 2032 n
rlabel metal5 119020 -35480 119120 -35380 1 PIX1999_IN
port 2033 n
rlabel metal5 520 -36980 620 -36880 1 PIX2000_IN
port 2034 n
rlabel metal2 -1500 -36760 -1500 -36715 3 ROW_SEL25
port 2035 e
rlabel metal5 2020 -36980 2120 -36880 1 PIX2001_IN
port 2036 n
rlabel metal5 3520 -36980 3620 -36880 1 PIX2002_IN
port 2037 n
rlabel metal5 5020 -36980 5120 -36880 1 PIX2003_IN
port 2038 n
rlabel metal5 6520 -36980 6620 -36880 1 PIX2004_IN
port 2039 n
rlabel metal5 8020 -36980 8120 -36880 1 PIX2005_IN
port 2040 n
rlabel metal5 9520 -36980 9620 -36880 1 PIX2006_IN
port 2041 n
rlabel metal5 11020 -36980 11120 -36880 1 PIX2007_IN
port 2042 n
rlabel metal5 12520 -36980 12620 -36880 1 PIX2008_IN
port 2043 n
rlabel metal5 14020 -36980 14120 -36880 1 PIX2009_IN
port 2044 n
rlabel metal5 15520 -36980 15620 -36880 1 PIX2010_IN
port 2045 n
rlabel metal5 17020 -36980 17120 -36880 1 PIX2011_IN
port 2046 n
rlabel metal5 18520 -36980 18620 -36880 1 PIX2012_IN
port 2047 n
rlabel metal5 20020 -36980 20120 -36880 1 PIX2013_IN
port 2048 n
rlabel metal5 21520 -36980 21620 -36880 1 PIX2014_IN
port 2049 n
rlabel metal5 23020 -36980 23120 -36880 1 PIX2015_IN
port 2050 n
rlabel metal5 24520 -36980 24620 -36880 1 PIX2016_IN
port 2051 n
rlabel metal5 26020 -36980 26120 -36880 1 PIX2017_IN
port 2052 n
rlabel metal5 27520 -36980 27620 -36880 1 PIX2018_IN
port 2053 n
rlabel metal5 29020 -36980 29120 -36880 1 PIX2019_IN
port 2054 n
rlabel metal5 30520 -36980 30620 -36880 1 PIX2020_IN
port 2055 n
rlabel metal5 32020 -36980 32120 -36880 1 PIX2021_IN
port 2056 n
rlabel metal5 33520 -36980 33620 -36880 1 PIX2022_IN
port 2057 n
rlabel metal5 35020 -36980 35120 -36880 1 PIX2023_IN
port 2058 n
rlabel metal5 36520 -36980 36620 -36880 1 PIX2024_IN
port 2059 n
rlabel metal5 38020 -36980 38120 -36880 1 PIX2025_IN
port 2060 n
rlabel metal5 39520 -36980 39620 -36880 1 PIX2026_IN
port 2061 n
rlabel metal5 41020 -36980 41120 -36880 1 PIX2027_IN
port 2062 n
rlabel metal5 42520 -36980 42620 -36880 1 PIX2028_IN
port 2063 n
rlabel metal5 44020 -36980 44120 -36880 1 PIX2029_IN
port 2064 n
rlabel metal5 45520 -36980 45620 -36880 1 PIX2030_IN
port 2065 n
rlabel metal5 47020 -36980 47120 -36880 1 PIX2031_IN
port 2066 n
rlabel metal5 48520 -36980 48620 -36880 1 PIX2032_IN
port 2067 n
rlabel metal5 50020 -36980 50120 -36880 1 PIX2033_IN
port 2068 n
rlabel metal5 51520 -36980 51620 -36880 1 PIX2034_IN
port 2069 n
rlabel metal5 53020 -36980 53120 -36880 1 PIX2035_IN
port 2070 n
rlabel metal5 54520 -36980 54620 -36880 1 PIX2036_IN
port 2071 n
rlabel metal5 56020 -36980 56120 -36880 1 PIX2037_IN
port 2072 n
rlabel metal5 57520 -36980 57620 -36880 1 PIX2038_IN
port 2073 n
rlabel metal5 59020 -36980 59120 -36880 1 PIX2039_IN
port 2074 n
rlabel metal5 60520 -36980 60620 -36880 1 PIX2040_IN
port 2075 n
rlabel metal5 62020 -36980 62120 -36880 1 PIX2041_IN
port 2076 n
rlabel metal5 63520 -36980 63620 -36880 1 PIX2042_IN
port 2077 n
rlabel metal5 65020 -36980 65120 -36880 1 PIX2043_IN
port 2078 n
rlabel metal5 66520 -36980 66620 -36880 1 PIX2044_IN
port 2079 n
rlabel metal5 68020 -36980 68120 -36880 1 PIX2045_IN
port 2080 n
rlabel metal5 69520 -36980 69620 -36880 1 PIX2046_IN
port 2081 n
rlabel metal5 71020 -36980 71120 -36880 1 PIX2047_IN
port 2082 n
rlabel metal5 72520 -36980 72620 -36880 1 PIX2048_IN
port 2083 n
rlabel metal5 74020 -36980 74120 -36880 1 PIX2049_IN
port 2084 n
rlabel metal5 75520 -36980 75620 -36880 1 PIX2050_IN
port 2085 n
rlabel metal5 77020 -36980 77120 -36880 1 PIX2051_IN
port 2086 n
rlabel metal5 78520 -36980 78620 -36880 1 PIX2052_IN
port 2087 n
rlabel metal5 80020 -36980 80120 -36880 1 PIX2053_IN
port 2088 n
rlabel metal5 81520 -36980 81620 -36880 1 PIX2054_IN
port 2089 n
rlabel metal5 83020 -36980 83120 -36880 1 PIX2055_IN
port 2090 n
rlabel metal5 84520 -36980 84620 -36880 1 PIX2056_IN
port 2091 n
rlabel metal5 86020 -36980 86120 -36880 1 PIX2057_IN
port 2092 n
rlabel metal5 87520 -36980 87620 -36880 1 PIX2058_IN
port 2093 n
rlabel metal5 89020 -36980 89120 -36880 1 PIX2059_IN
port 2094 n
rlabel metal5 90520 -36980 90620 -36880 1 PIX2060_IN
port 2095 n
rlabel metal5 92020 -36980 92120 -36880 1 PIX2061_IN
port 2096 n
rlabel metal5 93520 -36980 93620 -36880 1 PIX2062_IN
port 2097 n
rlabel metal5 95020 -36980 95120 -36880 1 PIX2063_IN
port 2098 n
rlabel metal5 96520 -36980 96620 -36880 1 PIX2064_IN
port 2099 n
rlabel metal5 98020 -36980 98120 -36880 1 PIX2065_IN
port 2100 n
rlabel metal5 99520 -36980 99620 -36880 1 PIX2066_IN
port 2101 n
rlabel metal5 101020 -36980 101120 -36880 1 PIX2067_IN
port 2102 n
rlabel metal5 102520 -36980 102620 -36880 1 PIX2068_IN
port 2103 n
rlabel metal5 104020 -36980 104120 -36880 1 PIX2069_IN
port 2104 n
rlabel metal5 105520 -36980 105620 -36880 1 PIX2070_IN
port 2105 n
rlabel metal5 107020 -36980 107120 -36880 1 PIX2071_IN
port 2106 n
rlabel metal5 108520 -36980 108620 -36880 1 PIX2072_IN
port 2107 n
rlabel metal5 110020 -36980 110120 -36880 1 PIX2073_IN
port 2108 n
rlabel metal5 111520 -36980 111620 -36880 1 PIX2074_IN
port 2109 n
rlabel metal5 113020 -36980 113120 -36880 1 PIX2075_IN
port 2110 n
rlabel metal5 114520 -36980 114620 -36880 1 PIX2076_IN
port 2111 n
rlabel metal5 116020 -36980 116120 -36880 1 PIX2077_IN
port 2112 n
rlabel metal5 117520 -36980 117620 -36880 1 PIX2078_IN
port 2113 n
rlabel metal5 119020 -36980 119120 -36880 1 PIX2079_IN
port 2114 n
rlabel metal5 520 -38480 620 -38380 1 PIX2080_IN
port 2115 n
rlabel metal2 -1500 -38260 -1500 -38215 3 ROW_SEL26
port 2116 e
rlabel metal5 2020 -38480 2120 -38380 1 PIX2081_IN
port 2117 n
rlabel metal5 3520 -38480 3620 -38380 1 PIX2082_IN
port 2118 n
rlabel metal5 5020 -38480 5120 -38380 1 PIX2083_IN
port 2119 n
rlabel metal5 6520 -38480 6620 -38380 1 PIX2084_IN
port 2120 n
rlabel metal5 8020 -38480 8120 -38380 1 PIX2085_IN
port 2121 n
rlabel metal5 9520 -38480 9620 -38380 1 PIX2086_IN
port 2122 n
rlabel metal5 11020 -38480 11120 -38380 1 PIX2087_IN
port 2123 n
rlabel metal5 12520 -38480 12620 -38380 1 PIX2088_IN
port 2124 n
rlabel metal5 14020 -38480 14120 -38380 1 PIX2089_IN
port 2125 n
rlabel metal5 15520 -38480 15620 -38380 1 PIX2090_IN
port 2126 n
rlabel metal5 17020 -38480 17120 -38380 1 PIX2091_IN
port 2127 n
rlabel metal5 18520 -38480 18620 -38380 1 PIX2092_IN
port 2128 n
rlabel metal5 20020 -38480 20120 -38380 1 PIX2093_IN
port 2129 n
rlabel metal5 21520 -38480 21620 -38380 1 PIX2094_IN
port 2130 n
rlabel metal5 23020 -38480 23120 -38380 1 PIX2095_IN
port 2131 n
rlabel metal5 24520 -38480 24620 -38380 1 PIX2096_IN
port 2132 n
rlabel metal5 26020 -38480 26120 -38380 1 PIX2097_IN
port 2133 n
rlabel metal5 27520 -38480 27620 -38380 1 PIX2098_IN
port 2134 n
rlabel metal5 29020 -38480 29120 -38380 1 PIX2099_IN
port 2135 n
rlabel metal5 30520 -38480 30620 -38380 1 PIX2100_IN
port 2136 n
rlabel metal5 32020 -38480 32120 -38380 1 PIX2101_IN
port 2137 n
rlabel metal5 33520 -38480 33620 -38380 1 PIX2102_IN
port 2138 n
rlabel metal5 35020 -38480 35120 -38380 1 PIX2103_IN
port 2139 n
rlabel metal5 36520 -38480 36620 -38380 1 PIX2104_IN
port 2140 n
rlabel metal5 38020 -38480 38120 -38380 1 PIX2105_IN
port 2141 n
rlabel metal5 39520 -38480 39620 -38380 1 PIX2106_IN
port 2142 n
rlabel metal5 41020 -38480 41120 -38380 1 PIX2107_IN
port 2143 n
rlabel metal5 42520 -38480 42620 -38380 1 PIX2108_IN
port 2144 n
rlabel metal5 44020 -38480 44120 -38380 1 PIX2109_IN
port 2145 n
rlabel metal5 45520 -38480 45620 -38380 1 PIX2110_IN
port 2146 n
rlabel metal5 47020 -38480 47120 -38380 1 PIX2111_IN
port 2147 n
rlabel metal5 48520 -38480 48620 -38380 1 PIX2112_IN
port 2148 n
rlabel metal5 50020 -38480 50120 -38380 1 PIX2113_IN
port 2149 n
rlabel metal5 51520 -38480 51620 -38380 1 PIX2114_IN
port 2150 n
rlabel metal5 53020 -38480 53120 -38380 1 PIX2115_IN
port 2151 n
rlabel metal5 54520 -38480 54620 -38380 1 PIX2116_IN
port 2152 n
rlabel metal5 56020 -38480 56120 -38380 1 PIX2117_IN
port 2153 n
rlabel metal5 57520 -38480 57620 -38380 1 PIX2118_IN
port 2154 n
rlabel metal5 59020 -38480 59120 -38380 1 PIX2119_IN
port 2155 n
rlabel metal5 60520 -38480 60620 -38380 1 PIX2120_IN
port 2156 n
rlabel metal5 62020 -38480 62120 -38380 1 PIX2121_IN
port 2157 n
rlabel metal5 63520 -38480 63620 -38380 1 PIX2122_IN
port 2158 n
rlabel metal5 65020 -38480 65120 -38380 1 PIX2123_IN
port 2159 n
rlabel metal5 66520 -38480 66620 -38380 1 PIX2124_IN
port 2160 n
rlabel metal5 68020 -38480 68120 -38380 1 PIX2125_IN
port 2161 n
rlabel metal5 69520 -38480 69620 -38380 1 PIX2126_IN
port 2162 n
rlabel metal5 71020 -38480 71120 -38380 1 PIX2127_IN
port 2163 n
rlabel metal5 72520 -38480 72620 -38380 1 PIX2128_IN
port 2164 n
rlabel metal5 74020 -38480 74120 -38380 1 PIX2129_IN
port 2165 n
rlabel metal5 75520 -38480 75620 -38380 1 PIX2130_IN
port 2166 n
rlabel metal5 77020 -38480 77120 -38380 1 PIX2131_IN
port 2167 n
rlabel metal5 78520 -38480 78620 -38380 1 PIX2132_IN
port 2168 n
rlabel metal5 80020 -38480 80120 -38380 1 PIX2133_IN
port 2169 n
rlabel metal5 81520 -38480 81620 -38380 1 PIX2134_IN
port 2170 n
rlabel metal5 83020 -38480 83120 -38380 1 PIX2135_IN
port 2171 n
rlabel metal5 84520 -38480 84620 -38380 1 PIX2136_IN
port 2172 n
rlabel metal5 86020 -38480 86120 -38380 1 PIX2137_IN
port 2173 n
rlabel metal5 87520 -38480 87620 -38380 1 PIX2138_IN
port 2174 n
rlabel metal5 89020 -38480 89120 -38380 1 PIX2139_IN
port 2175 n
rlabel metal5 90520 -38480 90620 -38380 1 PIX2140_IN
port 2176 n
rlabel metal5 92020 -38480 92120 -38380 1 PIX2141_IN
port 2177 n
rlabel metal5 93520 -38480 93620 -38380 1 PIX2142_IN
port 2178 n
rlabel metal5 95020 -38480 95120 -38380 1 PIX2143_IN
port 2179 n
rlabel metal5 96520 -38480 96620 -38380 1 PIX2144_IN
port 2180 n
rlabel metal5 98020 -38480 98120 -38380 1 PIX2145_IN
port 2181 n
rlabel metal5 99520 -38480 99620 -38380 1 PIX2146_IN
port 2182 n
rlabel metal5 101020 -38480 101120 -38380 1 PIX2147_IN
port 2183 n
rlabel metal5 102520 -38480 102620 -38380 1 PIX2148_IN
port 2184 n
rlabel metal5 104020 -38480 104120 -38380 1 PIX2149_IN
port 2185 n
rlabel metal5 105520 -38480 105620 -38380 1 PIX2150_IN
port 2186 n
rlabel metal5 107020 -38480 107120 -38380 1 PIX2151_IN
port 2187 n
rlabel metal5 108520 -38480 108620 -38380 1 PIX2152_IN
port 2188 n
rlabel metal5 110020 -38480 110120 -38380 1 PIX2153_IN
port 2189 n
rlabel metal5 111520 -38480 111620 -38380 1 PIX2154_IN
port 2190 n
rlabel metal5 113020 -38480 113120 -38380 1 PIX2155_IN
port 2191 n
rlabel metal5 114520 -38480 114620 -38380 1 PIX2156_IN
port 2192 n
rlabel metal5 116020 -38480 116120 -38380 1 PIX2157_IN
port 2193 n
rlabel metal5 117520 -38480 117620 -38380 1 PIX2158_IN
port 2194 n
rlabel metal5 119020 -38480 119120 -38380 1 PIX2159_IN
port 2195 n
rlabel metal5 520 -39980 620 -39880 1 PIX2160_IN
port 2196 n
rlabel metal2 -1500 -39760 -1500 -39715 3 ROW_SEL27
port 2197 e
rlabel metal5 2020 -39980 2120 -39880 1 PIX2161_IN
port 2198 n
rlabel metal5 3520 -39980 3620 -39880 1 PIX2162_IN
port 2199 n
rlabel metal5 5020 -39980 5120 -39880 1 PIX2163_IN
port 2200 n
rlabel metal5 6520 -39980 6620 -39880 1 PIX2164_IN
port 2201 n
rlabel metal5 8020 -39980 8120 -39880 1 PIX2165_IN
port 2202 n
rlabel metal5 9520 -39980 9620 -39880 1 PIX2166_IN
port 2203 n
rlabel metal5 11020 -39980 11120 -39880 1 PIX2167_IN
port 2204 n
rlabel metal5 12520 -39980 12620 -39880 1 PIX2168_IN
port 2205 n
rlabel metal5 14020 -39980 14120 -39880 1 PIX2169_IN
port 2206 n
rlabel metal5 15520 -39980 15620 -39880 1 PIX2170_IN
port 2207 n
rlabel metal5 17020 -39980 17120 -39880 1 PIX2171_IN
port 2208 n
rlabel metal5 18520 -39980 18620 -39880 1 PIX2172_IN
port 2209 n
rlabel metal5 20020 -39980 20120 -39880 1 PIX2173_IN
port 2210 n
rlabel metal5 21520 -39980 21620 -39880 1 PIX2174_IN
port 2211 n
rlabel metal5 23020 -39980 23120 -39880 1 PIX2175_IN
port 2212 n
rlabel metal5 24520 -39980 24620 -39880 1 PIX2176_IN
port 2213 n
rlabel metal5 26020 -39980 26120 -39880 1 PIX2177_IN
port 2214 n
rlabel metal5 27520 -39980 27620 -39880 1 PIX2178_IN
port 2215 n
rlabel metal5 29020 -39980 29120 -39880 1 PIX2179_IN
port 2216 n
rlabel metal5 30520 -39980 30620 -39880 1 PIX2180_IN
port 2217 n
rlabel metal5 32020 -39980 32120 -39880 1 PIX2181_IN
port 2218 n
rlabel metal5 33520 -39980 33620 -39880 1 PIX2182_IN
port 2219 n
rlabel metal5 35020 -39980 35120 -39880 1 PIX2183_IN
port 2220 n
rlabel metal5 36520 -39980 36620 -39880 1 PIX2184_IN
port 2221 n
rlabel metal5 38020 -39980 38120 -39880 1 PIX2185_IN
port 2222 n
rlabel metal5 39520 -39980 39620 -39880 1 PIX2186_IN
port 2223 n
rlabel metal5 41020 -39980 41120 -39880 1 PIX2187_IN
port 2224 n
rlabel metal5 42520 -39980 42620 -39880 1 PIX2188_IN
port 2225 n
rlabel metal5 44020 -39980 44120 -39880 1 PIX2189_IN
port 2226 n
rlabel metal5 45520 -39980 45620 -39880 1 PIX2190_IN
port 2227 n
rlabel metal5 47020 -39980 47120 -39880 1 PIX2191_IN
port 2228 n
rlabel metal5 48520 -39980 48620 -39880 1 PIX2192_IN
port 2229 n
rlabel metal5 50020 -39980 50120 -39880 1 PIX2193_IN
port 2230 n
rlabel metal5 51520 -39980 51620 -39880 1 PIX2194_IN
port 2231 n
rlabel metal5 53020 -39980 53120 -39880 1 PIX2195_IN
port 2232 n
rlabel metal5 54520 -39980 54620 -39880 1 PIX2196_IN
port 2233 n
rlabel metal5 56020 -39980 56120 -39880 1 PIX2197_IN
port 2234 n
rlabel metal5 57520 -39980 57620 -39880 1 PIX2198_IN
port 2235 n
rlabel metal5 59020 -39980 59120 -39880 1 PIX2199_IN
port 2236 n
rlabel metal5 60520 -39980 60620 -39880 1 PIX2200_IN
port 2237 n
rlabel metal5 62020 -39980 62120 -39880 1 PIX2201_IN
port 2238 n
rlabel metal5 63520 -39980 63620 -39880 1 PIX2202_IN
port 2239 n
rlabel metal5 65020 -39980 65120 -39880 1 PIX2203_IN
port 2240 n
rlabel metal5 66520 -39980 66620 -39880 1 PIX2204_IN
port 2241 n
rlabel metal5 68020 -39980 68120 -39880 1 PIX2205_IN
port 2242 n
rlabel metal5 69520 -39980 69620 -39880 1 PIX2206_IN
port 2243 n
rlabel metal5 71020 -39980 71120 -39880 1 PIX2207_IN
port 2244 n
rlabel metal5 72520 -39980 72620 -39880 1 PIX2208_IN
port 2245 n
rlabel metal5 74020 -39980 74120 -39880 1 PIX2209_IN
port 2246 n
rlabel metal5 75520 -39980 75620 -39880 1 PIX2210_IN
port 2247 n
rlabel metal5 77020 -39980 77120 -39880 1 PIX2211_IN
port 2248 n
rlabel metal5 78520 -39980 78620 -39880 1 PIX2212_IN
port 2249 n
rlabel metal5 80020 -39980 80120 -39880 1 PIX2213_IN
port 2250 n
rlabel metal5 81520 -39980 81620 -39880 1 PIX2214_IN
port 2251 n
rlabel metal5 83020 -39980 83120 -39880 1 PIX2215_IN
port 2252 n
rlabel metal5 84520 -39980 84620 -39880 1 PIX2216_IN
port 2253 n
rlabel metal5 86020 -39980 86120 -39880 1 PIX2217_IN
port 2254 n
rlabel metal5 87520 -39980 87620 -39880 1 PIX2218_IN
port 2255 n
rlabel metal5 89020 -39980 89120 -39880 1 PIX2219_IN
port 2256 n
rlabel metal5 90520 -39980 90620 -39880 1 PIX2220_IN
port 2257 n
rlabel metal5 92020 -39980 92120 -39880 1 PIX2221_IN
port 2258 n
rlabel metal5 93520 -39980 93620 -39880 1 PIX2222_IN
port 2259 n
rlabel metal5 95020 -39980 95120 -39880 1 PIX2223_IN
port 2260 n
rlabel metal5 96520 -39980 96620 -39880 1 PIX2224_IN
port 2261 n
rlabel metal5 98020 -39980 98120 -39880 1 PIX2225_IN
port 2262 n
rlabel metal5 99520 -39980 99620 -39880 1 PIX2226_IN
port 2263 n
rlabel metal5 101020 -39980 101120 -39880 1 PIX2227_IN
port 2264 n
rlabel metal5 102520 -39980 102620 -39880 1 PIX2228_IN
port 2265 n
rlabel metal5 104020 -39980 104120 -39880 1 PIX2229_IN
port 2266 n
rlabel metal5 105520 -39980 105620 -39880 1 PIX2230_IN
port 2267 n
rlabel metal5 107020 -39980 107120 -39880 1 PIX2231_IN
port 2268 n
rlabel metal5 108520 -39980 108620 -39880 1 PIX2232_IN
port 2269 n
rlabel metal5 110020 -39980 110120 -39880 1 PIX2233_IN
port 2270 n
rlabel metal5 111520 -39980 111620 -39880 1 PIX2234_IN
port 2271 n
rlabel metal5 113020 -39980 113120 -39880 1 PIX2235_IN
port 2272 n
rlabel metal5 114520 -39980 114620 -39880 1 PIX2236_IN
port 2273 n
rlabel metal5 116020 -39980 116120 -39880 1 PIX2237_IN
port 2274 n
rlabel metal5 117520 -39980 117620 -39880 1 PIX2238_IN
port 2275 n
rlabel metal5 119020 -39980 119120 -39880 1 PIX2239_IN
port 2276 n
rlabel metal5 520 -41480 620 -41380 1 PIX2240_IN
port 2277 n
rlabel metal2 -1500 -41260 -1500 -41215 3 ROW_SEL28
port 2278 e
rlabel metal5 2020 -41480 2120 -41380 1 PIX2241_IN
port 2279 n
rlabel metal5 3520 -41480 3620 -41380 1 PIX2242_IN
port 2280 n
rlabel metal5 5020 -41480 5120 -41380 1 PIX2243_IN
port 2281 n
rlabel metal5 6520 -41480 6620 -41380 1 PIX2244_IN
port 2282 n
rlabel metal5 8020 -41480 8120 -41380 1 PIX2245_IN
port 2283 n
rlabel metal5 9520 -41480 9620 -41380 1 PIX2246_IN
port 2284 n
rlabel metal5 11020 -41480 11120 -41380 1 PIX2247_IN
port 2285 n
rlabel metal5 12520 -41480 12620 -41380 1 PIX2248_IN
port 2286 n
rlabel metal5 14020 -41480 14120 -41380 1 PIX2249_IN
port 2287 n
rlabel metal5 15520 -41480 15620 -41380 1 PIX2250_IN
port 2288 n
rlabel metal5 17020 -41480 17120 -41380 1 PIX2251_IN
port 2289 n
rlabel metal5 18520 -41480 18620 -41380 1 PIX2252_IN
port 2290 n
rlabel metal5 20020 -41480 20120 -41380 1 PIX2253_IN
port 2291 n
rlabel metal5 21520 -41480 21620 -41380 1 PIX2254_IN
port 2292 n
rlabel metal5 23020 -41480 23120 -41380 1 PIX2255_IN
port 2293 n
rlabel metal5 24520 -41480 24620 -41380 1 PIX2256_IN
port 2294 n
rlabel metal5 26020 -41480 26120 -41380 1 PIX2257_IN
port 2295 n
rlabel metal5 27520 -41480 27620 -41380 1 PIX2258_IN
port 2296 n
rlabel metal5 29020 -41480 29120 -41380 1 PIX2259_IN
port 2297 n
rlabel metal5 30520 -41480 30620 -41380 1 PIX2260_IN
port 2298 n
rlabel metal5 32020 -41480 32120 -41380 1 PIX2261_IN
port 2299 n
rlabel metal5 33520 -41480 33620 -41380 1 PIX2262_IN
port 2300 n
rlabel metal5 35020 -41480 35120 -41380 1 PIX2263_IN
port 2301 n
rlabel metal5 36520 -41480 36620 -41380 1 PIX2264_IN
port 2302 n
rlabel metal5 38020 -41480 38120 -41380 1 PIX2265_IN
port 2303 n
rlabel metal5 39520 -41480 39620 -41380 1 PIX2266_IN
port 2304 n
rlabel metal5 41020 -41480 41120 -41380 1 PIX2267_IN
port 2305 n
rlabel metal5 42520 -41480 42620 -41380 1 PIX2268_IN
port 2306 n
rlabel metal5 44020 -41480 44120 -41380 1 PIX2269_IN
port 2307 n
rlabel metal5 45520 -41480 45620 -41380 1 PIX2270_IN
port 2308 n
rlabel metal5 47020 -41480 47120 -41380 1 PIX2271_IN
port 2309 n
rlabel metal5 48520 -41480 48620 -41380 1 PIX2272_IN
port 2310 n
rlabel metal5 50020 -41480 50120 -41380 1 PIX2273_IN
port 2311 n
rlabel metal5 51520 -41480 51620 -41380 1 PIX2274_IN
port 2312 n
rlabel metal5 53020 -41480 53120 -41380 1 PIX2275_IN
port 2313 n
rlabel metal5 54520 -41480 54620 -41380 1 PIX2276_IN
port 2314 n
rlabel metal5 56020 -41480 56120 -41380 1 PIX2277_IN
port 2315 n
rlabel metal5 57520 -41480 57620 -41380 1 PIX2278_IN
port 2316 n
rlabel metal5 59020 -41480 59120 -41380 1 PIX2279_IN
port 2317 n
rlabel metal5 60520 -41480 60620 -41380 1 PIX2280_IN
port 2318 n
rlabel metal5 62020 -41480 62120 -41380 1 PIX2281_IN
port 2319 n
rlabel metal5 63520 -41480 63620 -41380 1 PIX2282_IN
port 2320 n
rlabel metal5 65020 -41480 65120 -41380 1 PIX2283_IN
port 2321 n
rlabel metal5 66520 -41480 66620 -41380 1 PIX2284_IN
port 2322 n
rlabel metal5 68020 -41480 68120 -41380 1 PIX2285_IN
port 2323 n
rlabel metal5 69520 -41480 69620 -41380 1 PIX2286_IN
port 2324 n
rlabel metal5 71020 -41480 71120 -41380 1 PIX2287_IN
port 2325 n
rlabel metal5 72520 -41480 72620 -41380 1 PIX2288_IN
port 2326 n
rlabel metal5 74020 -41480 74120 -41380 1 PIX2289_IN
port 2327 n
rlabel metal5 75520 -41480 75620 -41380 1 PIX2290_IN
port 2328 n
rlabel metal5 77020 -41480 77120 -41380 1 PIX2291_IN
port 2329 n
rlabel metal5 78520 -41480 78620 -41380 1 PIX2292_IN
port 2330 n
rlabel metal5 80020 -41480 80120 -41380 1 PIX2293_IN
port 2331 n
rlabel metal5 81520 -41480 81620 -41380 1 PIX2294_IN
port 2332 n
rlabel metal5 83020 -41480 83120 -41380 1 PIX2295_IN
port 2333 n
rlabel metal5 84520 -41480 84620 -41380 1 PIX2296_IN
port 2334 n
rlabel metal5 86020 -41480 86120 -41380 1 PIX2297_IN
port 2335 n
rlabel metal5 87520 -41480 87620 -41380 1 PIX2298_IN
port 2336 n
rlabel metal5 89020 -41480 89120 -41380 1 PIX2299_IN
port 2337 n
rlabel metal5 90520 -41480 90620 -41380 1 PIX2300_IN
port 2338 n
rlabel metal5 92020 -41480 92120 -41380 1 PIX2301_IN
port 2339 n
rlabel metal5 93520 -41480 93620 -41380 1 PIX2302_IN
port 2340 n
rlabel metal5 95020 -41480 95120 -41380 1 PIX2303_IN
port 2341 n
rlabel metal5 96520 -41480 96620 -41380 1 PIX2304_IN
port 2342 n
rlabel metal5 98020 -41480 98120 -41380 1 PIX2305_IN
port 2343 n
rlabel metal5 99520 -41480 99620 -41380 1 PIX2306_IN
port 2344 n
rlabel metal5 101020 -41480 101120 -41380 1 PIX2307_IN
port 2345 n
rlabel metal5 102520 -41480 102620 -41380 1 PIX2308_IN
port 2346 n
rlabel metal5 104020 -41480 104120 -41380 1 PIX2309_IN
port 2347 n
rlabel metal5 105520 -41480 105620 -41380 1 PIX2310_IN
port 2348 n
rlabel metal5 107020 -41480 107120 -41380 1 PIX2311_IN
port 2349 n
rlabel metal5 108520 -41480 108620 -41380 1 PIX2312_IN
port 2350 n
rlabel metal5 110020 -41480 110120 -41380 1 PIX2313_IN
port 2351 n
rlabel metal5 111520 -41480 111620 -41380 1 PIX2314_IN
port 2352 n
rlabel metal5 113020 -41480 113120 -41380 1 PIX2315_IN
port 2353 n
rlabel metal5 114520 -41480 114620 -41380 1 PIX2316_IN
port 2354 n
rlabel metal5 116020 -41480 116120 -41380 1 PIX2317_IN
port 2355 n
rlabel metal5 117520 -41480 117620 -41380 1 PIX2318_IN
port 2356 n
rlabel metal5 119020 -41480 119120 -41380 1 PIX2319_IN
port 2357 n
rlabel metal5 520 -42980 620 -42880 1 PIX2320_IN
port 2358 n
rlabel metal2 -1500 -42760 -1500 -42715 3 ROW_SEL29
port 2359 e
rlabel metal5 2020 -42980 2120 -42880 1 PIX2321_IN
port 2360 n
rlabel metal5 3520 -42980 3620 -42880 1 PIX2322_IN
port 2361 n
rlabel metal5 5020 -42980 5120 -42880 1 PIX2323_IN
port 2362 n
rlabel metal5 6520 -42980 6620 -42880 1 PIX2324_IN
port 2363 n
rlabel metal5 8020 -42980 8120 -42880 1 PIX2325_IN
port 2364 n
rlabel metal5 9520 -42980 9620 -42880 1 PIX2326_IN
port 2365 n
rlabel metal5 11020 -42980 11120 -42880 1 PIX2327_IN
port 2366 n
rlabel metal5 12520 -42980 12620 -42880 1 PIX2328_IN
port 2367 n
rlabel metal5 14020 -42980 14120 -42880 1 PIX2329_IN
port 2368 n
rlabel metal5 15520 -42980 15620 -42880 1 PIX2330_IN
port 2369 n
rlabel metal5 17020 -42980 17120 -42880 1 PIX2331_IN
port 2370 n
rlabel metal5 18520 -42980 18620 -42880 1 PIX2332_IN
port 2371 n
rlabel metal5 20020 -42980 20120 -42880 1 PIX2333_IN
port 2372 n
rlabel metal5 21520 -42980 21620 -42880 1 PIX2334_IN
port 2373 n
rlabel metal5 23020 -42980 23120 -42880 1 PIX2335_IN
port 2374 n
rlabel metal5 24520 -42980 24620 -42880 1 PIX2336_IN
port 2375 n
rlabel metal5 26020 -42980 26120 -42880 1 PIX2337_IN
port 2376 n
rlabel metal5 27520 -42980 27620 -42880 1 PIX2338_IN
port 2377 n
rlabel metal5 29020 -42980 29120 -42880 1 PIX2339_IN
port 2378 n
rlabel metal5 30520 -42980 30620 -42880 1 PIX2340_IN
port 2379 n
rlabel metal5 32020 -42980 32120 -42880 1 PIX2341_IN
port 2380 n
rlabel metal5 33520 -42980 33620 -42880 1 PIX2342_IN
port 2381 n
rlabel metal5 35020 -42980 35120 -42880 1 PIX2343_IN
port 2382 n
rlabel metal5 36520 -42980 36620 -42880 1 PIX2344_IN
port 2383 n
rlabel metal5 38020 -42980 38120 -42880 1 PIX2345_IN
port 2384 n
rlabel metal5 39520 -42980 39620 -42880 1 PIX2346_IN
port 2385 n
rlabel metal5 41020 -42980 41120 -42880 1 PIX2347_IN
port 2386 n
rlabel metal5 42520 -42980 42620 -42880 1 PIX2348_IN
port 2387 n
rlabel metal5 44020 -42980 44120 -42880 1 PIX2349_IN
port 2388 n
rlabel metal5 45520 -42980 45620 -42880 1 PIX2350_IN
port 2389 n
rlabel metal5 47020 -42980 47120 -42880 1 PIX2351_IN
port 2390 n
rlabel metal5 48520 -42980 48620 -42880 1 PIX2352_IN
port 2391 n
rlabel metal5 50020 -42980 50120 -42880 1 PIX2353_IN
port 2392 n
rlabel metal5 51520 -42980 51620 -42880 1 PIX2354_IN
port 2393 n
rlabel metal5 53020 -42980 53120 -42880 1 PIX2355_IN
port 2394 n
rlabel metal5 54520 -42980 54620 -42880 1 PIX2356_IN
port 2395 n
rlabel metal5 56020 -42980 56120 -42880 1 PIX2357_IN
port 2396 n
rlabel metal5 57520 -42980 57620 -42880 1 PIX2358_IN
port 2397 n
rlabel metal5 59020 -42980 59120 -42880 1 PIX2359_IN
port 2398 n
rlabel metal5 60520 -42980 60620 -42880 1 PIX2360_IN
port 2399 n
rlabel metal5 62020 -42980 62120 -42880 1 PIX2361_IN
port 2400 n
rlabel metal5 63520 -42980 63620 -42880 1 PIX2362_IN
port 2401 n
rlabel metal5 65020 -42980 65120 -42880 1 PIX2363_IN
port 2402 n
rlabel metal5 66520 -42980 66620 -42880 1 PIX2364_IN
port 2403 n
rlabel metal5 68020 -42980 68120 -42880 1 PIX2365_IN
port 2404 n
rlabel metal5 69520 -42980 69620 -42880 1 PIX2366_IN
port 2405 n
rlabel metal5 71020 -42980 71120 -42880 1 PIX2367_IN
port 2406 n
rlabel metal5 72520 -42980 72620 -42880 1 PIX2368_IN
port 2407 n
rlabel metal5 74020 -42980 74120 -42880 1 PIX2369_IN
port 2408 n
rlabel metal5 75520 -42980 75620 -42880 1 PIX2370_IN
port 2409 n
rlabel metal5 77020 -42980 77120 -42880 1 PIX2371_IN
port 2410 n
rlabel metal5 78520 -42980 78620 -42880 1 PIX2372_IN
port 2411 n
rlabel metal5 80020 -42980 80120 -42880 1 PIX2373_IN
port 2412 n
rlabel metal5 81520 -42980 81620 -42880 1 PIX2374_IN
port 2413 n
rlabel metal5 83020 -42980 83120 -42880 1 PIX2375_IN
port 2414 n
rlabel metal5 84520 -42980 84620 -42880 1 PIX2376_IN
port 2415 n
rlabel metal5 86020 -42980 86120 -42880 1 PIX2377_IN
port 2416 n
rlabel metal5 87520 -42980 87620 -42880 1 PIX2378_IN
port 2417 n
rlabel metal5 89020 -42980 89120 -42880 1 PIX2379_IN
port 2418 n
rlabel metal5 90520 -42980 90620 -42880 1 PIX2380_IN
port 2419 n
rlabel metal5 92020 -42980 92120 -42880 1 PIX2381_IN
port 2420 n
rlabel metal5 93520 -42980 93620 -42880 1 PIX2382_IN
port 2421 n
rlabel metal5 95020 -42980 95120 -42880 1 PIX2383_IN
port 2422 n
rlabel metal5 96520 -42980 96620 -42880 1 PIX2384_IN
port 2423 n
rlabel metal5 98020 -42980 98120 -42880 1 PIX2385_IN
port 2424 n
rlabel metal5 99520 -42980 99620 -42880 1 PIX2386_IN
port 2425 n
rlabel metal5 101020 -42980 101120 -42880 1 PIX2387_IN
port 2426 n
rlabel metal5 102520 -42980 102620 -42880 1 PIX2388_IN
port 2427 n
rlabel metal5 104020 -42980 104120 -42880 1 PIX2389_IN
port 2428 n
rlabel metal5 105520 -42980 105620 -42880 1 PIX2390_IN
port 2429 n
rlabel metal5 107020 -42980 107120 -42880 1 PIX2391_IN
port 2430 n
rlabel metal5 108520 -42980 108620 -42880 1 PIX2392_IN
port 2431 n
rlabel metal5 110020 -42980 110120 -42880 1 PIX2393_IN
port 2432 n
rlabel metal5 111520 -42980 111620 -42880 1 PIX2394_IN
port 2433 n
rlabel metal5 113020 -42980 113120 -42880 1 PIX2395_IN
port 2434 n
rlabel metal5 114520 -42980 114620 -42880 1 PIX2396_IN
port 2435 n
rlabel metal5 116020 -42980 116120 -42880 1 PIX2397_IN
port 2436 n
rlabel metal5 117520 -42980 117620 -42880 1 PIX2398_IN
port 2437 n
rlabel metal5 119020 -42980 119120 -42880 1 PIX2399_IN
port 2438 n
rlabel metal5 520 -44480 620 -44380 1 PIX2400_IN
port 2439 n
rlabel metal2 -1500 -44260 -1500 -44215 3 ROW_SEL30
port 2440 e
rlabel metal5 2020 -44480 2120 -44380 1 PIX2401_IN
port 2441 n
rlabel metal5 3520 -44480 3620 -44380 1 PIX2402_IN
port 2442 n
rlabel metal5 5020 -44480 5120 -44380 1 PIX2403_IN
port 2443 n
rlabel metal5 6520 -44480 6620 -44380 1 PIX2404_IN
port 2444 n
rlabel metal5 8020 -44480 8120 -44380 1 PIX2405_IN
port 2445 n
rlabel metal5 9520 -44480 9620 -44380 1 PIX2406_IN
port 2446 n
rlabel metal5 11020 -44480 11120 -44380 1 PIX2407_IN
port 2447 n
rlabel metal5 12520 -44480 12620 -44380 1 PIX2408_IN
port 2448 n
rlabel metal5 14020 -44480 14120 -44380 1 PIX2409_IN
port 2449 n
rlabel metal5 15520 -44480 15620 -44380 1 PIX2410_IN
port 2450 n
rlabel metal5 17020 -44480 17120 -44380 1 PIX2411_IN
port 2451 n
rlabel metal5 18520 -44480 18620 -44380 1 PIX2412_IN
port 2452 n
rlabel metal5 20020 -44480 20120 -44380 1 PIX2413_IN
port 2453 n
rlabel metal5 21520 -44480 21620 -44380 1 PIX2414_IN
port 2454 n
rlabel metal5 23020 -44480 23120 -44380 1 PIX2415_IN
port 2455 n
rlabel metal5 24520 -44480 24620 -44380 1 PIX2416_IN
port 2456 n
rlabel metal5 26020 -44480 26120 -44380 1 PIX2417_IN
port 2457 n
rlabel metal5 27520 -44480 27620 -44380 1 PIX2418_IN
port 2458 n
rlabel metal5 29020 -44480 29120 -44380 1 PIX2419_IN
port 2459 n
rlabel metal5 30520 -44480 30620 -44380 1 PIX2420_IN
port 2460 n
rlabel metal5 32020 -44480 32120 -44380 1 PIX2421_IN
port 2461 n
rlabel metal5 33520 -44480 33620 -44380 1 PIX2422_IN
port 2462 n
rlabel metal5 35020 -44480 35120 -44380 1 PIX2423_IN
port 2463 n
rlabel metal5 36520 -44480 36620 -44380 1 PIX2424_IN
port 2464 n
rlabel metal5 38020 -44480 38120 -44380 1 PIX2425_IN
port 2465 n
rlabel metal5 39520 -44480 39620 -44380 1 PIX2426_IN
port 2466 n
rlabel metal5 41020 -44480 41120 -44380 1 PIX2427_IN
port 2467 n
rlabel metal5 42520 -44480 42620 -44380 1 PIX2428_IN
port 2468 n
rlabel metal5 44020 -44480 44120 -44380 1 PIX2429_IN
port 2469 n
rlabel metal5 45520 -44480 45620 -44380 1 PIX2430_IN
port 2470 n
rlabel metal5 47020 -44480 47120 -44380 1 PIX2431_IN
port 2471 n
rlabel metal5 48520 -44480 48620 -44380 1 PIX2432_IN
port 2472 n
rlabel metal5 50020 -44480 50120 -44380 1 PIX2433_IN
port 2473 n
rlabel metal5 51520 -44480 51620 -44380 1 PIX2434_IN
port 2474 n
rlabel metal5 53020 -44480 53120 -44380 1 PIX2435_IN
port 2475 n
rlabel metal5 54520 -44480 54620 -44380 1 PIX2436_IN
port 2476 n
rlabel metal5 56020 -44480 56120 -44380 1 PIX2437_IN
port 2477 n
rlabel metal5 57520 -44480 57620 -44380 1 PIX2438_IN
port 2478 n
rlabel metal5 59020 -44480 59120 -44380 1 PIX2439_IN
port 2479 n
rlabel metal5 60520 -44480 60620 -44380 1 PIX2440_IN
port 2480 n
rlabel metal5 62020 -44480 62120 -44380 1 PIX2441_IN
port 2481 n
rlabel metal5 63520 -44480 63620 -44380 1 PIX2442_IN
port 2482 n
rlabel metal5 65020 -44480 65120 -44380 1 PIX2443_IN
port 2483 n
rlabel metal5 66520 -44480 66620 -44380 1 PIX2444_IN
port 2484 n
rlabel metal5 68020 -44480 68120 -44380 1 PIX2445_IN
port 2485 n
rlabel metal5 69520 -44480 69620 -44380 1 PIX2446_IN
port 2486 n
rlabel metal5 71020 -44480 71120 -44380 1 PIX2447_IN
port 2487 n
rlabel metal5 72520 -44480 72620 -44380 1 PIX2448_IN
port 2488 n
rlabel metal5 74020 -44480 74120 -44380 1 PIX2449_IN
port 2489 n
rlabel metal5 75520 -44480 75620 -44380 1 PIX2450_IN
port 2490 n
rlabel metal5 77020 -44480 77120 -44380 1 PIX2451_IN
port 2491 n
rlabel metal5 78520 -44480 78620 -44380 1 PIX2452_IN
port 2492 n
rlabel metal5 80020 -44480 80120 -44380 1 PIX2453_IN
port 2493 n
rlabel metal5 81520 -44480 81620 -44380 1 PIX2454_IN
port 2494 n
rlabel metal5 83020 -44480 83120 -44380 1 PIX2455_IN
port 2495 n
rlabel metal5 84520 -44480 84620 -44380 1 PIX2456_IN
port 2496 n
rlabel metal5 86020 -44480 86120 -44380 1 PIX2457_IN
port 2497 n
rlabel metal5 87520 -44480 87620 -44380 1 PIX2458_IN
port 2498 n
rlabel metal5 89020 -44480 89120 -44380 1 PIX2459_IN
port 2499 n
rlabel metal5 90520 -44480 90620 -44380 1 PIX2460_IN
port 2500 n
rlabel metal5 92020 -44480 92120 -44380 1 PIX2461_IN
port 2501 n
rlabel metal5 93520 -44480 93620 -44380 1 PIX2462_IN
port 2502 n
rlabel metal5 95020 -44480 95120 -44380 1 PIX2463_IN
port 2503 n
rlabel metal5 96520 -44480 96620 -44380 1 PIX2464_IN
port 2504 n
rlabel metal5 98020 -44480 98120 -44380 1 PIX2465_IN
port 2505 n
rlabel metal5 99520 -44480 99620 -44380 1 PIX2466_IN
port 2506 n
rlabel metal5 101020 -44480 101120 -44380 1 PIX2467_IN
port 2507 n
rlabel metal5 102520 -44480 102620 -44380 1 PIX2468_IN
port 2508 n
rlabel metal5 104020 -44480 104120 -44380 1 PIX2469_IN
port 2509 n
rlabel metal5 105520 -44480 105620 -44380 1 PIX2470_IN
port 2510 n
rlabel metal5 107020 -44480 107120 -44380 1 PIX2471_IN
port 2511 n
rlabel metal5 108520 -44480 108620 -44380 1 PIX2472_IN
port 2512 n
rlabel metal5 110020 -44480 110120 -44380 1 PIX2473_IN
port 2513 n
rlabel metal5 111520 -44480 111620 -44380 1 PIX2474_IN
port 2514 n
rlabel metal5 113020 -44480 113120 -44380 1 PIX2475_IN
port 2515 n
rlabel metal5 114520 -44480 114620 -44380 1 PIX2476_IN
port 2516 n
rlabel metal5 116020 -44480 116120 -44380 1 PIX2477_IN
port 2517 n
rlabel metal5 117520 -44480 117620 -44380 1 PIX2478_IN
port 2518 n
rlabel metal5 119020 -44480 119120 -44380 1 PIX2479_IN
port 2519 n
rlabel metal5 520 -45980 620 -45880 1 PIX2480_IN
port 2520 n
rlabel metal2 -1500 -45760 -1500 -45715 3 ROW_SEL31
port 2521 e
rlabel metal5 2020 -45980 2120 -45880 1 PIX2481_IN
port 2522 n
rlabel metal5 3520 -45980 3620 -45880 1 PIX2482_IN
port 2523 n
rlabel metal5 5020 -45980 5120 -45880 1 PIX2483_IN
port 2524 n
rlabel metal5 6520 -45980 6620 -45880 1 PIX2484_IN
port 2525 n
rlabel metal5 8020 -45980 8120 -45880 1 PIX2485_IN
port 2526 n
rlabel metal5 9520 -45980 9620 -45880 1 PIX2486_IN
port 2527 n
rlabel metal5 11020 -45980 11120 -45880 1 PIX2487_IN
port 2528 n
rlabel metal5 12520 -45980 12620 -45880 1 PIX2488_IN
port 2529 n
rlabel metal5 14020 -45980 14120 -45880 1 PIX2489_IN
port 2530 n
rlabel metal5 15520 -45980 15620 -45880 1 PIX2490_IN
port 2531 n
rlabel metal5 17020 -45980 17120 -45880 1 PIX2491_IN
port 2532 n
rlabel metal5 18520 -45980 18620 -45880 1 PIX2492_IN
port 2533 n
rlabel metal5 20020 -45980 20120 -45880 1 PIX2493_IN
port 2534 n
rlabel metal5 21520 -45980 21620 -45880 1 PIX2494_IN
port 2535 n
rlabel metal5 23020 -45980 23120 -45880 1 PIX2495_IN
port 2536 n
rlabel metal5 24520 -45980 24620 -45880 1 PIX2496_IN
port 2537 n
rlabel metal5 26020 -45980 26120 -45880 1 PIX2497_IN
port 2538 n
rlabel metal5 27520 -45980 27620 -45880 1 PIX2498_IN
port 2539 n
rlabel metal5 29020 -45980 29120 -45880 1 PIX2499_IN
port 2540 n
rlabel metal5 30520 -45980 30620 -45880 1 PIX2500_IN
port 2541 n
rlabel metal5 32020 -45980 32120 -45880 1 PIX2501_IN
port 2542 n
rlabel metal5 33520 -45980 33620 -45880 1 PIX2502_IN
port 2543 n
rlabel metal5 35020 -45980 35120 -45880 1 PIX2503_IN
port 2544 n
rlabel metal5 36520 -45980 36620 -45880 1 PIX2504_IN
port 2545 n
rlabel metal5 38020 -45980 38120 -45880 1 PIX2505_IN
port 2546 n
rlabel metal5 39520 -45980 39620 -45880 1 PIX2506_IN
port 2547 n
rlabel metal5 41020 -45980 41120 -45880 1 PIX2507_IN
port 2548 n
rlabel metal5 42520 -45980 42620 -45880 1 PIX2508_IN
port 2549 n
rlabel metal5 44020 -45980 44120 -45880 1 PIX2509_IN
port 2550 n
rlabel metal5 45520 -45980 45620 -45880 1 PIX2510_IN
port 2551 n
rlabel metal5 47020 -45980 47120 -45880 1 PIX2511_IN
port 2552 n
rlabel metal5 48520 -45980 48620 -45880 1 PIX2512_IN
port 2553 n
rlabel metal5 50020 -45980 50120 -45880 1 PIX2513_IN
port 2554 n
rlabel metal5 51520 -45980 51620 -45880 1 PIX2514_IN
port 2555 n
rlabel metal5 53020 -45980 53120 -45880 1 PIX2515_IN
port 2556 n
rlabel metal5 54520 -45980 54620 -45880 1 PIX2516_IN
port 2557 n
rlabel metal5 56020 -45980 56120 -45880 1 PIX2517_IN
port 2558 n
rlabel metal5 57520 -45980 57620 -45880 1 PIX2518_IN
port 2559 n
rlabel metal5 59020 -45980 59120 -45880 1 PIX2519_IN
port 2560 n
rlabel metal5 60520 -45980 60620 -45880 1 PIX2520_IN
port 2561 n
rlabel metal5 62020 -45980 62120 -45880 1 PIX2521_IN
port 2562 n
rlabel metal5 63520 -45980 63620 -45880 1 PIX2522_IN
port 2563 n
rlabel metal5 65020 -45980 65120 -45880 1 PIX2523_IN
port 2564 n
rlabel metal5 66520 -45980 66620 -45880 1 PIX2524_IN
port 2565 n
rlabel metal5 68020 -45980 68120 -45880 1 PIX2525_IN
port 2566 n
rlabel metal5 69520 -45980 69620 -45880 1 PIX2526_IN
port 2567 n
rlabel metal5 71020 -45980 71120 -45880 1 PIX2527_IN
port 2568 n
rlabel metal5 72520 -45980 72620 -45880 1 PIX2528_IN
port 2569 n
rlabel metal5 74020 -45980 74120 -45880 1 PIX2529_IN
port 2570 n
rlabel metal5 75520 -45980 75620 -45880 1 PIX2530_IN
port 2571 n
rlabel metal5 77020 -45980 77120 -45880 1 PIX2531_IN
port 2572 n
rlabel metal5 78520 -45980 78620 -45880 1 PIX2532_IN
port 2573 n
rlabel metal5 80020 -45980 80120 -45880 1 PIX2533_IN
port 2574 n
rlabel metal5 81520 -45980 81620 -45880 1 PIX2534_IN
port 2575 n
rlabel metal5 83020 -45980 83120 -45880 1 PIX2535_IN
port 2576 n
rlabel metal5 84520 -45980 84620 -45880 1 PIX2536_IN
port 2577 n
rlabel metal5 86020 -45980 86120 -45880 1 PIX2537_IN
port 2578 n
rlabel metal5 87520 -45980 87620 -45880 1 PIX2538_IN
port 2579 n
rlabel metal5 89020 -45980 89120 -45880 1 PIX2539_IN
port 2580 n
rlabel metal5 90520 -45980 90620 -45880 1 PIX2540_IN
port 2581 n
rlabel metal5 92020 -45980 92120 -45880 1 PIX2541_IN
port 2582 n
rlabel metal5 93520 -45980 93620 -45880 1 PIX2542_IN
port 2583 n
rlabel metal5 95020 -45980 95120 -45880 1 PIX2543_IN
port 2584 n
rlabel metal5 96520 -45980 96620 -45880 1 PIX2544_IN
port 2585 n
rlabel metal5 98020 -45980 98120 -45880 1 PIX2545_IN
port 2586 n
rlabel metal5 99520 -45980 99620 -45880 1 PIX2546_IN
port 2587 n
rlabel metal5 101020 -45980 101120 -45880 1 PIX2547_IN
port 2588 n
rlabel metal5 102520 -45980 102620 -45880 1 PIX2548_IN
port 2589 n
rlabel metal5 104020 -45980 104120 -45880 1 PIX2549_IN
port 2590 n
rlabel metal5 105520 -45980 105620 -45880 1 PIX2550_IN
port 2591 n
rlabel metal5 107020 -45980 107120 -45880 1 PIX2551_IN
port 2592 n
rlabel metal5 108520 -45980 108620 -45880 1 PIX2552_IN
port 2593 n
rlabel metal5 110020 -45980 110120 -45880 1 PIX2553_IN
port 2594 n
rlabel metal5 111520 -45980 111620 -45880 1 PIX2554_IN
port 2595 n
rlabel metal5 113020 -45980 113120 -45880 1 PIX2555_IN
port 2596 n
rlabel metal5 114520 -45980 114620 -45880 1 PIX2556_IN
port 2597 n
rlabel metal5 116020 -45980 116120 -45880 1 PIX2557_IN
port 2598 n
rlabel metal5 117520 -45980 117620 -45880 1 PIX2558_IN
port 2599 n
rlabel metal5 119020 -45980 119120 -45880 1 PIX2559_IN
port 2600 n
rlabel metal5 520 -47480 620 -47380 1 PIX2560_IN
port 2601 n
rlabel metal2 -1500 -47260 -1500 -47215 3 ROW_SEL32
port 2602 e
rlabel metal5 2020 -47480 2120 -47380 1 PIX2561_IN
port 2603 n
rlabel metal5 3520 -47480 3620 -47380 1 PIX2562_IN
port 2604 n
rlabel metal5 5020 -47480 5120 -47380 1 PIX2563_IN
port 2605 n
rlabel metal5 6520 -47480 6620 -47380 1 PIX2564_IN
port 2606 n
rlabel metal5 8020 -47480 8120 -47380 1 PIX2565_IN
port 2607 n
rlabel metal5 9520 -47480 9620 -47380 1 PIX2566_IN
port 2608 n
rlabel metal5 11020 -47480 11120 -47380 1 PIX2567_IN
port 2609 n
rlabel metal5 12520 -47480 12620 -47380 1 PIX2568_IN
port 2610 n
rlabel metal5 14020 -47480 14120 -47380 1 PIX2569_IN
port 2611 n
rlabel metal5 15520 -47480 15620 -47380 1 PIX2570_IN
port 2612 n
rlabel metal5 17020 -47480 17120 -47380 1 PIX2571_IN
port 2613 n
rlabel metal5 18520 -47480 18620 -47380 1 PIX2572_IN
port 2614 n
rlabel metal5 20020 -47480 20120 -47380 1 PIX2573_IN
port 2615 n
rlabel metal5 21520 -47480 21620 -47380 1 PIX2574_IN
port 2616 n
rlabel metal5 23020 -47480 23120 -47380 1 PIX2575_IN
port 2617 n
rlabel metal5 24520 -47480 24620 -47380 1 PIX2576_IN
port 2618 n
rlabel metal5 26020 -47480 26120 -47380 1 PIX2577_IN
port 2619 n
rlabel metal5 27520 -47480 27620 -47380 1 PIX2578_IN
port 2620 n
rlabel metal5 29020 -47480 29120 -47380 1 PIX2579_IN
port 2621 n
rlabel metal5 30520 -47480 30620 -47380 1 PIX2580_IN
port 2622 n
rlabel metal5 32020 -47480 32120 -47380 1 PIX2581_IN
port 2623 n
rlabel metal5 33520 -47480 33620 -47380 1 PIX2582_IN
port 2624 n
rlabel metal5 35020 -47480 35120 -47380 1 PIX2583_IN
port 2625 n
rlabel metal5 36520 -47480 36620 -47380 1 PIX2584_IN
port 2626 n
rlabel metal5 38020 -47480 38120 -47380 1 PIX2585_IN
port 2627 n
rlabel metal5 39520 -47480 39620 -47380 1 PIX2586_IN
port 2628 n
rlabel metal5 41020 -47480 41120 -47380 1 PIX2587_IN
port 2629 n
rlabel metal5 42520 -47480 42620 -47380 1 PIX2588_IN
port 2630 n
rlabel metal5 44020 -47480 44120 -47380 1 PIX2589_IN
port 2631 n
rlabel metal5 45520 -47480 45620 -47380 1 PIX2590_IN
port 2632 n
rlabel metal5 47020 -47480 47120 -47380 1 PIX2591_IN
port 2633 n
rlabel metal5 48520 -47480 48620 -47380 1 PIX2592_IN
port 2634 n
rlabel metal5 50020 -47480 50120 -47380 1 PIX2593_IN
port 2635 n
rlabel metal5 51520 -47480 51620 -47380 1 PIX2594_IN
port 2636 n
rlabel metal5 53020 -47480 53120 -47380 1 PIX2595_IN
port 2637 n
rlabel metal5 54520 -47480 54620 -47380 1 PIX2596_IN
port 2638 n
rlabel metal5 56020 -47480 56120 -47380 1 PIX2597_IN
port 2639 n
rlabel metal5 57520 -47480 57620 -47380 1 PIX2598_IN
port 2640 n
rlabel metal5 59020 -47480 59120 -47380 1 PIX2599_IN
port 2641 n
rlabel metal5 60520 -47480 60620 -47380 1 PIX2600_IN
port 2642 n
rlabel metal5 62020 -47480 62120 -47380 1 PIX2601_IN
port 2643 n
rlabel metal5 63520 -47480 63620 -47380 1 PIX2602_IN
port 2644 n
rlabel metal5 65020 -47480 65120 -47380 1 PIX2603_IN
port 2645 n
rlabel metal5 66520 -47480 66620 -47380 1 PIX2604_IN
port 2646 n
rlabel metal5 68020 -47480 68120 -47380 1 PIX2605_IN
port 2647 n
rlabel metal5 69520 -47480 69620 -47380 1 PIX2606_IN
port 2648 n
rlabel metal5 71020 -47480 71120 -47380 1 PIX2607_IN
port 2649 n
rlabel metal5 72520 -47480 72620 -47380 1 PIX2608_IN
port 2650 n
rlabel metal5 74020 -47480 74120 -47380 1 PIX2609_IN
port 2651 n
rlabel metal5 75520 -47480 75620 -47380 1 PIX2610_IN
port 2652 n
rlabel metal5 77020 -47480 77120 -47380 1 PIX2611_IN
port 2653 n
rlabel metal5 78520 -47480 78620 -47380 1 PIX2612_IN
port 2654 n
rlabel metal5 80020 -47480 80120 -47380 1 PIX2613_IN
port 2655 n
rlabel metal5 81520 -47480 81620 -47380 1 PIX2614_IN
port 2656 n
rlabel metal5 83020 -47480 83120 -47380 1 PIX2615_IN
port 2657 n
rlabel metal5 84520 -47480 84620 -47380 1 PIX2616_IN
port 2658 n
rlabel metal5 86020 -47480 86120 -47380 1 PIX2617_IN
port 2659 n
rlabel metal5 87520 -47480 87620 -47380 1 PIX2618_IN
port 2660 n
rlabel metal5 89020 -47480 89120 -47380 1 PIX2619_IN
port 2661 n
rlabel metal5 90520 -47480 90620 -47380 1 PIX2620_IN
port 2662 n
rlabel metal5 92020 -47480 92120 -47380 1 PIX2621_IN
port 2663 n
rlabel metal5 93520 -47480 93620 -47380 1 PIX2622_IN
port 2664 n
rlabel metal5 95020 -47480 95120 -47380 1 PIX2623_IN
port 2665 n
rlabel metal5 96520 -47480 96620 -47380 1 PIX2624_IN
port 2666 n
rlabel metal5 98020 -47480 98120 -47380 1 PIX2625_IN
port 2667 n
rlabel metal5 99520 -47480 99620 -47380 1 PIX2626_IN
port 2668 n
rlabel metal5 101020 -47480 101120 -47380 1 PIX2627_IN
port 2669 n
rlabel metal5 102520 -47480 102620 -47380 1 PIX2628_IN
port 2670 n
rlabel metal5 104020 -47480 104120 -47380 1 PIX2629_IN
port 2671 n
rlabel metal5 105520 -47480 105620 -47380 1 PIX2630_IN
port 2672 n
rlabel metal5 107020 -47480 107120 -47380 1 PIX2631_IN
port 2673 n
rlabel metal5 108520 -47480 108620 -47380 1 PIX2632_IN
port 2674 n
rlabel metal5 110020 -47480 110120 -47380 1 PIX2633_IN
port 2675 n
rlabel metal5 111520 -47480 111620 -47380 1 PIX2634_IN
port 2676 n
rlabel metal5 113020 -47480 113120 -47380 1 PIX2635_IN
port 2677 n
rlabel metal5 114520 -47480 114620 -47380 1 PIX2636_IN
port 2678 n
rlabel metal5 116020 -47480 116120 -47380 1 PIX2637_IN
port 2679 n
rlabel metal5 117520 -47480 117620 -47380 1 PIX2638_IN
port 2680 n
rlabel metal5 119020 -47480 119120 -47380 1 PIX2639_IN
port 2681 n
rlabel metal5 520 -48980 620 -48880 1 PIX2640_IN
port 2682 n
rlabel metal2 -1500 -48760 -1500 -48715 3 ROW_SEL33
port 2683 e
rlabel metal5 2020 -48980 2120 -48880 1 PIX2641_IN
port 2684 n
rlabel metal5 3520 -48980 3620 -48880 1 PIX2642_IN
port 2685 n
rlabel metal5 5020 -48980 5120 -48880 1 PIX2643_IN
port 2686 n
rlabel metal5 6520 -48980 6620 -48880 1 PIX2644_IN
port 2687 n
rlabel metal5 8020 -48980 8120 -48880 1 PIX2645_IN
port 2688 n
rlabel metal5 9520 -48980 9620 -48880 1 PIX2646_IN
port 2689 n
rlabel metal5 11020 -48980 11120 -48880 1 PIX2647_IN
port 2690 n
rlabel metal5 12520 -48980 12620 -48880 1 PIX2648_IN
port 2691 n
rlabel metal5 14020 -48980 14120 -48880 1 PIX2649_IN
port 2692 n
rlabel metal5 15520 -48980 15620 -48880 1 PIX2650_IN
port 2693 n
rlabel metal5 17020 -48980 17120 -48880 1 PIX2651_IN
port 2694 n
rlabel metal5 18520 -48980 18620 -48880 1 PIX2652_IN
port 2695 n
rlabel metal5 20020 -48980 20120 -48880 1 PIX2653_IN
port 2696 n
rlabel metal5 21520 -48980 21620 -48880 1 PIX2654_IN
port 2697 n
rlabel metal5 23020 -48980 23120 -48880 1 PIX2655_IN
port 2698 n
rlabel metal5 24520 -48980 24620 -48880 1 PIX2656_IN
port 2699 n
rlabel metal5 26020 -48980 26120 -48880 1 PIX2657_IN
port 2700 n
rlabel metal5 27520 -48980 27620 -48880 1 PIX2658_IN
port 2701 n
rlabel metal5 29020 -48980 29120 -48880 1 PIX2659_IN
port 2702 n
rlabel metal5 30520 -48980 30620 -48880 1 PIX2660_IN
port 2703 n
rlabel metal5 32020 -48980 32120 -48880 1 PIX2661_IN
port 2704 n
rlabel metal5 33520 -48980 33620 -48880 1 PIX2662_IN
port 2705 n
rlabel metal5 35020 -48980 35120 -48880 1 PIX2663_IN
port 2706 n
rlabel metal5 36520 -48980 36620 -48880 1 PIX2664_IN
port 2707 n
rlabel metal5 38020 -48980 38120 -48880 1 PIX2665_IN
port 2708 n
rlabel metal5 39520 -48980 39620 -48880 1 PIX2666_IN
port 2709 n
rlabel metal5 41020 -48980 41120 -48880 1 PIX2667_IN
port 2710 n
rlabel metal5 42520 -48980 42620 -48880 1 PIX2668_IN
port 2711 n
rlabel metal5 44020 -48980 44120 -48880 1 PIX2669_IN
port 2712 n
rlabel metal5 45520 -48980 45620 -48880 1 PIX2670_IN
port 2713 n
rlabel metal5 47020 -48980 47120 -48880 1 PIX2671_IN
port 2714 n
rlabel metal5 48520 -48980 48620 -48880 1 PIX2672_IN
port 2715 n
rlabel metal5 50020 -48980 50120 -48880 1 PIX2673_IN
port 2716 n
rlabel metal5 51520 -48980 51620 -48880 1 PIX2674_IN
port 2717 n
rlabel metal5 53020 -48980 53120 -48880 1 PIX2675_IN
port 2718 n
rlabel metal5 54520 -48980 54620 -48880 1 PIX2676_IN
port 2719 n
rlabel metal5 56020 -48980 56120 -48880 1 PIX2677_IN
port 2720 n
rlabel metal5 57520 -48980 57620 -48880 1 PIX2678_IN
port 2721 n
rlabel metal5 59020 -48980 59120 -48880 1 PIX2679_IN
port 2722 n
rlabel metal5 60520 -48980 60620 -48880 1 PIX2680_IN
port 2723 n
rlabel metal5 62020 -48980 62120 -48880 1 PIX2681_IN
port 2724 n
rlabel metal5 63520 -48980 63620 -48880 1 PIX2682_IN
port 2725 n
rlabel metal5 65020 -48980 65120 -48880 1 PIX2683_IN
port 2726 n
rlabel metal5 66520 -48980 66620 -48880 1 PIX2684_IN
port 2727 n
rlabel metal5 68020 -48980 68120 -48880 1 PIX2685_IN
port 2728 n
rlabel metal5 69520 -48980 69620 -48880 1 PIX2686_IN
port 2729 n
rlabel metal5 71020 -48980 71120 -48880 1 PIX2687_IN
port 2730 n
rlabel metal5 72520 -48980 72620 -48880 1 PIX2688_IN
port 2731 n
rlabel metal5 74020 -48980 74120 -48880 1 PIX2689_IN
port 2732 n
rlabel metal5 75520 -48980 75620 -48880 1 PIX2690_IN
port 2733 n
rlabel metal5 77020 -48980 77120 -48880 1 PIX2691_IN
port 2734 n
rlabel metal5 78520 -48980 78620 -48880 1 PIX2692_IN
port 2735 n
rlabel metal5 80020 -48980 80120 -48880 1 PIX2693_IN
port 2736 n
rlabel metal5 81520 -48980 81620 -48880 1 PIX2694_IN
port 2737 n
rlabel metal5 83020 -48980 83120 -48880 1 PIX2695_IN
port 2738 n
rlabel metal5 84520 -48980 84620 -48880 1 PIX2696_IN
port 2739 n
rlabel metal5 86020 -48980 86120 -48880 1 PIX2697_IN
port 2740 n
rlabel metal5 87520 -48980 87620 -48880 1 PIX2698_IN
port 2741 n
rlabel metal5 89020 -48980 89120 -48880 1 PIX2699_IN
port 2742 n
rlabel metal5 90520 -48980 90620 -48880 1 PIX2700_IN
port 2743 n
rlabel metal5 92020 -48980 92120 -48880 1 PIX2701_IN
port 2744 n
rlabel metal5 93520 -48980 93620 -48880 1 PIX2702_IN
port 2745 n
rlabel metal5 95020 -48980 95120 -48880 1 PIX2703_IN
port 2746 n
rlabel metal5 96520 -48980 96620 -48880 1 PIX2704_IN
port 2747 n
rlabel metal5 98020 -48980 98120 -48880 1 PIX2705_IN
port 2748 n
rlabel metal5 99520 -48980 99620 -48880 1 PIX2706_IN
port 2749 n
rlabel metal5 101020 -48980 101120 -48880 1 PIX2707_IN
port 2750 n
rlabel metal5 102520 -48980 102620 -48880 1 PIX2708_IN
port 2751 n
rlabel metal5 104020 -48980 104120 -48880 1 PIX2709_IN
port 2752 n
rlabel metal5 105520 -48980 105620 -48880 1 PIX2710_IN
port 2753 n
rlabel metal5 107020 -48980 107120 -48880 1 PIX2711_IN
port 2754 n
rlabel metal5 108520 -48980 108620 -48880 1 PIX2712_IN
port 2755 n
rlabel metal5 110020 -48980 110120 -48880 1 PIX2713_IN
port 2756 n
rlabel metal5 111520 -48980 111620 -48880 1 PIX2714_IN
port 2757 n
rlabel metal5 113020 -48980 113120 -48880 1 PIX2715_IN
port 2758 n
rlabel metal5 114520 -48980 114620 -48880 1 PIX2716_IN
port 2759 n
rlabel metal5 116020 -48980 116120 -48880 1 PIX2717_IN
port 2760 n
rlabel metal5 117520 -48980 117620 -48880 1 PIX2718_IN
port 2761 n
rlabel metal5 119020 -48980 119120 -48880 1 PIX2719_IN
port 2762 n
rlabel metal5 520 -50480 620 -50380 1 PIX2720_IN
port 2763 n
rlabel metal2 -1500 -50260 -1500 -50215 3 ROW_SEL34
port 2764 e
rlabel metal5 2020 -50480 2120 -50380 1 PIX2721_IN
port 2765 n
rlabel metal5 3520 -50480 3620 -50380 1 PIX2722_IN
port 2766 n
rlabel metal5 5020 -50480 5120 -50380 1 PIX2723_IN
port 2767 n
rlabel metal5 6520 -50480 6620 -50380 1 PIX2724_IN
port 2768 n
rlabel metal5 8020 -50480 8120 -50380 1 PIX2725_IN
port 2769 n
rlabel metal5 9520 -50480 9620 -50380 1 PIX2726_IN
port 2770 n
rlabel metal5 11020 -50480 11120 -50380 1 PIX2727_IN
port 2771 n
rlabel metal5 12520 -50480 12620 -50380 1 PIX2728_IN
port 2772 n
rlabel metal5 14020 -50480 14120 -50380 1 PIX2729_IN
port 2773 n
rlabel metal5 15520 -50480 15620 -50380 1 PIX2730_IN
port 2774 n
rlabel metal5 17020 -50480 17120 -50380 1 PIX2731_IN
port 2775 n
rlabel metal5 18520 -50480 18620 -50380 1 PIX2732_IN
port 2776 n
rlabel metal5 20020 -50480 20120 -50380 1 PIX2733_IN
port 2777 n
rlabel metal5 21520 -50480 21620 -50380 1 PIX2734_IN
port 2778 n
rlabel metal5 23020 -50480 23120 -50380 1 PIX2735_IN
port 2779 n
rlabel metal5 24520 -50480 24620 -50380 1 PIX2736_IN
port 2780 n
rlabel metal5 26020 -50480 26120 -50380 1 PIX2737_IN
port 2781 n
rlabel metal5 27520 -50480 27620 -50380 1 PIX2738_IN
port 2782 n
rlabel metal5 29020 -50480 29120 -50380 1 PIX2739_IN
port 2783 n
rlabel metal5 30520 -50480 30620 -50380 1 PIX2740_IN
port 2784 n
rlabel metal5 32020 -50480 32120 -50380 1 PIX2741_IN
port 2785 n
rlabel metal5 33520 -50480 33620 -50380 1 PIX2742_IN
port 2786 n
rlabel metal5 35020 -50480 35120 -50380 1 PIX2743_IN
port 2787 n
rlabel metal5 36520 -50480 36620 -50380 1 PIX2744_IN
port 2788 n
rlabel metal5 38020 -50480 38120 -50380 1 PIX2745_IN
port 2789 n
rlabel metal5 39520 -50480 39620 -50380 1 PIX2746_IN
port 2790 n
rlabel metal5 41020 -50480 41120 -50380 1 PIX2747_IN
port 2791 n
rlabel metal5 42520 -50480 42620 -50380 1 PIX2748_IN
port 2792 n
rlabel metal5 44020 -50480 44120 -50380 1 PIX2749_IN
port 2793 n
rlabel metal5 45520 -50480 45620 -50380 1 PIX2750_IN
port 2794 n
rlabel metal5 47020 -50480 47120 -50380 1 PIX2751_IN
port 2795 n
rlabel metal5 48520 -50480 48620 -50380 1 PIX2752_IN
port 2796 n
rlabel metal5 50020 -50480 50120 -50380 1 PIX2753_IN
port 2797 n
rlabel metal5 51520 -50480 51620 -50380 1 PIX2754_IN
port 2798 n
rlabel metal5 53020 -50480 53120 -50380 1 PIX2755_IN
port 2799 n
rlabel metal5 54520 -50480 54620 -50380 1 PIX2756_IN
port 2800 n
rlabel metal5 56020 -50480 56120 -50380 1 PIX2757_IN
port 2801 n
rlabel metal5 57520 -50480 57620 -50380 1 PIX2758_IN
port 2802 n
rlabel metal5 59020 -50480 59120 -50380 1 PIX2759_IN
port 2803 n
rlabel metal5 60520 -50480 60620 -50380 1 PIX2760_IN
port 2804 n
rlabel metal5 62020 -50480 62120 -50380 1 PIX2761_IN
port 2805 n
rlabel metal5 63520 -50480 63620 -50380 1 PIX2762_IN
port 2806 n
rlabel metal5 65020 -50480 65120 -50380 1 PIX2763_IN
port 2807 n
rlabel metal5 66520 -50480 66620 -50380 1 PIX2764_IN
port 2808 n
rlabel metal5 68020 -50480 68120 -50380 1 PIX2765_IN
port 2809 n
rlabel metal5 69520 -50480 69620 -50380 1 PIX2766_IN
port 2810 n
rlabel metal5 71020 -50480 71120 -50380 1 PIX2767_IN
port 2811 n
rlabel metal5 72520 -50480 72620 -50380 1 PIX2768_IN
port 2812 n
rlabel metal5 74020 -50480 74120 -50380 1 PIX2769_IN
port 2813 n
rlabel metal5 75520 -50480 75620 -50380 1 PIX2770_IN
port 2814 n
rlabel metal5 77020 -50480 77120 -50380 1 PIX2771_IN
port 2815 n
rlabel metal5 78520 -50480 78620 -50380 1 PIX2772_IN
port 2816 n
rlabel metal5 80020 -50480 80120 -50380 1 PIX2773_IN
port 2817 n
rlabel metal5 81520 -50480 81620 -50380 1 PIX2774_IN
port 2818 n
rlabel metal5 83020 -50480 83120 -50380 1 PIX2775_IN
port 2819 n
rlabel metal5 84520 -50480 84620 -50380 1 PIX2776_IN
port 2820 n
rlabel metal5 86020 -50480 86120 -50380 1 PIX2777_IN
port 2821 n
rlabel metal5 87520 -50480 87620 -50380 1 PIX2778_IN
port 2822 n
rlabel metal5 89020 -50480 89120 -50380 1 PIX2779_IN
port 2823 n
rlabel metal5 90520 -50480 90620 -50380 1 PIX2780_IN
port 2824 n
rlabel metal5 92020 -50480 92120 -50380 1 PIX2781_IN
port 2825 n
rlabel metal5 93520 -50480 93620 -50380 1 PIX2782_IN
port 2826 n
rlabel metal5 95020 -50480 95120 -50380 1 PIX2783_IN
port 2827 n
rlabel metal5 96520 -50480 96620 -50380 1 PIX2784_IN
port 2828 n
rlabel metal5 98020 -50480 98120 -50380 1 PIX2785_IN
port 2829 n
rlabel metal5 99520 -50480 99620 -50380 1 PIX2786_IN
port 2830 n
rlabel metal5 101020 -50480 101120 -50380 1 PIX2787_IN
port 2831 n
rlabel metal5 102520 -50480 102620 -50380 1 PIX2788_IN
port 2832 n
rlabel metal5 104020 -50480 104120 -50380 1 PIX2789_IN
port 2833 n
rlabel metal5 105520 -50480 105620 -50380 1 PIX2790_IN
port 2834 n
rlabel metal5 107020 -50480 107120 -50380 1 PIX2791_IN
port 2835 n
rlabel metal5 108520 -50480 108620 -50380 1 PIX2792_IN
port 2836 n
rlabel metal5 110020 -50480 110120 -50380 1 PIX2793_IN
port 2837 n
rlabel metal5 111520 -50480 111620 -50380 1 PIX2794_IN
port 2838 n
rlabel metal5 113020 -50480 113120 -50380 1 PIX2795_IN
port 2839 n
rlabel metal5 114520 -50480 114620 -50380 1 PIX2796_IN
port 2840 n
rlabel metal5 116020 -50480 116120 -50380 1 PIX2797_IN
port 2841 n
rlabel metal5 117520 -50480 117620 -50380 1 PIX2798_IN
port 2842 n
rlabel metal5 119020 -50480 119120 -50380 1 PIX2799_IN
port 2843 n
rlabel metal5 520 -51980 620 -51880 1 PIX2800_IN
port 2844 n
rlabel metal2 -1500 -51760 -1500 -51715 3 ROW_SEL35
port 2845 e
rlabel metal5 2020 -51980 2120 -51880 1 PIX2801_IN
port 2846 n
rlabel metal5 3520 -51980 3620 -51880 1 PIX2802_IN
port 2847 n
rlabel metal5 5020 -51980 5120 -51880 1 PIX2803_IN
port 2848 n
rlabel metal5 6520 -51980 6620 -51880 1 PIX2804_IN
port 2849 n
rlabel metal5 8020 -51980 8120 -51880 1 PIX2805_IN
port 2850 n
rlabel metal5 9520 -51980 9620 -51880 1 PIX2806_IN
port 2851 n
rlabel metal5 11020 -51980 11120 -51880 1 PIX2807_IN
port 2852 n
rlabel metal5 12520 -51980 12620 -51880 1 PIX2808_IN
port 2853 n
rlabel metal5 14020 -51980 14120 -51880 1 PIX2809_IN
port 2854 n
rlabel metal5 15520 -51980 15620 -51880 1 PIX2810_IN
port 2855 n
rlabel metal5 17020 -51980 17120 -51880 1 PIX2811_IN
port 2856 n
rlabel metal5 18520 -51980 18620 -51880 1 PIX2812_IN
port 2857 n
rlabel metal5 20020 -51980 20120 -51880 1 PIX2813_IN
port 2858 n
rlabel metal5 21520 -51980 21620 -51880 1 PIX2814_IN
port 2859 n
rlabel metal5 23020 -51980 23120 -51880 1 PIX2815_IN
port 2860 n
rlabel metal5 24520 -51980 24620 -51880 1 PIX2816_IN
port 2861 n
rlabel metal5 26020 -51980 26120 -51880 1 PIX2817_IN
port 2862 n
rlabel metal5 27520 -51980 27620 -51880 1 PIX2818_IN
port 2863 n
rlabel metal5 29020 -51980 29120 -51880 1 PIX2819_IN
port 2864 n
rlabel metal5 30520 -51980 30620 -51880 1 PIX2820_IN
port 2865 n
rlabel metal5 32020 -51980 32120 -51880 1 PIX2821_IN
port 2866 n
rlabel metal5 33520 -51980 33620 -51880 1 PIX2822_IN
port 2867 n
rlabel metal5 35020 -51980 35120 -51880 1 PIX2823_IN
port 2868 n
rlabel metal5 36520 -51980 36620 -51880 1 PIX2824_IN
port 2869 n
rlabel metal5 38020 -51980 38120 -51880 1 PIX2825_IN
port 2870 n
rlabel metal5 39520 -51980 39620 -51880 1 PIX2826_IN
port 2871 n
rlabel metal5 41020 -51980 41120 -51880 1 PIX2827_IN
port 2872 n
rlabel metal5 42520 -51980 42620 -51880 1 PIX2828_IN
port 2873 n
rlabel metal5 44020 -51980 44120 -51880 1 PIX2829_IN
port 2874 n
rlabel metal5 45520 -51980 45620 -51880 1 PIX2830_IN
port 2875 n
rlabel metal5 47020 -51980 47120 -51880 1 PIX2831_IN
port 2876 n
rlabel metal5 48520 -51980 48620 -51880 1 PIX2832_IN
port 2877 n
rlabel metal5 50020 -51980 50120 -51880 1 PIX2833_IN
port 2878 n
rlabel metal5 51520 -51980 51620 -51880 1 PIX2834_IN
port 2879 n
rlabel metal5 53020 -51980 53120 -51880 1 PIX2835_IN
port 2880 n
rlabel metal5 54520 -51980 54620 -51880 1 PIX2836_IN
port 2881 n
rlabel metal5 56020 -51980 56120 -51880 1 PIX2837_IN
port 2882 n
rlabel metal5 57520 -51980 57620 -51880 1 PIX2838_IN
port 2883 n
rlabel metal5 59020 -51980 59120 -51880 1 PIX2839_IN
port 2884 n
rlabel metal5 60520 -51980 60620 -51880 1 PIX2840_IN
port 2885 n
rlabel metal5 62020 -51980 62120 -51880 1 PIX2841_IN
port 2886 n
rlabel metal5 63520 -51980 63620 -51880 1 PIX2842_IN
port 2887 n
rlabel metal5 65020 -51980 65120 -51880 1 PIX2843_IN
port 2888 n
rlabel metal5 66520 -51980 66620 -51880 1 PIX2844_IN
port 2889 n
rlabel metal5 68020 -51980 68120 -51880 1 PIX2845_IN
port 2890 n
rlabel metal5 69520 -51980 69620 -51880 1 PIX2846_IN
port 2891 n
rlabel metal5 71020 -51980 71120 -51880 1 PIX2847_IN
port 2892 n
rlabel metal5 72520 -51980 72620 -51880 1 PIX2848_IN
port 2893 n
rlabel metal5 74020 -51980 74120 -51880 1 PIX2849_IN
port 2894 n
rlabel metal5 75520 -51980 75620 -51880 1 PIX2850_IN
port 2895 n
rlabel metal5 77020 -51980 77120 -51880 1 PIX2851_IN
port 2896 n
rlabel metal5 78520 -51980 78620 -51880 1 PIX2852_IN
port 2897 n
rlabel metal5 80020 -51980 80120 -51880 1 PIX2853_IN
port 2898 n
rlabel metal5 81520 -51980 81620 -51880 1 PIX2854_IN
port 2899 n
rlabel metal5 83020 -51980 83120 -51880 1 PIX2855_IN
port 2900 n
rlabel metal5 84520 -51980 84620 -51880 1 PIX2856_IN
port 2901 n
rlabel metal5 86020 -51980 86120 -51880 1 PIX2857_IN
port 2902 n
rlabel metal5 87520 -51980 87620 -51880 1 PIX2858_IN
port 2903 n
rlabel metal5 89020 -51980 89120 -51880 1 PIX2859_IN
port 2904 n
rlabel metal5 90520 -51980 90620 -51880 1 PIX2860_IN
port 2905 n
rlabel metal5 92020 -51980 92120 -51880 1 PIX2861_IN
port 2906 n
rlabel metal5 93520 -51980 93620 -51880 1 PIX2862_IN
port 2907 n
rlabel metal5 95020 -51980 95120 -51880 1 PIX2863_IN
port 2908 n
rlabel metal5 96520 -51980 96620 -51880 1 PIX2864_IN
port 2909 n
rlabel metal5 98020 -51980 98120 -51880 1 PIX2865_IN
port 2910 n
rlabel metal5 99520 -51980 99620 -51880 1 PIX2866_IN
port 2911 n
rlabel metal5 101020 -51980 101120 -51880 1 PIX2867_IN
port 2912 n
rlabel metal5 102520 -51980 102620 -51880 1 PIX2868_IN
port 2913 n
rlabel metal5 104020 -51980 104120 -51880 1 PIX2869_IN
port 2914 n
rlabel metal5 105520 -51980 105620 -51880 1 PIX2870_IN
port 2915 n
rlabel metal5 107020 -51980 107120 -51880 1 PIX2871_IN
port 2916 n
rlabel metal5 108520 -51980 108620 -51880 1 PIX2872_IN
port 2917 n
rlabel metal5 110020 -51980 110120 -51880 1 PIX2873_IN
port 2918 n
rlabel metal5 111520 -51980 111620 -51880 1 PIX2874_IN
port 2919 n
rlabel metal5 113020 -51980 113120 -51880 1 PIX2875_IN
port 2920 n
rlabel metal5 114520 -51980 114620 -51880 1 PIX2876_IN
port 2921 n
rlabel metal5 116020 -51980 116120 -51880 1 PIX2877_IN
port 2922 n
rlabel metal5 117520 -51980 117620 -51880 1 PIX2878_IN
port 2923 n
rlabel metal5 119020 -51980 119120 -51880 1 PIX2879_IN
port 2924 n
rlabel metal5 520 -53480 620 -53380 1 PIX2880_IN
port 2925 n
rlabel metal2 -1500 -53260 -1500 -53215 3 ROW_SEL36
port 2926 e
rlabel metal5 2020 -53480 2120 -53380 1 PIX2881_IN
port 2927 n
rlabel metal5 3520 -53480 3620 -53380 1 PIX2882_IN
port 2928 n
rlabel metal5 5020 -53480 5120 -53380 1 PIX2883_IN
port 2929 n
rlabel metal5 6520 -53480 6620 -53380 1 PIX2884_IN
port 2930 n
rlabel metal5 8020 -53480 8120 -53380 1 PIX2885_IN
port 2931 n
rlabel metal5 9520 -53480 9620 -53380 1 PIX2886_IN
port 2932 n
rlabel metal5 11020 -53480 11120 -53380 1 PIX2887_IN
port 2933 n
rlabel metal5 12520 -53480 12620 -53380 1 PIX2888_IN
port 2934 n
rlabel metal5 14020 -53480 14120 -53380 1 PIX2889_IN
port 2935 n
rlabel metal5 15520 -53480 15620 -53380 1 PIX2890_IN
port 2936 n
rlabel metal5 17020 -53480 17120 -53380 1 PIX2891_IN
port 2937 n
rlabel metal5 18520 -53480 18620 -53380 1 PIX2892_IN
port 2938 n
rlabel metal5 20020 -53480 20120 -53380 1 PIX2893_IN
port 2939 n
rlabel metal5 21520 -53480 21620 -53380 1 PIX2894_IN
port 2940 n
rlabel metal5 23020 -53480 23120 -53380 1 PIX2895_IN
port 2941 n
rlabel metal5 24520 -53480 24620 -53380 1 PIX2896_IN
port 2942 n
rlabel metal5 26020 -53480 26120 -53380 1 PIX2897_IN
port 2943 n
rlabel metal5 27520 -53480 27620 -53380 1 PIX2898_IN
port 2944 n
rlabel metal5 29020 -53480 29120 -53380 1 PIX2899_IN
port 2945 n
rlabel metal5 30520 -53480 30620 -53380 1 PIX2900_IN
port 2946 n
rlabel metal5 32020 -53480 32120 -53380 1 PIX2901_IN
port 2947 n
rlabel metal5 33520 -53480 33620 -53380 1 PIX2902_IN
port 2948 n
rlabel metal5 35020 -53480 35120 -53380 1 PIX2903_IN
port 2949 n
rlabel metal5 36520 -53480 36620 -53380 1 PIX2904_IN
port 2950 n
rlabel metal5 38020 -53480 38120 -53380 1 PIX2905_IN
port 2951 n
rlabel metal5 39520 -53480 39620 -53380 1 PIX2906_IN
port 2952 n
rlabel metal5 41020 -53480 41120 -53380 1 PIX2907_IN
port 2953 n
rlabel metal5 42520 -53480 42620 -53380 1 PIX2908_IN
port 2954 n
rlabel metal5 44020 -53480 44120 -53380 1 PIX2909_IN
port 2955 n
rlabel metal5 45520 -53480 45620 -53380 1 PIX2910_IN
port 2956 n
rlabel metal5 47020 -53480 47120 -53380 1 PIX2911_IN
port 2957 n
rlabel metal5 48520 -53480 48620 -53380 1 PIX2912_IN
port 2958 n
rlabel metal5 50020 -53480 50120 -53380 1 PIX2913_IN
port 2959 n
rlabel metal5 51520 -53480 51620 -53380 1 PIX2914_IN
port 2960 n
rlabel metal5 53020 -53480 53120 -53380 1 PIX2915_IN
port 2961 n
rlabel metal5 54520 -53480 54620 -53380 1 PIX2916_IN
port 2962 n
rlabel metal5 56020 -53480 56120 -53380 1 PIX2917_IN
port 2963 n
rlabel metal5 57520 -53480 57620 -53380 1 PIX2918_IN
port 2964 n
rlabel metal5 59020 -53480 59120 -53380 1 PIX2919_IN
port 2965 n
rlabel metal5 60520 -53480 60620 -53380 1 PIX2920_IN
port 2966 n
rlabel metal5 62020 -53480 62120 -53380 1 PIX2921_IN
port 2967 n
rlabel metal5 63520 -53480 63620 -53380 1 PIX2922_IN
port 2968 n
rlabel metal5 65020 -53480 65120 -53380 1 PIX2923_IN
port 2969 n
rlabel metal5 66520 -53480 66620 -53380 1 PIX2924_IN
port 2970 n
rlabel metal5 68020 -53480 68120 -53380 1 PIX2925_IN
port 2971 n
rlabel metal5 69520 -53480 69620 -53380 1 PIX2926_IN
port 2972 n
rlabel metal5 71020 -53480 71120 -53380 1 PIX2927_IN
port 2973 n
rlabel metal5 72520 -53480 72620 -53380 1 PIX2928_IN
port 2974 n
rlabel metal5 74020 -53480 74120 -53380 1 PIX2929_IN
port 2975 n
rlabel metal5 75520 -53480 75620 -53380 1 PIX2930_IN
port 2976 n
rlabel metal5 77020 -53480 77120 -53380 1 PIX2931_IN
port 2977 n
rlabel metal5 78520 -53480 78620 -53380 1 PIX2932_IN
port 2978 n
rlabel metal5 80020 -53480 80120 -53380 1 PIX2933_IN
port 2979 n
rlabel metal5 81520 -53480 81620 -53380 1 PIX2934_IN
port 2980 n
rlabel metal5 83020 -53480 83120 -53380 1 PIX2935_IN
port 2981 n
rlabel metal5 84520 -53480 84620 -53380 1 PIX2936_IN
port 2982 n
rlabel metal5 86020 -53480 86120 -53380 1 PIX2937_IN
port 2983 n
rlabel metal5 87520 -53480 87620 -53380 1 PIX2938_IN
port 2984 n
rlabel metal5 89020 -53480 89120 -53380 1 PIX2939_IN
port 2985 n
rlabel metal5 90520 -53480 90620 -53380 1 PIX2940_IN
port 2986 n
rlabel metal5 92020 -53480 92120 -53380 1 PIX2941_IN
port 2987 n
rlabel metal5 93520 -53480 93620 -53380 1 PIX2942_IN
port 2988 n
rlabel metal5 95020 -53480 95120 -53380 1 PIX2943_IN
port 2989 n
rlabel metal5 96520 -53480 96620 -53380 1 PIX2944_IN
port 2990 n
rlabel metal5 98020 -53480 98120 -53380 1 PIX2945_IN
port 2991 n
rlabel metal5 99520 -53480 99620 -53380 1 PIX2946_IN
port 2992 n
rlabel metal5 101020 -53480 101120 -53380 1 PIX2947_IN
port 2993 n
rlabel metal5 102520 -53480 102620 -53380 1 PIX2948_IN
port 2994 n
rlabel metal5 104020 -53480 104120 -53380 1 PIX2949_IN
port 2995 n
rlabel metal5 105520 -53480 105620 -53380 1 PIX2950_IN
port 2996 n
rlabel metal5 107020 -53480 107120 -53380 1 PIX2951_IN
port 2997 n
rlabel metal5 108520 -53480 108620 -53380 1 PIX2952_IN
port 2998 n
rlabel metal5 110020 -53480 110120 -53380 1 PIX2953_IN
port 2999 n
rlabel metal5 111520 -53480 111620 -53380 1 PIX2954_IN
port 3000 n
rlabel metal5 113020 -53480 113120 -53380 1 PIX2955_IN
port 3001 n
rlabel metal5 114520 -53480 114620 -53380 1 PIX2956_IN
port 3002 n
rlabel metal5 116020 -53480 116120 -53380 1 PIX2957_IN
port 3003 n
rlabel metal5 117520 -53480 117620 -53380 1 PIX2958_IN
port 3004 n
rlabel metal5 119020 -53480 119120 -53380 1 PIX2959_IN
port 3005 n
rlabel metal5 520 -54980 620 -54880 1 PIX2960_IN
port 3006 n
rlabel metal2 -1500 -54760 -1500 -54715 3 ROW_SEL37
port 3007 e
rlabel metal5 2020 -54980 2120 -54880 1 PIX2961_IN
port 3008 n
rlabel metal5 3520 -54980 3620 -54880 1 PIX2962_IN
port 3009 n
rlabel metal5 5020 -54980 5120 -54880 1 PIX2963_IN
port 3010 n
rlabel metal5 6520 -54980 6620 -54880 1 PIX2964_IN
port 3011 n
rlabel metal5 8020 -54980 8120 -54880 1 PIX2965_IN
port 3012 n
rlabel metal5 9520 -54980 9620 -54880 1 PIX2966_IN
port 3013 n
rlabel metal5 11020 -54980 11120 -54880 1 PIX2967_IN
port 3014 n
rlabel metal5 12520 -54980 12620 -54880 1 PIX2968_IN
port 3015 n
rlabel metal5 14020 -54980 14120 -54880 1 PIX2969_IN
port 3016 n
rlabel metal5 15520 -54980 15620 -54880 1 PIX2970_IN
port 3017 n
rlabel metal5 17020 -54980 17120 -54880 1 PIX2971_IN
port 3018 n
rlabel metal5 18520 -54980 18620 -54880 1 PIX2972_IN
port 3019 n
rlabel metal5 20020 -54980 20120 -54880 1 PIX2973_IN
port 3020 n
rlabel metal5 21520 -54980 21620 -54880 1 PIX2974_IN
port 3021 n
rlabel metal5 23020 -54980 23120 -54880 1 PIX2975_IN
port 3022 n
rlabel metal5 24520 -54980 24620 -54880 1 PIX2976_IN
port 3023 n
rlabel metal5 26020 -54980 26120 -54880 1 PIX2977_IN
port 3024 n
rlabel metal5 27520 -54980 27620 -54880 1 PIX2978_IN
port 3025 n
rlabel metal5 29020 -54980 29120 -54880 1 PIX2979_IN
port 3026 n
rlabel metal5 30520 -54980 30620 -54880 1 PIX2980_IN
port 3027 n
rlabel metal5 32020 -54980 32120 -54880 1 PIX2981_IN
port 3028 n
rlabel metal5 33520 -54980 33620 -54880 1 PIX2982_IN
port 3029 n
rlabel metal5 35020 -54980 35120 -54880 1 PIX2983_IN
port 3030 n
rlabel metal5 36520 -54980 36620 -54880 1 PIX2984_IN
port 3031 n
rlabel metal5 38020 -54980 38120 -54880 1 PIX2985_IN
port 3032 n
rlabel metal5 39520 -54980 39620 -54880 1 PIX2986_IN
port 3033 n
rlabel metal5 41020 -54980 41120 -54880 1 PIX2987_IN
port 3034 n
rlabel metal5 42520 -54980 42620 -54880 1 PIX2988_IN
port 3035 n
rlabel metal5 44020 -54980 44120 -54880 1 PIX2989_IN
port 3036 n
rlabel metal5 45520 -54980 45620 -54880 1 PIX2990_IN
port 3037 n
rlabel metal5 47020 -54980 47120 -54880 1 PIX2991_IN
port 3038 n
rlabel metal5 48520 -54980 48620 -54880 1 PIX2992_IN
port 3039 n
rlabel metal5 50020 -54980 50120 -54880 1 PIX2993_IN
port 3040 n
rlabel metal5 51520 -54980 51620 -54880 1 PIX2994_IN
port 3041 n
rlabel metal5 53020 -54980 53120 -54880 1 PIX2995_IN
port 3042 n
rlabel metal5 54520 -54980 54620 -54880 1 PIX2996_IN
port 3043 n
rlabel metal5 56020 -54980 56120 -54880 1 PIX2997_IN
port 3044 n
rlabel metal5 57520 -54980 57620 -54880 1 PIX2998_IN
port 3045 n
rlabel metal5 59020 -54980 59120 -54880 1 PIX2999_IN
port 3046 n
rlabel metal5 60520 -54980 60620 -54880 1 PIX3000_IN
port 3047 n
rlabel metal5 62020 -54980 62120 -54880 1 PIX3001_IN
port 3048 n
rlabel metal5 63520 -54980 63620 -54880 1 PIX3002_IN
port 3049 n
rlabel metal5 65020 -54980 65120 -54880 1 PIX3003_IN
port 3050 n
rlabel metal5 66520 -54980 66620 -54880 1 PIX3004_IN
port 3051 n
rlabel metal5 68020 -54980 68120 -54880 1 PIX3005_IN
port 3052 n
rlabel metal5 69520 -54980 69620 -54880 1 PIX3006_IN
port 3053 n
rlabel metal5 71020 -54980 71120 -54880 1 PIX3007_IN
port 3054 n
rlabel metal5 72520 -54980 72620 -54880 1 PIX3008_IN
port 3055 n
rlabel metal5 74020 -54980 74120 -54880 1 PIX3009_IN
port 3056 n
rlabel metal5 75520 -54980 75620 -54880 1 PIX3010_IN
port 3057 n
rlabel metal5 77020 -54980 77120 -54880 1 PIX3011_IN
port 3058 n
rlabel metal5 78520 -54980 78620 -54880 1 PIX3012_IN
port 3059 n
rlabel metal5 80020 -54980 80120 -54880 1 PIX3013_IN
port 3060 n
rlabel metal5 81520 -54980 81620 -54880 1 PIX3014_IN
port 3061 n
rlabel metal5 83020 -54980 83120 -54880 1 PIX3015_IN
port 3062 n
rlabel metal5 84520 -54980 84620 -54880 1 PIX3016_IN
port 3063 n
rlabel metal5 86020 -54980 86120 -54880 1 PIX3017_IN
port 3064 n
rlabel metal5 87520 -54980 87620 -54880 1 PIX3018_IN
port 3065 n
rlabel metal5 89020 -54980 89120 -54880 1 PIX3019_IN
port 3066 n
rlabel metal5 90520 -54980 90620 -54880 1 PIX3020_IN
port 3067 n
rlabel metal5 92020 -54980 92120 -54880 1 PIX3021_IN
port 3068 n
rlabel metal5 93520 -54980 93620 -54880 1 PIX3022_IN
port 3069 n
rlabel metal5 95020 -54980 95120 -54880 1 PIX3023_IN
port 3070 n
rlabel metal5 96520 -54980 96620 -54880 1 PIX3024_IN
port 3071 n
rlabel metal5 98020 -54980 98120 -54880 1 PIX3025_IN
port 3072 n
rlabel metal5 99520 -54980 99620 -54880 1 PIX3026_IN
port 3073 n
rlabel metal5 101020 -54980 101120 -54880 1 PIX3027_IN
port 3074 n
rlabel metal5 102520 -54980 102620 -54880 1 PIX3028_IN
port 3075 n
rlabel metal5 104020 -54980 104120 -54880 1 PIX3029_IN
port 3076 n
rlabel metal5 105520 -54980 105620 -54880 1 PIX3030_IN
port 3077 n
rlabel metal5 107020 -54980 107120 -54880 1 PIX3031_IN
port 3078 n
rlabel metal5 108520 -54980 108620 -54880 1 PIX3032_IN
port 3079 n
rlabel metal5 110020 -54980 110120 -54880 1 PIX3033_IN
port 3080 n
rlabel metal5 111520 -54980 111620 -54880 1 PIX3034_IN
port 3081 n
rlabel metal5 113020 -54980 113120 -54880 1 PIX3035_IN
port 3082 n
rlabel metal5 114520 -54980 114620 -54880 1 PIX3036_IN
port 3083 n
rlabel metal5 116020 -54980 116120 -54880 1 PIX3037_IN
port 3084 n
rlabel metal5 117520 -54980 117620 -54880 1 PIX3038_IN
port 3085 n
rlabel metal5 119020 -54980 119120 -54880 1 PIX3039_IN
port 3086 n
rlabel metal5 520 -56480 620 -56380 1 PIX3040_IN
port 3087 n
rlabel metal2 -1500 -56260 -1500 -56215 3 ROW_SEL38
port 3088 e
rlabel metal5 2020 -56480 2120 -56380 1 PIX3041_IN
port 3089 n
rlabel metal5 3520 -56480 3620 -56380 1 PIX3042_IN
port 3090 n
rlabel metal5 5020 -56480 5120 -56380 1 PIX3043_IN
port 3091 n
rlabel metal5 6520 -56480 6620 -56380 1 PIX3044_IN
port 3092 n
rlabel metal5 8020 -56480 8120 -56380 1 PIX3045_IN
port 3093 n
rlabel metal5 9520 -56480 9620 -56380 1 PIX3046_IN
port 3094 n
rlabel metal5 11020 -56480 11120 -56380 1 PIX3047_IN
port 3095 n
rlabel metal5 12520 -56480 12620 -56380 1 PIX3048_IN
port 3096 n
rlabel metal5 14020 -56480 14120 -56380 1 PIX3049_IN
port 3097 n
rlabel metal5 15520 -56480 15620 -56380 1 PIX3050_IN
port 3098 n
rlabel metal5 17020 -56480 17120 -56380 1 PIX3051_IN
port 3099 n
rlabel metal5 18520 -56480 18620 -56380 1 PIX3052_IN
port 3100 n
rlabel metal5 20020 -56480 20120 -56380 1 PIX3053_IN
port 3101 n
rlabel metal5 21520 -56480 21620 -56380 1 PIX3054_IN
port 3102 n
rlabel metal5 23020 -56480 23120 -56380 1 PIX3055_IN
port 3103 n
rlabel metal5 24520 -56480 24620 -56380 1 PIX3056_IN
port 3104 n
rlabel metal5 26020 -56480 26120 -56380 1 PIX3057_IN
port 3105 n
rlabel metal5 27520 -56480 27620 -56380 1 PIX3058_IN
port 3106 n
rlabel metal5 29020 -56480 29120 -56380 1 PIX3059_IN
port 3107 n
rlabel metal5 30520 -56480 30620 -56380 1 PIX3060_IN
port 3108 n
rlabel metal5 32020 -56480 32120 -56380 1 PIX3061_IN
port 3109 n
rlabel metal5 33520 -56480 33620 -56380 1 PIX3062_IN
port 3110 n
rlabel metal5 35020 -56480 35120 -56380 1 PIX3063_IN
port 3111 n
rlabel metal5 36520 -56480 36620 -56380 1 PIX3064_IN
port 3112 n
rlabel metal5 38020 -56480 38120 -56380 1 PIX3065_IN
port 3113 n
rlabel metal5 39520 -56480 39620 -56380 1 PIX3066_IN
port 3114 n
rlabel metal5 41020 -56480 41120 -56380 1 PIX3067_IN
port 3115 n
rlabel metal5 42520 -56480 42620 -56380 1 PIX3068_IN
port 3116 n
rlabel metal5 44020 -56480 44120 -56380 1 PIX3069_IN
port 3117 n
rlabel metal5 45520 -56480 45620 -56380 1 PIX3070_IN
port 3118 n
rlabel metal5 47020 -56480 47120 -56380 1 PIX3071_IN
port 3119 n
rlabel metal5 48520 -56480 48620 -56380 1 PIX3072_IN
port 3120 n
rlabel metal5 50020 -56480 50120 -56380 1 PIX3073_IN
port 3121 n
rlabel metal5 51520 -56480 51620 -56380 1 PIX3074_IN
port 3122 n
rlabel metal5 53020 -56480 53120 -56380 1 PIX3075_IN
port 3123 n
rlabel metal5 54520 -56480 54620 -56380 1 PIX3076_IN
port 3124 n
rlabel metal5 56020 -56480 56120 -56380 1 PIX3077_IN
port 3125 n
rlabel metal5 57520 -56480 57620 -56380 1 PIX3078_IN
port 3126 n
rlabel metal5 59020 -56480 59120 -56380 1 PIX3079_IN
port 3127 n
rlabel metal5 60520 -56480 60620 -56380 1 PIX3080_IN
port 3128 n
rlabel metal5 62020 -56480 62120 -56380 1 PIX3081_IN
port 3129 n
rlabel metal5 63520 -56480 63620 -56380 1 PIX3082_IN
port 3130 n
rlabel metal5 65020 -56480 65120 -56380 1 PIX3083_IN
port 3131 n
rlabel metal5 66520 -56480 66620 -56380 1 PIX3084_IN
port 3132 n
rlabel metal5 68020 -56480 68120 -56380 1 PIX3085_IN
port 3133 n
rlabel metal5 69520 -56480 69620 -56380 1 PIX3086_IN
port 3134 n
rlabel metal5 71020 -56480 71120 -56380 1 PIX3087_IN
port 3135 n
rlabel metal5 72520 -56480 72620 -56380 1 PIX3088_IN
port 3136 n
rlabel metal5 74020 -56480 74120 -56380 1 PIX3089_IN
port 3137 n
rlabel metal5 75520 -56480 75620 -56380 1 PIX3090_IN
port 3138 n
rlabel metal5 77020 -56480 77120 -56380 1 PIX3091_IN
port 3139 n
rlabel metal5 78520 -56480 78620 -56380 1 PIX3092_IN
port 3140 n
rlabel metal5 80020 -56480 80120 -56380 1 PIX3093_IN
port 3141 n
rlabel metal5 81520 -56480 81620 -56380 1 PIX3094_IN
port 3142 n
rlabel metal5 83020 -56480 83120 -56380 1 PIX3095_IN
port 3143 n
rlabel metal5 84520 -56480 84620 -56380 1 PIX3096_IN
port 3144 n
rlabel metal5 86020 -56480 86120 -56380 1 PIX3097_IN
port 3145 n
rlabel metal5 87520 -56480 87620 -56380 1 PIX3098_IN
port 3146 n
rlabel metal5 89020 -56480 89120 -56380 1 PIX3099_IN
port 3147 n
rlabel metal5 90520 -56480 90620 -56380 1 PIX3100_IN
port 3148 n
rlabel metal5 92020 -56480 92120 -56380 1 PIX3101_IN
port 3149 n
rlabel metal5 93520 -56480 93620 -56380 1 PIX3102_IN
port 3150 n
rlabel metal5 95020 -56480 95120 -56380 1 PIX3103_IN
port 3151 n
rlabel metal5 96520 -56480 96620 -56380 1 PIX3104_IN
port 3152 n
rlabel metal5 98020 -56480 98120 -56380 1 PIX3105_IN
port 3153 n
rlabel metal5 99520 -56480 99620 -56380 1 PIX3106_IN
port 3154 n
rlabel metal5 101020 -56480 101120 -56380 1 PIX3107_IN
port 3155 n
rlabel metal5 102520 -56480 102620 -56380 1 PIX3108_IN
port 3156 n
rlabel metal5 104020 -56480 104120 -56380 1 PIX3109_IN
port 3157 n
rlabel metal5 105520 -56480 105620 -56380 1 PIX3110_IN
port 3158 n
rlabel metal5 107020 -56480 107120 -56380 1 PIX3111_IN
port 3159 n
rlabel metal5 108520 -56480 108620 -56380 1 PIX3112_IN
port 3160 n
rlabel metal5 110020 -56480 110120 -56380 1 PIX3113_IN
port 3161 n
rlabel metal5 111520 -56480 111620 -56380 1 PIX3114_IN
port 3162 n
rlabel metal5 113020 -56480 113120 -56380 1 PIX3115_IN
port 3163 n
rlabel metal5 114520 -56480 114620 -56380 1 PIX3116_IN
port 3164 n
rlabel metal5 116020 -56480 116120 -56380 1 PIX3117_IN
port 3165 n
rlabel metal5 117520 -56480 117620 -56380 1 PIX3118_IN
port 3166 n
rlabel metal5 119020 -56480 119120 -56380 1 PIX3119_IN
port 3167 n
rlabel metal5 520 -57980 620 -57880 1 PIX3120_IN
port 3168 n
rlabel metal2 -1500 -57760 -1500 -57715 3 ROW_SEL39
port 3169 e
rlabel metal5 2020 -57980 2120 -57880 1 PIX3121_IN
port 3170 n
rlabel metal5 3520 -57980 3620 -57880 1 PIX3122_IN
port 3171 n
rlabel metal5 5020 -57980 5120 -57880 1 PIX3123_IN
port 3172 n
rlabel metal5 6520 -57980 6620 -57880 1 PIX3124_IN
port 3173 n
rlabel metal5 8020 -57980 8120 -57880 1 PIX3125_IN
port 3174 n
rlabel metal5 9520 -57980 9620 -57880 1 PIX3126_IN
port 3175 n
rlabel metal5 11020 -57980 11120 -57880 1 PIX3127_IN
port 3176 n
rlabel metal5 12520 -57980 12620 -57880 1 PIX3128_IN
port 3177 n
rlabel metal5 14020 -57980 14120 -57880 1 PIX3129_IN
port 3178 n
rlabel metal5 15520 -57980 15620 -57880 1 PIX3130_IN
port 3179 n
rlabel metal5 17020 -57980 17120 -57880 1 PIX3131_IN
port 3180 n
rlabel metal5 18520 -57980 18620 -57880 1 PIX3132_IN
port 3181 n
rlabel metal5 20020 -57980 20120 -57880 1 PIX3133_IN
port 3182 n
rlabel metal5 21520 -57980 21620 -57880 1 PIX3134_IN
port 3183 n
rlabel metal5 23020 -57980 23120 -57880 1 PIX3135_IN
port 3184 n
rlabel metal5 24520 -57980 24620 -57880 1 PIX3136_IN
port 3185 n
rlabel metal5 26020 -57980 26120 -57880 1 PIX3137_IN
port 3186 n
rlabel metal5 27520 -57980 27620 -57880 1 PIX3138_IN
port 3187 n
rlabel metal5 29020 -57980 29120 -57880 1 PIX3139_IN
port 3188 n
rlabel metal5 30520 -57980 30620 -57880 1 PIX3140_IN
port 3189 n
rlabel metal5 32020 -57980 32120 -57880 1 PIX3141_IN
port 3190 n
rlabel metal5 33520 -57980 33620 -57880 1 PIX3142_IN
port 3191 n
rlabel metal5 35020 -57980 35120 -57880 1 PIX3143_IN
port 3192 n
rlabel metal5 36520 -57980 36620 -57880 1 PIX3144_IN
port 3193 n
rlabel metal5 38020 -57980 38120 -57880 1 PIX3145_IN
port 3194 n
rlabel metal5 39520 -57980 39620 -57880 1 PIX3146_IN
port 3195 n
rlabel metal5 41020 -57980 41120 -57880 1 PIX3147_IN
port 3196 n
rlabel metal5 42520 -57980 42620 -57880 1 PIX3148_IN
port 3197 n
rlabel metal5 44020 -57980 44120 -57880 1 PIX3149_IN
port 3198 n
rlabel metal5 45520 -57980 45620 -57880 1 PIX3150_IN
port 3199 n
rlabel metal5 47020 -57980 47120 -57880 1 PIX3151_IN
port 3200 n
rlabel metal5 48520 -57980 48620 -57880 1 PIX3152_IN
port 3201 n
rlabel metal5 50020 -57980 50120 -57880 1 PIX3153_IN
port 3202 n
rlabel metal5 51520 -57980 51620 -57880 1 PIX3154_IN
port 3203 n
rlabel metal5 53020 -57980 53120 -57880 1 PIX3155_IN
port 3204 n
rlabel metal5 54520 -57980 54620 -57880 1 PIX3156_IN
port 3205 n
rlabel metal5 56020 -57980 56120 -57880 1 PIX3157_IN
port 3206 n
rlabel metal5 57520 -57980 57620 -57880 1 PIX3158_IN
port 3207 n
rlabel metal5 59020 -57980 59120 -57880 1 PIX3159_IN
port 3208 n
rlabel metal5 60520 -57980 60620 -57880 1 PIX3160_IN
port 3209 n
rlabel metal5 62020 -57980 62120 -57880 1 PIX3161_IN
port 3210 n
rlabel metal5 63520 -57980 63620 -57880 1 PIX3162_IN
port 3211 n
rlabel metal5 65020 -57980 65120 -57880 1 PIX3163_IN
port 3212 n
rlabel metal5 66520 -57980 66620 -57880 1 PIX3164_IN
port 3213 n
rlabel metal5 68020 -57980 68120 -57880 1 PIX3165_IN
port 3214 n
rlabel metal5 69520 -57980 69620 -57880 1 PIX3166_IN
port 3215 n
rlabel metal5 71020 -57980 71120 -57880 1 PIX3167_IN
port 3216 n
rlabel metal5 72520 -57980 72620 -57880 1 PIX3168_IN
port 3217 n
rlabel metal5 74020 -57980 74120 -57880 1 PIX3169_IN
port 3218 n
rlabel metal5 75520 -57980 75620 -57880 1 PIX3170_IN
port 3219 n
rlabel metal5 77020 -57980 77120 -57880 1 PIX3171_IN
port 3220 n
rlabel metal5 78520 -57980 78620 -57880 1 PIX3172_IN
port 3221 n
rlabel metal5 80020 -57980 80120 -57880 1 PIX3173_IN
port 3222 n
rlabel metal5 81520 -57980 81620 -57880 1 PIX3174_IN
port 3223 n
rlabel metal5 83020 -57980 83120 -57880 1 PIX3175_IN
port 3224 n
rlabel metal5 84520 -57980 84620 -57880 1 PIX3176_IN
port 3225 n
rlabel metal5 86020 -57980 86120 -57880 1 PIX3177_IN
port 3226 n
rlabel metal5 87520 -57980 87620 -57880 1 PIX3178_IN
port 3227 n
rlabel metal5 89020 -57980 89120 -57880 1 PIX3179_IN
port 3228 n
rlabel metal5 90520 -57980 90620 -57880 1 PIX3180_IN
port 3229 n
rlabel metal5 92020 -57980 92120 -57880 1 PIX3181_IN
port 3230 n
rlabel metal5 93520 -57980 93620 -57880 1 PIX3182_IN
port 3231 n
rlabel metal5 95020 -57980 95120 -57880 1 PIX3183_IN
port 3232 n
rlabel metal5 96520 -57980 96620 -57880 1 PIX3184_IN
port 3233 n
rlabel metal5 98020 -57980 98120 -57880 1 PIX3185_IN
port 3234 n
rlabel metal5 99520 -57980 99620 -57880 1 PIX3186_IN
port 3235 n
rlabel metal5 101020 -57980 101120 -57880 1 PIX3187_IN
port 3236 n
rlabel metal5 102520 -57980 102620 -57880 1 PIX3188_IN
port 3237 n
rlabel metal5 104020 -57980 104120 -57880 1 PIX3189_IN
port 3238 n
rlabel metal5 105520 -57980 105620 -57880 1 PIX3190_IN
port 3239 n
rlabel metal5 107020 -57980 107120 -57880 1 PIX3191_IN
port 3240 n
rlabel metal5 108520 -57980 108620 -57880 1 PIX3192_IN
port 3241 n
rlabel metal5 110020 -57980 110120 -57880 1 PIX3193_IN
port 3242 n
rlabel metal5 111520 -57980 111620 -57880 1 PIX3194_IN
port 3243 n
rlabel metal5 113020 -57980 113120 -57880 1 PIX3195_IN
port 3244 n
rlabel metal5 114520 -57980 114620 -57880 1 PIX3196_IN
port 3245 n
rlabel metal5 116020 -57980 116120 -57880 1 PIX3197_IN
port 3246 n
rlabel metal5 117520 -57980 117620 -57880 1 PIX3198_IN
port 3247 n
rlabel metal5 119020 -57980 119120 -57880 1 PIX3199_IN
port 3248 n
rlabel metal5 520 -59480 620 -59380 1 PIX3200_IN
port 3249 n
rlabel metal2 -1500 -59260 -1500 -59215 3 ROW_SEL40
port 3250 e
rlabel metal5 2020 -59480 2120 -59380 1 PIX3201_IN
port 3251 n
rlabel metal5 3520 -59480 3620 -59380 1 PIX3202_IN
port 3252 n
rlabel metal5 5020 -59480 5120 -59380 1 PIX3203_IN
port 3253 n
rlabel metal5 6520 -59480 6620 -59380 1 PIX3204_IN
port 3254 n
rlabel metal5 8020 -59480 8120 -59380 1 PIX3205_IN
port 3255 n
rlabel metal5 9520 -59480 9620 -59380 1 PIX3206_IN
port 3256 n
rlabel metal5 11020 -59480 11120 -59380 1 PIX3207_IN
port 3257 n
rlabel metal5 12520 -59480 12620 -59380 1 PIX3208_IN
port 3258 n
rlabel metal5 14020 -59480 14120 -59380 1 PIX3209_IN
port 3259 n
rlabel metal5 15520 -59480 15620 -59380 1 PIX3210_IN
port 3260 n
rlabel metal5 17020 -59480 17120 -59380 1 PIX3211_IN
port 3261 n
rlabel metal5 18520 -59480 18620 -59380 1 PIX3212_IN
port 3262 n
rlabel metal5 20020 -59480 20120 -59380 1 PIX3213_IN
port 3263 n
rlabel metal5 21520 -59480 21620 -59380 1 PIX3214_IN
port 3264 n
rlabel metal5 23020 -59480 23120 -59380 1 PIX3215_IN
port 3265 n
rlabel metal5 24520 -59480 24620 -59380 1 PIX3216_IN
port 3266 n
rlabel metal5 26020 -59480 26120 -59380 1 PIX3217_IN
port 3267 n
rlabel metal5 27520 -59480 27620 -59380 1 PIX3218_IN
port 3268 n
rlabel metal5 29020 -59480 29120 -59380 1 PIX3219_IN
port 3269 n
rlabel metal5 30520 -59480 30620 -59380 1 PIX3220_IN
port 3270 n
rlabel metal5 32020 -59480 32120 -59380 1 PIX3221_IN
port 3271 n
rlabel metal5 33520 -59480 33620 -59380 1 PIX3222_IN
port 3272 n
rlabel metal5 35020 -59480 35120 -59380 1 PIX3223_IN
port 3273 n
rlabel metal5 36520 -59480 36620 -59380 1 PIX3224_IN
port 3274 n
rlabel metal5 38020 -59480 38120 -59380 1 PIX3225_IN
port 3275 n
rlabel metal5 39520 -59480 39620 -59380 1 PIX3226_IN
port 3276 n
rlabel metal5 41020 -59480 41120 -59380 1 PIX3227_IN
port 3277 n
rlabel metal5 42520 -59480 42620 -59380 1 PIX3228_IN
port 3278 n
rlabel metal5 44020 -59480 44120 -59380 1 PIX3229_IN
port 3279 n
rlabel metal5 45520 -59480 45620 -59380 1 PIX3230_IN
port 3280 n
rlabel metal5 47020 -59480 47120 -59380 1 PIX3231_IN
port 3281 n
rlabel metal5 48520 -59480 48620 -59380 1 PIX3232_IN
port 3282 n
rlabel metal5 50020 -59480 50120 -59380 1 PIX3233_IN
port 3283 n
rlabel metal5 51520 -59480 51620 -59380 1 PIX3234_IN
port 3284 n
rlabel metal5 53020 -59480 53120 -59380 1 PIX3235_IN
port 3285 n
rlabel metal5 54520 -59480 54620 -59380 1 PIX3236_IN
port 3286 n
rlabel metal5 56020 -59480 56120 -59380 1 PIX3237_IN
port 3287 n
rlabel metal5 57520 -59480 57620 -59380 1 PIX3238_IN
port 3288 n
rlabel metal5 59020 -59480 59120 -59380 1 PIX3239_IN
port 3289 n
rlabel metal5 60520 -59480 60620 -59380 1 PIX3240_IN
port 3290 n
rlabel metal5 62020 -59480 62120 -59380 1 PIX3241_IN
port 3291 n
rlabel metal5 63520 -59480 63620 -59380 1 PIX3242_IN
port 3292 n
rlabel metal5 65020 -59480 65120 -59380 1 PIX3243_IN
port 3293 n
rlabel metal5 66520 -59480 66620 -59380 1 PIX3244_IN
port 3294 n
rlabel metal5 68020 -59480 68120 -59380 1 PIX3245_IN
port 3295 n
rlabel metal5 69520 -59480 69620 -59380 1 PIX3246_IN
port 3296 n
rlabel metal5 71020 -59480 71120 -59380 1 PIX3247_IN
port 3297 n
rlabel metal5 72520 -59480 72620 -59380 1 PIX3248_IN
port 3298 n
rlabel metal5 74020 -59480 74120 -59380 1 PIX3249_IN
port 3299 n
rlabel metal5 75520 -59480 75620 -59380 1 PIX3250_IN
port 3300 n
rlabel metal5 77020 -59480 77120 -59380 1 PIX3251_IN
port 3301 n
rlabel metal5 78520 -59480 78620 -59380 1 PIX3252_IN
port 3302 n
rlabel metal5 80020 -59480 80120 -59380 1 PIX3253_IN
port 3303 n
rlabel metal5 81520 -59480 81620 -59380 1 PIX3254_IN
port 3304 n
rlabel metal5 83020 -59480 83120 -59380 1 PIX3255_IN
port 3305 n
rlabel metal5 84520 -59480 84620 -59380 1 PIX3256_IN
port 3306 n
rlabel metal5 86020 -59480 86120 -59380 1 PIX3257_IN
port 3307 n
rlabel metal5 87520 -59480 87620 -59380 1 PIX3258_IN
port 3308 n
rlabel metal5 89020 -59480 89120 -59380 1 PIX3259_IN
port 3309 n
rlabel metal5 90520 -59480 90620 -59380 1 PIX3260_IN
port 3310 n
rlabel metal5 92020 -59480 92120 -59380 1 PIX3261_IN
port 3311 n
rlabel metal5 93520 -59480 93620 -59380 1 PIX3262_IN
port 3312 n
rlabel metal5 95020 -59480 95120 -59380 1 PIX3263_IN
port 3313 n
rlabel metal5 96520 -59480 96620 -59380 1 PIX3264_IN
port 3314 n
rlabel metal5 98020 -59480 98120 -59380 1 PIX3265_IN
port 3315 n
rlabel metal5 99520 -59480 99620 -59380 1 PIX3266_IN
port 3316 n
rlabel metal5 101020 -59480 101120 -59380 1 PIX3267_IN
port 3317 n
rlabel metal5 102520 -59480 102620 -59380 1 PIX3268_IN
port 3318 n
rlabel metal5 104020 -59480 104120 -59380 1 PIX3269_IN
port 3319 n
rlabel metal5 105520 -59480 105620 -59380 1 PIX3270_IN
port 3320 n
rlabel metal5 107020 -59480 107120 -59380 1 PIX3271_IN
port 3321 n
rlabel metal5 108520 -59480 108620 -59380 1 PIX3272_IN
port 3322 n
rlabel metal5 110020 -59480 110120 -59380 1 PIX3273_IN
port 3323 n
rlabel metal5 111520 -59480 111620 -59380 1 PIX3274_IN
port 3324 n
rlabel metal5 113020 -59480 113120 -59380 1 PIX3275_IN
port 3325 n
rlabel metal5 114520 -59480 114620 -59380 1 PIX3276_IN
port 3326 n
rlabel metal5 116020 -59480 116120 -59380 1 PIX3277_IN
port 3327 n
rlabel metal5 117520 -59480 117620 -59380 1 PIX3278_IN
port 3328 n
rlabel metal5 119020 -59480 119120 -59380 1 PIX3279_IN
port 3329 n
rlabel metal5 520 -60980 620 -60880 1 PIX3280_IN
port 3330 n
rlabel metal2 -1500 -60760 -1500 -60715 3 ROW_SEL41
port 3331 e
rlabel metal5 2020 -60980 2120 -60880 1 PIX3281_IN
port 3332 n
rlabel metal5 3520 -60980 3620 -60880 1 PIX3282_IN
port 3333 n
rlabel metal5 5020 -60980 5120 -60880 1 PIX3283_IN
port 3334 n
rlabel metal5 6520 -60980 6620 -60880 1 PIX3284_IN
port 3335 n
rlabel metal5 8020 -60980 8120 -60880 1 PIX3285_IN
port 3336 n
rlabel metal5 9520 -60980 9620 -60880 1 PIX3286_IN
port 3337 n
rlabel metal5 11020 -60980 11120 -60880 1 PIX3287_IN
port 3338 n
rlabel metal5 12520 -60980 12620 -60880 1 PIX3288_IN
port 3339 n
rlabel metal5 14020 -60980 14120 -60880 1 PIX3289_IN
port 3340 n
rlabel metal5 15520 -60980 15620 -60880 1 PIX3290_IN
port 3341 n
rlabel metal5 17020 -60980 17120 -60880 1 PIX3291_IN
port 3342 n
rlabel metal5 18520 -60980 18620 -60880 1 PIX3292_IN
port 3343 n
rlabel metal5 20020 -60980 20120 -60880 1 PIX3293_IN
port 3344 n
rlabel metal5 21520 -60980 21620 -60880 1 PIX3294_IN
port 3345 n
rlabel metal5 23020 -60980 23120 -60880 1 PIX3295_IN
port 3346 n
rlabel metal5 24520 -60980 24620 -60880 1 PIX3296_IN
port 3347 n
rlabel metal5 26020 -60980 26120 -60880 1 PIX3297_IN
port 3348 n
rlabel metal5 27520 -60980 27620 -60880 1 PIX3298_IN
port 3349 n
rlabel metal5 29020 -60980 29120 -60880 1 PIX3299_IN
port 3350 n
rlabel metal5 30520 -60980 30620 -60880 1 PIX3300_IN
port 3351 n
rlabel metal5 32020 -60980 32120 -60880 1 PIX3301_IN
port 3352 n
rlabel metal5 33520 -60980 33620 -60880 1 PIX3302_IN
port 3353 n
rlabel metal5 35020 -60980 35120 -60880 1 PIX3303_IN
port 3354 n
rlabel metal5 36520 -60980 36620 -60880 1 PIX3304_IN
port 3355 n
rlabel metal5 38020 -60980 38120 -60880 1 PIX3305_IN
port 3356 n
rlabel metal5 39520 -60980 39620 -60880 1 PIX3306_IN
port 3357 n
rlabel metal5 41020 -60980 41120 -60880 1 PIX3307_IN
port 3358 n
rlabel metal5 42520 -60980 42620 -60880 1 PIX3308_IN
port 3359 n
rlabel metal5 44020 -60980 44120 -60880 1 PIX3309_IN
port 3360 n
rlabel metal5 45520 -60980 45620 -60880 1 PIX3310_IN
port 3361 n
rlabel metal5 47020 -60980 47120 -60880 1 PIX3311_IN
port 3362 n
rlabel metal5 48520 -60980 48620 -60880 1 PIX3312_IN
port 3363 n
rlabel metal5 50020 -60980 50120 -60880 1 PIX3313_IN
port 3364 n
rlabel metal5 51520 -60980 51620 -60880 1 PIX3314_IN
port 3365 n
rlabel metal5 53020 -60980 53120 -60880 1 PIX3315_IN
port 3366 n
rlabel metal5 54520 -60980 54620 -60880 1 PIX3316_IN
port 3367 n
rlabel metal5 56020 -60980 56120 -60880 1 PIX3317_IN
port 3368 n
rlabel metal5 57520 -60980 57620 -60880 1 PIX3318_IN
port 3369 n
rlabel metal5 59020 -60980 59120 -60880 1 PIX3319_IN
port 3370 n
rlabel metal5 60520 -60980 60620 -60880 1 PIX3320_IN
port 3371 n
rlabel metal5 62020 -60980 62120 -60880 1 PIX3321_IN
port 3372 n
rlabel metal5 63520 -60980 63620 -60880 1 PIX3322_IN
port 3373 n
rlabel metal5 65020 -60980 65120 -60880 1 PIX3323_IN
port 3374 n
rlabel metal5 66520 -60980 66620 -60880 1 PIX3324_IN
port 3375 n
rlabel metal5 68020 -60980 68120 -60880 1 PIX3325_IN
port 3376 n
rlabel metal5 69520 -60980 69620 -60880 1 PIX3326_IN
port 3377 n
rlabel metal5 71020 -60980 71120 -60880 1 PIX3327_IN
port 3378 n
rlabel metal5 72520 -60980 72620 -60880 1 PIX3328_IN
port 3379 n
rlabel metal5 74020 -60980 74120 -60880 1 PIX3329_IN
port 3380 n
rlabel metal5 75520 -60980 75620 -60880 1 PIX3330_IN
port 3381 n
rlabel metal5 77020 -60980 77120 -60880 1 PIX3331_IN
port 3382 n
rlabel metal5 78520 -60980 78620 -60880 1 PIX3332_IN
port 3383 n
rlabel metal5 80020 -60980 80120 -60880 1 PIX3333_IN
port 3384 n
rlabel metal5 81520 -60980 81620 -60880 1 PIX3334_IN
port 3385 n
rlabel metal5 83020 -60980 83120 -60880 1 PIX3335_IN
port 3386 n
rlabel metal5 84520 -60980 84620 -60880 1 PIX3336_IN
port 3387 n
rlabel metal5 86020 -60980 86120 -60880 1 PIX3337_IN
port 3388 n
rlabel metal5 87520 -60980 87620 -60880 1 PIX3338_IN
port 3389 n
rlabel metal5 89020 -60980 89120 -60880 1 PIX3339_IN
port 3390 n
rlabel metal5 90520 -60980 90620 -60880 1 PIX3340_IN
port 3391 n
rlabel metal5 92020 -60980 92120 -60880 1 PIX3341_IN
port 3392 n
rlabel metal5 93520 -60980 93620 -60880 1 PIX3342_IN
port 3393 n
rlabel metal5 95020 -60980 95120 -60880 1 PIX3343_IN
port 3394 n
rlabel metal5 96520 -60980 96620 -60880 1 PIX3344_IN
port 3395 n
rlabel metal5 98020 -60980 98120 -60880 1 PIX3345_IN
port 3396 n
rlabel metal5 99520 -60980 99620 -60880 1 PIX3346_IN
port 3397 n
rlabel metal5 101020 -60980 101120 -60880 1 PIX3347_IN
port 3398 n
rlabel metal5 102520 -60980 102620 -60880 1 PIX3348_IN
port 3399 n
rlabel metal5 104020 -60980 104120 -60880 1 PIX3349_IN
port 3400 n
rlabel metal5 105520 -60980 105620 -60880 1 PIX3350_IN
port 3401 n
rlabel metal5 107020 -60980 107120 -60880 1 PIX3351_IN
port 3402 n
rlabel metal5 108520 -60980 108620 -60880 1 PIX3352_IN
port 3403 n
rlabel metal5 110020 -60980 110120 -60880 1 PIX3353_IN
port 3404 n
rlabel metal5 111520 -60980 111620 -60880 1 PIX3354_IN
port 3405 n
rlabel metal5 113020 -60980 113120 -60880 1 PIX3355_IN
port 3406 n
rlabel metal5 114520 -60980 114620 -60880 1 PIX3356_IN
port 3407 n
rlabel metal5 116020 -60980 116120 -60880 1 PIX3357_IN
port 3408 n
rlabel metal5 117520 -60980 117620 -60880 1 PIX3358_IN
port 3409 n
rlabel metal5 119020 -60980 119120 -60880 1 PIX3359_IN
port 3410 n
rlabel metal5 520 -62480 620 -62380 1 PIX3360_IN
port 3411 n
rlabel metal2 -1500 -62260 -1500 -62215 3 ROW_SEL42
port 3412 e
rlabel metal5 2020 -62480 2120 -62380 1 PIX3361_IN
port 3413 n
rlabel metal5 3520 -62480 3620 -62380 1 PIX3362_IN
port 3414 n
rlabel metal5 5020 -62480 5120 -62380 1 PIX3363_IN
port 3415 n
rlabel metal5 6520 -62480 6620 -62380 1 PIX3364_IN
port 3416 n
rlabel metal5 8020 -62480 8120 -62380 1 PIX3365_IN
port 3417 n
rlabel metal5 9520 -62480 9620 -62380 1 PIX3366_IN
port 3418 n
rlabel metal5 11020 -62480 11120 -62380 1 PIX3367_IN
port 3419 n
rlabel metal5 12520 -62480 12620 -62380 1 PIX3368_IN
port 3420 n
rlabel metal5 14020 -62480 14120 -62380 1 PIX3369_IN
port 3421 n
rlabel metal5 15520 -62480 15620 -62380 1 PIX3370_IN
port 3422 n
rlabel metal5 17020 -62480 17120 -62380 1 PIX3371_IN
port 3423 n
rlabel metal5 18520 -62480 18620 -62380 1 PIX3372_IN
port 3424 n
rlabel metal5 20020 -62480 20120 -62380 1 PIX3373_IN
port 3425 n
rlabel metal5 21520 -62480 21620 -62380 1 PIX3374_IN
port 3426 n
rlabel metal5 23020 -62480 23120 -62380 1 PIX3375_IN
port 3427 n
rlabel metal5 24520 -62480 24620 -62380 1 PIX3376_IN
port 3428 n
rlabel metal5 26020 -62480 26120 -62380 1 PIX3377_IN
port 3429 n
rlabel metal5 27520 -62480 27620 -62380 1 PIX3378_IN
port 3430 n
rlabel metal5 29020 -62480 29120 -62380 1 PIX3379_IN
port 3431 n
rlabel metal5 30520 -62480 30620 -62380 1 PIX3380_IN
port 3432 n
rlabel metal5 32020 -62480 32120 -62380 1 PIX3381_IN
port 3433 n
rlabel metal5 33520 -62480 33620 -62380 1 PIX3382_IN
port 3434 n
rlabel metal5 35020 -62480 35120 -62380 1 PIX3383_IN
port 3435 n
rlabel metal5 36520 -62480 36620 -62380 1 PIX3384_IN
port 3436 n
rlabel metal5 38020 -62480 38120 -62380 1 PIX3385_IN
port 3437 n
rlabel metal5 39520 -62480 39620 -62380 1 PIX3386_IN
port 3438 n
rlabel metal5 41020 -62480 41120 -62380 1 PIX3387_IN
port 3439 n
rlabel metal5 42520 -62480 42620 -62380 1 PIX3388_IN
port 3440 n
rlabel metal5 44020 -62480 44120 -62380 1 PIX3389_IN
port 3441 n
rlabel metal5 45520 -62480 45620 -62380 1 PIX3390_IN
port 3442 n
rlabel metal5 47020 -62480 47120 -62380 1 PIX3391_IN
port 3443 n
rlabel metal5 48520 -62480 48620 -62380 1 PIX3392_IN
port 3444 n
rlabel metal5 50020 -62480 50120 -62380 1 PIX3393_IN
port 3445 n
rlabel metal5 51520 -62480 51620 -62380 1 PIX3394_IN
port 3446 n
rlabel metal5 53020 -62480 53120 -62380 1 PIX3395_IN
port 3447 n
rlabel metal5 54520 -62480 54620 -62380 1 PIX3396_IN
port 3448 n
rlabel metal5 56020 -62480 56120 -62380 1 PIX3397_IN
port 3449 n
rlabel metal5 57520 -62480 57620 -62380 1 PIX3398_IN
port 3450 n
rlabel metal5 59020 -62480 59120 -62380 1 PIX3399_IN
port 3451 n
rlabel metal5 60520 -62480 60620 -62380 1 PIX3400_IN
port 3452 n
rlabel metal5 62020 -62480 62120 -62380 1 PIX3401_IN
port 3453 n
rlabel metal5 63520 -62480 63620 -62380 1 PIX3402_IN
port 3454 n
rlabel metal5 65020 -62480 65120 -62380 1 PIX3403_IN
port 3455 n
rlabel metal5 66520 -62480 66620 -62380 1 PIX3404_IN
port 3456 n
rlabel metal5 68020 -62480 68120 -62380 1 PIX3405_IN
port 3457 n
rlabel metal5 69520 -62480 69620 -62380 1 PIX3406_IN
port 3458 n
rlabel metal5 71020 -62480 71120 -62380 1 PIX3407_IN
port 3459 n
rlabel metal5 72520 -62480 72620 -62380 1 PIX3408_IN
port 3460 n
rlabel metal5 74020 -62480 74120 -62380 1 PIX3409_IN
port 3461 n
rlabel metal5 75520 -62480 75620 -62380 1 PIX3410_IN
port 3462 n
rlabel metal5 77020 -62480 77120 -62380 1 PIX3411_IN
port 3463 n
rlabel metal5 78520 -62480 78620 -62380 1 PIX3412_IN
port 3464 n
rlabel metal5 80020 -62480 80120 -62380 1 PIX3413_IN
port 3465 n
rlabel metal5 81520 -62480 81620 -62380 1 PIX3414_IN
port 3466 n
rlabel metal5 83020 -62480 83120 -62380 1 PIX3415_IN
port 3467 n
rlabel metal5 84520 -62480 84620 -62380 1 PIX3416_IN
port 3468 n
rlabel metal5 86020 -62480 86120 -62380 1 PIX3417_IN
port 3469 n
rlabel metal5 87520 -62480 87620 -62380 1 PIX3418_IN
port 3470 n
rlabel metal5 89020 -62480 89120 -62380 1 PIX3419_IN
port 3471 n
rlabel metal5 90520 -62480 90620 -62380 1 PIX3420_IN
port 3472 n
rlabel metal5 92020 -62480 92120 -62380 1 PIX3421_IN
port 3473 n
rlabel metal5 93520 -62480 93620 -62380 1 PIX3422_IN
port 3474 n
rlabel metal5 95020 -62480 95120 -62380 1 PIX3423_IN
port 3475 n
rlabel metal5 96520 -62480 96620 -62380 1 PIX3424_IN
port 3476 n
rlabel metal5 98020 -62480 98120 -62380 1 PIX3425_IN
port 3477 n
rlabel metal5 99520 -62480 99620 -62380 1 PIX3426_IN
port 3478 n
rlabel metal5 101020 -62480 101120 -62380 1 PIX3427_IN
port 3479 n
rlabel metal5 102520 -62480 102620 -62380 1 PIX3428_IN
port 3480 n
rlabel metal5 104020 -62480 104120 -62380 1 PIX3429_IN
port 3481 n
rlabel metal5 105520 -62480 105620 -62380 1 PIX3430_IN
port 3482 n
rlabel metal5 107020 -62480 107120 -62380 1 PIX3431_IN
port 3483 n
rlabel metal5 108520 -62480 108620 -62380 1 PIX3432_IN
port 3484 n
rlabel metal5 110020 -62480 110120 -62380 1 PIX3433_IN
port 3485 n
rlabel metal5 111520 -62480 111620 -62380 1 PIX3434_IN
port 3486 n
rlabel metal5 113020 -62480 113120 -62380 1 PIX3435_IN
port 3487 n
rlabel metal5 114520 -62480 114620 -62380 1 PIX3436_IN
port 3488 n
rlabel metal5 116020 -62480 116120 -62380 1 PIX3437_IN
port 3489 n
rlabel metal5 117520 -62480 117620 -62380 1 PIX3438_IN
port 3490 n
rlabel metal5 119020 -62480 119120 -62380 1 PIX3439_IN
port 3491 n
rlabel metal5 520 -63980 620 -63880 1 PIX3440_IN
port 3492 n
rlabel metal2 -1500 -63760 -1500 -63715 3 ROW_SEL43
port 3493 e
rlabel metal5 2020 -63980 2120 -63880 1 PIX3441_IN
port 3494 n
rlabel metal5 3520 -63980 3620 -63880 1 PIX3442_IN
port 3495 n
rlabel metal5 5020 -63980 5120 -63880 1 PIX3443_IN
port 3496 n
rlabel metal5 6520 -63980 6620 -63880 1 PIX3444_IN
port 3497 n
rlabel metal5 8020 -63980 8120 -63880 1 PIX3445_IN
port 3498 n
rlabel metal5 9520 -63980 9620 -63880 1 PIX3446_IN
port 3499 n
rlabel metal5 11020 -63980 11120 -63880 1 PIX3447_IN
port 3500 n
rlabel metal5 12520 -63980 12620 -63880 1 PIX3448_IN
port 3501 n
rlabel metal5 14020 -63980 14120 -63880 1 PIX3449_IN
port 3502 n
rlabel metal5 15520 -63980 15620 -63880 1 PIX3450_IN
port 3503 n
rlabel metal5 17020 -63980 17120 -63880 1 PIX3451_IN
port 3504 n
rlabel metal5 18520 -63980 18620 -63880 1 PIX3452_IN
port 3505 n
rlabel metal5 20020 -63980 20120 -63880 1 PIX3453_IN
port 3506 n
rlabel metal5 21520 -63980 21620 -63880 1 PIX3454_IN
port 3507 n
rlabel metal5 23020 -63980 23120 -63880 1 PIX3455_IN
port 3508 n
rlabel metal5 24520 -63980 24620 -63880 1 PIX3456_IN
port 3509 n
rlabel metal5 26020 -63980 26120 -63880 1 PIX3457_IN
port 3510 n
rlabel metal5 27520 -63980 27620 -63880 1 PIX3458_IN
port 3511 n
rlabel metal5 29020 -63980 29120 -63880 1 PIX3459_IN
port 3512 n
rlabel metal5 30520 -63980 30620 -63880 1 PIX3460_IN
port 3513 n
rlabel metal5 32020 -63980 32120 -63880 1 PIX3461_IN
port 3514 n
rlabel metal5 33520 -63980 33620 -63880 1 PIX3462_IN
port 3515 n
rlabel metal5 35020 -63980 35120 -63880 1 PIX3463_IN
port 3516 n
rlabel metal5 36520 -63980 36620 -63880 1 PIX3464_IN
port 3517 n
rlabel metal5 38020 -63980 38120 -63880 1 PIX3465_IN
port 3518 n
rlabel metal5 39520 -63980 39620 -63880 1 PIX3466_IN
port 3519 n
rlabel metal5 41020 -63980 41120 -63880 1 PIX3467_IN
port 3520 n
rlabel metal5 42520 -63980 42620 -63880 1 PIX3468_IN
port 3521 n
rlabel metal5 44020 -63980 44120 -63880 1 PIX3469_IN
port 3522 n
rlabel metal5 45520 -63980 45620 -63880 1 PIX3470_IN
port 3523 n
rlabel metal5 47020 -63980 47120 -63880 1 PIX3471_IN
port 3524 n
rlabel metal5 48520 -63980 48620 -63880 1 PIX3472_IN
port 3525 n
rlabel metal5 50020 -63980 50120 -63880 1 PIX3473_IN
port 3526 n
rlabel metal5 51520 -63980 51620 -63880 1 PIX3474_IN
port 3527 n
rlabel metal5 53020 -63980 53120 -63880 1 PIX3475_IN
port 3528 n
rlabel metal5 54520 -63980 54620 -63880 1 PIX3476_IN
port 3529 n
rlabel metal5 56020 -63980 56120 -63880 1 PIX3477_IN
port 3530 n
rlabel metal5 57520 -63980 57620 -63880 1 PIX3478_IN
port 3531 n
rlabel metal5 59020 -63980 59120 -63880 1 PIX3479_IN
port 3532 n
rlabel metal5 60520 -63980 60620 -63880 1 PIX3480_IN
port 3533 n
rlabel metal5 62020 -63980 62120 -63880 1 PIX3481_IN
port 3534 n
rlabel metal5 63520 -63980 63620 -63880 1 PIX3482_IN
port 3535 n
rlabel metal5 65020 -63980 65120 -63880 1 PIX3483_IN
port 3536 n
rlabel metal5 66520 -63980 66620 -63880 1 PIX3484_IN
port 3537 n
rlabel metal5 68020 -63980 68120 -63880 1 PIX3485_IN
port 3538 n
rlabel metal5 69520 -63980 69620 -63880 1 PIX3486_IN
port 3539 n
rlabel metal5 71020 -63980 71120 -63880 1 PIX3487_IN
port 3540 n
rlabel metal5 72520 -63980 72620 -63880 1 PIX3488_IN
port 3541 n
rlabel metal5 74020 -63980 74120 -63880 1 PIX3489_IN
port 3542 n
rlabel metal5 75520 -63980 75620 -63880 1 PIX3490_IN
port 3543 n
rlabel metal5 77020 -63980 77120 -63880 1 PIX3491_IN
port 3544 n
rlabel metal5 78520 -63980 78620 -63880 1 PIX3492_IN
port 3545 n
rlabel metal5 80020 -63980 80120 -63880 1 PIX3493_IN
port 3546 n
rlabel metal5 81520 -63980 81620 -63880 1 PIX3494_IN
port 3547 n
rlabel metal5 83020 -63980 83120 -63880 1 PIX3495_IN
port 3548 n
rlabel metal5 84520 -63980 84620 -63880 1 PIX3496_IN
port 3549 n
rlabel metal5 86020 -63980 86120 -63880 1 PIX3497_IN
port 3550 n
rlabel metal5 87520 -63980 87620 -63880 1 PIX3498_IN
port 3551 n
rlabel metal5 89020 -63980 89120 -63880 1 PIX3499_IN
port 3552 n
rlabel metal5 90520 -63980 90620 -63880 1 PIX3500_IN
port 3553 n
rlabel metal5 92020 -63980 92120 -63880 1 PIX3501_IN
port 3554 n
rlabel metal5 93520 -63980 93620 -63880 1 PIX3502_IN
port 3555 n
rlabel metal5 95020 -63980 95120 -63880 1 PIX3503_IN
port 3556 n
rlabel metal5 96520 -63980 96620 -63880 1 PIX3504_IN
port 3557 n
rlabel metal5 98020 -63980 98120 -63880 1 PIX3505_IN
port 3558 n
rlabel metal5 99520 -63980 99620 -63880 1 PIX3506_IN
port 3559 n
rlabel metal5 101020 -63980 101120 -63880 1 PIX3507_IN
port 3560 n
rlabel metal5 102520 -63980 102620 -63880 1 PIX3508_IN
port 3561 n
rlabel metal5 104020 -63980 104120 -63880 1 PIX3509_IN
port 3562 n
rlabel metal5 105520 -63980 105620 -63880 1 PIX3510_IN
port 3563 n
rlabel metal5 107020 -63980 107120 -63880 1 PIX3511_IN
port 3564 n
rlabel metal5 108520 -63980 108620 -63880 1 PIX3512_IN
port 3565 n
rlabel metal5 110020 -63980 110120 -63880 1 PIX3513_IN
port 3566 n
rlabel metal5 111520 -63980 111620 -63880 1 PIX3514_IN
port 3567 n
rlabel metal5 113020 -63980 113120 -63880 1 PIX3515_IN
port 3568 n
rlabel metal5 114520 -63980 114620 -63880 1 PIX3516_IN
port 3569 n
rlabel metal5 116020 -63980 116120 -63880 1 PIX3517_IN
port 3570 n
rlabel metal5 117520 -63980 117620 -63880 1 PIX3518_IN
port 3571 n
rlabel metal5 119020 -63980 119120 -63880 1 PIX3519_IN
port 3572 n
rlabel metal5 520 -65480 620 -65380 1 PIX3520_IN
port 3573 n
rlabel metal2 -1500 -65260 -1500 -65215 3 ROW_SEL44
port 3574 e
rlabel metal5 2020 -65480 2120 -65380 1 PIX3521_IN
port 3575 n
rlabel metal5 3520 -65480 3620 -65380 1 PIX3522_IN
port 3576 n
rlabel metal5 5020 -65480 5120 -65380 1 PIX3523_IN
port 3577 n
rlabel metal5 6520 -65480 6620 -65380 1 PIX3524_IN
port 3578 n
rlabel metal5 8020 -65480 8120 -65380 1 PIX3525_IN
port 3579 n
rlabel metal5 9520 -65480 9620 -65380 1 PIX3526_IN
port 3580 n
rlabel metal5 11020 -65480 11120 -65380 1 PIX3527_IN
port 3581 n
rlabel metal5 12520 -65480 12620 -65380 1 PIX3528_IN
port 3582 n
rlabel metal5 14020 -65480 14120 -65380 1 PIX3529_IN
port 3583 n
rlabel metal5 15520 -65480 15620 -65380 1 PIX3530_IN
port 3584 n
rlabel metal5 17020 -65480 17120 -65380 1 PIX3531_IN
port 3585 n
rlabel metal5 18520 -65480 18620 -65380 1 PIX3532_IN
port 3586 n
rlabel metal5 20020 -65480 20120 -65380 1 PIX3533_IN
port 3587 n
rlabel metal5 21520 -65480 21620 -65380 1 PIX3534_IN
port 3588 n
rlabel metal5 23020 -65480 23120 -65380 1 PIX3535_IN
port 3589 n
rlabel metal5 24520 -65480 24620 -65380 1 PIX3536_IN
port 3590 n
rlabel metal5 26020 -65480 26120 -65380 1 PIX3537_IN
port 3591 n
rlabel metal5 27520 -65480 27620 -65380 1 PIX3538_IN
port 3592 n
rlabel metal5 29020 -65480 29120 -65380 1 PIX3539_IN
port 3593 n
rlabel metal5 30520 -65480 30620 -65380 1 PIX3540_IN
port 3594 n
rlabel metal5 32020 -65480 32120 -65380 1 PIX3541_IN
port 3595 n
rlabel metal5 33520 -65480 33620 -65380 1 PIX3542_IN
port 3596 n
rlabel metal5 35020 -65480 35120 -65380 1 PIX3543_IN
port 3597 n
rlabel metal5 36520 -65480 36620 -65380 1 PIX3544_IN
port 3598 n
rlabel metal5 38020 -65480 38120 -65380 1 PIX3545_IN
port 3599 n
rlabel metal5 39520 -65480 39620 -65380 1 PIX3546_IN
port 3600 n
rlabel metal5 41020 -65480 41120 -65380 1 PIX3547_IN
port 3601 n
rlabel metal5 42520 -65480 42620 -65380 1 PIX3548_IN
port 3602 n
rlabel metal5 44020 -65480 44120 -65380 1 PIX3549_IN
port 3603 n
rlabel metal5 45520 -65480 45620 -65380 1 PIX3550_IN
port 3604 n
rlabel metal5 47020 -65480 47120 -65380 1 PIX3551_IN
port 3605 n
rlabel metal5 48520 -65480 48620 -65380 1 PIX3552_IN
port 3606 n
rlabel metal5 50020 -65480 50120 -65380 1 PIX3553_IN
port 3607 n
rlabel metal5 51520 -65480 51620 -65380 1 PIX3554_IN
port 3608 n
rlabel metal5 53020 -65480 53120 -65380 1 PIX3555_IN
port 3609 n
rlabel metal5 54520 -65480 54620 -65380 1 PIX3556_IN
port 3610 n
rlabel metal5 56020 -65480 56120 -65380 1 PIX3557_IN
port 3611 n
rlabel metal5 57520 -65480 57620 -65380 1 PIX3558_IN
port 3612 n
rlabel metal5 59020 -65480 59120 -65380 1 PIX3559_IN
port 3613 n
rlabel metal5 60520 -65480 60620 -65380 1 PIX3560_IN
port 3614 n
rlabel metal5 62020 -65480 62120 -65380 1 PIX3561_IN
port 3615 n
rlabel metal5 63520 -65480 63620 -65380 1 PIX3562_IN
port 3616 n
rlabel metal5 65020 -65480 65120 -65380 1 PIX3563_IN
port 3617 n
rlabel metal5 66520 -65480 66620 -65380 1 PIX3564_IN
port 3618 n
rlabel metal5 68020 -65480 68120 -65380 1 PIX3565_IN
port 3619 n
rlabel metal5 69520 -65480 69620 -65380 1 PIX3566_IN
port 3620 n
rlabel metal5 71020 -65480 71120 -65380 1 PIX3567_IN
port 3621 n
rlabel metal5 72520 -65480 72620 -65380 1 PIX3568_IN
port 3622 n
rlabel metal5 74020 -65480 74120 -65380 1 PIX3569_IN
port 3623 n
rlabel metal5 75520 -65480 75620 -65380 1 PIX3570_IN
port 3624 n
rlabel metal5 77020 -65480 77120 -65380 1 PIX3571_IN
port 3625 n
rlabel metal5 78520 -65480 78620 -65380 1 PIX3572_IN
port 3626 n
rlabel metal5 80020 -65480 80120 -65380 1 PIX3573_IN
port 3627 n
rlabel metal5 81520 -65480 81620 -65380 1 PIX3574_IN
port 3628 n
rlabel metal5 83020 -65480 83120 -65380 1 PIX3575_IN
port 3629 n
rlabel metal5 84520 -65480 84620 -65380 1 PIX3576_IN
port 3630 n
rlabel metal5 86020 -65480 86120 -65380 1 PIX3577_IN
port 3631 n
rlabel metal5 87520 -65480 87620 -65380 1 PIX3578_IN
port 3632 n
rlabel metal5 89020 -65480 89120 -65380 1 PIX3579_IN
port 3633 n
rlabel metal5 90520 -65480 90620 -65380 1 PIX3580_IN
port 3634 n
rlabel metal5 92020 -65480 92120 -65380 1 PIX3581_IN
port 3635 n
rlabel metal5 93520 -65480 93620 -65380 1 PIX3582_IN
port 3636 n
rlabel metal5 95020 -65480 95120 -65380 1 PIX3583_IN
port 3637 n
rlabel metal5 96520 -65480 96620 -65380 1 PIX3584_IN
port 3638 n
rlabel metal5 98020 -65480 98120 -65380 1 PIX3585_IN
port 3639 n
rlabel metal5 99520 -65480 99620 -65380 1 PIX3586_IN
port 3640 n
rlabel metal5 101020 -65480 101120 -65380 1 PIX3587_IN
port 3641 n
rlabel metal5 102520 -65480 102620 -65380 1 PIX3588_IN
port 3642 n
rlabel metal5 104020 -65480 104120 -65380 1 PIX3589_IN
port 3643 n
rlabel metal5 105520 -65480 105620 -65380 1 PIX3590_IN
port 3644 n
rlabel metal5 107020 -65480 107120 -65380 1 PIX3591_IN
port 3645 n
rlabel metal5 108520 -65480 108620 -65380 1 PIX3592_IN
port 3646 n
rlabel metal5 110020 -65480 110120 -65380 1 PIX3593_IN
port 3647 n
rlabel metal5 111520 -65480 111620 -65380 1 PIX3594_IN
port 3648 n
rlabel metal5 113020 -65480 113120 -65380 1 PIX3595_IN
port 3649 n
rlabel metal5 114520 -65480 114620 -65380 1 PIX3596_IN
port 3650 n
rlabel metal5 116020 -65480 116120 -65380 1 PIX3597_IN
port 3651 n
rlabel metal5 117520 -65480 117620 -65380 1 PIX3598_IN
port 3652 n
rlabel metal5 119020 -65480 119120 -65380 1 PIX3599_IN
port 3653 n
rlabel metal5 520 -66980 620 -66880 1 PIX3600_IN
port 3654 n
rlabel metal2 -1500 -66760 -1500 -66715 3 ROW_SEL45
port 3655 e
rlabel metal5 2020 -66980 2120 -66880 1 PIX3601_IN
port 3656 n
rlabel metal5 3520 -66980 3620 -66880 1 PIX3602_IN
port 3657 n
rlabel metal5 5020 -66980 5120 -66880 1 PIX3603_IN
port 3658 n
rlabel metal5 6520 -66980 6620 -66880 1 PIX3604_IN
port 3659 n
rlabel metal5 8020 -66980 8120 -66880 1 PIX3605_IN
port 3660 n
rlabel metal5 9520 -66980 9620 -66880 1 PIX3606_IN
port 3661 n
rlabel metal5 11020 -66980 11120 -66880 1 PIX3607_IN
port 3662 n
rlabel metal5 12520 -66980 12620 -66880 1 PIX3608_IN
port 3663 n
rlabel metal5 14020 -66980 14120 -66880 1 PIX3609_IN
port 3664 n
rlabel metal5 15520 -66980 15620 -66880 1 PIX3610_IN
port 3665 n
rlabel metal5 17020 -66980 17120 -66880 1 PIX3611_IN
port 3666 n
rlabel metal5 18520 -66980 18620 -66880 1 PIX3612_IN
port 3667 n
rlabel metal5 20020 -66980 20120 -66880 1 PIX3613_IN
port 3668 n
rlabel metal5 21520 -66980 21620 -66880 1 PIX3614_IN
port 3669 n
rlabel metal5 23020 -66980 23120 -66880 1 PIX3615_IN
port 3670 n
rlabel metal5 24520 -66980 24620 -66880 1 PIX3616_IN
port 3671 n
rlabel metal5 26020 -66980 26120 -66880 1 PIX3617_IN
port 3672 n
rlabel metal5 27520 -66980 27620 -66880 1 PIX3618_IN
port 3673 n
rlabel metal5 29020 -66980 29120 -66880 1 PIX3619_IN
port 3674 n
rlabel metal5 30520 -66980 30620 -66880 1 PIX3620_IN
port 3675 n
rlabel metal5 32020 -66980 32120 -66880 1 PIX3621_IN
port 3676 n
rlabel metal5 33520 -66980 33620 -66880 1 PIX3622_IN
port 3677 n
rlabel metal5 35020 -66980 35120 -66880 1 PIX3623_IN
port 3678 n
rlabel metal5 36520 -66980 36620 -66880 1 PIX3624_IN
port 3679 n
rlabel metal5 38020 -66980 38120 -66880 1 PIX3625_IN
port 3680 n
rlabel metal5 39520 -66980 39620 -66880 1 PIX3626_IN
port 3681 n
rlabel metal5 41020 -66980 41120 -66880 1 PIX3627_IN
port 3682 n
rlabel metal5 42520 -66980 42620 -66880 1 PIX3628_IN
port 3683 n
rlabel metal5 44020 -66980 44120 -66880 1 PIX3629_IN
port 3684 n
rlabel metal5 45520 -66980 45620 -66880 1 PIX3630_IN
port 3685 n
rlabel metal5 47020 -66980 47120 -66880 1 PIX3631_IN
port 3686 n
rlabel metal5 48520 -66980 48620 -66880 1 PIX3632_IN
port 3687 n
rlabel metal5 50020 -66980 50120 -66880 1 PIX3633_IN
port 3688 n
rlabel metal5 51520 -66980 51620 -66880 1 PIX3634_IN
port 3689 n
rlabel metal5 53020 -66980 53120 -66880 1 PIX3635_IN
port 3690 n
rlabel metal5 54520 -66980 54620 -66880 1 PIX3636_IN
port 3691 n
rlabel metal5 56020 -66980 56120 -66880 1 PIX3637_IN
port 3692 n
rlabel metal5 57520 -66980 57620 -66880 1 PIX3638_IN
port 3693 n
rlabel metal5 59020 -66980 59120 -66880 1 PIX3639_IN
port 3694 n
rlabel metal5 60520 -66980 60620 -66880 1 PIX3640_IN
port 3695 n
rlabel metal5 62020 -66980 62120 -66880 1 PIX3641_IN
port 3696 n
rlabel metal5 63520 -66980 63620 -66880 1 PIX3642_IN
port 3697 n
rlabel metal5 65020 -66980 65120 -66880 1 PIX3643_IN
port 3698 n
rlabel metal5 66520 -66980 66620 -66880 1 PIX3644_IN
port 3699 n
rlabel metal5 68020 -66980 68120 -66880 1 PIX3645_IN
port 3700 n
rlabel metal5 69520 -66980 69620 -66880 1 PIX3646_IN
port 3701 n
rlabel metal5 71020 -66980 71120 -66880 1 PIX3647_IN
port 3702 n
rlabel metal5 72520 -66980 72620 -66880 1 PIX3648_IN
port 3703 n
rlabel metal5 74020 -66980 74120 -66880 1 PIX3649_IN
port 3704 n
rlabel metal5 75520 -66980 75620 -66880 1 PIX3650_IN
port 3705 n
rlabel metal5 77020 -66980 77120 -66880 1 PIX3651_IN
port 3706 n
rlabel metal5 78520 -66980 78620 -66880 1 PIX3652_IN
port 3707 n
rlabel metal5 80020 -66980 80120 -66880 1 PIX3653_IN
port 3708 n
rlabel metal5 81520 -66980 81620 -66880 1 PIX3654_IN
port 3709 n
rlabel metal5 83020 -66980 83120 -66880 1 PIX3655_IN
port 3710 n
rlabel metal5 84520 -66980 84620 -66880 1 PIX3656_IN
port 3711 n
rlabel metal5 86020 -66980 86120 -66880 1 PIX3657_IN
port 3712 n
rlabel metal5 87520 -66980 87620 -66880 1 PIX3658_IN
port 3713 n
rlabel metal5 89020 -66980 89120 -66880 1 PIX3659_IN
port 3714 n
rlabel metal5 90520 -66980 90620 -66880 1 PIX3660_IN
port 3715 n
rlabel metal5 92020 -66980 92120 -66880 1 PIX3661_IN
port 3716 n
rlabel metal5 93520 -66980 93620 -66880 1 PIX3662_IN
port 3717 n
rlabel metal5 95020 -66980 95120 -66880 1 PIX3663_IN
port 3718 n
rlabel metal5 96520 -66980 96620 -66880 1 PIX3664_IN
port 3719 n
rlabel metal5 98020 -66980 98120 -66880 1 PIX3665_IN
port 3720 n
rlabel metal5 99520 -66980 99620 -66880 1 PIX3666_IN
port 3721 n
rlabel metal5 101020 -66980 101120 -66880 1 PIX3667_IN
port 3722 n
rlabel metal5 102520 -66980 102620 -66880 1 PIX3668_IN
port 3723 n
rlabel metal5 104020 -66980 104120 -66880 1 PIX3669_IN
port 3724 n
rlabel metal5 105520 -66980 105620 -66880 1 PIX3670_IN
port 3725 n
rlabel metal5 107020 -66980 107120 -66880 1 PIX3671_IN
port 3726 n
rlabel metal5 108520 -66980 108620 -66880 1 PIX3672_IN
port 3727 n
rlabel metal5 110020 -66980 110120 -66880 1 PIX3673_IN
port 3728 n
rlabel metal5 111520 -66980 111620 -66880 1 PIX3674_IN
port 3729 n
rlabel metal5 113020 -66980 113120 -66880 1 PIX3675_IN
port 3730 n
rlabel metal5 114520 -66980 114620 -66880 1 PIX3676_IN
port 3731 n
rlabel metal5 116020 -66980 116120 -66880 1 PIX3677_IN
port 3732 n
rlabel metal5 117520 -66980 117620 -66880 1 PIX3678_IN
port 3733 n
rlabel metal5 119020 -66980 119120 -66880 1 PIX3679_IN
port 3734 n
rlabel metal5 520 -68480 620 -68380 1 PIX3680_IN
port 3735 n
rlabel metal2 -1500 -68260 -1500 -68215 3 ROW_SEL46
port 3736 e
rlabel metal5 2020 -68480 2120 -68380 1 PIX3681_IN
port 3737 n
rlabel metal5 3520 -68480 3620 -68380 1 PIX3682_IN
port 3738 n
rlabel metal5 5020 -68480 5120 -68380 1 PIX3683_IN
port 3739 n
rlabel metal5 6520 -68480 6620 -68380 1 PIX3684_IN
port 3740 n
rlabel metal5 8020 -68480 8120 -68380 1 PIX3685_IN
port 3741 n
rlabel metal5 9520 -68480 9620 -68380 1 PIX3686_IN
port 3742 n
rlabel metal5 11020 -68480 11120 -68380 1 PIX3687_IN
port 3743 n
rlabel metal5 12520 -68480 12620 -68380 1 PIX3688_IN
port 3744 n
rlabel metal5 14020 -68480 14120 -68380 1 PIX3689_IN
port 3745 n
rlabel metal5 15520 -68480 15620 -68380 1 PIX3690_IN
port 3746 n
rlabel metal5 17020 -68480 17120 -68380 1 PIX3691_IN
port 3747 n
rlabel metal5 18520 -68480 18620 -68380 1 PIX3692_IN
port 3748 n
rlabel metal5 20020 -68480 20120 -68380 1 PIX3693_IN
port 3749 n
rlabel metal5 21520 -68480 21620 -68380 1 PIX3694_IN
port 3750 n
rlabel metal5 23020 -68480 23120 -68380 1 PIX3695_IN
port 3751 n
rlabel metal5 24520 -68480 24620 -68380 1 PIX3696_IN
port 3752 n
rlabel metal5 26020 -68480 26120 -68380 1 PIX3697_IN
port 3753 n
rlabel metal5 27520 -68480 27620 -68380 1 PIX3698_IN
port 3754 n
rlabel metal5 29020 -68480 29120 -68380 1 PIX3699_IN
port 3755 n
rlabel metal5 30520 -68480 30620 -68380 1 PIX3700_IN
port 3756 n
rlabel metal5 32020 -68480 32120 -68380 1 PIX3701_IN
port 3757 n
rlabel metal5 33520 -68480 33620 -68380 1 PIX3702_IN
port 3758 n
rlabel metal5 35020 -68480 35120 -68380 1 PIX3703_IN
port 3759 n
rlabel metal5 36520 -68480 36620 -68380 1 PIX3704_IN
port 3760 n
rlabel metal5 38020 -68480 38120 -68380 1 PIX3705_IN
port 3761 n
rlabel metal5 39520 -68480 39620 -68380 1 PIX3706_IN
port 3762 n
rlabel metal5 41020 -68480 41120 -68380 1 PIX3707_IN
port 3763 n
rlabel metal5 42520 -68480 42620 -68380 1 PIX3708_IN
port 3764 n
rlabel metal5 44020 -68480 44120 -68380 1 PIX3709_IN
port 3765 n
rlabel metal5 45520 -68480 45620 -68380 1 PIX3710_IN
port 3766 n
rlabel metal5 47020 -68480 47120 -68380 1 PIX3711_IN
port 3767 n
rlabel metal5 48520 -68480 48620 -68380 1 PIX3712_IN
port 3768 n
rlabel metal5 50020 -68480 50120 -68380 1 PIX3713_IN
port 3769 n
rlabel metal5 51520 -68480 51620 -68380 1 PIX3714_IN
port 3770 n
rlabel metal5 53020 -68480 53120 -68380 1 PIX3715_IN
port 3771 n
rlabel metal5 54520 -68480 54620 -68380 1 PIX3716_IN
port 3772 n
rlabel metal5 56020 -68480 56120 -68380 1 PIX3717_IN
port 3773 n
rlabel metal5 57520 -68480 57620 -68380 1 PIX3718_IN
port 3774 n
rlabel metal5 59020 -68480 59120 -68380 1 PIX3719_IN
port 3775 n
rlabel metal5 60520 -68480 60620 -68380 1 PIX3720_IN
port 3776 n
rlabel metal5 62020 -68480 62120 -68380 1 PIX3721_IN
port 3777 n
rlabel metal5 63520 -68480 63620 -68380 1 PIX3722_IN
port 3778 n
rlabel metal5 65020 -68480 65120 -68380 1 PIX3723_IN
port 3779 n
rlabel metal5 66520 -68480 66620 -68380 1 PIX3724_IN
port 3780 n
rlabel metal5 68020 -68480 68120 -68380 1 PIX3725_IN
port 3781 n
rlabel metal5 69520 -68480 69620 -68380 1 PIX3726_IN
port 3782 n
rlabel metal5 71020 -68480 71120 -68380 1 PIX3727_IN
port 3783 n
rlabel metal5 72520 -68480 72620 -68380 1 PIX3728_IN
port 3784 n
rlabel metal5 74020 -68480 74120 -68380 1 PIX3729_IN
port 3785 n
rlabel metal5 75520 -68480 75620 -68380 1 PIX3730_IN
port 3786 n
rlabel metal5 77020 -68480 77120 -68380 1 PIX3731_IN
port 3787 n
rlabel metal5 78520 -68480 78620 -68380 1 PIX3732_IN
port 3788 n
rlabel metal5 80020 -68480 80120 -68380 1 PIX3733_IN
port 3789 n
rlabel metal5 81520 -68480 81620 -68380 1 PIX3734_IN
port 3790 n
rlabel metal5 83020 -68480 83120 -68380 1 PIX3735_IN
port 3791 n
rlabel metal5 84520 -68480 84620 -68380 1 PIX3736_IN
port 3792 n
rlabel metal5 86020 -68480 86120 -68380 1 PIX3737_IN
port 3793 n
rlabel metal5 87520 -68480 87620 -68380 1 PIX3738_IN
port 3794 n
rlabel metal5 89020 -68480 89120 -68380 1 PIX3739_IN
port 3795 n
rlabel metal5 90520 -68480 90620 -68380 1 PIX3740_IN
port 3796 n
rlabel metal5 92020 -68480 92120 -68380 1 PIX3741_IN
port 3797 n
rlabel metal5 93520 -68480 93620 -68380 1 PIX3742_IN
port 3798 n
rlabel metal5 95020 -68480 95120 -68380 1 PIX3743_IN
port 3799 n
rlabel metal5 96520 -68480 96620 -68380 1 PIX3744_IN
port 3800 n
rlabel metal5 98020 -68480 98120 -68380 1 PIX3745_IN
port 3801 n
rlabel metal5 99520 -68480 99620 -68380 1 PIX3746_IN
port 3802 n
rlabel metal5 101020 -68480 101120 -68380 1 PIX3747_IN
port 3803 n
rlabel metal5 102520 -68480 102620 -68380 1 PIX3748_IN
port 3804 n
rlabel metal5 104020 -68480 104120 -68380 1 PIX3749_IN
port 3805 n
rlabel metal5 105520 -68480 105620 -68380 1 PIX3750_IN
port 3806 n
rlabel metal5 107020 -68480 107120 -68380 1 PIX3751_IN
port 3807 n
rlabel metal5 108520 -68480 108620 -68380 1 PIX3752_IN
port 3808 n
rlabel metal5 110020 -68480 110120 -68380 1 PIX3753_IN
port 3809 n
rlabel metal5 111520 -68480 111620 -68380 1 PIX3754_IN
port 3810 n
rlabel metal5 113020 -68480 113120 -68380 1 PIX3755_IN
port 3811 n
rlabel metal5 114520 -68480 114620 -68380 1 PIX3756_IN
port 3812 n
rlabel metal5 116020 -68480 116120 -68380 1 PIX3757_IN
port 3813 n
rlabel metal5 117520 -68480 117620 -68380 1 PIX3758_IN
port 3814 n
rlabel metal5 119020 -68480 119120 -68380 1 PIX3759_IN
port 3815 n
rlabel metal5 520 -69980 620 -69880 1 PIX3760_IN
port 3816 n
rlabel metal2 -1500 -69760 -1500 -69715 3 ROW_SEL47
port 3817 e
rlabel metal5 2020 -69980 2120 -69880 1 PIX3761_IN
port 3818 n
rlabel metal5 3520 -69980 3620 -69880 1 PIX3762_IN
port 3819 n
rlabel metal5 5020 -69980 5120 -69880 1 PIX3763_IN
port 3820 n
rlabel metal5 6520 -69980 6620 -69880 1 PIX3764_IN
port 3821 n
rlabel metal5 8020 -69980 8120 -69880 1 PIX3765_IN
port 3822 n
rlabel metal5 9520 -69980 9620 -69880 1 PIX3766_IN
port 3823 n
rlabel metal5 11020 -69980 11120 -69880 1 PIX3767_IN
port 3824 n
rlabel metal5 12520 -69980 12620 -69880 1 PIX3768_IN
port 3825 n
rlabel metal5 14020 -69980 14120 -69880 1 PIX3769_IN
port 3826 n
rlabel metal5 15520 -69980 15620 -69880 1 PIX3770_IN
port 3827 n
rlabel metal5 17020 -69980 17120 -69880 1 PIX3771_IN
port 3828 n
rlabel metal5 18520 -69980 18620 -69880 1 PIX3772_IN
port 3829 n
rlabel metal5 20020 -69980 20120 -69880 1 PIX3773_IN
port 3830 n
rlabel metal5 21520 -69980 21620 -69880 1 PIX3774_IN
port 3831 n
rlabel metal5 23020 -69980 23120 -69880 1 PIX3775_IN
port 3832 n
rlabel metal5 24520 -69980 24620 -69880 1 PIX3776_IN
port 3833 n
rlabel metal5 26020 -69980 26120 -69880 1 PIX3777_IN
port 3834 n
rlabel metal5 27520 -69980 27620 -69880 1 PIX3778_IN
port 3835 n
rlabel metal5 29020 -69980 29120 -69880 1 PIX3779_IN
port 3836 n
rlabel metal5 30520 -69980 30620 -69880 1 PIX3780_IN
port 3837 n
rlabel metal5 32020 -69980 32120 -69880 1 PIX3781_IN
port 3838 n
rlabel metal5 33520 -69980 33620 -69880 1 PIX3782_IN
port 3839 n
rlabel metal5 35020 -69980 35120 -69880 1 PIX3783_IN
port 3840 n
rlabel metal5 36520 -69980 36620 -69880 1 PIX3784_IN
port 3841 n
rlabel metal5 38020 -69980 38120 -69880 1 PIX3785_IN
port 3842 n
rlabel metal5 39520 -69980 39620 -69880 1 PIX3786_IN
port 3843 n
rlabel metal5 41020 -69980 41120 -69880 1 PIX3787_IN
port 3844 n
rlabel metal5 42520 -69980 42620 -69880 1 PIX3788_IN
port 3845 n
rlabel metal5 44020 -69980 44120 -69880 1 PIX3789_IN
port 3846 n
rlabel metal5 45520 -69980 45620 -69880 1 PIX3790_IN
port 3847 n
rlabel metal5 47020 -69980 47120 -69880 1 PIX3791_IN
port 3848 n
rlabel metal5 48520 -69980 48620 -69880 1 PIX3792_IN
port 3849 n
rlabel metal5 50020 -69980 50120 -69880 1 PIX3793_IN
port 3850 n
rlabel metal5 51520 -69980 51620 -69880 1 PIX3794_IN
port 3851 n
rlabel metal5 53020 -69980 53120 -69880 1 PIX3795_IN
port 3852 n
rlabel metal5 54520 -69980 54620 -69880 1 PIX3796_IN
port 3853 n
rlabel metal5 56020 -69980 56120 -69880 1 PIX3797_IN
port 3854 n
rlabel metal5 57520 -69980 57620 -69880 1 PIX3798_IN
port 3855 n
rlabel metal5 59020 -69980 59120 -69880 1 PIX3799_IN
port 3856 n
rlabel metal5 60520 -69980 60620 -69880 1 PIX3800_IN
port 3857 n
rlabel metal5 62020 -69980 62120 -69880 1 PIX3801_IN
port 3858 n
rlabel metal5 63520 -69980 63620 -69880 1 PIX3802_IN
port 3859 n
rlabel metal5 65020 -69980 65120 -69880 1 PIX3803_IN
port 3860 n
rlabel metal5 66520 -69980 66620 -69880 1 PIX3804_IN
port 3861 n
rlabel metal5 68020 -69980 68120 -69880 1 PIX3805_IN
port 3862 n
rlabel metal5 69520 -69980 69620 -69880 1 PIX3806_IN
port 3863 n
rlabel metal5 71020 -69980 71120 -69880 1 PIX3807_IN
port 3864 n
rlabel metal5 72520 -69980 72620 -69880 1 PIX3808_IN
port 3865 n
rlabel metal5 74020 -69980 74120 -69880 1 PIX3809_IN
port 3866 n
rlabel metal5 75520 -69980 75620 -69880 1 PIX3810_IN
port 3867 n
rlabel metal5 77020 -69980 77120 -69880 1 PIX3811_IN
port 3868 n
rlabel metal5 78520 -69980 78620 -69880 1 PIX3812_IN
port 3869 n
rlabel metal5 80020 -69980 80120 -69880 1 PIX3813_IN
port 3870 n
rlabel metal5 81520 -69980 81620 -69880 1 PIX3814_IN
port 3871 n
rlabel metal5 83020 -69980 83120 -69880 1 PIX3815_IN
port 3872 n
rlabel metal5 84520 -69980 84620 -69880 1 PIX3816_IN
port 3873 n
rlabel metal5 86020 -69980 86120 -69880 1 PIX3817_IN
port 3874 n
rlabel metal5 87520 -69980 87620 -69880 1 PIX3818_IN
port 3875 n
rlabel metal5 89020 -69980 89120 -69880 1 PIX3819_IN
port 3876 n
rlabel metal5 90520 -69980 90620 -69880 1 PIX3820_IN
port 3877 n
rlabel metal5 92020 -69980 92120 -69880 1 PIX3821_IN
port 3878 n
rlabel metal5 93520 -69980 93620 -69880 1 PIX3822_IN
port 3879 n
rlabel metal5 95020 -69980 95120 -69880 1 PIX3823_IN
port 3880 n
rlabel metal5 96520 -69980 96620 -69880 1 PIX3824_IN
port 3881 n
rlabel metal5 98020 -69980 98120 -69880 1 PIX3825_IN
port 3882 n
rlabel metal5 99520 -69980 99620 -69880 1 PIX3826_IN
port 3883 n
rlabel metal5 101020 -69980 101120 -69880 1 PIX3827_IN
port 3884 n
rlabel metal5 102520 -69980 102620 -69880 1 PIX3828_IN
port 3885 n
rlabel metal5 104020 -69980 104120 -69880 1 PIX3829_IN
port 3886 n
rlabel metal5 105520 -69980 105620 -69880 1 PIX3830_IN
port 3887 n
rlabel metal5 107020 -69980 107120 -69880 1 PIX3831_IN
port 3888 n
rlabel metal5 108520 -69980 108620 -69880 1 PIX3832_IN
port 3889 n
rlabel metal5 110020 -69980 110120 -69880 1 PIX3833_IN
port 3890 n
rlabel metal5 111520 -69980 111620 -69880 1 PIX3834_IN
port 3891 n
rlabel metal5 113020 -69980 113120 -69880 1 PIX3835_IN
port 3892 n
rlabel metal5 114520 -69980 114620 -69880 1 PIX3836_IN
port 3893 n
rlabel metal5 116020 -69980 116120 -69880 1 PIX3837_IN
port 3894 n
rlabel metal5 117520 -69980 117620 -69880 1 PIX3838_IN
port 3895 n
rlabel metal5 119020 -69980 119120 -69880 1 PIX3839_IN
port 3896 n
rlabel metal5 520 -71480 620 -71380 1 PIX3840_IN
port 3897 n
rlabel metal2 -1500 -71260 -1500 -71215 3 ROW_SEL48
port 3898 e
rlabel metal5 2020 -71480 2120 -71380 1 PIX3841_IN
port 3899 n
rlabel metal5 3520 -71480 3620 -71380 1 PIX3842_IN
port 3900 n
rlabel metal5 5020 -71480 5120 -71380 1 PIX3843_IN
port 3901 n
rlabel metal5 6520 -71480 6620 -71380 1 PIX3844_IN
port 3902 n
rlabel metal5 8020 -71480 8120 -71380 1 PIX3845_IN
port 3903 n
rlabel metal5 9520 -71480 9620 -71380 1 PIX3846_IN
port 3904 n
rlabel metal5 11020 -71480 11120 -71380 1 PIX3847_IN
port 3905 n
rlabel metal5 12520 -71480 12620 -71380 1 PIX3848_IN
port 3906 n
rlabel metal5 14020 -71480 14120 -71380 1 PIX3849_IN
port 3907 n
rlabel metal5 15520 -71480 15620 -71380 1 PIX3850_IN
port 3908 n
rlabel metal5 17020 -71480 17120 -71380 1 PIX3851_IN
port 3909 n
rlabel metal5 18520 -71480 18620 -71380 1 PIX3852_IN
port 3910 n
rlabel metal5 20020 -71480 20120 -71380 1 PIX3853_IN
port 3911 n
rlabel metal5 21520 -71480 21620 -71380 1 PIX3854_IN
port 3912 n
rlabel metal5 23020 -71480 23120 -71380 1 PIX3855_IN
port 3913 n
rlabel metal5 24520 -71480 24620 -71380 1 PIX3856_IN
port 3914 n
rlabel metal5 26020 -71480 26120 -71380 1 PIX3857_IN
port 3915 n
rlabel metal5 27520 -71480 27620 -71380 1 PIX3858_IN
port 3916 n
rlabel metal5 29020 -71480 29120 -71380 1 PIX3859_IN
port 3917 n
rlabel metal5 30520 -71480 30620 -71380 1 PIX3860_IN
port 3918 n
rlabel metal5 32020 -71480 32120 -71380 1 PIX3861_IN
port 3919 n
rlabel metal5 33520 -71480 33620 -71380 1 PIX3862_IN
port 3920 n
rlabel metal5 35020 -71480 35120 -71380 1 PIX3863_IN
port 3921 n
rlabel metal5 36520 -71480 36620 -71380 1 PIX3864_IN
port 3922 n
rlabel metal5 38020 -71480 38120 -71380 1 PIX3865_IN
port 3923 n
rlabel metal5 39520 -71480 39620 -71380 1 PIX3866_IN
port 3924 n
rlabel metal5 41020 -71480 41120 -71380 1 PIX3867_IN
port 3925 n
rlabel metal5 42520 -71480 42620 -71380 1 PIX3868_IN
port 3926 n
rlabel metal5 44020 -71480 44120 -71380 1 PIX3869_IN
port 3927 n
rlabel metal5 45520 -71480 45620 -71380 1 PIX3870_IN
port 3928 n
rlabel metal5 47020 -71480 47120 -71380 1 PIX3871_IN
port 3929 n
rlabel metal5 48520 -71480 48620 -71380 1 PIX3872_IN
port 3930 n
rlabel metal5 50020 -71480 50120 -71380 1 PIX3873_IN
port 3931 n
rlabel metal5 51520 -71480 51620 -71380 1 PIX3874_IN
port 3932 n
rlabel metal5 53020 -71480 53120 -71380 1 PIX3875_IN
port 3933 n
rlabel metal5 54520 -71480 54620 -71380 1 PIX3876_IN
port 3934 n
rlabel metal5 56020 -71480 56120 -71380 1 PIX3877_IN
port 3935 n
rlabel metal5 57520 -71480 57620 -71380 1 PIX3878_IN
port 3936 n
rlabel metal5 59020 -71480 59120 -71380 1 PIX3879_IN
port 3937 n
rlabel metal5 60520 -71480 60620 -71380 1 PIX3880_IN
port 3938 n
rlabel metal5 62020 -71480 62120 -71380 1 PIX3881_IN
port 3939 n
rlabel metal5 63520 -71480 63620 -71380 1 PIX3882_IN
port 3940 n
rlabel metal5 65020 -71480 65120 -71380 1 PIX3883_IN
port 3941 n
rlabel metal5 66520 -71480 66620 -71380 1 PIX3884_IN
port 3942 n
rlabel metal5 68020 -71480 68120 -71380 1 PIX3885_IN
port 3943 n
rlabel metal5 69520 -71480 69620 -71380 1 PIX3886_IN
port 3944 n
rlabel metal5 71020 -71480 71120 -71380 1 PIX3887_IN
port 3945 n
rlabel metal5 72520 -71480 72620 -71380 1 PIX3888_IN
port 3946 n
rlabel metal5 74020 -71480 74120 -71380 1 PIX3889_IN
port 3947 n
rlabel metal5 75520 -71480 75620 -71380 1 PIX3890_IN
port 3948 n
rlabel metal5 77020 -71480 77120 -71380 1 PIX3891_IN
port 3949 n
rlabel metal5 78520 -71480 78620 -71380 1 PIX3892_IN
port 3950 n
rlabel metal5 80020 -71480 80120 -71380 1 PIX3893_IN
port 3951 n
rlabel metal5 81520 -71480 81620 -71380 1 PIX3894_IN
port 3952 n
rlabel metal5 83020 -71480 83120 -71380 1 PIX3895_IN
port 3953 n
rlabel metal5 84520 -71480 84620 -71380 1 PIX3896_IN
port 3954 n
rlabel metal5 86020 -71480 86120 -71380 1 PIX3897_IN
port 3955 n
rlabel metal5 87520 -71480 87620 -71380 1 PIX3898_IN
port 3956 n
rlabel metal5 89020 -71480 89120 -71380 1 PIX3899_IN
port 3957 n
rlabel metal5 90520 -71480 90620 -71380 1 PIX3900_IN
port 3958 n
rlabel metal5 92020 -71480 92120 -71380 1 PIX3901_IN
port 3959 n
rlabel metal5 93520 -71480 93620 -71380 1 PIX3902_IN
port 3960 n
rlabel metal5 95020 -71480 95120 -71380 1 PIX3903_IN
port 3961 n
rlabel metal5 96520 -71480 96620 -71380 1 PIX3904_IN
port 3962 n
rlabel metal5 98020 -71480 98120 -71380 1 PIX3905_IN
port 3963 n
rlabel metal5 99520 -71480 99620 -71380 1 PIX3906_IN
port 3964 n
rlabel metal5 101020 -71480 101120 -71380 1 PIX3907_IN
port 3965 n
rlabel metal5 102520 -71480 102620 -71380 1 PIX3908_IN
port 3966 n
rlabel metal5 104020 -71480 104120 -71380 1 PIX3909_IN
port 3967 n
rlabel metal5 105520 -71480 105620 -71380 1 PIX3910_IN
port 3968 n
rlabel metal5 107020 -71480 107120 -71380 1 PIX3911_IN
port 3969 n
rlabel metal5 108520 -71480 108620 -71380 1 PIX3912_IN
port 3970 n
rlabel metal5 110020 -71480 110120 -71380 1 PIX3913_IN
port 3971 n
rlabel metal5 111520 -71480 111620 -71380 1 PIX3914_IN
port 3972 n
rlabel metal5 113020 -71480 113120 -71380 1 PIX3915_IN
port 3973 n
rlabel metal5 114520 -71480 114620 -71380 1 PIX3916_IN
port 3974 n
rlabel metal5 116020 -71480 116120 -71380 1 PIX3917_IN
port 3975 n
rlabel metal5 117520 -71480 117620 -71380 1 PIX3918_IN
port 3976 n
rlabel metal5 119020 -71480 119120 -71380 1 PIX3919_IN
port 3977 n
rlabel metal5 520 -72980 620 -72880 1 PIX3920_IN
port 3978 n
rlabel metal2 -1500 -72760 -1500 -72715 3 ROW_SEL49
port 3979 e
rlabel metal5 2020 -72980 2120 -72880 1 PIX3921_IN
port 3980 n
rlabel metal5 3520 -72980 3620 -72880 1 PIX3922_IN
port 3981 n
rlabel metal5 5020 -72980 5120 -72880 1 PIX3923_IN
port 3982 n
rlabel metal5 6520 -72980 6620 -72880 1 PIX3924_IN
port 3983 n
rlabel metal5 8020 -72980 8120 -72880 1 PIX3925_IN
port 3984 n
rlabel metal5 9520 -72980 9620 -72880 1 PIX3926_IN
port 3985 n
rlabel metal5 11020 -72980 11120 -72880 1 PIX3927_IN
port 3986 n
rlabel metal5 12520 -72980 12620 -72880 1 PIX3928_IN
port 3987 n
rlabel metal5 14020 -72980 14120 -72880 1 PIX3929_IN
port 3988 n
rlabel metal5 15520 -72980 15620 -72880 1 PIX3930_IN
port 3989 n
rlabel metal5 17020 -72980 17120 -72880 1 PIX3931_IN
port 3990 n
rlabel metal5 18520 -72980 18620 -72880 1 PIX3932_IN
port 3991 n
rlabel metal5 20020 -72980 20120 -72880 1 PIX3933_IN
port 3992 n
rlabel metal5 21520 -72980 21620 -72880 1 PIX3934_IN
port 3993 n
rlabel metal5 23020 -72980 23120 -72880 1 PIX3935_IN
port 3994 n
rlabel metal5 24520 -72980 24620 -72880 1 PIX3936_IN
port 3995 n
rlabel metal5 26020 -72980 26120 -72880 1 PIX3937_IN
port 3996 n
rlabel metal5 27520 -72980 27620 -72880 1 PIX3938_IN
port 3997 n
rlabel metal5 29020 -72980 29120 -72880 1 PIX3939_IN
port 3998 n
rlabel metal5 30520 -72980 30620 -72880 1 PIX3940_IN
port 3999 n
rlabel metal5 32020 -72980 32120 -72880 1 PIX3941_IN
port 4000 n
rlabel metal5 33520 -72980 33620 -72880 1 PIX3942_IN
port 4001 n
rlabel metal5 35020 -72980 35120 -72880 1 PIX3943_IN
port 4002 n
rlabel metal5 36520 -72980 36620 -72880 1 PIX3944_IN
port 4003 n
rlabel metal5 38020 -72980 38120 -72880 1 PIX3945_IN
port 4004 n
rlabel metal5 39520 -72980 39620 -72880 1 PIX3946_IN
port 4005 n
rlabel metal5 41020 -72980 41120 -72880 1 PIX3947_IN
port 4006 n
rlabel metal5 42520 -72980 42620 -72880 1 PIX3948_IN
port 4007 n
rlabel metal5 44020 -72980 44120 -72880 1 PIX3949_IN
port 4008 n
rlabel metal5 45520 -72980 45620 -72880 1 PIX3950_IN
port 4009 n
rlabel metal5 47020 -72980 47120 -72880 1 PIX3951_IN
port 4010 n
rlabel metal5 48520 -72980 48620 -72880 1 PIX3952_IN
port 4011 n
rlabel metal5 50020 -72980 50120 -72880 1 PIX3953_IN
port 4012 n
rlabel metal5 51520 -72980 51620 -72880 1 PIX3954_IN
port 4013 n
rlabel metal5 53020 -72980 53120 -72880 1 PIX3955_IN
port 4014 n
rlabel metal5 54520 -72980 54620 -72880 1 PIX3956_IN
port 4015 n
rlabel metal5 56020 -72980 56120 -72880 1 PIX3957_IN
port 4016 n
rlabel metal5 57520 -72980 57620 -72880 1 PIX3958_IN
port 4017 n
rlabel metal5 59020 -72980 59120 -72880 1 PIX3959_IN
port 4018 n
rlabel metal5 60520 -72980 60620 -72880 1 PIX3960_IN
port 4019 n
rlabel metal5 62020 -72980 62120 -72880 1 PIX3961_IN
port 4020 n
rlabel metal5 63520 -72980 63620 -72880 1 PIX3962_IN
port 4021 n
rlabel metal5 65020 -72980 65120 -72880 1 PIX3963_IN
port 4022 n
rlabel metal5 66520 -72980 66620 -72880 1 PIX3964_IN
port 4023 n
rlabel metal5 68020 -72980 68120 -72880 1 PIX3965_IN
port 4024 n
rlabel metal5 69520 -72980 69620 -72880 1 PIX3966_IN
port 4025 n
rlabel metal5 71020 -72980 71120 -72880 1 PIX3967_IN
port 4026 n
rlabel metal5 72520 -72980 72620 -72880 1 PIX3968_IN
port 4027 n
rlabel metal5 74020 -72980 74120 -72880 1 PIX3969_IN
port 4028 n
rlabel metal5 75520 -72980 75620 -72880 1 PIX3970_IN
port 4029 n
rlabel metal5 77020 -72980 77120 -72880 1 PIX3971_IN
port 4030 n
rlabel metal5 78520 -72980 78620 -72880 1 PIX3972_IN
port 4031 n
rlabel metal5 80020 -72980 80120 -72880 1 PIX3973_IN
port 4032 n
rlabel metal5 81520 -72980 81620 -72880 1 PIX3974_IN
port 4033 n
rlabel metal5 83020 -72980 83120 -72880 1 PIX3975_IN
port 4034 n
rlabel metal5 84520 -72980 84620 -72880 1 PIX3976_IN
port 4035 n
rlabel metal5 86020 -72980 86120 -72880 1 PIX3977_IN
port 4036 n
rlabel metal5 87520 -72980 87620 -72880 1 PIX3978_IN
port 4037 n
rlabel metal5 89020 -72980 89120 -72880 1 PIX3979_IN
port 4038 n
rlabel metal5 90520 -72980 90620 -72880 1 PIX3980_IN
port 4039 n
rlabel metal5 92020 -72980 92120 -72880 1 PIX3981_IN
port 4040 n
rlabel metal5 93520 -72980 93620 -72880 1 PIX3982_IN
port 4041 n
rlabel metal5 95020 -72980 95120 -72880 1 PIX3983_IN
port 4042 n
rlabel metal5 96520 -72980 96620 -72880 1 PIX3984_IN
port 4043 n
rlabel metal5 98020 -72980 98120 -72880 1 PIX3985_IN
port 4044 n
rlabel metal5 99520 -72980 99620 -72880 1 PIX3986_IN
port 4045 n
rlabel metal5 101020 -72980 101120 -72880 1 PIX3987_IN
port 4046 n
rlabel metal5 102520 -72980 102620 -72880 1 PIX3988_IN
port 4047 n
rlabel metal5 104020 -72980 104120 -72880 1 PIX3989_IN
port 4048 n
rlabel metal5 105520 -72980 105620 -72880 1 PIX3990_IN
port 4049 n
rlabel metal5 107020 -72980 107120 -72880 1 PIX3991_IN
port 4050 n
rlabel metal5 108520 -72980 108620 -72880 1 PIX3992_IN
port 4051 n
rlabel metal5 110020 -72980 110120 -72880 1 PIX3993_IN
port 4052 n
rlabel metal5 111520 -72980 111620 -72880 1 PIX3994_IN
port 4053 n
rlabel metal5 113020 -72980 113120 -72880 1 PIX3995_IN
port 4054 n
rlabel metal5 114520 -72980 114620 -72880 1 PIX3996_IN
port 4055 n
rlabel metal5 116020 -72980 116120 -72880 1 PIX3997_IN
port 4056 n
rlabel metal5 117520 -72980 117620 -72880 1 PIX3998_IN
port 4057 n
rlabel metal5 119020 -72980 119120 -72880 1 PIX3999_IN
port 4058 n
rlabel metal5 520 -74480 620 -74380 1 PIX4000_IN
port 4059 n
rlabel metal2 -1500 -74260 -1500 -74215 3 ROW_SEL50
port 4060 e
rlabel metal5 2020 -74480 2120 -74380 1 PIX4001_IN
port 4061 n
rlabel metal5 3520 -74480 3620 -74380 1 PIX4002_IN
port 4062 n
rlabel metal5 5020 -74480 5120 -74380 1 PIX4003_IN
port 4063 n
rlabel metal5 6520 -74480 6620 -74380 1 PIX4004_IN
port 4064 n
rlabel metal5 8020 -74480 8120 -74380 1 PIX4005_IN
port 4065 n
rlabel metal5 9520 -74480 9620 -74380 1 PIX4006_IN
port 4066 n
rlabel metal5 11020 -74480 11120 -74380 1 PIX4007_IN
port 4067 n
rlabel metal5 12520 -74480 12620 -74380 1 PIX4008_IN
port 4068 n
rlabel metal5 14020 -74480 14120 -74380 1 PIX4009_IN
port 4069 n
rlabel metal5 15520 -74480 15620 -74380 1 PIX4010_IN
port 4070 n
rlabel metal5 17020 -74480 17120 -74380 1 PIX4011_IN
port 4071 n
rlabel metal5 18520 -74480 18620 -74380 1 PIX4012_IN
port 4072 n
rlabel metal5 20020 -74480 20120 -74380 1 PIX4013_IN
port 4073 n
rlabel metal5 21520 -74480 21620 -74380 1 PIX4014_IN
port 4074 n
rlabel metal5 23020 -74480 23120 -74380 1 PIX4015_IN
port 4075 n
rlabel metal5 24520 -74480 24620 -74380 1 PIX4016_IN
port 4076 n
rlabel metal5 26020 -74480 26120 -74380 1 PIX4017_IN
port 4077 n
rlabel metal5 27520 -74480 27620 -74380 1 PIX4018_IN
port 4078 n
rlabel metal5 29020 -74480 29120 -74380 1 PIX4019_IN
port 4079 n
rlabel metal5 30520 -74480 30620 -74380 1 PIX4020_IN
port 4080 n
rlabel metal5 32020 -74480 32120 -74380 1 PIX4021_IN
port 4081 n
rlabel metal5 33520 -74480 33620 -74380 1 PIX4022_IN
port 4082 n
rlabel metal5 35020 -74480 35120 -74380 1 PIX4023_IN
port 4083 n
rlabel metal5 36520 -74480 36620 -74380 1 PIX4024_IN
port 4084 n
rlabel metal5 38020 -74480 38120 -74380 1 PIX4025_IN
port 4085 n
rlabel metal5 39520 -74480 39620 -74380 1 PIX4026_IN
port 4086 n
rlabel metal5 41020 -74480 41120 -74380 1 PIX4027_IN
port 4087 n
rlabel metal5 42520 -74480 42620 -74380 1 PIX4028_IN
port 4088 n
rlabel metal5 44020 -74480 44120 -74380 1 PIX4029_IN
port 4089 n
rlabel metal5 45520 -74480 45620 -74380 1 PIX4030_IN
port 4090 n
rlabel metal5 47020 -74480 47120 -74380 1 PIX4031_IN
port 4091 n
rlabel metal5 48520 -74480 48620 -74380 1 PIX4032_IN
port 4092 n
rlabel metal5 50020 -74480 50120 -74380 1 PIX4033_IN
port 4093 n
rlabel metal5 51520 -74480 51620 -74380 1 PIX4034_IN
port 4094 n
rlabel metal5 53020 -74480 53120 -74380 1 PIX4035_IN
port 4095 n
rlabel metal5 54520 -74480 54620 -74380 1 PIX4036_IN
port 4096 n
rlabel metal5 56020 -74480 56120 -74380 1 PIX4037_IN
port 4097 n
rlabel metal5 57520 -74480 57620 -74380 1 PIX4038_IN
port 4098 n
rlabel metal5 59020 -74480 59120 -74380 1 PIX4039_IN
port 4099 n
rlabel metal5 60520 -74480 60620 -74380 1 PIX4040_IN
port 4100 n
rlabel metal5 62020 -74480 62120 -74380 1 PIX4041_IN
port 4101 n
rlabel metal5 63520 -74480 63620 -74380 1 PIX4042_IN
port 4102 n
rlabel metal5 65020 -74480 65120 -74380 1 PIX4043_IN
port 4103 n
rlabel metal5 66520 -74480 66620 -74380 1 PIX4044_IN
port 4104 n
rlabel metal5 68020 -74480 68120 -74380 1 PIX4045_IN
port 4105 n
rlabel metal5 69520 -74480 69620 -74380 1 PIX4046_IN
port 4106 n
rlabel metal5 71020 -74480 71120 -74380 1 PIX4047_IN
port 4107 n
rlabel metal5 72520 -74480 72620 -74380 1 PIX4048_IN
port 4108 n
rlabel metal5 74020 -74480 74120 -74380 1 PIX4049_IN
port 4109 n
rlabel metal5 75520 -74480 75620 -74380 1 PIX4050_IN
port 4110 n
rlabel metal5 77020 -74480 77120 -74380 1 PIX4051_IN
port 4111 n
rlabel metal5 78520 -74480 78620 -74380 1 PIX4052_IN
port 4112 n
rlabel metal5 80020 -74480 80120 -74380 1 PIX4053_IN
port 4113 n
rlabel metal5 81520 -74480 81620 -74380 1 PIX4054_IN
port 4114 n
rlabel metal5 83020 -74480 83120 -74380 1 PIX4055_IN
port 4115 n
rlabel metal5 84520 -74480 84620 -74380 1 PIX4056_IN
port 4116 n
rlabel metal5 86020 -74480 86120 -74380 1 PIX4057_IN
port 4117 n
rlabel metal5 87520 -74480 87620 -74380 1 PIX4058_IN
port 4118 n
rlabel metal5 89020 -74480 89120 -74380 1 PIX4059_IN
port 4119 n
rlabel metal5 90520 -74480 90620 -74380 1 PIX4060_IN
port 4120 n
rlabel metal5 92020 -74480 92120 -74380 1 PIX4061_IN
port 4121 n
rlabel metal5 93520 -74480 93620 -74380 1 PIX4062_IN
port 4122 n
rlabel metal5 95020 -74480 95120 -74380 1 PIX4063_IN
port 4123 n
rlabel metal5 96520 -74480 96620 -74380 1 PIX4064_IN
port 4124 n
rlabel metal5 98020 -74480 98120 -74380 1 PIX4065_IN
port 4125 n
rlabel metal5 99520 -74480 99620 -74380 1 PIX4066_IN
port 4126 n
rlabel metal5 101020 -74480 101120 -74380 1 PIX4067_IN
port 4127 n
rlabel metal5 102520 -74480 102620 -74380 1 PIX4068_IN
port 4128 n
rlabel metal5 104020 -74480 104120 -74380 1 PIX4069_IN
port 4129 n
rlabel metal5 105520 -74480 105620 -74380 1 PIX4070_IN
port 4130 n
rlabel metal5 107020 -74480 107120 -74380 1 PIX4071_IN
port 4131 n
rlabel metal5 108520 -74480 108620 -74380 1 PIX4072_IN
port 4132 n
rlabel metal5 110020 -74480 110120 -74380 1 PIX4073_IN
port 4133 n
rlabel metal5 111520 -74480 111620 -74380 1 PIX4074_IN
port 4134 n
rlabel metal5 113020 -74480 113120 -74380 1 PIX4075_IN
port 4135 n
rlabel metal5 114520 -74480 114620 -74380 1 PIX4076_IN
port 4136 n
rlabel metal5 116020 -74480 116120 -74380 1 PIX4077_IN
port 4137 n
rlabel metal5 117520 -74480 117620 -74380 1 PIX4078_IN
port 4138 n
rlabel metal5 119020 -74480 119120 -74380 1 PIX4079_IN
port 4139 n
rlabel metal5 520 -75980 620 -75880 1 PIX4080_IN
port 4140 n
rlabel metal2 -1500 -75760 -1500 -75715 3 ROW_SEL51
port 4141 e
rlabel metal5 2020 -75980 2120 -75880 1 PIX4081_IN
port 4142 n
rlabel metal5 3520 -75980 3620 -75880 1 PIX4082_IN
port 4143 n
rlabel metal5 5020 -75980 5120 -75880 1 PIX4083_IN
port 4144 n
rlabel metal5 6520 -75980 6620 -75880 1 PIX4084_IN
port 4145 n
rlabel metal5 8020 -75980 8120 -75880 1 PIX4085_IN
port 4146 n
rlabel metal5 9520 -75980 9620 -75880 1 PIX4086_IN
port 4147 n
rlabel metal5 11020 -75980 11120 -75880 1 PIX4087_IN
port 4148 n
rlabel metal5 12520 -75980 12620 -75880 1 PIX4088_IN
port 4149 n
rlabel metal5 14020 -75980 14120 -75880 1 PIX4089_IN
port 4150 n
rlabel metal5 15520 -75980 15620 -75880 1 PIX4090_IN
port 4151 n
rlabel metal5 17020 -75980 17120 -75880 1 PIX4091_IN
port 4152 n
rlabel metal5 18520 -75980 18620 -75880 1 PIX4092_IN
port 4153 n
rlabel metal5 20020 -75980 20120 -75880 1 PIX4093_IN
port 4154 n
rlabel metal5 21520 -75980 21620 -75880 1 PIX4094_IN
port 4155 n
rlabel metal5 23020 -75980 23120 -75880 1 PIX4095_IN
port 4156 n
rlabel metal5 24520 -75980 24620 -75880 1 PIX4096_IN
port 4157 n
rlabel metal5 26020 -75980 26120 -75880 1 PIX4097_IN
port 4158 n
rlabel metal5 27520 -75980 27620 -75880 1 PIX4098_IN
port 4159 n
rlabel metal5 29020 -75980 29120 -75880 1 PIX4099_IN
port 4160 n
rlabel metal5 30520 -75980 30620 -75880 1 PIX4100_IN
port 4161 n
rlabel metal5 32020 -75980 32120 -75880 1 PIX4101_IN
port 4162 n
rlabel metal5 33520 -75980 33620 -75880 1 PIX4102_IN
port 4163 n
rlabel metal5 35020 -75980 35120 -75880 1 PIX4103_IN
port 4164 n
rlabel metal5 36520 -75980 36620 -75880 1 PIX4104_IN
port 4165 n
rlabel metal5 38020 -75980 38120 -75880 1 PIX4105_IN
port 4166 n
rlabel metal5 39520 -75980 39620 -75880 1 PIX4106_IN
port 4167 n
rlabel metal5 41020 -75980 41120 -75880 1 PIX4107_IN
port 4168 n
rlabel metal5 42520 -75980 42620 -75880 1 PIX4108_IN
port 4169 n
rlabel metal5 44020 -75980 44120 -75880 1 PIX4109_IN
port 4170 n
rlabel metal5 45520 -75980 45620 -75880 1 PIX4110_IN
port 4171 n
rlabel metal5 47020 -75980 47120 -75880 1 PIX4111_IN
port 4172 n
rlabel metal5 48520 -75980 48620 -75880 1 PIX4112_IN
port 4173 n
rlabel metal5 50020 -75980 50120 -75880 1 PIX4113_IN
port 4174 n
rlabel metal5 51520 -75980 51620 -75880 1 PIX4114_IN
port 4175 n
rlabel metal5 53020 -75980 53120 -75880 1 PIX4115_IN
port 4176 n
rlabel metal5 54520 -75980 54620 -75880 1 PIX4116_IN
port 4177 n
rlabel metal5 56020 -75980 56120 -75880 1 PIX4117_IN
port 4178 n
rlabel metal5 57520 -75980 57620 -75880 1 PIX4118_IN
port 4179 n
rlabel metal5 59020 -75980 59120 -75880 1 PIX4119_IN
port 4180 n
rlabel metal5 60520 -75980 60620 -75880 1 PIX4120_IN
port 4181 n
rlabel metal5 62020 -75980 62120 -75880 1 PIX4121_IN
port 4182 n
rlabel metal5 63520 -75980 63620 -75880 1 PIX4122_IN
port 4183 n
rlabel metal5 65020 -75980 65120 -75880 1 PIX4123_IN
port 4184 n
rlabel metal5 66520 -75980 66620 -75880 1 PIX4124_IN
port 4185 n
rlabel metal5 68020 -75980 68120 -75880 1 PIX4125_IN
port 4186 n
rlabel metal5 69520 -75980 69620 -75880 1 PIX4126_IN
port 4187 n
rlabel metal5 71020 -75980 71120 -75880 1 PIX4127_IN
port 4188 n
rlabel metal5 72520 -75980 72620 -75880 1 PIX4128_IN
port 4189 n
rlabel metal5 74020 -75980 74120 -75880 1 PIX4129_IN
port 4190 n
rlabel metal5 75520 -75980 75620 -75880 1 PIX4130_IN
port 4191 n
rlabel metal5 77020 -75980 77120 -75880 1 PIX4131_IN
port 4192 n
rlabel metal5 78520 -75980 78620 -75880 1 PIX4132_IN
port 4193 n
rlabel metal5 80020 -75980 80120 -75880 1 PIX4133_IN
port 4194 n
rlabel metal5 81520 -75980 81620 -75880 1 PIX4134_IN
port 4195 n
rlabel metal5 83020 -75980 83120 -75880 1 PIX4135_IN
port 4196 n
rlabel metal5 84520 -75980 84620 -75880 1 PIX4136_IN
port 4197 n
rlabel metal5 86020 -75980 86120 -75880 1 PIX4137_IN
port 4198 n
rlabel metal5 87520 -75980 87620 -75880 1 PIX4138_IN
port 4199 n
rlabel metal5 89020 -75980 89120 -75880 1 PIX4139_IN
port 4200 n
rlabel metal5 90520 -75980 90620 -75880 1 PIX4140_IN
port 4201 n
rlabel metal5 92020 -75980 92120 -75880 1 PIX4141_IN
port 4202 n
rlabel metal5 93520 -75980 93620 -75880 1 PIX4142_IN
port 4203 n
rlabel metal5 95020 -75980 95120 -75880 1 PIX4143_IN
port 4204 n
rlabel metal5 96520 -75980 96620 -75880 1 PIX4144_IN
port 4205 n
rlabel metal5 98020 -75980 98120 -75880 1 PIX4145_IN
port 4206 n
rlabel metal5 99520 -75980 99620 -75880 1 PIX4146_IN
port 4207 n
rlabel metal5 101020 -75980 101120 -75880 1 PIX4147_IN
port 4208 n
rlabel metal5 102520 -75980 102620 -75880 1 PIX4148_IN
port 4209 n
rlabel metal5 104020 -75980 104120 -75880 1 PIX4149_IN
port 4210 n
rlabel metal5 105520 -75980 105620 -75880 1 PIX4150_IN
port 4211 n
rlabel metal5 107020 -75980 107120 -75880 1 PIX4151_IN
port 4212 n
rlabel metal5 108520 -75980 108620 -75880 1 PIX4152_IN
port 4213 n
rlabel metal5 110020 -75980 110120 -75880 1 PIX4153_IN
port 4214 n
rlabel metal5 111520 -75980 111620 -75880 1 PIX4154_IN
port 4215 n
rlabel metal5 113020 -75980 113120 -75880 1 PIX4155_IN
port 4216 n
rlabel metal5 114520 -75980 114620 -75880 1 PIX4156_IN
port 4217 n
rlabel metal5 116020 -75980 116120 -75880 1 PIX4157_IN
port 4218 n
rlabel metal5 117520 -75980 117620 -75880 1 PIX4158_IN
port 4219 n
rlabel metal5 119020 -75980 119120 -75880 1 PIX4159_IN
port 4220 n
rlabel metal5 520 -77480 620 -77380 1 PIX4160_IN
port 4221 n
rlabel metal2 -1500 -77260 -1500 -77215 3 ROW_SEL52
port 4222 e
rlabel metal5 2020 -77480 2120 -77380 1 PIX4161_IN
port 4223 n
rlabel metal5 3520 -77480 3620 -77380 1 PIX4162_IN
port 4224 n
rlabel metal5 5020 -77480 5120 -77380 1 PIX4163_IN
port 4225 n
rlabel metal5 6520 -77480 6620 -77380 1 PIX4164_IN
port 4226 n
rlabel metal5 8020 -77480 8120 -77380 1 PIX4165_IN
port 4227 n
rlabel metal5 9520 -77480 9620 -77380 1 PIX4166_IN
port 4228 n
rlabel metal5 11020 -77480 11120 -77380 1 PIX4167_IN
port 4229 n
rlabel metal5 12520 -77480 12620 -77380 1 PIX4168_IN
port 4230 n
rlabel metal5 14020 -77480 14120 -77380 1 PIX4169_IN
port 4231 n
rlabel metal5 15520 -77480 15620 -77380 1 PIX4170_IN
port 4232 n
rlabel metal5 17020 -77480 17120 -77380 1 PIX4171_IN
port 4233 n
rlabel metal5 18520 -77480 18620 -77380 1 PIX4172_IN
port 4234 n
rlabel metal5 20020 -77480 20120 -77380 1 PIX4173_IN
port 4235 n
rlabel metal5 21520 -77480 21620 -77380 1 PIX4174_IN
port 4236 n
rlabel metal5 23020 -77480 23120 -77380 1 PIX4175_IN
port 4237 n
rlabel metal5 24520 -77480 24620 -77380 1 PIX4176_IN
port 4238 n
rlabel metal5 26020 -77480 26120 -77380 1 PIX4177_IN
port 4239 n
rlabel metal5 27520 -77480 27620 -77380 1 PIX4178_IN
port 4240 n
rlabel metal5 29020 -77480 29120 -77380 1 PIX4179_IN
port 4241 n
rlabel metal5 30520 -77480 30620 -77380 1 PIX4180_IN
port 4242 n
rlabel metal5 32020 -77480 32120 -77380 1 PIX4181_IN
port 4243 n
rlabel metal5 33520 -77480 33620 -77380 1 PIX4182_IN
port 4244 n
rlabel metal5 35020 -77480 35120 -77380 1 PIX4183_IN
port 4245 n
rlabel metal5 36520 -77480 36620 -77380 1 PIX4184_IN
port 4246 n
rlabel metal5 38020 -77480 38120 -77380 1 PIX4185_IN
port 4247 n
rlabel metal5 39520 -77480 39620 -77380 1 PIX4186_IN
port 4248 n
rlabel metal5 41020 -77480 41120 -77380 1 PIX4187_IN
port 4249 n
rlabel metal5 42520 -77480 42620 -77380 1 PIX4188_IN
port 4250 n
rlabel metal5 44020 -77480 44120 -77380 1 PIX4189_IN
port 4251 n
rlabel metal5 45520 -77480 45620 -77380 1 PIX4190_IN
port 4252 n
rlabel metal5 47020 -77480 47120 -77380 1 PIX4191_IN
port 4253 n
rlabel metal5 48520 -77480 48620 -77380 1 PIX4192_IN
port 4254 n
rlabel metal5 50020 -77480 50120 -77380 1 PIX4193_IN
port 4255 n
rlabel metal5 51520 -77480 51620 -77380 1 PIX4194_IN
port 4256 n
rlabel metal5 53020 -77480 53120 -77380 1 PIX4195_IN
port 4257 n
rlabel metal5 54520 -77480 54620 -77380 1 PIX4196_IN
port 4258 n
rlabel metal5 56020 -77480 56120 -77380 1 PIX4197_IN
port 4259 n
rlabel metal5 57520 -77480 57620 -77380 1 PIX4198_IN
port 4260 n
rlabel metal5 59020 -77480 59120 -77380 1 PIX4199_IN
port 4261 n
rlabel metal5 60520 -77480 60620 -77380 1 PIX4200_IN
port 4262 n
rlabel metal5 62020 -77480 62120 -77380 1 PIX4201_IN
port 4263 n
rlabel metal5 63520 -77480 63620 -77380 1 PIX4202_IN
port 4264 n
rlabel metal5 65020 -77480 65120 -77380 1 PIX4203_IN
port 4265 n
rlabel metal5 66520 -77480 66620 -77380 1 PIX4204_IN
port 4266 n
rlabel metal5 68020 -77480 68120 -77380 1 PIX4205_IN
port 4267 n
rlabel metal5 69520 -77480 69620 -77380 1 PIX4206_IN
port 4268 n
rlabel metal5 71020 -77480 71120 -77380 1 PIX4207_IN
port 4269 n
rlabel metal5 72520 -77480 72620 -77380 1 PIX4208_IN
port 4270 n
rlabel metal5 74020 -77480 74120 -77380 1 PIX4209_IN
port 4271 n
rlabel metal5 75520 -77480 75620 -77380 1 PIX4210_IN
port 4272 n
rlabel metal5 77020 -77480 77120 -77380 1 PIX4211_IN
port 4273 n
rlabel metal5 78520 -77480 78620 -77380 1 PIX4212_IN
port 4274 n
rlabel metal5 80020 -77480 80120 -77380 1 PIX4213_IN
port 4275 n
rlabel metal5 81520 -77480 81620 -77380 1 PIX4214_IN
port 4276 n
rlabel metal5 83020 -77480 83120 -77380 1 PIX4215_IN
port 4277 n
rlabel metal5 84520 -77480 84620 -77380 1 PIX4216_IN
port 4278 n
rlabel metal5 86020 -77480 86120 -77380 1 PIX4217_IN
port 4279 n
rlabel metal5 87520 -77480 87620 -77380 1 PIX4218_IN
port 4280 n
rlabel metal5 89020 -77480 89120 -77380 1 PIX4219_IN
port 4281 n
rlabel metal5 90520 -77480 90620 -77380 1 PIX4220_IN
port 4282 n
rlabel metal5 92020 -77480 92120 -77380 1 PIX4221_IN
port 4283 n
rlabel metal5 93520 -77480 93620 -77380 1 PIX4222_IN
port 4284 n
rlabel metal5 95020 -77480 95120 -77380 1 PIX4223_IN
port 4285 n
rlabel metal5 96520 -77480 96620 -77380 1 PIX4224_IN
port 4286 n
rlabel metal5 98020 -77480 98120 -77380 1 PIX4225_IN
port 4287 n
rlabel metal5 99520 -77480 99620 -77380 1 PIX4226_IN
port 4288 n
rlabel metal5 101020 -77480 101120 -77380 1 PIX4227_IN
port 4289 n
rlabel metal5 102520 -77480 102620 -77380 1 PIX4228_IN
port 4290 n
rlabel metal5 104020 -77480 104120 -77380 1 PIX4229_IN
port 4291 n
rlabel metal5 105520 -77480 105620 -77380 1 PIX4230_IN
port 4292 n
rlabel metal5 107020 -77480 107120 -77380 1 PIX4231_IN
port 4293 n
rlabel metal5 108520 -77480 108620 -77380 1 PIX4232_IN
port 4294 n
rlabel metal5 110020 -77480 110120 -77380 1 PIX4233_IN
port 4295 n
rlabel metal5 111520 -77480 111620 -77380 1 PIX4234_IN
port 4296 n
rlabel metal5 113020 -77480 113120 -77380 1 PIX4235_IN
port 4297 n
rlabel metal5 114520 -77480 114620 -77380 1 PIX4236_IN
port 4298 n
rlabel metal5 116020 -77480 116120 -77380 1 PIX4237_IN
port 4299 n
rlabel metal5 117520 -77480 117620 -77380 1 PIX4238_IN
port 4300 n
rlabel metal5 119020 -77480 119120 -77380 1 PIX4239_IN
port 4301 n
rlabel metal5 520 -78980 620 -78880 1 PIX4240_IN
port 4302 n
rlabel metal2 -1500 -78760 -1500 -78715 3 ROW_SEL53
port 4303 e
rlabel metal5 2020 -78980 2120 -78880 1 PIX4241_IN
port 4304 n
rlabel metal5 3520 -78980 3620 -78880 1 PIX4242_IN
port 4305 n
rlabel metal5 5020 -78980 5120 -78880 1 PIX4243_IN
port 4306 n
rlabel metal5 6520 -78980 6620 -78880 1 PIX4244_IN
port 4307 n
rlabel metal5 8020 -78980 8120 -78880 1 PIX4245_IN
port 4308 n
rlabel metal5 9520 -78980 9620 -78880 1 PIX4246_IN
port 4309 n
rlabel metal5 11020 -78980 11120 -78880 1 PIX4247_IN
port 4310 n
rlabel metal5 12520 -78980 12620 -78880 1 PIX4248_IN
port 4311 n
rlabel metal5 14020 -78980 14120 -78880 1 PIX4249_IN
port 4312 n
rlabel metal5 15520 -78980 15620 -78880 1 PIX4250_IN
port 4313 n
rlabel metal5 17020 -78980 17120 -78880 1 PIX4251_IN
port 4314 n
rlabel metal5 18520 -78980 18620 -78880 1 PIX4252_IN
port 4315 n
rlabel metal5 20020 -78980 20120 -78880 1 PIX4253_IN
port 4316 n
rlabel metal5 21520 -78980 21620 -78880 1 PIX4254_IN
port 4317 n
rlabel metal5 23020 -78980 23120 -78880 1 PIX4255_IN
port 4318 n
rlabel metal5 24520 -78980 24620 -78880 1 PIX4256_IN
port 4319 n
rlabel metal5 26020 -78980 26120 -78880 1 PIX4257_IN
port 4320 n
rlabel metal5 27520 -78980 27620 -78880 1 PIX4258_IN
port 4321 n
rlabel metal5 29020 -78980 29120 -78880 1 PIX4259_IN
port 4322 n
rlabel metal5 30520 -78980 30620 -78880 1 PIX4260_IN
port 4323 n
rlabel metal5 32020 -78980 32120 -78880 1 PIX4261_IN
port 4324 n
rlabel metal5 33520 -78980 33620 -78880 1 PIX4262_IN
port 4325 n
rlabel metal5 35020 -78980 35120 -78880 1 PIX4263_IN
port 4326 n
rlabel metal5 36520 -78980 36620 -78880 1 PIX4264_IN
port 4327 n
rlabel metal5 38020 -78980 38120 -78880 1 PIX4265_IN
port 4328 n
rlabel metal5 39520 -78980 39620 -78880 1 PIX4266_IN
port 4329 n
rlabel metal5 41020 -78980 41120 -78880 1 PIX4267_IN
port 4330 n
rlabel metal5 42520 -78980 42620 -78880 1 PIX4268_IN
port 4331 n
rlabel metal5 44020 -78980 44120 -78880 1 PIX4269_IN
port 4332 n
rlabel metal5 45520 -78980 45620 -78880 1 PIX4270_IN
port 4333 n
rlabel metal5 47020 -78980 47120 -78880 1 PIX4271_IN
port 4334 n
rlabel metal5 48520 -78980 48620 -78880 1 PIX4272_IN
port 4335 n
rlabel metal5 50020 -78980 50120 -78880 1 PIX4273_IN
port 4336 n
rlabel metal5 51520 -78980 51620 -78880 1 PIX4274_IN
port 4337 n
rlabel metal5 53020 -78980 53120 -78880 1 PIX4275_IN
port 4338 n
rlabel metal5 54520 -78980 54620 -78880 1 PIX4276_IN
port 4339 n
rlabel metal5 56020 -78980 56120 -78880 1 PIX4277_IN
port 4340 n
rlabel metal5 57520 -78980 57620 -78880 1 PIX4278_IN
port 4341 n
rlabel metal5 59020 -78980 59120 -78880 1 PIX4279_IN
port 4342 n
rlabel metal5 60520 -78980 60620 -78880 1 PIX4280_IN
port 4343 n
rlabel metal5 62020 -78980 62120 -78880 1 PIX4281_IN
port 4344 n
rlabel metal5 63520 -78980 63620 -78880 1 PIX4282_IN
port 4345 n
rlabel metal5 65020 -78980 65120 -78880 1 PIX4283_IN
port 4346 n
rlabel metal5 66520 -78980 66620 -78880 1 PIX4284_IN
port 4347 n
rlabel metal5 68020 -78980 68120 -78880 1 PIX4285_IN
port 4348 n
rlabel metal5 69520 -78980 69620 -78880 1 PIX4286_IN
port 4349 n
rlabel metal5 71020 -78980 71120 -78880 1 PIX4287_IN
port 4350 n
rlabel metal5 72520 -78980 72620 -78880 1 PIX4288_IN
port 4351 n
rlabel metal5 74020 -78980 74120 -78880 1 PIX4289_IN
port 4352 n
rlabel metal5 75520 -78980 75620 -78880 1 PIX4290_IN
port 4353 n
rlabel metal5 77020 -78980 77120 -78880 1 PIX4291_IN
port 4354 n
rlabel metal5 78520 -78980 78620 -78880 1 PIX4292_IN
port 4355 n
rlabel metal5 80020 -78980 80120 -78880 1 PIX4293_IN
port 4356 n
rlabel metal5 81520 -78980 81620 -78880 1 PIX4294_IN
port 4357 n
rlabel metal5 83020 -78980 83120 -78880 1 PIX4295_IN
port 4358 n
rlabel metal5 84520 -78980 84620 -78880 1 PIX4296_IN
port 4359 n
rlabel metal5 86020 -78980 86120 -78880 1 PIX4297_IN
port 4360 n
rlabel metal5 87520 -78980 87620 -78880 1 PIX4298_IN
port 4361 n
rlabel metal5 89020 -78980 89120 -78880 1 PIX4299_IN
port 4362 n
rlabel metal5 90520 -78980 90620 -78880 1 PIX4300_IN
port 4363 n
rlabel metal5 92020 -78980 92120 -78880 1 PIX4301_IN
port 4364 n
rlabel metal5 93520 -78980 93620 -78880 1 PIX4302_IN
port 4365 n
rlabel metal5 95020 -78980 95120 -78880 1 PIX4303_IN
port 4366 n
rlabel metal5 96520 -78980 96620 -78880 1 PIX4304_IN
port 4367 n
rlabel metal5 98020 -78980 98120 -78880 1 PIX4305_IN
port 4368 n
rlabel metal5 99520 -78980 99620 -78880 1 PIX4306_IN
port 4369 n
rlabel metal5 101020 -78980 101120 -78880 1 PIX4307_IN
port 4370 n
rlabel metal5 102520 -78980 102620 -78880 1 PIX4308_IN
port 4371 n
rlabel metal5 104020 -78980 104120 -78880 1 PIX4309_IN
port 4372 n
rlabel metal5 105520 -78980 105620 -78880 1 PIX4310_IN
port 4373 n
rlabel metal5 107020 -78980 107120 -78880 1 PIX4311_IN
port 4374 n
rlabel metal5 108520 -78980 108620 -78880 1 PIX4312_IN
port 4375 n
rlabel metal5 110020 -78980 110120 -78880 1 PIX4313_IN
port 4376 n
rlabel metal5 111520 -78980 111620 -78880 1 PIX4314_IN
port 4377 n
rlabel metal5 113020 -78980 113120 -78880 1 PIX4315_IN
port 4378 n
rlabel metal5 114520 -78980 114620 -78880 1 PIX4316_IN
port 4379 n
rlabel metal5 116020 -78980 116120 -78880 1 PIX4317_IN
port 4380 n
rlabel metal5 117520 -78980 117620 -78880 1 PIX4318_IN
port 4381 n
rlabel metal5 119020 -78980 119120 -78880 1 PIX4319_IN
port 4382 n
rlabel metal5 520 -80480 620 -80380 1 PIX4320_IN
port 4383 n
rlabel metal2 -1500 -80260 -1500 -80215 3 ROW_SEL54
port 4384 e
rlabel metal5 2020 -80480 2120 -80380 1 PIX4321_IN
port 4385 n
rlabel metal5 3520 -80480 3620 -80380 1 PIX4322_IN
port 4386 n
rlabel metal5 5020 -80480 5120 -80380 1 PIX4323_IN
port 4387 n
rlabel metal5 6520 -80480 6620 -80380 1 PIX4324_IN
port 4388 n
rlabel metal5 8020 -80480 8120 -80380 1 PIX4325_IN
port 4389 n
rlabel metal5 9520 -80480 9620 -80380 1 PIX4326_IN
port 4390 n
rlabel metal5 11020 -80480 11120 -80380 1 PIX4327_IN
port 4391 n
rlabel metal5 12520 -80480 12620 -80380 1 PIX4328_IN
port 4392 n
rlabel metal5 14020 -80480 14120 -80380 1 PIX4329_IN
port 4393 n
rlabel metal5 15520 -80480 15620 -80380 1 PIX4330_IN
port 4394 n
rlabel metal5 17020 -80480 17120 -80380 1 PIX4331_IN
port 4395 n
rlabel metal5 18520 -80480 18620 -80380 1 PIX4332_IN
port 4396 n
rlabel metal5 20020 -80480 20120 -80380 1 PIX4333_IN
port 4397 n
rlabel metal5 21520 -80480 21620 -80380 1 PIX4334_IN
port 4398 n
rlabel metal5 23020 -80480 23120 -80380 1 PIX4335_IN
port 4399 n
rlabel metal5 24520 -80480 24620 -80380 1 PIX4336_IN
port 4400 n
rlabel metal5 26020 -80480 26120 -80380 1 PIX4337_IN
port 4401 n
rlabel metal5 27520 -80480 27620 -80380 1 PIX4338_IN
port 4402 n
rlabel metal5 29020 -80480 29120 -80380 1 PIX4339_IN
port 4403 n
rlabel metal5 30520 -80480 30620 -80380 1 PIX4340_IN
port 4404 n
rlabel metal5 32020 -80480 32120 -80380 1 PIX4341_IN
port 4405 n
rlabel metal5 33520 -80480 33620 -80380 1 PIX4342_IN
port 4406 n
rlabel metal5 35020 -80480 35120 -80380 1 PIX4343_IN
port 4407 n
rlabel metal5 36520 -80480 36620 -80380 1 PIX4344_IN
port 4408 n
rlabel metal5 38020 -80480 38120 -80380 1 PIX4345_IN
port 4409 n
rlabel metal5 39520 -80480 39620 -80380 1 PIX4346_IN
port 4410 n
rlabel metal5 41020 -80480 41120 -80380 1 PIX4347_IN
port 4411 n
rlabel metal5 42520 -80480 42620 -80380 1 PIX4348_IN
port 4412 n
rlabel metal5 44020 -80480 44120 -80380 1 PIX4349_IN
port 4413 n
rlabel metal5 45520 -80480 45620 -80380 1 PIX4350_IN
port 4414 n
rlabel metal5 47020 -80480 47120 -80380 1 PIX4351_IN
port 4415 n
rlabel metal5 48520 -80480 48620 -80380 1 PIX4352_IN
port 4416 n
rlabel metal5 50020 -80480 50120 -80380 1 PIX4353_IN
port 4417 n
rlabel metal5 51520 -80480 51620 -80380 1 PIX4354_IN
port 4418 n
rlabel metal5 53020 -80480 53120 -80380 1 PIX4355_IN
port 4419 n
rlabel metal5 54520 -80480 54620 -80380 1 PIX4356_IN
port 4420 n
rlabel metal5 56020 -80480 56120 -80380 1 PIX4357_IN
port 4421 n
rlabel metal5 57520 -80480 57620 -80380 1 PIX4358_IN
port 4422 n
rlabel metal5 59020 -80480 59120 -80380 1 PIX4359_IN
port 4423 n
rlabel metal5 60520 -80480 60620 -80380 1 PIX4360_IN
port 4424 n
rlabel metal5 62020 -80480 62120 -80380 1 PIX4361_IN
port 4425 n
rlabel metal5 63520 -80480 63620 -80380 1 PIX4362_IN
port 4426 n
rlabel metal5 65020 -80480 65120 -80380 1 PIX4363_IN
port 4427 n
rlabel metal5 66520 -80480 66620 -80380 1 PIX4364_IN
port 4428 n
rlabel metal5 68020 -80480 68120 -80380 1 PIX4365_IN
port 4429 n
rlabel metal5 69520 -80480 69620 -80380 1 PIX4366_IN
port 4430 n
rlabel metal5 71020 -80480 71120 -80380 1 PIX4367_IN
port 4431 n
rlabel metal5 72520 -80480 72620 -80380 1 PIX4368_IN
port 4432 n
rlabel metal5 74020 -80480 74120 -80380 1 PIX4369_IN
port 4433 n
rlabel metal5 75520 -80480 75620 -80380 1 PIX4370_IN
port 4434 n
rlabel metal5 77020 -80480 77120 -80380 1 PIX4371_IN
port 4435 n
rlabel metal5 78520 -80480 78620 -80380 1 PIX4372_IN
port 4436 n
rlabel metal5 80020 -80480 80120 -80380 1 PIX4373_IN
port 4437 n
rlabel metal5 81520 -80480 81620 -80380 1 PIX4374_IN
port 4438 n
rlabel metal5 83020 -80480 83120 -80380 1 PIX4375_IN
port 4439 n
rlabel metal5 84520 -80480 84620 -80380 1 PIX4376_IN
port 4440 n
rlabel metal5 86020 -80480 86120 -80380 1 PIX4377_IN
port 4441 n
rlabel metal5 87520 -80480 87620 -80380 1 PIX4378_IN
port 4442 n
rlabel metal5 89020 -80480 89120 -80380 1 PIX4379_IN
port 4443 n
rlabel metal5 90520 -80480 90620 -80380 1 PIX4380_IN
port 4444 n
rlabel metal5 92020 -80480 92120 -80380 1 PIX4381_IN
port 4445 n
rlabel metal5 93520 -80480 93620 -80380 1 PIX4382_IN
port 4446 n
rlabel metal5 95020 -80480 95120 -80380 1 PIX4383_IN
port 4447 n
rlabel metal5 96520 -80480 96620 -80380 1 PIX4384_IN
port 4448 n
rlabel metal5 98020 -80480 98120 -80380 1 PIX4385_IN
port 4449 n
rlabel metal5 99520 -80480 99620 -80380 1 PIX4386_IN
port 4450 n
rlabel metal5 101020 -80480 101120 -80380 1 PIX4387_IN
port 4451 n
rlabel metal5 102520 -80480 102620 -80380 1 PIX4388_IN
port 4452 n
rlabel metal5 104020 -80480 104120 -80380 1 PIX4389_IN
port 4453 n
rlabel metal5 105520 -80480 105620 -80380 1 PIX4390_IN
port 4454 n
rlabel metal5 107020 -80480 107120 -80380 1 PIX4391_IN
port 4455 n
rlabel metal5 108520 -80480 108620 -80380 1 PIX4392_IN
port 4456 n
rlabel metal5 110020 -80480 110120 -80380 1 PIX4393_IN
port 4457 n
rlabel metal5 111520 -80480 111620 -80380 1 PIX4394_IN
port 4458 n
rlabel metal5 113020 -80480 113120 -80380 1 PIX4395_IN
port 4459 n
rlabel metal5 114520 -80480 114620 -80380 1 PIX4396_IN
port 4460 n
rlabel metal5 116020 -80480 116120 -80380 1 PIX4397_IN
port 4461 n
rlabel metal5 117520 -80480 117620 -80380 1 PIX4398_IN
port 4462 n
rlabel metal5 119020 -80480 119120 -80380 1 PIX4399_IN
port 4463 n
rlabel metal5 520 -81980 620 -81880 1 PIX4400_IN
port 4464 n
rlabel metal2 -1500 -81760 -1500 -81715 3 ROW_SEL55
port 4465 e
rlabel metal5 2020 -81980 2120 -81880 1 PIX4401_IN
port 4466 n
rlabel metal5 3520 -81980 3620 -81880 1 PIX4402_IN
port 4467 n
rlabel metal5 5020 -81980 5120 -81880 1 PIX4403_IN
port 4468 n
rlabel metal5 6520 -81980 6620 -81880 1 PIX4404_IN
port 4469 n
rlabel metal5 8020 -81980 8120 -81880 1 PIX4405_IN
port 4470 n
rlabel metal5 9520 -81980 9620 -81880 1 PIX4406_IN
port 4471 n
rlabel metal5 11020 -81980 11120 -81880 1 PIX4407_IN
port 4472 n
rlabel metal5 12520 -81980 12620 -81880 1 PIX4408_IN
port 4473 n
rlabel metal5 14020 -81980 14120 -81880 1 PIX4409_IN
port 4474 n
rlabel metal5 15520 -81980 15620 -81880 1 PIX4410_IN
port 4475 n
rlabel metal5 17020 -81980 17120 -81880 1 PIX4411_IN
port 4476 n
rlabel metal5 18520 -81980 18620 -81880 1 PIX4412_IN
port 4477 n
rlabel metal5 20020 -81980 20120 -81880 1 PIX4413_IN
port 4478 n
rlabel metal5 21520 -81980 21620 -81880 1 PIX4414_IN
port 4479 n
rlabel metal5 23020 -81980 23120 -81880 1 PIX4415_IN
port 4480 n
rlabel metal5 24520 -81980 24620 -81880 1 PIX4416_IN
port 4481 n
rlabel metal5 26020 -81980 26120 -81880 1 PIX4417_IN
port 4482 n
rlabel metal5 27520 -81980 27620 -81880 1 PIX4418_IN
port 4483 n
rlabel metal5 29020 -81980 29120 -81880 1 PIX4419_IN
port 4484 n
rlabel metal5 30520 -81980 30620 -81880 1 PIX4420_IN
port 4485 n
rlabel metal5 32020 -81980 32120 -81880 1 PIX4421_IN
port 4486 n
rlabel metal5 33520 -81980 33620 -81880 1 PIX4422_IN
port 4487 n
rlabel metal5 35020 -81980 35120 -81880 1 PIX4423_IN
port 4488 n
rlabel metal5 36520 -81980 36620 -81880 1 PIX4424_IN
port 4489 n
rlabel metal5 38020 -81980 38120 -81880 1 PIX4425_IN
port 4490 n
rlabel metal5 39520 -81980 39620 -81880 1 PIX4426_IN
port 4491 n
rlabel metal5 41020 -81980 41120 -81880 1 PIX4427_IN
port 4492 n
rlabel metal5 42520 -81980 42620 -81880 1 PIX4428_IN
port 4493 n
rlabel metal5 44020 -81980 44120 -81880 1 PIX4429_IN
port 4494 n
rlabel metal5 45520 -81980 45620 -81880 1 PIX4430_IN
port 4495 n
rlabel metal5 47020 -81980 47120 -81880 1 PIX4431_IN
port 4496 n
rlabel metal5 48520 -81980 48620 -81880 1 PIX4432_IN
port 4497 n
rlabel metal5 50020 -81980 50120 -81880 1 PIX4433_IN
port 4498 n
rlabel metal5 51520 -81980 51620 -81880 1 PIX4434_IN
port 4499 n
rlabel metal5 53020 -81980 53120 -81880 1 PIX4435_IN
port 4500 n
rlabel metal5 54520 -81980 54620 -81880 1 PIX4436_IN
port 4501 n
rlabel metal5 56020 -81980 56120 -81880 1 PIX4437_IN
port 4502 n
rlabel metal5 57520 -81980 57620 -81880 1 PIX4438_IN
port 4503 n
rlabel metal5 59020 -81980 59120 -81880 1 PIX4439_IN
port 4504 n
rlabel metal5 60520 -81980 60620 -81880 1 PIX4440_IN
port 4505 n
rlabel metal5 62020 -81980 62120 -81880 1 PIX4441_IN
port 4506 n
rlabel metal5 63520 -81980 63620 -81880 1 PIX4442_IN
port 4507 n
rlabel metal5 65020 -81980 65120 -81880 1 PIX4443_IN
port 4508 n
rlabel metal5 66520 -81980 66620 -81880 1 PIX4444_IN
port 4509 n
rlabel metal5 68020 -81980 68120 -81880 1 PIX4445_IN
port 4510 n
rlabel metal5 69520 -81980 69620 -81880 1 PIX4446_IN
port 4511 n
rlabel metal5 71020 -81980 71120 -81880 1 PIX4447_IN
port 4512 n
rlabel metal5 72520 -81980 72620 -81880 1 PIX4448_IN
port 4513 n
rlabel metal5 74020 -81980 74120 -81880 1 PIX4449_IN
port 4514 n
rlabel metal5 75520 -81980 75620 -81880 1 PIX4450_IN
port 4515 n
rlabel metal5 77020 -81980 77120 -81880 1 PIX4451_IN
port 4516 n
rlabel metal5 78520 -81980 78620 -81880 1 PIX4452_IN
port 4517 n
rlabel metal5 80020 -81980 80120 -81880 1 PIX4453_IN
port 4518 n
rlabel metal5 81520 -81980 81620 -81880 1 PIX4454_IN
port 4519 n
rlabel metal5 83020 -81980 83120 -81880 1 PIX4455_IN
port 4520 n
rlabel metal5 84520 -81980 84620 -81880 1 PIX4456_IN
port 4521 n
rlabel metal5 86020 -81980 86120 -81880 1 PIX4457_IN
port 4522 n
rlabel metal5 87520 -81980 87620 -81880 1 PIX4458_IN
port 4523 n
rlabel metal5 89020 -81980 89120 -81880 1 PIX4459_IN
port 4524 n
rlabel metal5 90520 -81980 90620 -81880 1 PIX4460_IN
port 4525 n
rlabel metal5 92020 -81980 92120 -81880 1 PIX4461_IN
port 4526 n
rlabel metal5 93520 -81980 93620 -81880 1 PIX4462_IN
port 4527 n
rlabel metal5 95020 -81980 95120 -81880 1 PIX4463_IN
port 4528 n
rlabel metal5 96520 -81980 96620 -81880 1 PIX4464_IN
port 4529 n
rlabel metal5 98020 -81980 98120 -81880 1 PIX4465_IN
port 4530 n
rlabel metal5 99520 -81980 99620 -81880 1 PIX4466_IN
port 4531 n
rlabel metal5 101020 -81980 101120 -81880 1 PIX4467_IN
port 4532 n
rlabel metal5 102520 -81980 102620 -81880 1 PIX4468_IN
port 4533 n
rlabel metal5 104020 -81980 104120 -81880 1 PIX4469_IN
port 4534 n
rlabel metal5 105520 -81980 105620 -81880 1 PIX4470_IN
port 4535 n
rlabel metal5 107020 -81980 107120 -81880 1 PIX4471_IN
port 4536 n
rlabel metal5 108520 -81980 108620 -81880 1 PIX4472_IN
port 4537 n
rlabel metal5 110020 -81980 110120 -81880 1 PIX4473_IN
port 4538 n
rlabel metal5 111520 -81980 111620 -81880 1 PIX4474_IN
port 4539 n
rlabel metal5 113020 -81980 113120 -81880 1 PIX4475_IN
port 4540 n
rlabel metal5 114520 -81980 114620 -81880 1 PIX4476_IN
port 4541 n
rlabel metal5 116020 -81980 116120 -81880 1 PIX4477_IN
port 4542 n
rlabel metal5 117520 -81980 117620 -81880 1 PIX4478_IN
port 4543 n
rlabel metal5 119020 -81980 119120 -81880 1 PIX4479_IN
port 4544 n
rlabel metal5 520 -83480 620 -83380 1 PIX4480_IN
port 4545 n
rlabel metal2 -1500 -83260 -1500 -83215 3 ROW_SEL56
port 4546 e
rlabel metal5 2020 -83480 2120 -83380 1 PIX4481_IN
port 4547 n
rlabel metal5 3520 -83480 3620 -83380 1 PIX4482_IN
port 4548 n
rlabel metal5 5020 -83480 5120 -83380 1 PIX4483_IN
port 4549 n
rlabel metal5 6520 -83480 6620 -83380 1 PIX4484_IN
port 4550 n
rlabel metal5 8020 -83480 8120 -83380 1 PIX4485_IN
port 4551 n
rlabel metal5 9520 -83480 9620 -83380 1 PIX4486_IN
port 4552 n
rlabel metal5 11020 -83480 11120 -83380 1 PIX4487_IN
port 4553 n
rlabel metal5 12520 -83480 12620 -83380 1 PIX4488_IN
port 4554 n
rlabel metal5 14020 -83480 14120 -83380 1 PIX4489_IN
port 4555 n
rlabel metal5 15520 -83480 15620 -83380 1 PIX4490_IN
port 4556 n
rlabel metal5 17020 -83480 17120 -83380 1 PIX4491_IN
port 4557 n
rlabel metal5 18520 -83480 18620 -83380 1 PIX4492_IN
port 4558 n
rlabel metal5 20020 -83480 20120 -83380 1 PIX4493_IN
port 4559 n
rlabel metal5 21520 -83480 21620 -83380 1 PIX4494_IN
port 4560 n
rlabel metal5 23020 -83480 23120 -83380 1 PIX4495_IN
port 4561 n
rlabel metal5 24520 -83480 24620 -83380 1 PIX4496_IN
port 4562 n
rlabel metal5 26020 -83480 26120 -83380 1 PIX4497_IN
port 4563 n
rlabel metal5 27520 -83480 27620 -83380 1 PIX4498_IN
port 4564 n
rlabel metal5 29020 -83480 29120 -83380 1 PIX4499_IN
port 4565 n
rlabel metal5 30520 -83480 30620 -83380 1 PIX4500_IN
port 4566 n
rlabel metal5 32020 -83480 32120 -83380 1 PIX4501_IN
port 4567 n
rlabel metal5 33520 -83480 33620 -83380 1 PIX4502_IN
port 4568 n
rlabel metal5 35020 -83480 35120 -83380 1 PIX4503_IN
port 4569 n
rlabel metal5 36520 -83480 36620 -83380 1 PIX4504_IN
port 4570 n
rlabel metal5 38020 -83480 38120 -83380 1 PIX4505_IN
port 4571 n
rlabel metal5 39520 -83480 39620 -83380 1 PIX4506_IN
port 4572 n
rlabel metal5 41020 -83480 41120 -83380 1 PIX4507_IN
port 4573 n
rlabel metal5 42520 -83480 42620 -83380 1 PIX4508_IN
port 4574 n
rlabel metal5 44020 -83480 44120 -83380 1 PIX4509_IN
port 4575 n
rlabel metal5 45520 -83480 45620 -83380 1 PIX4510_IN
port 4576 n
rlabel metal5 47020 -83480 47120 -83380 1 PIX4511_IN
port 4577 n
rlabel metal5 48520 -83480 48620 -83380 1 PIX4512_IN
port 4578 n
rlabel metal5 50020 -83480 50120 -83380 1 PIX4513_IN
port 4579 n
rlabel metal5 51520 -83480 51620 -83380 1 PIX4514_IN
port 4580 n
rlabel metal5 53020 -83480 53120 -83380 1 PIX4515_IN
port 4581 n
rlabel metal5 54520 -83480 54620 -83380 1 PIX4516_IN
port 4582 n
rlabel metal5 56020 -83480 56120 -83380 1 PIX4517_IN
port 4583 n
rlabel metal5 57520 -83480 57620 -83380 1 PIX4518_IN
port 4584 n
rlabel metal5 59020 -83480 59120 -83380 1 PIX4519_IN
port 4585 n
rlabel metal5 60520 -83480 60620 -83380 1 PIX4520_IN
port 4586 n
rlabel metal5 62020 -83480 62120 -83380 1 PIX4521_IN
port 4587 n
rlabel metal5 63520 -83480 63620 -83380 1 PIX4522_IN
port 4588 n
rlabel metal5 65020 -83480 65120 -83380 1 PIX4523_IN
port 4589 n
rlabel metal5 66520 -83480 66620 -83380 1 PIX4524_IN
port 4590 n
rlabel metal5 68020 -83480 68120 -83380 1 PIX4525_IN
port 4591 n
rlabel metal5 69520 -83480 69620 -83380 1 PIX4526_IN
port 4592 n
rlabel metal5 71020 -83480 71120 -83380 1 PIX4527_IN
port 4593 n
rlabel metal5 72520 -83480 72620 -83380 1 PIX4528_IN
port 4594 n
rlabel metal5 74020 -83480 74120 -83380 1 PIX4529_IN
port 4595 n
rlabel metal5 75520 -83480 75620 -83380 1 PIX4530_IN
port 4596 n
rlabel metal5 77020 -83480 77120 -83380 1 PIX4531_IN
port 4597 n
rlabel metal5 78520 -83480 78620 -83380 1 PIX4532_IN
port 4598 n
rlabel metal5 80020 -83480 80120 -83380 1 PIX4533_IN
port 4599 n
rlabel metal5 81520 -83480 81620 -83380 1 PIX4534_IN
port 4600 n
rlabel metal5 83020 -83480 83120 -83380 1 PIX4535_IN
port 4601 n
rlabel metal5 84520 -83480 84620 -83380 1 PIX4536_IN
port 4602 n
rlabel metal5 86020 -83480 86120 -83380 1 PIX4537_IN
port 4603 n
rlabel metal5 87520 -83480 87620 -83380 1 PIX4538_IN
port 4604 n
rlabel metal5 89020 -83480 89120 -83380 1 PIX4539_IN
port 4605 n
rlabel metal5 90520 -83480 90620 -83380 1 PIX4540_IN
port 4606 n
rlabel metal5 92020 -83480 92120 -83380 1 PIX4541_IN
port 4607 n
rlabel metal5 93520 -83480 93620 -83380 1 PIX4542_IN
port 4608 n
rlabel metal5 95020 -83480 95120 -83380 1 PIX4543_IN
port 4609 n
rlabel metal5 96520 -83480 96620 -83380 1 PIX4544_IN
port 4610 n
rlabel metal5 98020 -83480 98120 -83380 1 PIX4545_IN
port 4611 n
rlabel metal5 99520 -83480 99620 -83380 1 PIX4546_IN
port 4612 n
rlabel metal5 101020 -83480 101120 -83380 1 PIX4547_IN
port 4613 n
rlabel metal5 102520 -83480 102620 -83380 1 PIX4548_IN
port 4614 n
rlabel metal5 104020 -83480 104120 -83380 1 PIX4549_IN
port 4615 n
rlabel metal5 105520 -83480 105620 -83380 1 PIX4550_IN
port 4616 n
rlabel metal5 107020 -83480 107120 -83380 1 PIX4551_IN
port 4617 n
rlabel metal5 108520 -83480 108620 -83380 1 PIX4552_IN
port 4618 n
rlabel metal5 110020 -83480 110120 -83380 1 PIX4553_IN
port 4619 n
rlabel metal5 111520 -83480 111620 -83380 1 PIX4554_IN
port 4620 n
rlabel metal5 113020 -83480 113120 -83380 1 PIX4555_IN
port 4621 n
rlabel metal5 114520 -83480 114620 -83380 1 PIX4556_IN
port 4622 n
rlabel metal5 116020 -83480 116120 -83380 1 PIX4557_IN
port 4623 n
rlabel metal5 117520 -83480 117620 -83380 1 PIX4558_IN
port 4624 n
rlabel metal5 119020 -83480 119120 -83380 1 PIX4559_IN
port 4625 n
rlabel metal5 520 -84980 620 -84880 1 PIX4560_IN
port 4626 n
rlabel metal2 -1500 -84760 -1500 -84715 3 ROW_SEL57
port 4627 e
rlabel metal5 2020 -84980 2120 -84880 1 PIX4561_IN
port 4628 n
rlabel metal5 3520 -84980 3620 -84880 1 PIX4562_IN
port 4629 n
rlabel metal5 5020 -84980 5120 -84880 1 PIX4563_IN
port 4630 n
rlabel metal5 6520 -84980 6620 -84880 1 PIX4564_IN
port 4631 n
rlabel metal5 8020 -84980 8120 -84880 1 PIX4565_IN
port 4632 n
rlabel metal5 9520 -84980 9620 -84880 1 PIX4566_IN
port 4633 n
rlabel metal5 11020 -84980 11120 -84880 1 PIX4567_IN
port 4634 n
rlabel metal5 12520 -84980 12620 -84880 1 PIX4568_IN
port 4635 n
rlabel metal5 14020 -84980 14120 -84880 1 PIX4569_IN
port 4636 n
rlabel metal5 15520 -84980 15620 -84880 1 PIX4570_IN
port 4637 n
rlabel metal5 17020 -84980 17120 -84880 1 PIX4571_IN
port 4638 n
rlabel metal5 18520 -84980 18620 -84880 1 PIX4572_IN
port 4639 n
rlabel metal5 20020 -84980 20120 -84880 1 PIX4573_IN
port 4640 n
rlabel metal5 21520 -84980 21620 -84880 1 PIX4574_IN
port 4641 n
rlabel metal5 23020 -84980 23120 -84880 1 PIX4575_IN
port 4642 n
rlabel metal5 24520 -84980 24620 -84880 1 PIX4576_IN
port 4643 n
rlabel metal5 26020 -84980 26120 -84880 1 PIX4577_IN
port 4644 n
rlabel metal5 27520 -84980 27620 -84880 1 PIX4578_IN
port 4645 n
rlabel metal5 29020 -84980 29120 -84880 1 PIX4579_IN
port 4646 n
rlabel metal5 30520 -84980 30620 -84880 1 PIX4580_IN
port 4647 n
rlabel metal5 32020 -84980 32120 -84880 1 PIX4581_IN
port 4648 n
rlabel metal5 33520 -84980 33620 -84880 1 PIX4582_IN
port 4649 n
rlabel metal5 35020 -84980 35120 -84880 1 PIX4583_IN
port 4650 n
rlabel metal5 36520 -84980 36620 -84880 1 PIX4584_IN
port 4651 n
rlabel metal5 38020 -84980 38120 -84880 1 PIX4585_IN
port 4652 n
rlabel metal5 39520 -84980 39620 -84880 1 PIX4586_IN
port 4653 n
rlabel metal5 41020 -84980 41120 -84880 1 PIX4587_IN
port 4654 n
rlabel metal5 42520 -84980 42620 -84880 1 PIX4588_IN
port 4655 n
rlabel metal5 44020 -84980 44120 -84880 1 PIX4589_IN
port 4656 n
rlabel metal5 45520 -84980 45620 -84880 1 PIX4590_IN
port 4657 n
rlabel metal5 47020 -84980 47120 -84880 1 PIX4591_IN
port 4658 n
rlabel metal5 48520 -84980 48620 -84880 1 PIX4592_IN
port 4659 n
rlabel metal5 50020 -84980 50120 -84880 1 PIX4593_IN
port 4660 n
rlabel metal5 51520 -84980 51620 -84880 1 PIX4594_IN
port 4661 n
rlabel metal5 53020 -84980 53120 -84880 1 PIX4595_IN
port 4662 n
rlabel metal5 54520 -84980 54620 -84880 1 PIX4596_IN
port 4663 n
rlabel metal5 56020 -84980 56120 -84880 1 PIX4597_IN
port 4664 n
rlabel metal5 57520 -84980 57620 -84880 1 PIX4598_IN
port 4665 n
rlabel metal5 59020 -84980 59120 -84880 1 PIX4599_IN
port 4666 n
rlabel metal5 60520 -84980 60620 -84880 1 PIX4600_IN
port 4667 n
rlabel metal5 62020 -84980 62120 -84880 1 PIX4601_IN
port 4668 n
rlabel metal5 63520 -84980 63620 -84880 1 PIX4602_IN
port 4669 n
rlabel metal5 65020 -84980 65120 -84880 1 PIX4603_IN
port 4670 n
rlabel metal5 66520 -84980 66620 -84880 1 PIX4604_IN
port 4671 n
rlabel metal5 68020 -84980 68120 -84880 1 PIX4605_IN
port 4672 n
rlabel metal5 69520 -84980 69620 -84880 1 PIX4606_IN
port 4673 n
rlabel metal5 71020 -84980 71120 -84880 1 PIX4607_IN
port 4674 n
rlabel metal5 72520 -84980 72620 -84880 1 PIX4608_IN
port 4675 n
rlabel metal5 74020 -84980 74120 -84880 1 PIX4609_IN
port 4676 n
rlabel metal5 75520 -84980 75620 -84880 1 PIX4610_IN
port 4677 n
rlabel metal5 77020 -84980 77120 -84880 1 PIX4611_IN
port 4678 n
rlabel metal5 78520 -84980 78620 -84880 1 PIX4612_IN
port 4679 n
rlabel metal5 80020 -84980 80120 -84880 1 PIX4613_IN
port 4680 n
rlabel metal5 81520 -84980 81620 -84880 1 PIX4614_IN
port 4681 n
rlabel metal5 83020 -84980 83120 -84880 1 PIX4615_IN
port 4682 n
rlabel metal5 84520 -84980 84620 -84880 1 PIX4616_IN
port 4683 n
rlabel metal5 86020 -84980 86120 -84880 1 PIX4617_IN
port 4684 n
rlabel metal5 87520 -84980 87620 -84880 1 PIX4618_IN
port 4685 n
rlabel metal5 89020 -84980 89120 -84880 1 PIX4619_IN
port 4686 n
rlabel metal5 90520 -84980 90620 -84880 1 PIX4620_IN
port 4687 n
rlabel metal5 92020 -84980 92120 -84880 1 PIX4621_IN
port 4688 n
rlabel metal5 93520 -84980 93620 -84880 1 PIX4622_IN
port 4689 n
rlabel metal5 95020 -84980 95120 -84880 1 PIX4623_IN
port 4690 n
rlabel metal5 96520 -84980 96620 -84880 1 PIX4624_IN
port 4691 n
rlabel metal5 98020 -84980 98120 -84880 1 PIX4625_IN
port 4692 n
rlabel metal5 99520 -84980 99620 -84880 1 PIX4626_IN
port 4693 n
rlabel metal5 101020 -84980 101120 -84880 1 PIX4627_IN
port 4694 n
rlabel metal5 102520 -84980 102620 -84880 1 PIX4628_IN
port 4695 n
rlabel metal5 104020 -84980 104120 -84880 1 PIX4629_IN
port 4696 n
rlabel metal5 105520 -84980 105620 -84880 1 PIX4630_IN
port 4697 n
rlabel metal5 107020 -84980 107120 -84880 1 PIX4631_IN
port 4698 n
rlabel metal5 108520 -84980 108620 -84880 1 PIX4632_IN
port 4699 n
rlabel metal5 110020 -84980 110120 -84880 1 PIX4633_IN
port 4700 n
rlabel metal5 111520 -84980 111620 -84880 1 PIX4634_IN
port 4701 n
rlabel metal5 113020 -84980 113120 -84880 1 PIX4635_IN
port 4702 n
rlabel metal5 114520 -84980 114620 -84880 1 PIX4636_IN
port 4703 n
rlabel metal5 116020 -84980 116120 -84880 1 PIX4637_IN
port 4704 n
rlabel metal5 117520 -84980 117620 -84880 1 PIX4638_IN
port 4705 n
rlabel metal5 119020 -84980 119120 -84880 1 PIX4639_IN
port 4706 n
rlabel metal5 520 -86480 620 -86380 1 PIX4640_IN
port 4707 n
rlabel metal2 -1500 -86260 -1500 -86215 3 ROW_SEL58
port 4708 e
rlabel metal5 2020 -86480 2120 -86380 1 PIX4641_IN
port 4709 n
rlabel metal5 3520 -86480 3620 -86380 1 PIX4642_IN
port 4710 n
rlabel metal5 5020 -86480 5120 -86380 1 PIX4643_IN
port 4711 n
rlabel metal5 6520 -86480 6620 -86380 1 PIX4644_IN
port 4712 n
rlabel metal5 8020 -86480 8120 -86380 1 PIX4645_IN
port 4713 n
rlabel metal5 9520 -86480 9620 -86380 1 PIX4646_IN
port 4714 n
rlabel metal5 11020 -86480 11120 -86380 1 PIX4647_IN
port 4715 n
rlabel metal5 12520 -86480 12620 -86380 1 PIX4648_IN
port 4716 n
rlabel metal5 14020 -86480 14120 -86380 1 PIX4649_IN
port 4717 n
rlabel metal5 15520 -86480 15620 -86380 1 PIX4650_IN
port 4718 n
rlabel metal5 17020 -86480 17120 -86380 1 PIX4651_IN
port 4719 n
rlabel metal5 18520 -86480 18620 -86380 1 PIX4652_IN
port 4720 n
rlabel metal5 20020 -86480 20120 -86380 1 PIX4653_IN
port 4721 n
rlabel metal5 21520 -86480 21620 -86380 1 PIX4654_IN
port 4722 n
rlabel metal5 23020 -86480 23120 -86380 1 PIX4655_IN
port 4723 n
rlabel metal5 24520 -86480 24620 -86380 1 PIX4656_IN
port 4724 n
rlabel metal5 26020 -86480 26120 -86380 1 PIX4657_IN
port 4725 n
rlabel metal5 27520 -86480 27620 -86380 1 PIX4658_IN
port 4726 n
rlabel metal5 29020 -86480 29120 -86380 1 PIX4659_IN
port 4727 n
rlabel metal5 30520 -86480 30620 -86380 1 PIX4660_IN
port 4728 n
rlabel metal5 32020 -86480 32120 -86380 1 PIX4661_IN
port 4729 n
rlabel metal5 33520 -86480 33620 -86380 1 PIX4662_IN
port 4730 n
rlabel metal5 35020 -86480 35120 -86380 1 PIX4663_IN
port 4731 n
rlabel metal5 36520 -86480 36620 -86380 1 PIX4664_IN
port 4732 n
rlabel metal5 38020 -86480 38120 -86380 1 PIX4665_IN
port 4733 n
rlabel metal5 39520 -86480 39620 -86380 1 PIX4666_IN
port 4734 n
rlabel metal5 41020 -86480 41120 -86380 1 PIX4667_IN
port 4735 n
rlabel metal5 42520 -86480 42620 -86380 1 PIX4668_IN
port 4736 n
rlabel metal5 44020 -86480 44120 -86380 1 PIX4669_IN
port 4737 n
rlabel metal5 45520 -86480 45620 -86380 1 PIX4670_IN
port 4738 n
rlabel metal5 47020 -86480 47120 -86380 1 PIX4671_IN
port 4739 n
rlabel metal5 48520 -86480 48620 -86380 1 PIX4672_IN
port 4740 n
rlabel metal5 50020 -86480 50120 -86380 1 PIX4673_IN
port 4741 n
rlabel metal5 51520 -86480 51620 -86380 1 PIX4674_IN
port 4742 n
rlabel metal5 53020 -86480 53120 -86380 1 PIX4675_IN
port 4743 n
rlabel metal5 54520 -86480 54620 -86380 1 PIX4676_IN
port 4744 n
rlabel metal5 56020 -86480 56120 -86380 1 PIX4677_IN
port 4745 n
rlabel metal5 57520 -86480 57620 -86380 1 PIX4678_IN
port 4746 n
rlabel metal5 59020 -86480 59120 -86380 1 PIX4679_IN
port 4747 n
rlabel metal5 60520 -86480 60620 -86380 1 PIX4680_IN
port 4748 n
rlabel metal5 62020 -86480 62120 -86380 1 PIX4681_IN
port 4749 n
rlabel metal5 63520 -86480 63620 -86380 1 PIX4682_IN
port 4750 n
rlabel metal5 65020 -86480 65120 -86380 1 PIX4683_IN
port 4751 n
rlabel metal5 66520 -86480 66620 -86380 1 PIX4684_IN
port 4752 n
rlabel metal5 68020 -86480 68120 -86380 1 PIX4685_IN
port 4753 n
rlabel metal5 69520 -86480 69620 -86380 1 PIX4686_IN
port 4754 n
rlabel metal5 71020 -86480 71120 -86380 1 PIX4687_IN
port 4755 n
rlabel metal5 72520 -86480 72620 -86380 1 PIX4688_IN
port 4756 n
rlabel metal5 74020 -86480 74120 -86380 1 PIX4689_IN
port 4757 n
rlabel metal5 75520 -86480 75620 -86380 1 PIX4690_IN
port 4758 n
rlabel metal5 77020 -86480 77120 -86380 1 PIX4691_IN
port 4759 n
rlabel metal5 78520 -86480 78620 -86380 1 PIX4692_IN
port 4760 n
rlabel metal5 80020 -86480 80120 -86380 1 PIX4693_IN
port 4761 n
rlabel metal5 81520 -86480 81620 -86380 1 PIX4694_IN
port 4762 n
rlabel metal5 83020 -86480 83120 -86380 1 PIX4695_IN
port 4763 n
rlabel metal5 84520 -86480 84620 -86380 1 PIX4696_IN
port 4764 n
rlabel metal5 86020 -86480 86120 -86380 1 PIX4697_IN
port 4765 n
rlabel metal5 87520 -86480 87620 -86380 1 PIX4698_IN
port 4766 n
rlabel metal5 89020 -86480 89120 -86380 1 PIX4699_IN
port 4767 n
rlabel metal5 90520 -86480 90620 -86380 1 PIX4700_IN
port 4768 n
rlabel metal5 92020 -86480 92120 -86380 1 PIX4701_IN
port 4769 n
rlabel metal5 93520 -86480 93620 -86380 1 PIX4702_IN
port 4770 n
rlabel metal5 95020 -86480 95120 -86380 1 PIX4703_IN
port 4771 n
rlabel metal5 96520 -86480 96620 -86380 1 PIX4704_IN
port 4772 n
rlabel metal5 98020 -86480 98120 -86380 1 PIX4705_IN
port 4773 n
rlabel metal5 99520 -86480 99620 -86380 1 PIX4706_IN
port 4774 n
rlabel metal5 101020 -86480 101120 -86380 1 PIX4707_IN
port 4775 n
rlabel metal5 102520 -86480 102620 -86380 1 PIX4708_IN
port 4776 n
rlabel metal5 104020 -86480 104120 -86380 1 PIX4709_IN
port 4777 n
rlabel metal5 105520 -86480 105620 -86380 1 PIX4710_IN
port 4778 n
rlabel metal5 107020 -86480 107120 -86380 1 PIX4711_IN
port 4779 n
rlabel metal5 108520 -86480 108620 -86380 1 PIX4712_IN
port 4780 n
rlabel metal5 110020 -86480 110120 -86380 1 PIX4713_IN
port 4781 n
rlabel metal5 111520 -86480 111620 -86380 1 PIX4714_IN
port 4782 n
rlabel metal5 113020 -86480 113120 -86380 1 PIX4715_IN
port 4783 n
rlabel metal5 114520 -86480 114620 -86380 1 PIX4716_IN
port 4784 n
rlabel metal5 116020 -86480 116120 -86380 1 PIX4717_IN
port 4785 n
rlabel metal5 117520 -86480 117620 -86380 1 PIX4718_IN
port 4786 n
rlabel metal5 119020 -86480 119120 -86380 1 PIX4719_IN
port 4787 n
rlabel metal5 520 -87980 620 -87880 1 PIX4720_IN
port 4788 n
rlabel metal2 -1500 -87760 -1500 -87715 3 ROW_SEL59
port 4789 e
rlabel metal5 2020 -87980 2120 -87880 1 PIX4721_IN
port 4790 n
rlabel metal5 3520 -87980 3620 -87880 1 PIX4722_IN
port 4791 n
rlabel metal5 5020 -87980 5120 -87880 1 PIX4723_IN
port 4792 n
rlabel metal5 6520 -87980 6620 -87880 1 PIX4724_IN
port 4793 n
rlabel metal5 8020 -87980 8120 -87880 1 PIX4725_IN
port 4794 n
rlabel metal5 9520 -87980 9620 -87880 1 PIX4726_IN
port 4795 n
rlabel metal5 11020 -87980 11120 -87880 1 PIX4727_IN
port 4796 n
rlabel metal5 12520 -87980 12620 -87880 1 PIX4728_IN
port 4797 n
rlabel metal5 14020 -87980 14120 -87880 1 PIX4729_IN
port 4798 n
rlabel metal5 15520 -87980 15620 -87880 1 PIX4730_IN
port 4799 n
rlabel metal5 17020 -87980 17120 -87880 1 PIX4731_IN
port 4800 n
rlabel metal5 18520 -87980 18620 -87880 1 PIX4732_IN
port 4801 n
rlabel metal5 20020 -87980 20120 -87880 1 PIX4733_IN
port 4802 n
rlabel metal5 21520 -87980 21620 -87880 1 PIX4734_IN
port 4803 n
rlabel metal5 23020 -87980 23120 -87880 1 PIX4735_IN
port 4804 n
rlabel metal5 24520 -87980 24620 -87880 1 PIX4736_IN
port 4805 n
rlabel metal5 26020 -87980 26120 -87880 1 PIX4737_IN
port 4806 n
rlabel metal5 27520 -87980 27620 -87880 1 PIX4738_IN
port 4807 n
rlabel metal5 29020 -87980 29120 -87880 1 PIX4739_IN
port 4808 n
rlabel metal5 30520 -87980 30620 -87880 1 PIX4740_IN
port 4809 n
rlabel metal5 32020 -87980 32120 -87880 1 PIX4741_IN
port 4810 n
rlabel metal5 33520 -87980 33620 -87880 1 PIX4742_IN
port 4811 n
rlabel metal5 35020 -87980 35120 -87880 1 PIX4743_IN
port 4812 n
rlabel metal5 36520 -87980 36620 -87880 1 PIX4744_IN
port 4813 n
rlabel metal5 38020 -87980 38120 -87880 1 PIX4745_IN
port 4814 n
rlabel metal5 39520 -87980 39620 -87880 1 PIX4746_IN
port 4815 n
rlabel metal5 41020 -87980 41120 -87880 1 PIX4747_IN
port 4816 n
rlabel metal5 42520 -87980 42620 -87880 1 PIX4748_IN
port 4817 n
rlabel metal5 44020 -87980 44120 -87880 1 PIX4749_IN
port 4818 n
rlabel metal5 45520 -87980 45620 -87880 1 PIX4750_IN
port 4819 n
rlabel metal5 47020 -87980 47120 -87880 1 PIX4751_IN
port 4820 n
rlabel metal5 48520 -87980 48620 -87880 1 PIX4752_IN
port 4821 n
rlabel metal5 50020 -87980 50120 -87880 1 PIX4753_IN
port 4822 n
rlabel metal5 51520 -87980 51620 -87880 1 PIX4754_IN
port 4823 n
rlabel metal5 53020 -87980 53120 -87880 1 PIX4755_IN
port 4824 n
rlabel metal5 54520 -87980 54620 -87880 1 PIX4756_IN
port 4825 n
rlabel metal5 56020 -87980 56120 -87880 1 PIX4757_IN
port 4826 n
rlabel metal5 57520 -87980 57620 -87880 1 PIX4758_IN
port 4827 n
rlabel metal5 59020 -87980 59120 -87880 1 PIX4759_IN
port 4828 n
rlabel metal5 60520 -87980 60620 -87880 1 PIX4760_IN
port 4829 n
rlabel metal5 62020 -87980 62120 -87880 1 PIX4761_IN
port 4830 n
rlabel metal5 63520 -87980 63620 -87880 1 PIX4762_IN
port 4831 n
rlabel metal5 65020 -87980 65120 -87880 1 PIX4763_IN
port 4832 n
rlabel metal5 66520 -87980 66620 -87880 1 PIX4764_IN
port 4833 n
rlabel metal5 68020 -87980 68120 -87880 1 PIX4765_IN
port 4834 n
rlabel metal5 69520 -87980 69620 -87880 1 PIX4766_IN
port 4835 n
rlabel metal5 71020 -87980 71120 -87880 1 PIX4767_IN
port 4836 n
rlabel metal5 72520 -87980 72620 -87880 1 PIX4768_IN
port 4837 n
rlabel metal5 74020 -87980 74120 -87880 1 PIX4769_IN
port 4838 n
rlabel metal5 75520 -87980 75620 -87880 1 PIX4770_IN
port 4839 n
rlabel metal5 77020 -87980 77120 -87880 1 PIX4771_IN
port 4840 n
rlabel metal5 78520 -87980 78620 -87880 1 PIX4772_IN
port 4841 n
rlabel metal5 80020 -87980 80120 -87880 1 PIX4773_IN
port 4842 n
rlabel metal5 81520 -87980 81620 -87880 1 PIX4774_IN
port 4843 n
rlabel metal5 83020 -87980 83120 -87880 1 PIX4775_IN
port 4844 n
rlabel metal5 84520 -87980 84620 -87880 1 PIX4776_IN
port 4845 n
rlabel metal5 86020 -87980 86120 -87880 1 PIX4777_IN
port 4846 n
rlabel metal5 87520 -87980 87620 -87880 1 PIX4778_IN
port 4847 n
rlabel metal5 89020 -87980 89120 -87880 1 PIX4779_IN
port 4848 n
rlabel metal5 90520 -87980 90620 -87880 1 PIX4780_IN
port 4849 n
rlabel metal5 92020 -87980 92120 -87880 1 PIX4781_IN
port 4850 n
rlabel metal5 93520 -87980 93620 -87880 1 PIX4782_IN
port 4851 n
rlabel metal5 95020 -87980 95120 -87880 1 PIX4783_IN
port 4852 n
rlabel metal5 96520 -87980 96620 -87880 1 PIX4784_IN
port 4853 n
rlabel metal5 98020 -87980 98120 -87880 1 PIX4785_IN
port 4854 n
rlabel metal5 99520 -87980 99620 -87880 1 PIX4786_IN
port 4855 n
rlabel metal5 101020 -87980 101120 -87880 1 PIX4787_IN
port 4856 n
rlabel metal5 102520 -87980 102620 -87880 1 PIX4788_IN
port 4857 n
rlabel metal5 104020 -87980 104120 -87880 1 PIX4789_IN
port 4858 n
rlabel metal5 105520 -87980 105620 -87880 1 PIX4790_IN
port 4859 n
rlabel metal5 107020 -87980 107120 -87880 1 PIX4791_IN
port 4860 n
rlabel metal5 108520 -87980 108620 -87880 1 PIX4792_IN
port 4861 n
rlabel metal5 110020 -87980 110120 -87880 1 PIX4793_IN
port 4862 n
rlabel metal5 111520 -87980 111620 -87880 1 PIX4794_IN
port 4863 n
rlabel metal5 113020 -87980 113120 -87880 1 PIX4795_IN
port 4864 n
rlabel metal5 114520 -87980 114620 -87880 1 PIX4796_IN
port 4865 n
rlabel metal5 116020 -87980 116120 -87880 1 PIX4797_IN
port 4866 n
rlabel metal5 117520 -87980 117620 -87880 1 PIX4798_IN
port 4867 n
rlabel metal5 119020 -87980 119120 -87880 1 PIX4799_IN
port 4868 n
rlabel metal5 520 -89480 620 -89380 1 PIX4800_IN
port 4869 n
rlabel metal2 -1500 -89260 -1500 -89215 3 ROW_SEL60
port 4870 e
rlabel metal5 2020 -89480 2120 -89380 1 PIX4801_IN
port 4871 n
rlabel metal5 3520 -89480 3620 -89380 1 PIX4802_IN
port 4872 n
rlabel metal5 5020 -89480 5120 -89380 1 PIX4803_IN
port 4873 n
rlabel metal5 6520 -89480 6620 -89380 1 PIX4804_IN
port 4874 n
rlabel metal5 8020 -89480 8120 -89380 1 PIX4805_IN
port 4875 n
rlabel metal5 9520 -89480 9620 -89380 1 PIX4806_IN
port 4876 n
rlabel metal5 11020 -89480 11120 -89380 1 PIX4807_IN
port 4877 n
rlabel metal5 12520 -89480 12620 -89380 1 PIX4808_IN
port 4878 n
rlabel metal5 14020 -89480 14120 -89380 1 PIX4809_IN
port 4879 n
rlabel metal5 15520 -89480 15620 -89380 1 PIX4810_IN
port 4880 n
rlabel metal5 17020 -89480 17120 -89380 1 PIX4811_IN
port 4881 n
rlabel metal5 18520 -89480 18620 -89380 1 PIX4812_IN
port 4882 n
rlabel metal5 20020 -89480 20120 -89380 1 PIX4813_IN
port 4883 n
rlabel metal5 21520 -89480 21620 -89380 1 PIX4814_IN
port 4884 n
rlabel metal5 23020 -89480 23120 -89380 1 PIX4815_IN
port 4885 n
rlabel metal5 24520 -89480 24620 -89380 1 PIX4816_IN
port 4886 n
rlabel metal5 26020 -89480 26120 -89380 1 PIX4817_IN
port 4887 n
rlabel metal5 27520 -89480 27620 -89380 1 PIX4818_IN
port 4888 n
rlabel metal5 29020 -89480 29120 -89380 1 PIX4819_IN
port 4889 n
rlabel metal5 30520 -89480 30620 -89380 1 PIX4820_IN
port 4890 n
rlabel metal5 32020 -89480 32120 -89380 1 PIX4821_IN
port 4891 n
rlabel metal5 33520 -89480 33620 -89380 1 PIX4822_IN
port 4892 n
rlabel metal5 35020 -89480 35120 -89380 1 PIX4823_IN
port 4893 n
rlabel metal5 36520 -89480 36620 -89380 1 PIX4824_IN
port 4894 n
rlabel metal5 38020 -89480 38120 -89380 1 PIX4825_IN
port 4895 n
rlabel metal5 39520 -89480 39620 -89380 1 PIX4826_IN
port 4896 n
rlabel metal5 41020 -89480 41120 -89380 1 PIX4827_IN
port 4897 n
rlabel metal5 42520 -89480 42620 -89380 1 PIX4828_IN
port 4898 n
rlabel metal5 44020 -89480 44120 -89380 1 PIX4829_IN
port 4899 n
rlabel metal5 45520 -89480 45620 -89380 1 PIX4830_IN
port 4900 n
rlabel metal5 47020 -89480 47120 -89380 1 PIX4831_IN
port 4901 n
rlabel metal5 48520 -89480 48620 -89380 1 PIX4832_IN
port 4902 n
rlabel metal5 50020 -89480 50120 -89380 1 PIX4833_IN
port 4903 n
rlabel metal5 51520 -89480 51620 -89380 1 PIX4834_IN
port 4904 n
rlabel metal5 53020 -89480 53120 -89380 1 PIX4835_IN
port 4905 n
rlabel metal5 54520 -89480 54620 -89380 1 PIX4836_IN
port 4906 n
rlabel metal5 56020 -89480 56120 -89380 1 PIX4837_IN
port 4907 n
rlabel metal5 57520 -89480 57620 -89380 1 PIX4838_IN
port 4908 n
rlabel metal5 59020 -89480 59120 -89380 1 PIX4839_IN
port 4909 n
rlabel metal5 60520 -89480 60620 -89380 1 PIX4840_IN
port 4910 n
rlabel metal5 62020 -89480 62120 -89380 1 PIX4841_IN
port 4911 n
rlabel metal5 63520 -89480 63620 -89380 1 PIX4842_IN
port 4912 n
rlabel metal5 65020 -89480 65120 -89380 1 PIX4843_IN
port 4913 n
rlabel metal5 66520 -89480 66620 -89380 1 PIX4844_IN
port 4914 n
rlabel metal5 68020 -89480 68120 -89380 1 PIX4845_IN
port 4915 n
rlabel metal5 69520 -89480 69620 -89380 1 PIX4846_IN
port 4916 n
rlabel metal5 71020 -89480 71120 -89380 1 PIX4847_IN
port 4917 n
rlabel metal5 72520 -89480 72620 -89380 1 PIX4848_IN
port 4918 n
rlabel metal5 74020 -89480 74120 -89380 1 PIX4849_IN
port 4919 n
rlabel metal5 75520 -89480 75620 -89380 1 PIX4850_IN
port 4920 n
rlabel metal5 77020 -89480 77120 -89380 1 PIX4851_IN
port 4921 n
rlabel metal5 78520 -89480 78620 -89380 1 PIX4852_IN
port 4922 n
rlabel metal5 80020 -89480 80120 -89380 1 PIX4853_IN
port 4923 n
rlabel metal5 81520 -89480 81620 -89380 1 PIX4854_IN
port 4924 n
rlabel metal5 83020 -89480 83120 -89380 1 PIX4855_IN
port 4925 n
rlabel metal5 84520 -89480 84620 -89380 1 PIX4856_IN
port 4926 n
rlabel metal5 86020 -89480 86120 -89380 1 PIX4857_IN
port 4927 n
rlabel metal5 87520 -89480 87620 -89380 1 PIX4858_IN
port 4928 n
rlabel metal5 89020 -89480 89120 -89380 1 PIX4859_IN
port 4929 n
rlabel metal5 90520 -89480 90620 -89380 1 PIX4860_IN
port 4930 n
rlabel metal5 92020 -89480 92120 -89380 1 PIX4861_IN
port 4931 n
rlabel metal5 93520 -89480 93620 -89380 1 PIX4862_IN
port 4932 n
rlabel metal5 95020 -89480 95120 -89380 1 PIX4863_IN
port 4933 n
rlabel metal5 96520 -89480 96620 -89380 1 PIX4864_IN
port 4934 n
rlabel metal5 98020 -89480 98120 -89380 1 PIX4865_IN
port 4935 n
rlabel metal5 99520 -89480 99620 -89380 1 PIX4866_IN
port 4936 n
rlabel metal5 101020 -89480 101120 -89380 1 PIX4867_IN
port 4937 n
rlabel metal5 102520 -89480 102620 -89380 1 PIX4868_IN
port 4938 n
rlabel metal5 104020 -89480 104120 -89380 1 PIX4869_IN
port 4939 n
rlabel metal5 105520 -89480 105620 -89380 1 PIX4870_IN
port 4940 n
rlabel metal5 107020 -89480 107120 -89380 1 PIX4871_IN
port 4941 n
rlabel metal5 108520 -89480 108620 -89380 1 PIX4872_IN
port 4942 n
rlabel metal5 110020 -89480 110120 -89380 1 PIX4873_IN
port 4943 n
rlabel metal5 111520 -89480 111620 -89380 1 PIX4874_IN
port 4944 n
rlabel metal5 113020 -89480 113120 -89380 1 PIX4875_IN
port 4945 n
rlabel metal5 114520 -89480 114620 -89380 1 PIX4876_IN
port 4946 n
rlabel metal5 116020 -89480 116120 -89380 1 PIX4877_IN
port 4947 n
rlabel metal5 117520 -89480 117620 -89380 1 PIX4878_IN
port 4948 n
rlabel metal5 119020 -89480 119120 -89380 1 PIX4879_IN
port 4949 n
rlabel metal5 520 -90980 620 -90880 1 PIX4880_IN
port 4950 n
rlabel metal2 -1500 -90760 -1500 -90715 3 ROW_SEL61
port 4951 e
rlabel metal5 2020 -90980 2120 -90880 1 PIX4881_IN
port 4952 n
rlabel metal5 3520 -90980 3620 -90880 1 PIX4882_IN
port 4953 n
rlabel metal5 5020 -90980 5120 -90880 1 PIX4883_IN
port 4954 n
rlabel metal5 6520 -90980 6620 -90880 1 PIX4884_IN
port 4955 n
rlabel metal5 8020 -90980 8120 -90880 1 PIX4885_IN
port 4956 n
rlabel metal5 9520 -90980 9620 -90880 1 PIX4886_IN
port 4957 n
rlabel metal5 11020 -90980 11120 -90880 1 PIX4887_IN
port 4958 n
rlabel metal5 12520 -90980 12620 -90880 1 PIX4888_IN
port 4959 n
rlabel metal5 14020 -90980 14120 -90880 1 PIX4889_IN
port 4960 n
rlabel metal5 15520 -90980 15620 -90880 1 PIX4890_IN
port 4961 n
rlabel metal5 17020 -90980 17120 -90880 1 PIX4891_IN
port 4962 n
rlabel metal5 18520 -90980 18620 -90880 1 PIX4892_IN
port 4963 n
rlabel metal5 20020 -90980 20120 -90880 1 PIX4893_IN
port 4964 n
rlabel metal5 21520 -90980 21620 -90880 1 PIX4894_IN
port 4965 n
rlabel metal5 23020 -90980 23120 -90880 1 PIX4895_IN
port 4966 n
rlabel metal5 24520 -90980 24620 -90880 1 PIX4896_IN
port 4967 n
rlabel metal5 26020 -90980 26120 -90880 1 PIX4897_IN
port 4968 n
rlabel metal5 27520 -90980 27620 -90880 1 PIX4898_IN
port 4969 n
rlabel metal5 29020 -90980 29120 -90880 1 PIX4899_IN
port 4970 n
rlabel metal5 30520 -90980 30620 -90880 1 PIX4900_IN
port 4971 n
rlabel metal5 32020 -90980 32120 -90880 1 PIX4901_IN
port 4972 n
rlabel metal5 33520 -90980 33620 -90880 1 PIX4902_IN
port 4973 n
rlabel metal5 35020 -90980 35120 -90880 1 PIX4903_IN
port 4974 n
rlabel metal5 36520 -90980 36620 -90880 1 PIX4904_IN
port 4975 n
rlabel metal5 38020 -90980 38120 -90880 1 PIX4905_IN
port 4976 n
rlabel metal5 39520 -90980 39620 -90880 1 PIX4906_IN
port 4977 n
rlabel metal5 41020 -90980 41120 -90880 1 PIX4907_IN
port 4978 n
rlabel metal5 42520 -90980 42620 -90880 1 PIX4908_IN
port 4979 n
rlabel metal5 44020 -90980 44120 -90880 1 PIX4909_IN
port 4980 n
rlabel metal5 45520 -90980 45620 -90880 1 PIX4910_IN
port 4981 n
rlabel metal5 47020 -90980 47120 -90880 1 PIX4911_IN
port 4982 n
rlabel metal5 48520 -90980 48620 -90880 1 PIX4912_IN
port 4983 n
rlabel metal5 50020 -90980 50120 -90880 1 PIX4913_IN
port 4984 n
rlabel metal5 51520 -90980 51620 -90880 1 PIX4914_IN
port 4985 n
rlabel metal5 53020 -90980 53120 -90880 1 PIX4915_IN
port 4986 n
rlabel metal5 54520 -90980 54620 -90880 1 PIX4916_IN
port 4987 n
rlabel metal5 56020 -90980 56120 -90880 1 PIX4917_IN
port 4988 n
rlabel metal5 57520 -90980 57620 -90880 1 PIX4918_IN
port 4989 n
rlabel metal5 59020 -90980 59120 -90880 1 PIX4919_IN
port 4990 n
rlabel metal5 60520 -90980 60620 -90880 1 PIX4920_IN
port 4991 n
rlabel metal5 62020 -90980 62120 -90880 1 PIX4921_IN
port 4992 n
rlabel metal5 63520 -90980 63620 -90880 1 PIX4922_IN
port 4993 n
rlabel metal5 65020 -90980 65120 -90880 1 PIX4923_IN
port 4994 n
rlabel metal5 66520 -90980 66620 -90880 1 PIX4924_IN
port 4995 n
rlabel metal5 68020 -90980 68120 -90880 1 PIX4925_IN
port 4996 n
rlabel metal5 69520 -90980 69620 -90880 1 PIX4926_IN
port 4997 n
rlabel metal5 71020 -90980 71120 -90880 1 PIX4927_IN
port 4998 n
rlabel metal5 72520 -90980 72620 -90880 1 PIX4928_IN
port 4999 n
rlabel metal5 74020 -90980 74120 -90880 1 PIX4929_IN
port 5000 n
rlabel metal5 75520 -90980 75620 -90880 1 PIX4930_IN
port 5001 n
rlabel metal5 77020 -90980 77120 -90880 1 PIX4931_IN
port 5002 n
rlabel metal5 78520 -90980 78620 -90880 1 PIX4932_IN
port 5003 n
rlabel metal5 80020 -90980 80120 -90880 1 PIX4933_IN
port 5004 n
rlabel metal5 81520 -90980 81620 -90880 1 PIX4934_IN
port 5005 n
rlabel metal5 83020 -90980 83120 -90880 1 PIX4935_IN
port 5006 n
rlabel metal5 84520 -90980 84620 -90880 1 PIX4936_IN
port 5007 n
rlabel metal5 86020 -90980 86120 -90880 1 PIX4937_IN
port 5008 n
rlabel metal5 87520 -90980 87620 -90880 1 PIX4938_IN
port 5009 n
rlabel metal5 89020 -90980 89120 -90880 1 PIX4939_IN
port 5010 n
rlabel metal5 90520 -90980 90620 -90880 1 PIX4940_IN
port 5011 n
rlabel metal5 92020 -90980 92120 -90880 1 PIX4941_IN
port 5012 n
rlabel metal5 93520 -90980 93620 -90880 1 PIX4942_IN
port 5013 n
rlabel metal5 95020 -90980 95120 -90880 1 PIX4943_IN
port 5014 n
rlabel metal5 96520 -90980 96620 -90880 1 PIX4944_IN
port 5015 n
rlabel metal5 98020 -90980 98120 -90880 1 PIX4945_IN
port 5016 n
rlabel metal5 99520 -90980 99620 -90880 1 PIX4946_IN
port 5017 n
rlabel metal5 101020 -90980 101120 -90880 1 PIX4947_IN
port 5018 n
rlabel metal5 102520 -90980 102620 -90880 1 PIX4948_IN
port 5019 n
rlabel metal5 104020 -90980 104120 -90880 1 PIX4949_IN
port 5020 n
rlabel metal5 105520 -90980 105620 -90880 1 PIX4950_IN
port 5021 n
rlabel metal5 107020 -90980 107120 -90880 1 PIX4951_IN
port 5022 n
rlabel metal5 108520 -90980 108620 -90880 1 PIX4952_IN
port 5023 n
rlabel metal5 110020 -90980 110120 -90880 1 PIX4953_IN
port 5024 n
rlabel metal5 111520 -90980 111620 -90880 1 PIX4954_IN
port 5025 n
rlabel metal5 113020 -90980 113120 -90880 1 PIX4955_IN
port 5026 n
rlabel metal5 114520 -90980 114620 -90880 1 PIX4956_IN
port 5027 n
rlabel metal5 116020 -90980 116120 -90880 1 PIX4957_IN
port 5028 n
rlabel metal5 117520 -90980 117620 -90880 1 PIX4958_IN
port 5029 n
rlabel metal5 119020 -90980 119120 -90880 1 PIX4959_IN
port 5030 n
rlabel metal5 520 -92480 620 -92380 1 PIX4960_IN
port 5031 n
rlabel metal2 -1500 -92260 -1500 -92215 3 ROW_SEL62
port 5032 e
rlabel metal5 2020 -92480 2120 -92380 1 PIX4961_IN
port 5033 n
rlabel metal5 3520 -92480 3620 -92380 1 PIX4962_IN
port 5034 n
rlabel metal5 5020 -92480 5120 -92380 1 PIX4963_IN
port 5035 n
rlabel metal5 6520 -92480 6620 -92380 1 PIX4964_IN
port 5036 n
rlabel metal5 8020 -92480 8120 -92380 1 PIX4965_IN
port 5037 n
rlabel metal5 9520 -92480 9620 -92380 1 PIX4966_IN
port 5038 n
rlabel metal5 11020 -92480 11120 -92380 1 PIX4967_IN
port 5039 n
rlabel metal5 12520 -92480 12620 -92380 1 PIX4968_IN
port 5040 n
rlabel metal5 14020 -92480 14120 -92380 1 PIX4969_IN
port 5041 n
rlabel metal5 15520 -92480 15620 -92380 1 PIX4970_IN
port 5042 n
rlabel metal5 17020 -92480 17120 -92380 1 PIX4971_IN
port 5043 n
rlabel metal5 18520 -92480 18620 -92380 1 PIX4972_IN
port 5044 n
rlabel metal5 20020 -92480 20120 -92380 1 PIX4973_IN
port 5045 n
rlabel metal5 21520 -92480 21620 -92380 1 PIX4974_IN
port 5046 n
rlabel metal5 23020 -92480 23120 -92380 1 PIX4975_IN
port 5047 n
rlabel metal5 24520 -92480 24620 -92380 1 PIX4976_IN
port 5048 n
rlabel metal5 26020 -92480 26120 -92380 1 PIX4977_IN
port 5049 n
rlabel metal5 27520 -92480 27620 -92380 1 PIX4978_IN
port 5050 n
rlabel metal5 29020 -92480 29120 -92380 1 PIX4979_IN
port 5051 n
rlabel metal5 30520 -92480 30620 -92380 1 PIX4980_IN
port 5052 n
rlabel metal5 32020 -92480 32120 -92380 1 PIX4981_IN
port 5053 n
rlabel metal5 33520 -92480 33620 -92380 1 PIX4982_IN
port 5054 n
rlabel metal5 35020 -92480 35120 -92380 1 PIX4983_IN
port 5055 n
rlabel metal5 36520 -92480 36620 -92380 1 PIX4984_IN
port 5056 n
rlabel metal5 38020 -92480 38120 -92380 1 PIX4985_IN
port 5057 n
rlabel metal5 39520 -92480 39620 -92380 1 PIX4986_IN
port 5058 n
rlabel metal5 41020 -92480 41120 -92380 1 PIX4987_IN
port 5059 n
rlabel metal5 42520 -92480 42620 -92380 1 PIX4988_IN
port 5060 n
rlabel metal5 44020 -92480 44120 -92380 1 PIX4989_IN
port 5061 n
rlabel metal5 45520 -92480 45620 -92380 1 PIX4990_IN
port 5062 n
rlabel metal5 47020 -92480 47120 -92380 1 PIX4991_IN
port 5063 n
rlabel metal5 48520 -92480 48620 -92380 1 PIX4992_IN
port 5064 n
rlabel metal5 50020 -92480 50120 -92380 1 PIX4993_IN
port 5065 n
rlabel metal5 51520 -92480 51620 -92380 1 PIX4994_IN
port 5066 n
rlabel metal5 53020 -92480 53120 -92380 1 PIX4995_IN
port 5067 n
rlabel metal5 54520 -92480 54620 -92380 1 PIX4996_IN
port 5068 n
rlabel metal5 56020 -92480 56120 -92380 1 PIX4997_IN
port 5069 n
rlabel metal5 57520 -92480 57620 -92380 1 PIX4998_IN
port 5070 n
rlabel metal5 59020 -92480 59120 -92380 1 PIX4999_IN
port 5071 n
rlabel metal5 60520 -92480 60620 -92380 1 PIX5000_IN
port 5072 n
rlabel metal5 62020 -92480 62120 -92380 1 PIX5001_IN
port 5073 n
rlabel metal5 63520 -92480 63620 -92380 1 PIX5002_IN
port 5074 n
rlabel metal5 65020 -92480 65120 -92380 1 PIX5003_IN
port 5075 n
rlabel metal5 66520 -92480 66620 -92380 1 PIX5004_IN
port 5076 n
rlabel metal5 68020 -92480 68120 -92380 1 PIX5005_IN
port 5077 n
rlabel metal5 69520 -92480 69620 -92380 1 PIX5006_IN
port 5078 n
rlabel metal5 71020 -92480 71120 -92380 1 PIX5007_IN
port 5079 n
rlabel metal5 72520 -92480 72620 -92380 1 PIX5008_IN
port 5080 n
rlabel metal5 74020 -92480 74120 -92380 1 PIX5009_IN
port 5081 n
rlabel metal5 75520 -92480 75620 -92380 1 PIX5010_IN
port 5082 n
rlabel metal5 77020 -92480 77120 -92380 1 PIX5011_IN
port 5083 n
rlabel metal5 78520 -92480 78620 -92380 1 PIX5012_IN
port 5084 n
rlabel metal5 80020 -92480 80120 -92380 1 PIX5013_IN
port 5085 n
rlabel metal5 81520 -92480 81620 -92380 1 PIX5014_IN
port 5086 n
rlabel metal5 83020 -92480 83120 -92380 1 PIX5015_IN
port 5087 n
rlabel metal5 84520 -92480 84620 -92380 1 PIX5016_IN
port 5088 n
rlabel metal5 86020 -92480 86120 -92380 1 PIX5017_IN
port 5089 n
rlabel metal5 87520 -92480 87620 -92380 1 PIX5018_IN
port 5090 n
rlabel metal5 89020 -92480 89120 -92380 1 PIX5019_IN
port 5091 n
rlabel metal5 90520 -92480 90620 -92380 1 PIX5020_IN
port 5092 n
rlabel metal5 92020 -92480 92120 -92380 1 PIX5021_IN
port 5093 n
rlabel metal5 93520 -92480 93620 -92380 1 PIX5022_IN
port 5094 n
rlabel metal5 95020 -92480 95120 -92380 1 PIX5023_IN
port 5095 n
rlabel metal5 96520 -92480 96620 -92380 1 PIX5024_IN
port 5096 n
rlabel metal5 98020 -92480 98120 -92380 1 PIX5025_IN
port 5097 n
rlabel metal5 99520 -92480 99620 -92380 1 PIX5026_IN
port 5098 n
rlabel metal5 101020 -92480 101120 -92380 1 PIX5027_IN
port 5099 n
rlabel metal5 102520 -92480 102620 -92380 1 PIX5028_IN
port 5100 n
rlabel metal5 104020 -92480 104120 -92380 1 PIX5029_IN
port 5101 n
rlabel metal5 105520 -92480 105620 -92380 1 PIX5030_IN
port 5102 n
rlabel metal5 107020 -92480 107120 -92380 1 PIX5031_IN
port 5103 n
rlabel metal5 108520 -92480 108620 -92380 1 PIX5032_IN
port 5104 n
rlabel metal5 110020 -92480 110120 -92380 1 PIX5033_IN
port 5105 n
rlabel metal5 111520 -92480 111620 -92380 1 PIX5034_IN
port 5106 n
rlabel metal5 113020 -92480 113120 -92380 1 PIX5035_IN
port 5107 n
rlabel metal5 114520 -92480 114620 -92380 1 PIX5036_IN
port 5108 n
rlabel metal5 116020 -92480 116120 -92380 1 PIX5037_IN
port 5109 n
rlabel metal5 117520 -92480 117620 -92380 1 PIX5038_IN
port 5110 n
rlabel metal5 119020 -92480 119120 -92380 1 PIX5039_IN
port 5111 n
rlabel metal5 520 -93980 620 -93880 1 PIX5040_IN
port 5112 n
rlabel metal2 -1500 -93760 -1500 -93715 3 ROW_SEL63
port 5113 e
rlabel metal5 2020 -93980 2120 -93880 1 PIX5041_IN
port 5114 n
rlabel metal5 3520 -93980 3620 -93880 1 PIX5042_IN
port 5115 n
rlabel metal5 5020 -93980 5120 -93880 1 PIX5043_IN
port 5116 n
rlabel metal5 6520 -93980 6620 -93880 1 PIX5044_IN
port 5117 n
rlabel metal5 8020 -93980 8120 -93880 1 PIX5045_IN
port 5118 n
rlabel metal5 9520 -93980 9620 -93880 1 PIX5046_IN
port 5119 n
rlabel metal5 11020 -93980 11120 -93880 1 PIX5047_IN
port 5120 n
rlabel metal5 12520 -93980 12620 -93880 1 PIX5048_IN
port 5121 n
rlabel metal5 14020 -93980 14120 -93880 1 PIX5049_IN
port 5122 n
rlabel metal5 15520 -93980 15620 -93880 1 PIX5050_IN
port 5123 n
rlabel metal5 17020 -93980 17120 -93880 1 PIX5051_IN
port 5124 n
rlabel metal5 18520 -93980 18620 -93880 1 PIX5052_IN
port 5125 n
rlabel metal5 20020 -93980 20120 -93880 1 PIX5053_IN
port 5126 n
rlabel metal5 21520 -93980 21620 -93880 1 PIX5054_IN
port 5127 n
rlabel metal5 23020 -93980 23120 -93880 1 PIX5055_IN
port 5128 n
rlabel metal5 24520 -93980 24620 -93880 1 PIX5056_IN
port 5129 n
rlabel metal5 26020 -93980 26120 -93880 1 PIX5057_IN
port 5130 n
rlabel metal5 27520 -93980 27620 -93880 1 PIX5058_IN
port 5131 n
rlabel metal5 29020 -93980 29120 -93880 1 PIX5059_IN
port 5132 n
rlabel metal5 30520 -93980 30620 -93880 1 PIX5060_IN
port 5133 n
rlabel metal5 32020 -93980 32120 -93880 1 PIX5061_IN
port 5134 n
rlabel metal5 33520 -93980 33620 -93880 1 PIX5062_IN
port 5135 n
rlabel metal5 35020 -93980 35120 -93880 1 PIX5063_IN
port 5136 n
rlabel metal5 36520 -93980 36620 -93880 1 PIX5064_IN
port 5137 n
rlabel metal5 38020 -93980 38120 -93880 1 PIX5065_IN
port 5138 n
rlabel metal5 39520 -93980 39620 -93880 1 PIX5066_IN
port 5139 n
rlabel metal5 41020 -93980 41120 -93880 1 PIX5067_IN
port 5140 n
rlabel metal5 42520 -93980 42620 -93880 1 PIX5068_IN
port 5141 n
rlabel metal5 44020 -93980 44120 -93880 1 PIX5069_IN
port 5142 n
rlabel metal5 45520 -93980 45620 -93880 1 PIX5070_IN
port 5143 n
rlabel metal5 47020 -93980 47120 -93880 1 PIX5071_IN
port 5144 n
rlabel metal5 48520 -93980 48620 -93880 1 PIX5072_IN
port 5145 n
rlabel metal5 50020 -93980 50120 -93880 1 PIX5073_IN
port 5146 n
rlabel metal5 51520 -93980 51620 -93880 1 PIX5074_IN
port 5147 n
rlabel metal5 53020 -93980 53120 -93880 1 PIX5075_IN
port 5148 n
rlabel metal5 54520 -93980 54620 -93880 1 PIX5076_IN
port 5149 n
rlabel metal5 56020 -93980 56120 -93880 1 PIX5077_IN
port 5150 n
rlabel metal5 57520 -93980 57620 -93880 1 PIX5078_IN
port 5151 n
rlabel metal5 59020 -93980 59120 -93880 1 PIX5079_IN
port 5152 n
rlabel metal5 60520 -93980 60620 -93880 1 PIX5080_IN
port 5153 n
rlabel metal5 62020 -93980 62120 -93880 1 PIX5081_IN
port 5154 n
rlabel metal5 63520 -93980 63620 -93880 1 PIX5082_IN
port 5155 n
rlabel metal5 65020 -93980 65120 -93880 1 PIX5083_IN
port 5156 n
rlabel metal5 66520 -93980 66620 -93880 1 PIX5084_IN
port 5157 n
rlabel metal5 68020 -93980 68120 -93880 1 PIX5085_IN
port 5158 n
rlabel metal5 69520 -93980 69620 -93880 1 PIX5086_IN
port 5159 n
rlabel metal5 71020 -93980 71120 -93880 1 PIX5087_IN
port 5160 n
rlabel metal5 72520 -93980 72620 -93880 1 PIX5088_IN
port 5161 n
rlabel metal5 74020 -93980 74120 -93880 1 PIX5089_IN
port 5162 n
rlabel metal5 75520 -93980 75620 -93880 1 PIX5090_IN
port 5163 n
rlabel metal5 77020 -93980 77120 -93880 1 PIX5091_IN
port 5164 n
rlabel metal5 78520 -93980 78620 -93880 1 PIX5092_IN
port 5165 n
rlabel metal5 80020 -93980 80120 -93880 1 PIX5093_IN
port 5166 n
rlabel metal5 81520 -93980 81620 -93880 1 PIX5094_IN
port 5167 n
rlabel metal5 83020 -93980 83120 -93880 1 PIX5095_IN
port 5168 n
rlabel metal5 84520 -93980 84620 -93880 1 PIX5096_IN
port 5169 n
rlabel metal5 86020 -93980 86120 -93880 1 PIX5097_IN
port 5170 n
rlabel metal5 87520 -93980 87620 -93880 1 PIX5098_IN
port 5171 n
rlabel metal5 89020 -93980 89120 -93880 1 PIX5099_IN
port 5172 n
rlabel metal5 90520 -93980 90620 -93880 1 PIX5100_IN
port 5173 n
rlabel metal5 92020 -93980 92120 -93880 1 PIX5101_IN
port 5174 n
rlabel metal5 93520 -93980 93620 -93880 1 PIX5102_IN
port 5175 n
rlabel metal5 95020 -93980 95120 -93880 1 PIX5103_IN
port 5176 n
rlabel metal5 96520 -93980 96620 -93880 1 PIX5104_IN
port 5177 n
rlabel metal5 98020 -93980 98120 -93880 1 PIX5105_IN
port 5178 n
rlabel metal5 99520 -93980 99620 -93880 1 PIX5106_IN
port 5179 n
rlabel metal5 101020 -93980 101120 -93880 1 PIX5107_IN
port 5180 n
rlabel metal5 102520 -93980 102620 -93880 1 PIX5108_IN
port 5181 n
rlabel metal5 104020 -93980 104120 -93880 1 PIX5109_IN
port 5182 n
rlabel metal5 105520 -93980 105620 -93880 1 PIX5110_IN
port 5183 n
rlabel metal5 107020 -93980 107120 -93880 1 PIX5111_IN
port 5184 n
rlabel metal5 108520 -93980 108620 -93880 1 PIX5112_IN
port 5185 n
rlabel metal5 110020 -93980 110120 -93880 1 PIX5113_IN
port 5186 n
rlabel metal5 111520 -93980 111620 -93880 1 PIX5114_IN
port 5187 n
rlabel metal5 113020 -93980 113120 -93880 1 PIX5115_IN
port 5188 n
rlabel metal5 114520 -93980 114620 -93880 1 PIX5116_IN
port 5189 n
rlabel metal5 116020 -93980 116120 -93880 1 PIX5117_IN
port 5190 n
rlabel metal5 117520 -93980 117620 -93880 1 PIX5118_IN
port 5191 n
rlabel metal5 119020 -93980 119120 -93880 1 PIX5119_IN
port 5192 n
rlabel metal5 520 -95480 620 -95380 1 PIX5120_IN
port 5193 n
rlabel metal2 -1500 -95260 -1500 -95215 3 ROW_SEL64
port 5194 e
rlabel metal5 2020 -95480 2120 -95380 1 PIX5121_IN
port 5195 n
rlabel metal5 3520 -95480 3620 -95380 1 PIX5122_IN
port 5196 n
rlabel metal5 5020 -95480 5120 -95380 1 PIX5123_IN
port 5197 n
rlabel metal5 6520 -95480 6620 -95380 1 PIX5124_IN
port 5198 n
rlabel metal5 8020 -95480 8120 -95380 1 PIX5125_IN
port 5199 n
rlabel metal5 9520 -95480 9620 -95380 1 PIX5126_IN
port 5200 n
rlabel metal5 11020 -95480 11120 -95380 1 PIX5127_IN
port 5201 n
rlabel metal5 12520 -95480 12620 -95380 1 PIX5128_IN
port 5202 n
rlabel metal5 14020 -95480 14120 -95380 1 PIX5129_IN
port 5203 n
rlabel metal5 15520 -95480 15620 -95380 1 PIX5130_IN
port 5204 n
rlabel metal5 17020 -95480 17120 -95380 1 PIX5131_IN
port 5205 n
rlabel metal5 18520 -95480 18620 -95380 1 PIX5132_IN
port 5206 n
rlabel metal5 20020 -95480 20120 -95380 1 PIX5133_IN
port 5207 n
rlabel metal5 21520 -95480 21620 -95380 1 PIX5134_IN
port 5208 n
rlabel metal5 23020 -95480 23120 -95380 1 PIX5135_IN
port 5209 n
rlabel metal5 24520 -95480 24620 -95380 1 PIX5136_IN
port 5210 n
rlabel metal5 26020 -95480 26120 -95380 1 PIX5137_IN
port 5211 n
rlabel metal5 27520 -95480 27620 -95380 1 PIX5138_IN
port 5212 n
rlabel metal5 29020 -95480 29120 -95380 1 PIX5139_IN
port 5213 n
rlabel metal5 30520 -95480 30620 -95380 1 PIX5140_IN
port 5214 n
rlabel metal5 32020 -95480 32120 -95380 1 PIX5141_IN
port 5215 n
rlabel metal5 33520 -95480 33620 -95380 1 PIX5142_IN
port 5216 n
rlabel metal5 35020 -95480 35120 -95380 1 PIX5143_IN
port 5217 n
rlabel metal5 36520 -95480 36620 -95380 1 PIX5144_IN
port 5218 n
rlabel metal5 38020 -95480 38120 -95380 1 PIX5145_IN
port 5219 n
rlabel metal5 39520 -95480 39620 -95380 1 PIX5146_IN
port 5220 n
rlabel metal5 41020 -95480 41120 -95380 1 PIX5147_IN
port 5221 n
rlabel metal5 42520 -95480 42620 -95380 1 PIX5148_IN
port 5222 n
rlabel metal5 44020 -95480 44120 -95380 1 PIX5149_IN
port 5223 n
rlabel metal5 45520 -95480 45620 -95380 1 PIX5150_IN
port 5224 n
rlabel metal5 47020 -95480 47120 -95380 1 PIX5151_IN
port 5225 n
rlabel metal5 48520 -95480 48620 -95380 1 PIX5152_IN
port 5226 n
rlabel metal5 50020 -95480 50120 -95380 1 PIX5153_IN
port 5227 n
rlabel metal5 51520 -95480 51620 -95380 1 PIX5154_IN
port 5228 n
rlabel metal5 53020 -95480 53120 -95380 1 PIX5155_IN
port 5229 n
rlabel metal5 54520 -95480 54620 -95380 1 PIX5156_IN
port 5230 n
rlabel metal5 56020 -95480 56120 -95380 1 PIX5157_IN
port 5231 n
rlabel metal5 57520 -95480 57620 -95380 1 PIX5158_IN
port 5232 n
rlabel metal5 59020 -95480 59120 -95380 1 PIX5159_IN
port 5233 n
rlabel metal5 60520 -95480 60620 -95380 1 PIX5160_IN
port 5234 n
rlabel metal5 62020 -95480 62120 -95380 1 PIX5161_IN
port 5235 n
rlabel metal5 63520 -95480 63620 -95380 1 PIX5162_IN
port 5236 n
rlabel metal5 65020 -95480 65120 -95380 1 PIX5163_IN
port 5237 n
rlabel metal5 66520 -95480 66620 -95380 1 PIX5164_IN
port 5238 n
rlabel metal5 68020 -95480 68120 -95380 1 PIX5165_IN
port 5239 n
rlabel metal5 69520 -95480 69620 -95380 1 PIX5166_IN
port 5240 n
rlabel metal5 71020 -95480 71120 -95380 1 PIX5167_IN
port 5241 n
rlabel metal5 72520 -95480 72620 -95380 1 PIX5168_IN
port 5242 n
rlabel metal5 74020 -95480 74120 -95380 1 PIX5169_IN
port 5243 n
rlabel metal5 75520 -95480 75620 -95380 1 PIX5170_IN
port 5244 n
rlabel metal5 77020 -95480 77120 -95380 1 PIX5171_IN
port 5245 n
rlabel metal5 78520 -95480 78620 -95380 1 PIX5172_IN
port 5246 n
rlabel metal5 80020 -95480 80120 -95380 1 PIX5173_IN
port 5247 n
rlabel metal5 81520 -95480 81620 -95380 1 PIX5174_IN
port 5248 n
rlabel metal5 83020 -95480 83120 -95380 1 PIX5175_IN
port 5249 n
rlabel metal5 84520 -95480 84620 -95380 1 PIX5176_IN
port 5250 n
rlabel metal5 86020 -95480 86120 -95380 1 PIX5177_IN
port 5251 n
rlabel metal5 87520 -95480 87620 -95380 1 PIX5178_IN
port 5252 n
rlabel metal5 89020 -95480 89120 -95380 1 PIX5179_IN
port 5253 n
rlabel metal5 90520 -95480 90620 -95380 1 PIX5180_IN
port 5254 n
rlabel metal5 92020 -95480 92120 -95380 1 PIX5181_IN
port 5255 n
rlabel metal5 93520 -95480 93620 -95380 1 PIX5182_IN
port 5256 n
rlabel metal5 95020 -95480 95120 -95380 1 PIX5183_IN
port 5257 n
rlabel metal5 96520 -95480 96620 -95380 1 PIX5184_IN
port 5258 n
rlabel metal5 98020 -95480 98120 -95380 1 PIX5185_IN
port 5259 n
rlabel metal5 99520 -95480 99620 -95380 1 PIX5186_IN
port 5260 n
rlabel metal5 101020 -95480 101120 -95380 1 PIX5187_IN
port 5261 n
rlabel metal5 102520 -95480 102620 -95380 1 PIX5188_IN
port 5262 n
rlabel metal5 104020 -95480 104120 -95380 1 PIX5189_IN
port 5263 n
rlabel metal5 105520 -95480 105620 -95380 1 PIX5190_IN
port 5264 n
rlabel metal5 107020 -95480 107120 -95380 1 PIX5191_IN
port 5265 n
rlabel metal5 108520 -95480 108620 -95380 1 PIX5192_IN
port 5266 n
rlabel metal5 110020 -95480 110120 -95380 1 PIX5193_IN
port 5267 n
rlabel metal5 111520 -95480 111620 -95380 1 PIX5194_IN
port 5268 n
rlabel metal5 113020 -95480 113120 -95380 1 PIX5195_IN
port 5269 n
rlabel metal5 114520 -95480 114620 -95380 1 PIX5196_IN
port 5270 n
rlabel metal5 116020 -95480 116120 -95380 1 PIX5197_IN
port 5271 n
rlabel metal5 117520 -95480 117620 -95380 1 PIX5198_IN
port 5272 n
rlabel metal5 119020 -95480 119120 -95380 1 PIX5199_IN
port 5273 n
rlabel metal5 520 -96980 620 -96880 1 PIX5200_IN
port 5274 n
rlabel metal2 -1500 -96760 -1500 -96715 3 ROW_SEL65
port 5275 e
rlabel metal5 2020 -96980 2120 -96880 1 PIX5201_IN
port 5276 n
rlabel metal5 3520 -96980 3620 -96880 1 PIX5202_IN
port 5277 n
rlabel metal5 5020 -96980 5120 -96880 1 PIX5203_IN
port 5278 n
rlabel metal5 6520 -96980 6620 -96880 1 PIX5204_IN
port 5279 n
rlabel metal5 8020 -96980 8120 -96880 1 PIX5205_IN
port 5280 n
rlabel metal5 9520 -96980 9620 -96880 1 PIX5206_IN
port 5281 n
rlabel metal5 11020 -96980 11120 -96880 1 PIX5207_IN
port 5282 n
rlabel metal5 12520 -96980 12620 -96880 1 PIX5208_IN
port 5283 n
rlabel metal5 14020 -96980 14120 -96880 1 PIX5209_IN
port 5284 n
rlabel metal5 15520 -96980 15620 -96880 1 PIX5210_IN
port 5285 n
rlabel metal5 17020 -96980 17120 -96880 1 PIX5211_IN
port 5286 n
rlabel metal5 18520 -96980 18620 -96880 1 PIX5212_IN
port 5287 n
rlabel metal5 20020 -96980 20120 -96880 1 PIX5213_IN
port 5288 n
rlabel metal5 21520 -96980 21620 -96880 1 PIX5214_IN
port 5289 n
rlabel metal5 23020 -96980 23120 -96880 1 PIX5215_IN
port 5290 n
rlabel metal5 24520 -96980 24620 -96880 1 PIX5216_IN
port 5291 n
rlabel metal5 26020 -96980 26120 -96880 1 PIX5217_IN
port 5292 n
rlabel metal5 27520 -96980 27620 -96880 1 PIX5218_IN
port 5293 n
rlabel metal5 29020 -96980 29120 -96880 1 PIX5219_IN
port 5294 n
rlabel metal5 30520 -96980 30620 -96880 1 PIX5220_IN
port 5295 n
rlabel metal5 32020 -96980 32120 -96880 1 PIX5221_IN
port 5296 n
rlabel metal5 33520 -96980 33620 -96880 1 PIX5222_IN
port 5297 n
rlabel metal5 35020 -96980 35120 -96880 1 PIX5223_IN
port 5298 n
rlabel metal5 36520 -96980 36620 -96880 1 PIX5224_IN
port 5299 n
rlabel metal5 38020 -96980 38120 -96880 1 PIX5225_IN
port 5300 n
rlabel metal5 39520 -96980 39620 -96880 1 PIX5226_IN
port 5301 n
rlabel metal5 41020 -96980 41120 -96880 1 PIX5227_IN
port 5302 n
rlabel metal5 42520 -96980 42620 -96880 1 PIX5228_IN
port 5303 n
rlabel metal5 44020 -96980 44120 -96880 1 PIX5229_IN
port 5304 n
rlabel metal5 45520 -96980 45620 -96880 1 PIX5230_IN
port 5305 n
rlabel metal5 47020 -96980 47120 -96880 1 PIX5231_IN
port 5306 n
rlabel metal5 48520 -96980 48620 -96880 1 PIX5232_IN
port 5307 n
rlabel metal5 50020 -96980 50120 -96880 1 PIX5233_IN
port 5308 n
rlabel metal5 51520 -96980 51620 -96880 1 PIX5234_IN
port 5309 n
rlabel metal5 53020 -96980 53120 -96880 1 PIX5235_IN
port 5310 n
rlabel metal5 54520 -96980 54620 -96880 1 PIX5236_IN
port 5311 n
rlabel metal5 56020 -96980 56120 -96880 1 PIX5237_IN
port 5312 n
rlabel metal5 57520 -96980 57620 -96880 1 PIX5238_IN
port 5313 n
rlabel metal5 59020 -96980 59120 -96880 1 PIX5239_IN
port 5314 n
rlabel metal5 60520 -96980 60620 -96880 1 PIX5240_IN
port 5315 n
rlabel metal5 62020 -96980 62120 -96880 1 PIX5241_IN
port 5316 n
rlabel metal5 63520 -96980 63620 -96880 1 PIX5242_IN
port 5317 n
rlabel metal5 65020 -96980 65120 -96880 1 PIX5243_IN
port 5318 n
rlabel metal5 66520 -96980 66620 -96880 1 PIX5244_IN
port 5319 n
rlabel metal5 68020 -96980 68120 -96880 1 PIX5245_IN
port 5320 n
rlabel metal5 69520 -96980 69620 -96880 1 PIX5246_IN
port 5321 n
rlabel metal5 71020 -96980 71120 -96880 1 PIX5247_IN
port 5322 n
rlabel metal5 72520 -96980 72620 -96880 1 PIX5248_IN
port 5323 n
rlabel metal5 74020 -96980 74120 -96880 1 PIX5249_IN
port 5324 n
rlabel metal5 75520 -96980 75620 -96880 1 PIX5250_IN
port 5325 n
rlabel metal5 77020 -96980 77120 -96880 1 PIX5251_IN
port 5326 n
rlabel metal5 78520 -96980 78620 -96880 1 PIX5252_IN
port 5327 n
rlabel metal5 80020 -96980 80120 -96880 1 PIX5253_IN
port 5328 n
rlabel metal5 81520 -96980 81620 -96880 1 PIX5254_IN
port 5329 n
rlabel metal5 83020 -96980 83120 -96880 1 PIX5255_IN
port 5330 n
rlabel metal5 84520 -96980 84620 -96880 1 PIX5256_IN
port 5331 n
rlabel metal5 86020 -96980 86120 -96880 1 PIX5257_IN
port 5332 n
rlabel metal5 87520 -96980 87620 -96880 1 PIX5258_IN
port 5333 n
rlabel metal5 89020 -96980 89120 -96880 1 PIX5259_IN
port 5334 n
rlabel metal5 90520 -96980 90620 -96880 1 PIX5260_IN
port 5335 n
rlabel metal5 92020 -96980 92120 -96880 1 PIX5261_IN
port 5336 n
rlabel metal5 93520 -96980 93620 -96880 1 PIX5262_IN
port 5337 n
rlabel metal5 95020 -96980 95120 -96880 1 PIX5263_IN
port 5338 n
rlabel metal5 96520 -96980 96620 -96880 1 PIX5264_IN
port 5339 n
rlabel metal5 98020 -96980 98120 -96880 1 PIX5265_IN
port 5340 n
rlabel metal5 99520 -96980 99620 -96880 1 PIX5266_IN
port 5341 n
rlabel metal5 101020 -96980 101120 -96880 1 PIX5267_IN
port 5342 n
rlabel metal5 102520 -96980 102620 -96880 1 PIX5268_IN
port 5343 n
rlabel metal5 104020 -96980 104120 -96880 1 PIX5269_IN
port 5344 n
rlabel metal5 105520 -96980 105620 -96880 1 PIX5270_IN
port 5345 n
rlabel metal5 107020 -96980 107120 -96880 1 PIX5271_IN
port 5346 n
rlabel metal5 108520 -96980 108620 -96880 1 PIX5272_IN
port 5347 n
rlabel metal5 110020 -96980 110120 -96880 1 PIX5273_IN
port 5348 n
rlabel metal5 111520 -96980 111620 -96880 1 PIX5274_IN
port 5349 n
rlabel metal5 113020 -96980 113120 -96880 1 PIX5275_IN
port 5350 n
rlabel metal5 114520 -96980 114620 -96880 1 PIX5276_IN
port 5351 n
rlabel metal5 116020 -96980 116120 -96880 1 PIX5277_IN
port 5352 n
rlabel metal5 117520 -96980 117620 -96880 1 PIX5278_IN
port 5353 n
rlabel metal5 119020 -96980 119120 -96880 1 PIX5279_IN
port 5354 n
rlabel metal5 520 -98480 620 -98380 1 PIX5280_IN
port 5355 n
rlabel metal2 -1500 -98260 -1500 -98215 3 ROW_SEL66
port 5356 e
rlabel metal5 2020 -98480 2120 -98380 1 PIX5281_IN
port 5357 n
rlabel metal5 3520 -98480 3620 -98380 1 PIX5282_IN
port 5358 n
rlabel metal5 5020 -98480 5120 -98380 1 PIX5283_IN
port 5359 n
rlabel metal5 6520 -98480 6620 -98380 1 PIX5284_IN
port 5360 n
rlabel metal5 8020 -98480 8120 -98380 1 PIX5285_IN
port 5361 n
rlabel metal5 9520 -98480 9620 -98380 1 PIX5286_IN
port 5362 n
rlabel metal5 11020 -98480 11120 -98380 1 PIX5287_IN
port 5363 n
rlabel metal5 12520 -98480 12620 -98380 1 PIX5288_IN
port 5364 n
rlabel metal5 14020 -98480 14120 -98380 1 PIX5289_IN
port 5365 n
rlabel metal5 15520 -98480 15620 -98380 1 PIX5290_IN
port 5366 n
rlabel metal5 17020 -98480 17120 -98380 1 PIX5291_IN
port 5367 n
rlabel metal5 18520 -98480 18620 -98380 1 PIX5292_IN
port 5368 n
rlabel metal5 20020 -98480 20120 -98380 1 PIX5293_IN
port 5369 n
rlabel metal5 21520 -98480 21620 -98380 1 PIX5294_IN
port 5370 n
rlabel metal5 23020 -98480 23120 -98380 1 PIX5295_IN
port 5371 n
rlabel metal5 24520 -98480 24620 -98380 1 PIX5296_IN
port 5372 n
rlabel metal5 26020 -98480 26120 -98380 1 PIX5297_IN
port 5373 n
rlabel metal5 27520 -98480 27620 -98380 1 PIX5298_IN
port 5374 n
rlabel metal5 29020 -98480 29120 -98380 1 PIX5299_IN
port 5375 n
rlabel metal5 30520 -98480 30620 -98380 1 PIX5300_IN
port 5376 n
rlabel metal5 32020 -98480 32120 -98380 1 PIX5301_IN
port 5377 n
rlabel metal5 33520 -98480 33620 -98380 1 PIX5302_IN
port 5378 n
rlabel metal5 35020 -98480 35120 -98380 1 PIX5303_IN
port 5379 n
rlabel metal5 36520 -98480 36620 -98380 1 PIX5304_IN
port 5380 n
rlabel metal5 38020 -98480 38120 -98380 1 PIX5305_IN
port 5381 n
rlabel metal5 39520 -98480 39620 -98380 1 PIX5306_IN
port 5382 n
rlabel metal5 41020 -98480 41120 -98380 1 PIX5307_IN
port 5383 n
rlabel metal5 42520 -98480 42620 -98380 1 PIX5308_IN
port 5384 n
rlabel metal5 44020 -98480 44120 -98380 1 PIX5309_IN
port 5385 n
rlabel metal5 45520 -98480 45620 -98380 1 PIX5310_IN
port 5386 n
rlabel metal5 47020 -98480 47120 -98380 1 PIX5311_IN
port 5387 n
rlabel metal5 48520 -98480 48620 -98380 1 PIX5312_IN
port 5388 n
rlabel metal5 50020 -98480 50120 -98380 1 PIX5313_IN
port 5389 n
rlabel metal5 51520 -98480 51620 -98380 1 PIX5314_IN
port 5390 n
rlabel metal5 53020 -98480 53120 -98380 1 PIX5315_IN
port 5391 n
rlabel metal5 54520 -98480 54620 -98380 1 PIX5316_IN
port 5392 n
rlabel metal5 56020 -98480 56120 -98380 1 PIX5317_IN
port 5393 n
rlabel metal5 57520 -98480 57620 -98380 1 PIX5318_IN
port 5394 n
rlabel metal5 59020 -98480 59120 -98380 1 PIX5319_IN
port 5395 n
rlabel metal5 60520 -98480 60620 -98380 1 PIX5320_IN
port 5396 n
rlabel metal5 62020 -98480 62120 -98380 1 PIX5321_IN
port 5397 n
rlabel metal5 63520 -98480 63620 -98380 1 PIX5322_IN
port 5398 n
rlabel metal5 65020 -98480 65120 -98380 1 PIX5323_IN
port 5399 n
rlabel metal5 66520 -98480 66620 -98380 1 PIX5324_IN
port 5400 n
rlabel metal5 68020 -98480 68120 -98380 1 PIX5325_IN
port 5401 n
rlabel metal5 69520 -98480 69620 -98380 1 PIX5326_IN
port 5402 n
rlabel metal5 71020 -98480 71120 -98380 1 PIX5327_IN
port 5403 n
rlabel metal5 72520 -98480 72620 -98380 1 PIX5328_IN
port 5404 n
rlabel metal5 74020 -98480 74120 -98380 1 PIX5329_IN
port 5405 n
rlabel metal5 75520 -98480 75620 -98380 1 PIX5330_IN
port 5406 n
rlabel metal5 77020 -98480 77120 -98380 1 PIX5331_IN
port 5407 n
rlabel metal5 78520 -98480 78620 -98380 1 PIX5332_IN
port 5408 n
rlabel metal5 80020 -98480 80120 -98380 1 PIX5333_IN
port 5409 n
rlabel metal5 81520 -98480 81620 -98380 1 PIX5334_IN
port 5410 n
rlabel metal5 83020 -98480 83120 -98380 1 PIX5335_IN
port 5411 n
rlabel metal5 84520 -98480 84620 -98380 1 PIX5336_IN
port 5412 n
rlabel metal5 86020 -98480 86120 -98380 1 PIX5337_IN
port 5413 n
rlabel metal5 87520 -98480 87620 -98380 1 PIX5338_IN
port 5414 n
rlabel metal5 89020 -98480 89120 -98380 1 PIX5339_IN
port 5415 n
rlabel metal5 90520 -98480 90620 -98380 1 PIX5340_IN
port 5416 n
rlabel metal5 92020 -98480 92120 -98380 1 PIX5341_IN
port 5417 n
rlabel metal5 93520 -98480 93620 -98380 1 PIX5342_IN
port 5418 n
rlabel metal5 95020 -98480 95120 -98380 1 PIX5343_IN
port 5419 n
rlabel metal5 96520 -98480 96620 -98380 1 PIX5344_IN
port 5420 n
rlabel metal5 98020 -98480 98120 -98380 1 PIX5345_IN
port 5421 n
rlabel metal5 99520 -98480 99620 -98380 1 PIX5346_IN
port 5422 n
rlabel metal5 101020 -98480 101120 -98380 1 PIX5347_IN
port 5423 n
rlabel metal5 102520 -98480 102620 -98380 1 PIX5348_IN
port 5424 n
rlabel metal5 104020 -98480 104120 -98380 1 PIX5349_IN
port 5425 n
rlabel metal5 105520 -98480 105620 -98380 1 PIX5350_IN
port 5426 n
rlabel metal5 107020 -98480 107120 -98380 1 PIX5351_IN
port 5427 n
rlabel metal5 108520 -98480 108620 -98380 1 PIX5352_IN
port 5428 n
rlabel metal5 110020 -98480 110120 -98380 1 PIX5353_IN
port 5429 n
rlabel metal5 111520 -98480 111620 -98380 1 PIX5354_IN
port 5430 n
rlabel metal5 113020 -98480 113120 -98380 1 PIX5355_IN
port 5431 n
rlabel metal5 114520 -98480 114620 -98380 1 PIX5356_IN
port 5432 n
rlabel metal5 116020 -98480 116120 -98380 1 PIX5357_IN
port 5433 n
rlabel metal5 117520 -98480 117620 -98380 1 PIX5358_IN
port 5434 n
rlabel metal5 119020 -98480 119120 -98380 1 PIX5359_IN
port 5435 n
rlabel metal5 520 -99980 620 -99880 1 PIX5360_IN
port 5436 n
rlabel metal2 -1500 -99760 -1500 -99715 3 ROW_SEL67
port 5437 e
rlabel metal5 2020 -99980 2120 -99880 1 PIX5361_IN
port 5438 n
rlabel metal5 3520 -99980 3620 -99880 1 PIX5362_IN
port 5439 n
rlabel metal5 5020 -99980 5120 -99880 1 PIX5363_IN
port 5440 n
rlabel metal5 6520 -99980 6620 -99880 1 PIX5364_IN
port 5441 n
rlabel metal5 8020 -99980 8120 -99880 1 PIX5365_IN
port 5442 n
rlabel metal5 9520 -99980 9620 -99880 1 PIX5366_IN
port 5443 n
rlabel metal5 11020 -99980 11120 -99880 1 PIX5367_IN
port 5444 n
rlabel metal5 12520 -99980 12620 -99880 1 PIX5368_IN
port 5445 n
rlabel metal5 14020 -99980 14120 -99880 1 PIX5369_IN
port 5446 n
rlabel metal5 15520 -99980 15620 -99880 1 PIX5370_IN
port 5447 n
rlabel metal5 17020 -99980 17120 -99880 1 PIX5371_IN
port 5448 n
rlabel metal5 18520 -99980 18620 -99880 1 PIX5372_IN
port 5449 n
rlabel metal5 20020 -99980 20120 -99880 1 PIX5373_IN
port 5450 n
rlabel metal5 21520 -99980 21620 -99880 1 PIX5374_IN
port 5451 n
rlabel metal5 23020 -99980 23120 -99880 1 PIX5375_IN
port 5452 n
rlabel metal5 24520 -99980 24620 -99880 1 PIX5376_IN
port 5453 n
rlabel metal5 26020 -99980 26120 -99880 1 PIX5377_IN
port 5454 n
rlabel metal5 27520 -99980 27620 -99880 1 PIX5378_IN
port 5455 n
rlabel metal5 29020 -99980 29120 -99880 1 PIX5379_IN
port 5456 n
rlabel metal5 30520 -99980 30620 -99880 1 PIX5380_IN
port 5457 n
rlabel metal5 32020 -99980 32120 -99880 1 PIX5381_IN
port 5458 n
rlabel metal5 33520 -99980 33620 -99880 1 PIX5382_IN
port 5459 n
rlabel metal5 35020 -99980 35120 -99880 1 PIX5383_IN
port 5460 n
rlabel metal5 36520 -99980 36620 -99880 1 PIX5384_IN
port 5461 n
rlabel metal5 38020 -99980 38120 -99880 1 PIX5385_IN
port 5462 n
rlabel metal5 39520 -99980 39620 -99880 1 PIX5386_IN
port 5463 n
rlabel metal5 41020 -99980 41120 -99880 1 PIX5387_IN
port 5464 n
rlabel metal5 42520 -99980 42620 -99880 1 PIX5388_IN
port 5465 n
rlabel metal5 44020 -99980 44120 -99880 1 PIX5389_IN
port 5466 n
rlabel metal5 45520 -99980 45620 -99880 1 PIX5390_IN
port 5467 n
rlabel metal5 47020 -99980 47120 -99880 1 PIX5391_IN
port 5468 n
rlabel metal5 48520 -99980 48620 -99880 1 PIX5392_IN
port 5469 n
rlabel metal5 50020 -99980 50120 -99880 1 PIX5393_IN
port 5470 n
rlabel metal5 51520 -99980 51620 -99880 1 PIX5394_IN
port 5471 n
rlabel metal5 53020 -99980 53120 -99880 1 PIX5395_IN
port 5472 n
rlabel metal5 54520 -99980 54620 -99880 1 PIX5396_IN
port 5473 n
rlabel metal5 56020 -99980 56120 -99880 1 PIX5397_IN
port 5474 n
rlabel metal5 57520 -99980 57620 -99880 1 PIX5398_IN
port 5475 n
rlabel metal5 59020 -99980 59120 -99880 1 PIX5399_IN
port 5476 n
rlabel metal5 60520 -99980 60620 -99880 1 PIX5400_IN
port 5477 n
rlabel metal5 62020 -99980 62120 -99880 1 PIX5401_IN
port 5478 n
rlabel metal5 63520 -99980 63620 -99880 1 PIX5402_IN
port 5479 n
rlabel metal5 65020 -99980 65120 -99880 1 PIX5403_IN
port 5480 n
rlabel metal5 66520 -99980 66620 -99880 1 PIX5404_IN
port 5481 n
rlabel metal5 68020 -99980 68120 -99880 1 PIX5405_IN
port 5482 n
rlabel metal5 69520 -99980 69620 -99880 1 PIX5406_IN
port 5483 n
rlabel metal5 71020 -99980 71120 -99880 1 PIX5407_IN
port 5484 n
rlabel metal5 72520 -99980 72620 -99880 1 PIX5408_IN
port 5485 n
rlabel metal5 74020 -99980 74120 -99880 1 PIX5409_IN
port 5486 n
rlabel metal5 75520 -99980 75620 -99880 1 PIX5410_IN
port 5487 n
rlabel metal5 77020 -99980 77120 -99880 1 PIX5411_IN
port 5488 n
rlabel metal5 78520 -99980 78620 -99880 1 PIX5412_IN
port 5489 n
rlabel metal5 80020 -99980 80120 -99880 1 PIX5413_IN
port 5490 n
rlabel metal5 81520 -99980 81620 -99880 1 PIX5414_IN
port 5491 n
rlabel metal5 83020 -99980 83120 -99880 1 PIX5415_IN
port 5492 n
rlabel metal5 84520 -99980 84620 -99880 1 PIX5416_IN
port 5493 n
rlabel metal5 86020 -99980 86120 -99880 1 PIX5417_IN
port 5494 n
rlabel metal5 87520 -99980 87620 -99880 1 PIX5418_IN
port 5495 n
rlabel metal5 89020 -99980 89120 -99880 1 PIX5419_IN
port 5496 n
rlabel metal5 90520 -99980 90620 -99880 1 PIX5420_IN
port 5497 n
rlabel metal5 92020 -99980 92120 -99880 1 PIX5421_IN
port 5498 n
rlabel metal5 93520 -99980 93620 -99880 1 PIX5422_IN
port 5499 n
rlabel metal5 95020 -99980 95120 -99880 1 PIX5423_IN
port 5500 n
rlabel metal5 96520 -99980 96620 -99880 1 PIX5424_IN
port 5501 n
rlabel metal5 98020 -99980 98120 -99880 1 PIX5425_IN
port 5502 n
rlabel metal5 99520 -99980 99620 -99880 1 PIX5426_IN
port 5503 n
rlabel metal5 101020 -99980 101120 -99880 1 PIX5427_IN
port 5504 n
rlabel metal5 102520 -99980 102620 -99880 1 PIX5428_IN
port 5505 n
rlabel metal5 104020 -99980 104120 -99880 1 PIX5429_IN
port 5506 n
rlabel metal5 105520 -99980 105620 -99880 1 PIX5430_IN
port 5507 n
rlabel metal5 107020 -99980 107120 -99880 1 PIX5431_IN
port 5508 n
rlabel metal5 108520 -99980 108620 -99880 1 PIX5432_IN
port 5509 n
rlabel metal5 110020 -99980 110120 -99880 1 PIX5433_IN
port 5510 n
rlabel metal5 111520 -99980 111620 -99880 1 PIX5434_IN
port 5511 n
rlabel metal5 113020 -99980 113120 -99880 1 PIX5435_IN
port 5512 n
rlabel metal5 114520 -99980 114620 -99880 1 PIX5436_IN
port 5513 n
rlabel metal5 116020 -99980 116120 -99880 1 PIX5437_IN
port 5514 n
rlabel metal5 117520 -99980 117620 -99880 1 PIX5438_IN
port 5515 n
rlabel metal5 119020 -99980 119120 -99880 1 PIX5439_IN
port 5516 n
rlabel metal5 520 -101480 620 -101380 1 PIX5440_IN
port 5517 n
rlabel metal2 -1500 -101260 -1500 -101215 3 ROW_SEL68
port 5518 e
rlabel metal5 2020 -101480 2120 -101380 1 PIX5441_IN
port 5519 n
rlabel metal5 3520 -101480 3620 -101380 1 PIX5442_IN
port 5520 n
rlabel metal5 5020 -101480 5120 -101380 1 PIX5443_IN
port 5521 n
rlabel metal5 6520 -101480 6620 -101380 1 PIX5444_IN
port 5522 n
rlabel metal5 8020 -101480 8120 -101380 1 PIX5445_IN
port 5523 n
rlabel metal5 9520 -101480 9620 -101380 1 PIX5446_IN
port 5524 n
rlabel metal5 11020 -101480 11120 -101380 1 PIX5447_IN
port 5525 n
rlabel metal5 12520 -101480 12620 -101380 1 PIX5448_IN
port 5526 n
rlabel metal5 14020 -101480 14120 -101380 1 PIX5449_IN
port 5527 n
rlabel metal5 15520 -101480 15620 -101380 1 PIX5450_IN
port 5528 n
rlabel metal5 17020 -101480 17120 -101380 1 PIX5451_IN
port 5529 n
rlabel metal5 18520 -101480 18620 -101380 1 PIX5452_IN
port 5530 n
rlabel metal5 20020 -101480 20120 -101380 1 PIX5453_IN
port 5531 n
rlabel metal5 21520 -101480 21620 -101380 1 PIX5454_IN
port 5532 n
rlabel metal5 23020 -101480 23120 -101380 1 PIX5455_IN
port 5533 n
rlabel metal5 24520 -101480 24620 -101380 1 PIX5456_IN
port 5534 n
rlabel metal5 26020 -101480 26120 -101380 1 PIX5457_IN
port 5535 n
rlabel metal5 27520 -101480 27620 -101380 1 PIX5458_IN
port 5536 n
rlabel metal5 29020 -101480 29120 -101380 1 PIX5459_IN
port 5537 n
rlabel metal5 30520 -101480 30620 -101380 1 PIX5460_IN
port 5538 n
rlabel metal5 32020 -101480 32120 -101380 1 PIX5461_IN
port 5539 n
rlabel metal5 33520 -101480 33620 -101380 1 PIX5462_IN
port 5540 n
rlabel metal5 35020 -101480 35120 -101380 1 PIX5463_IN
port 5541 n
rlabel metal5 36520 -101480 36620 -101380 1 PIX5464_IN
port 5542 n
rlabel metal5 38020 -101480 38120 -101380 1 PIX5465_IN
port 5543 n
rlabel metal5 39520 -101480 39620 -101380 1 PIX5466_IN
port 5544 n
rlabel metal5 41020 -101480 41120 -101380 1 PIX5467_IN
port 5545 n
rlabel metal5 42520 -101480 42620 -101380 1 PIX5468_IN
port 5546 n
rlabel metal5 44020 -101480 44120 -101380 1 PIX5469_IN
port 5547 n
rlabel metal5 45520 -101480 45620 -101380 1 PIX5470_IN
port 5548 n
rlabel metal5 47020 -101480 47120 -101380 1 PIX5471_IN
port 5549 n
rlabel metal5 48520 -101480 48620 -101380 1 PIX5472_IN
port 5550 n
rlabel metal5 50020 -101480 50120 -101380 1 PIX5473_IN
port 5551 n
rlabel metal5 51520 -101480 51620 -101380 1 PIX5474_IN
port 5552 n
rlabel metal5 53020 -101480 53120 -101380 1 PIX5475_IN
port 5553 n
rlabel metal5 54520 -101480 54620 -101380 1 PIX5476_IN
port 5554 n
rlabel metal5 56020 -101480 56120 -101380 1 PIX5477_IN
port 5555 n
rlabel metal5 57520 -101480 57620 -101380 1 PIX5478_IN
port 5556 n
rlabel metal5 59020 -101480 59120 -101380 1 PIX5479_IN
port 5557 n
rlabel metal5 60520 -101480 60620 -101380 1 PIX5480_IN
port 5558 n
rlabel metal5 62020 -101480 62120 -101380 1 PIX5481_IN
port 5559 n
rlabel metal5 63520 -101480 63620 -101380 1 PIX5482_IN
port 5560 n
rlabel metal5 65020 -101480 65120 -101380 1 PIX5483_IN
port 5561 n
rlabel metal5 66520 -101480 66620 -101380 1 PIX5484_IN
port 5562 n
rlabel metal5 68020 -101480 68120 -101380 1 PIX5485_IN
port 5563 n
rlabel metal5 69520 -101480 69620 -101380 1 PIX5486_IN
port 5564 n
rlabel metal5 71020 -101480 71120 -101380 1 PIX5487_IN
port 5565 n
rlabel metal5 72520 -101480 72620 -101380 1 PIX5488_IN
port 5566 n
rlabel metal5 74020 -101480 74120 -101380 1 PIX5489_IN
port 5567 n
rlabel metal5 75520 -101480 75620 -101380 1 PIX5490_IN
port 5568 n
rlabel metal5 77020 -101480 77120 -101380 1 PIX5491_IN
port 5569 n
rlabel metal5 78520 -101480 78620 -101380 1 PIX5492_IN
port 5570 n
rlabel metal5 80020 -101480 80120 -101380 1 PIX5493_IN
port 5571 n
rlabel metal5 81520 -101480 81620 -101380 1 PIX5494_IN
port 5572 n
rlabel metal5 83020 -101480 83120 -101380 1 PIX5495_IN
port 5573 n
rlabel metal5 84520 -101480 84620 -101380 1 PIX5496_IN
port 5574 n
rlabel metal5 86020 -101480 86120 -101380 1 PIX5497_IN
port 5575 n
rlabel metal5 87520 -101480 87620 -101380 1 PIX5498_IN
port 5576 n
rlabel metal5 89020 -101480 89120 -101380 1 PIX5499_IN
port 5577 n
rlabel metal5 90520 -101480 90620 -101380 1 PIX5500_IN
port 5578 n
rlabel metal5 92020 -101480 92120 -101380 1 PIX5501_IN
port 5579 n
rlabel metal5 93520 -101480 93620 -101380 1 PIX5502_IN
port 5580 n
rlabel metal5 95020 -101480 95120 -101380 1 PIX5503_IN
port 5581 n
rlabel metal5 96520 -101480 96620 -101380 1 PIX5504_IN
port 5582 n
rlabel metal5 98020 -101480 98120 -101380 1 PIX5505_IN
port 5583 n
rlabel metal5 99520 -101480 99620 -101380 1 PIX5506_IN
port 5584 n
rlabel metal5 101020 -101480 101120 -101380 1 PIX5507_IN
port 5585 n
rlabel metal5 102520 -101480 102620 -101380 1 PIX5508_IN
port 5586 n
rlabel metal5 104020 -101480 104120 -101380 1 PIX5509_IN
port 5587 n
rlabel metal5 105520 -101480 105620 -101380 1 PIX5510_IN
port 5588 n
rlabel metal5 107020 -101480 107120 -101380 1 PIX5511_IN
port 5589 n
rlabel metal5 108520 -101480 108620 -101380 1 PIX5512_IN
port 5590 n
rlabel metal5 110020 -101480 110120 -101380 1 PIX5513_IN
port 5591 n
rlabel metal5 111520 -101480 111620 -101380 1 PIX5514_IN
port 5592 n
rlabel metal5 113020 -101480 113120 -101380 1 PIX5515_IN
port 5593 n
rlabel metal5 114520 -101480 114620 -101380 1 PIX5516_IN
port 5594 n
rlabel metal5 116020 -101480 116120 -101380 1 PIX5517_IN
port 5595 n
rlabel metal5 117520 -101480 117620 -101380 1 PIX5518_IN
port 5596 n
rlabel metal5 119020 -101480 119120 -101380 1 PIX5519_IN
port 5597 n
rlabel metal5 520 -102980 620 -102880 1 PIX5520_IN
port 5598 n
rlabel metal2 -1500 -102760 -1500 -102715 3 ROW_SEL69
port 5599 e
rlabel metal5 2020 -102980 2120 -102880 1 PIX5521_IN
port 5600 n
rlabel metal5 3520 -102980 3620 -102880 1 PIX5522_IN
port 5601 n
rlabel metal5 5020 -102980 5120 -102880 1 PIX5523_IN
port 5602 n
rlabel metal5 6520 -102980 6620 -102880 1 PIX5524_IN
port 5603 n
rlabel metal5 8020 -102980 8120 -102880 1 PIX5525_IN
port 5604 n
rlabel metal5 9520 -102980 9620 -102880 1 PIX5526_IN
port 5605 n
rlabel metal5 11020 -102980 11120 -102880 1 PIX5527_IN
port 5606 n
rlabel metal5 12520 -102980 12620 -102880 1 PIX5528_IN
port 5607 n
rlabel metal5 14020 -102980 14120 -102880 1 PIX5529_IN
port 5608 n
rlabel metal5 15520 -102980 15620 -102880 1 PIX5530_IN
port 5609 n
rlabel metal5 17020 -102980 17120 -102880 1 PIX5531_IN
port 5610 n
rlabel metal5 18520 -102980 18620 -102880 1 PIX5532_IN
port 5611 n
rlabel metal5 20020 -102980 20120 -102880 1 PIX5533_IN
port 5612 n
rlabel metal5 21520 -102980 21620 -102880 1 PIX5534_IN
port 5613 n
rlabel metal5 23020 -102980 23120 -102880 1 PIX5535_IN
port 5614 n
rlabel metal5 24520 -102980 24620 -102880 1 PIX5536_IN
port 5615 n
rlabel metal5 26020 -102980 26120 -102880 1 PIX5537_IN
port 5616 n
rlabel metal5 27520 -102980 27620 -102880 1 PIX5538_IN
port 5617 n
rlabel metal5 29020 -102980 29120 -102880 1 PIX5539_IN
port 5618 n
rlabel metal5 30520 -102980 30620 -102880 1 PIX5540_IN
port 5619 n
rlabel metal5 32020 -102980 32120 -102880 1 PIX5541_IN
port 5620 n
rlabel metal5 33520 -102980 33620 -102880 1 PIX5542_IN
port 5621 n
rlabel metal5 35020 -102980 35120 -102880 1 PIX5543_IN
port 5622 n
rlabel metal5 36520 -102980 36620 -102880 1 PIX5544_IN
port 5623 n
rlabel metal5 38020 -102980 38120 -102880 1 PIX5545_IN
port 5624 n
rlabel metal5 39520 -102980 39620 -102880 1 PIX5546_IN
port 5625 n
rlabel metal5 41020 -102980 41120 -102880 1 PIX5547_IN
port 5626 n
rlabel metal5 42520 -102980 42620 -102880 1 PIX5548_IN
port 5627 n
rlabel metal5 44020 -102980 44120 -102880 1 PIX5549_IN
port 5628 n
rlabel metal5 45520 -102980 45620 -102880 1 PIX5550_IN
port 5629 n
rlabel metal5 47020 -102980 47120 -102880 1 PIX5551_IN
port 5630 n
rlabel metal5 48520 -102980 48620 -102880 1 PIX5552_IN
port 5631 n
rlabel metal5 50020 -102980 50120 -102880 1 PIX5553_IN
port 5632 n
rlabel metal5 51520 -102980 51620 -102880 1 PIX5554_IN
port 5633 n
rlabel metal5 53020 -102980 53120 -102880 1 PIX5555_IN
port 5634 n
rlabel metal5 54520 -102980 54620 -102880 1 PIX5556_IN
port 5635 n
rlabel metal5 56020 -102980 56120 -102880 1 PIX5557_IN
port 5636 n
rlabel metal5 57520 -102980 57620 -102880 1 PIX5558_IN
port 5637 n
rlabel metal5 59020 -102980 59120 -102880 1 PIX5559_IN
port 5638 n
rlabel metal5 60520 -102980 60620 -102880 1 PIX5560_IN
port 5639 n
rlabel metal5 62020 -102980 62120 -102880 1 PIX5561_IN
port 5640 n
rlabel metal5 63520 -102980 63620 -102880 1 PIX5562_IN
port 5641 n
rlabel metal5 65020 -102980 65120 -102880 1 PIX5563_IN
port 5642 n
rlabel metal5 66520 -102980 66620 -102880 1 PIX5564_IN
port 5643 n
rlabel metal5 68020 -102980 68120 -102880 1 PIX5565_IN
port 5644 n
rlabel metal5 69520 -102980 69620 -102880 1 PIX5566_IN
port 5645 n
rlabel metal5 71020 -102980 71120 -102880 1 PIX5567_IN
port 5646 n
rlabel metal5 72520 -102980 72620 -102880 1 PIX5568_IN
port 5647 n
rlabel metal5 74020 -102980 74120 -102880 1 PIX5569_IN
port 5648 n
rlabel metal5 75520 -102980 75620 -102880 1 PIX5570_IN
port 5649 n
rlabel metal5 77020 -102980 77120 -102880 1 PIX5571_IN
port 5650 n
rlabel metal5 78520 -102980 78620 -102880 1 PIX5572_IN
port 5651 n
rlabel metal5 80020 -102980 80120 -102880 1 PIX5573_IN
port 5652 n
rlabel metal5 81520 -102980 81620 -102880 1 PIX5574_IN
port 5653 n
rlabel metal5 83020 -102980 83120 -102880 1 PIX5575_IN
port 5654 n
rlabel metal5 84520 -102980 84620 -102880 1 PIX5576_IN
port 5655 n
rlabel metal5 86020 -102980 86120 -102880 1 PIX5577_IN
port 5656 n
rlabel metal5 87520 -102980 87620 -102880 1 PIX5578_IN
port 5657 n
rlabel metal5 89020 -102980 89120 -102880 1 PIX5579_IN
port 5658 n
rlabel metal5 90520 -102980 90620 -102880 1 PIX5580_IN
port 5659 n
rlabel metal5 92020 -102980 92120 -102880 1 PIX5581_IN
port 5660 n
rlabel metal5 93520 -102980 93620 -102880 1 PIX5582_IN
port 5661 n
rlabel metal5 95020 -102980 95120 -102880 1 PIX5583_IN
port 5662 n
rlabel metal5 96520 -102980 96620 -102880 1 PIX5584_IN
port 5663 n
rlabel metal5 98020 -102980 98120 -102880 1 PIX5585_IN
port 5664 n
rlabel metal5 99520 -102980 99620 -102880 1 PIX5586_IN
port 5665 n
rlabel metal5 101020 -102980 101120 -102880 1 PIX5587_IN
port 5666 n
rlabel metal5 102520 -102980 102620 -102880 1 PIX5588_IN
port 5667 n
rlabel metal5 104020 -102980 104120 -102880 1 PIX5589_IN
port 5668 n
rlabel metal5 105520 -102980 105620 -102880 1 PIX5590_IN
port 5669 n
rlabel metal5 107020 -102980 107120 -102880 1 PIX5591_IN
port 5670 n
rlabel metal5 108520 -102980 108620 -102880 1 PIX5592_IN
port 5671 n
rlabel metal5 110020 -102980 110120 -102880 1 PIX5593_IN
port 5672 n
rlabel metal5 111520 -102980 111620 -102880 1 PIX5594_IN
port 5673 n
rlabel metal5 113020 -102980 113120 -102880 1 PIX5595_IN
port 5674 n
rlabel metal5 114520 -102980 114620 -102880 1 PIX5596_IN
port 5675 n
rlabel metal5 116020 -102980 116120 -102880 1 PIX5597_IN
port 5676 n
rlabel metal5 117520 -102980 117620 -102880 1 PIX5598_IN
port 5677 n
rlabel metal5 119020 -102980 119120 -102880 1 PIX5599_IN
port 5678 n
rlabel metal5 520 -104480 620 -104380 1 PIX5600_IN
port 5679 n
rlabel metal2 -1500 -104260 -1500 -104215 3 ROW_SEL70
port 5680 e
rlabel metal5 2020 -104480 2120 -104380 1 PIX5601_IN
port 5681 n
rlabel metal5 3520 -104480 3620 -104380 1 PIX5602_IN
port 5682 n
rlabel metal5 5020 -104480 5120 -104380 1 PIX5603_IN
port 5683 n
rlabel metal5 6520 -104480 6620 -104380 1 PIX5604_IN
port 5684 n
rlabel metal5 8020 -104480 8120 -104380 1 PIX5605_IN
port 5685 n
rlabel metal5 9520 -104480 9620 -104380 1 PIX5606_IN
port 5686 n
rlabel metal5 11020 -104480 11120 -104380 1 PIX5607_IN
port 5687 n
rlabel metal5 12520 -104480 12620 -104380 1 PIX5608_IN
port 5688 n
rlabel metal5 14020 -104480 14120 -104380 1 PIX5609_IN
port 5689 n
rlabel metal5 15520 -104480 15620 -104380 1 PIX5610_IN
port 5690 n
rlabel metal5 17020 -104480 17120 -104380 1 PIX5611_IN
port 5691 n
rlabel metal5 18520 -104480 18620 -104380 1 PIX5612_IN
port 5692 n
rlabel metal5 20020 -104480 20120 -104380 1 PIX5613_IN
port 5693 n
rlabel metal5 21520 -104480 21620 -104380 1 PIX5614_IN
port 5694 n
rlabel metal5 23020 -104480 23120 -104380 1 PIX5615_IN
port 5695 n
rlabel metal5 24520 -104480 24620 -104380 1 PIX5616_IN
port 5696 n
rlabel metal5 26020 -104480 26120 -104380 1 PIX5617_IN
port 5697 n
rlabel metal5 27520 -104480 27620 -104380 1 PIX5618_IN
port 5698 n
rlabel metal5 29020 -104480 29120 -104380 1 PIX5619_IN
port 5699 n
rlabel metal5 30520 -104480 30620 -104380 1 PIX5620_IN
port 5700 n
rlabel metal5 32020 -104480 32120 -104380 1 PIX5621_IN
port 5701 n
rlabel metal5 33520 -104480 33620 -104380 1 PIX5622_IN
port 5702 n
rlabel metal5 35020 -104480 35120 -104380 1 PIX5623_IN
port 5703 n
rlabel metal5 36520 -104480 36620 -104380 1 PIX5624_IN
port 5704 n
rlabel metal5 38020 -104480 38120 -104380 1 PIX5625_IN
port 5705 n
rlabel metal5 39520 -104480 39620 -104380 1 PIX5626_IN
port 5706 n
rlabel metal5 41020 -104480 41120 -104380 1 PIX5627_IN
port 5707 n
rlabel metal5 42520 -104480 42620 -104380 1 PIX5628_IN
port 5708 n
rlabel metal5 44020 -104480 44120 -104380 1 PIX5629_IN
port 5709 n
rlabel metal5 45520 -104480 45620 -104380 1 PIX5630_IN
port 5710 n
rlabel metal5 47020 -104480 47120 -104380 1 PIX5631_IN
port 5711 n
rlabel metal5 48520 -104480 48620 -104380 1 PIX5632_IN
port 5712 n
rlabel metal5 50020 -104480 50120 -104380 1 PIX5633_IN
port 5713 n
rlabel metal5 51520 -104480 51620 -104380 1 PIX5634_IN
port 5714 n
rlabel metal5 53020 -104480 53120 -104380 1 PIX5635_IN
port 5715 n
rlabel metal5 54520 -104480 54620 -104380 1 PIX5636_IN
port 5716 n
rlabel metal5 56020 -104480 56120 -104380 1 PIX5637_IN
port 5717 n
rlabel metal5 57520 -104480 57620 -104380 1 PIX5638_IN
port 5718 n
rlabel metal5 59020 -104480 59120 -104380 1 PIX5639_IN
port 5719 n
rlabel metal5 60520 -104480 60620 -104380 1 PIX5640_IN
port 5720 n
rlabel metal5 62020 -104480 62120 -104380 1 PIX5641_IN
port 5721 n
rlabel metal5 63520 -104480 63620 -104380 1 PIX5642_IN
port 5722 n
rlabel metal5 65020 -104480 65120 -104380 1 PIX5643_IN
port 5723 n
rlabel metal5 66520 -104480 66620 -104380 1 PIX5644_IN
port 5724 n
rlabel metal5 68020 -104480 68120 -104380 1 PIX5645_IN
port 5725 n
rlabel metal5 69520 -104480 69620 -104380 1 PIX5646_IN
port 5726 n
rlabel metal5 71020 -104480 71120 -104380 1 PIX5647_IN
port 5727 n
rlabel metal5 72520 -104480 72620 -104380 1 PIX5648_IN
port 5728 n
rlabel metal5 74020 -104480 74120 -104380 1 PIX5649_IN
port 5729 n
rlabel metal5 75520 -104480 75620 -104380 1 PIX5650_IN
port 5730 n
rlabel metal5 77020 -104480 77120 -104380 1 PIX5651_IN
port 5731 n
rlabel metal5 78520 -104480 78620 -104380 1 PIX5652_IN
port 5732 n
rlabel metal5 80020 -104480 80120 -104380 1 PIX5653_IN
port 5733 n
rlabel metal5 81520 -104480 81620 -104380 1 PIX5654_IN
port 5734 n
rlabel metal5 83020 -104480 83120 -104380 1 PIX5655_IN
port 5735 n
rlabel metal5 84520 -104480 84620 -104380 1 PIX5656_IN
port 5736 n
rlabel metal5 86020 -104480 86120 -104380 1 PIX5657_IN
port 5737 n
rlabel metal5 87520 -104480 87620 -104380 1 PIX5658_IN
port 5738 n
rlabel metal5 89020 -104480 89120 -104380 1 PIX5659_IN
port 5739 n
rlabel metal5 90520 -104480 90620 -104380 1 PIX5660_IN
port 5740 n
rlabel metal5 92020 -104480 92120 -104380 1 PIX5661_IN
port 5741 n
rlabel metal5 93520 -104480 93620 -104380 1 PIX5662_IN
port 5742 n
rlabel metal5 95020 -104480 95120 -104380 1 PIX5663_IN
port 5743 n
rlabel metal5 96520 -104480 96620 -104380 1 PIX5664_IN
port 5744 n
rlabel metal5 98020 -104480 98120 -104380 1 PIX5665_IN
port 5745 n
rlabel metal5 99520 -104480 99620 -104380 1 PIX5666_IN
port 5746 n
rlabel metal5 101020 -104480 101120 -104380 1 PIX5667_IN
port 5747 n
rlabel metal5 102520 -104480 102620 -104380 1 PIX5668_IN
port 5748 n
rlabel metal5 104020 -104480 104120 -104380 1 PIX5669_IN
port 5749 n
rlabel metal5 105520 -104480 105620 -104380 1 PIX5670_IN
port 5750 n
rlabel metal5 107020 -104480 107120 -104380 1 PIX5671_IN
port 5751 n
rlabel metal5 108520 -104480 108620 -104380 1 PIX5672_IN
port 5752 n
rlabel metal5 110020 -104480 110120 -104380 1 PIX5673_IN
port 5753 n
rlabel metal5 111520 -104480 111620 -104380 1 PIX5674_IN
port 5754 n
rlabel metal5 113020 -104480 113120 -104380 1 PIX5675_IN
port 5755 n
rlabel metal5 114520 -104480 114620 -104380 1 PIX5676_IN
port 5756 n
rlabel metal5 116020 -104480 116120 -104380 1 PIX5677_IN
port 5757 n
rlabel metal5 117520 -104480 117620 -104380 1 PIX5678_IN
port 5758 n
rlabel metal5 119020 -104480 119120 -104380 1 PIX5679_IN
port 5759 n
rlabel metal5 520 -105980 620 -105880 1 PIX5680_IN
port 5760 n
rlabel metal2 -1500 -105760 -1500 -105715 3 ROW_SEL71
port 5761 e
rlabel metal5 2020 -105980 2120 -105880 1 PIX5681_IN
port 5762 n
rlabel metal5 3520 -105980 3620 -105880 1 PIX5682_IN
port 5763 n
rlabel metal5 5020 -105980 5120 -105880 1 PIX5683_IN
port 5764 n
rlabel metal5 6520 -105980 6620 -105880 1 PIX5684_IN
port 5765 n
rlabel metal5 8020 -105980 8120 -105880 1 PIX5685_IN
port 5766 n
rlabel metal5 9520 -105980 9620 -105880 1 PIX5686_IN
port 5767 n
rlabel metal5 11020 -105980 11120 -105880 1 PIX5687_IN
port 5768 n
rlabel metal5 12520 -105980 12620 -105880 1 PIX5688_IN
port 5769 n
rlabel metal5 14020 -105980 14120 -105880 1 PIX5689_IN
port 5770 n
rlabel metal5 15520 -105980 15620 -105880 1 PIX5690_IN
port 5771 n
rlabel metal5 17020 -105980 17120 -105880 1 PIX5691_IN
port 5772 n
rlabel metal5 18520 -105980 18620 -105880 1 PIX5692_IN
port 5773 n
rlabel metal5 20020 -105980 20120 -105880 1 PIX5693_IN
port 5774 n
rlabel metal5 21520 -105980 21620 -105880 1 PIX5694_IN
port 5775 n
rlabel metal5 23020 -105980 23120 -105880 1 PIX5695_IN
port 5776 n
rlabel metal5 24520 -105980 24620 -105880 1 PIX5696_IN
port 5777 n
rlabel metal5 26020 -105980 26120 -105880 1 PIX5697_IN
port 5778 n
rlabel metal5 27520 -105980 27620 -105880 1 PIX5698_IN
port 5779 n
rlabel metal5 29020 -105980 29120 -105880 1 PIX5699_IN
port 5780 n
rlabel metal5 30520 -105980 30620 -105880 1 PIX5700_IN
port 5781 n
rlabel metal5 32020 -105980 32120 -105880 1 PIX5701_IN
port 5782 n
rlabel metal5 33520 -105980 33620 -105880 1 PIX5702_IN
port 5783 n
rlabel metal5 35020 -105980 35120 -105880 1 PIX5703_IN
port 5784 n
rlabel metal5 36520 -105980 36620 -105880 1 PIX5704_IN
port 5785 n
rlabel metal5 38020 -105980 38120 -105880 1 PIX5705_IN
port 5786 n
rlabel metal5 39520 -105980 39620 -105880 1 PIX5706_IN
port 5787 n
rlabel metal5 41020 -105980 41120 -105880 1 PIX5707_IN
port 5788 n
rlabel metal5 42520 -105980 42620 -105880 1 PIX5708_IN
port 5789 n
rlabel metal5 44020 -105980 44120 -105880 1 PIX5709_IN
port 5790 n
rlabel metal5 45520 -105980 45620 -105880 1 PIX5710_IN
port 5791 n
rlabel metal5 47020 -105980 47120 -105880 1 PIX5711_IN
port 5792 n
rlabel metal5 48520 -105980 48620 -105880 1 PIX5712_IN
port 5793 n
rlabel metal5 50020 -105980 50120 -105880 1 PIX5713_IN
port 5794 n
rlabel metal5 51520 -105980 51620 -105880 1 PIX5714_IN
port 5795 n
rlabel metal5 53020 -105980 53120 -105880 1 PIX5715_IN
port 5796 n
rlabel metal5 54520 -105980 54620 -105880 1 PIX5716_IN
port 5797 n
rlabel metal5 56020 -105980 56120 -105880 1 PIX5717_IN
port 5798 n
rlabel metal5 57520 -105980 57620 -105880 1 PIX5718_IN
port 5799 n
rlabel metal5 59020 -105980 59120 -105880 1 PIX5719_IN
port 5800 n
rlabel metal5 60520 -105980 60620 -105880 1 PIX5720_IN
port 5801 n
rlabel metal5 62020 -105980 62120 -105880 1 PIX5721_IN
port 5802 n
rlabel metal5 63520 -105980 63620 -105880 1 PIX5722_IN
port 5803 n
rlabel metal5 65020 -105980 65120 -105880 1 PIX5723_IN
port 5804 n
rlabel metal5 66520 -105980 66620 -105880 1 PIX5724_IN
port 5805 n
rlabel metal5 68020 -105980 68120 -105880 1 PIX5725_IN
port 5806 n
rlabel metal5 69520 -105980 69620 -105880 1 PIX5726_IN
port 5807 n
rlabel metal5 71020 -105980 71120 -105880 1 PIX5727_IN
port 5808 n
rlabel metal5 72520 -105980 72620 -105880 1 PIX5728_IN
port 5809 n
rlabel metal5 74020 -105980 74120 -105880 1 PIX5729_IN
port 5810 n
rlabel metal5 75520 -105980 75620 -105880 1 PIX5730_IN
port 5811 n
rlabel metal5 77020 -105980 77120 -105880 1 PIX5731_IN
port 5812 n
rlabel metal5 78520 -105980 78620 -105880 1 PIX5732_IN
port 5813 n
rlabel metal5 80020 -105980 80120 -105880 1 PIX5733_IN
port 5814 n
rlabel metal5 81520 -105980 81620 -105880 1 PIX5734_IN
port 5815 n
rlabel metal5 83020 -105980 83120 -105880 1 PIX5735_IN
port 5816 n
rlabel metal5 84520 -105980 84620 -105880 1 PIX5736_IN
port 5817 n
rlabel metal5 86020 -105980 86120 -105880 1 PIX5737_IN
port 5818 n
rlabel metal5 87520 -105980 87620 -105880 1 PIX5738_IN
port 5819 n
rlabel metal5 89020 -105980 89120 -105880 1 PIX5739_IN
port 5820 n
rlabel metal5 90520 -105980 90620 -105880 1 PIX5740_IN
port 5821 n
rlabel metal5 92020 -105980 92120 -105880 1 PIX5741_IN
port 5822 n
rlabel metal5 93520 -105980 93620 -105880 1 PIX5742_IN
port 5823 n
rlabel metal5 95020 -105980 95120 -105880 1 PIX5743_IN
port 5824 n
rlabel metal5 96520 -105980 96620 -105880 1 PIX5744_IN
port 5825 n
rlabel metal5 98020 -105980 98120 -105880 1 PIX5745_IN
port 5826 n
rlabel metal5 99520 -105980 99620 -105880 1 PIX5746_IN
port 5827 n
rlabel metal5 101020 -105980 101120 -105880 1 PIX5747_IN
port 5828 n
rlabel metal5 102520 -105980 102620 -105880 1 PIX5748_IN
port 5829 n
rlabel metal5 104020 -105980 104120 -105880 1 PIX5749_IN
port 5830 n
rlabel metal5 105520 -105980 105620 -105880 1 PIX5750_IN
port 5831 n
rlabel metal5 107020 -105980 107120 -105880 1 PIX5751_IN
port 5832 n
rlabel metal5 108520 -105980 108620 -105880 1 PIX5752_IN
port 5833 n
rlabel metal5 110020 -105980 110120 -105880 1 PIX5753_IN
port 5834 n
rlabel metal5 111520 -105980 111620 -105880 1 PIX5754_IN
port 5835 n
rlabel metal5 113020 -105980 113120 -105880 1 PIX5755_IN
port 5836 n
rlabel metal5 114520 -105980 114620 -105880 1 PIX5756_IN
port 5837 n
rlabel metal5 116020 -105980 116120 -105880 1 PIX5757_IN
port 5838 n
rlabel metal5 117520 -105980 117620 -105880 1 PIX5758_IN
port 5839 n
rlabel metal5 119020 -105980 119120 -105880 1 PIX5759_IN
port 5840 n
rlabel metal5 520 -107480 620 -107380 1 PIX5760_IN
port 5841 n
rlabel metal2 -1500 -107260 -1500 -107215 3 ROW_SEL72
port 5842 e
rlabel metal5 2020 -107480 2120 -107380 1 PIX5761_IN
port 5843 n
rlabel metal5 3520 -107480 3620 -107380 1 PIX5762_IN
port 5844 n
rlabel metal5 5020 -107480 5120 -107380 1 PIX5763_IN
port 5845 n
rlabel metal5 6520 -107480 6620 -107380 1 PIX5764_IN
port 5846 n
rlabel metal5 8020 -107480 8120 -107380 1 PIX5765_IN
port 5847 n
rlabel metal5 9520 -107480 9620 -107380 1 PIX5766_IN
port 5848 n
rlabel metal5 11020 -107480 11120 -107380 1 PIX5767_IN
port 5849 n
rlabel metal5 12520 -107480 12620 -107380 1 PIX5768_IN
port 5850 n
rlabel metal5 14020 -107480 14120 -107380 1 PIX5769_IN
port 5851 n
rlabel metal5 15520 -107480 15620 -107380 1 PIX5770_IN
port 5852 n
rlabel metal5 17020 -107480 17120 -107380 1 PIX5771_IN
port 5853 n
rlabel metal5 18520 -107480 18620 -107380 1 PIX5772_IN
port 5854 n
rlabel metal5 20020 -107480 20120 -107380 1 PIX5773_IN
port 5855 n
rlabel metal5 21520 -107480 21620 -107380 1 PIX5774_IN
port 5856 n
rlabel metal5 23020 -107480 23120 -107380 1 PIX5775_IN
port 5857 n
rlabel metal5 24520 -107480 24620 -107380 1 PIX5776_IN
port 5858 n
rlabel metal5 26020 -107480 26120 -107380 1 PIX5777_IN
port 5859 n
rlabel metal5 27520 -107480 27620 -107380 1 PIX5778_IN
port 5860 n
rlabel metal5 29020 -107480 29120 -107380 1 PIX5779_IN
port 5861 n
rlabel metal5 30520 -107480 30620 -107380 1 PIX5780_IN
port 5862 n
rlabel metal5 32020 -107480 32120 -107380 1 PIX5781_IN
port 5863 n
rlabel metal5 33520 -107480 33620 -107380 1 PIX5782_IN
port 5864 n
rlabel metal5 35020 -107480 35120 -107380 1 PIX5783_IN
port 5865 n
rlabel metal5 36520 -107480 36620 -107380 1 PIX5784_IN
port 5866 n
rlabel metal5 38020 -107480 38120 -107380 1 PIX5785_IN
port 5867 n
rlabel metal5 39520 -107480 39620 -107380 1 PIX5786_IN
port 5868 n
rlabel metal5 41020 -107480 41120 -107380 1 PIX5787_IN
port 5869 n
rlabel metal5 42520 -107480 42620 -107380 1 PIX5788_IN
port 5870 n
rlabel metal5 44020 -107480 44120 -107380 1 PIX5789_IN
port 5871 n
rlabel metal5 45520 -107480 45620 -107380 1 PIX5790_IN
port 5872 n
rlabel metal5 47020 -107480 47120 -107380 1 PIX5791_IN
port 5873 n
rlabel metal5 48520 -107480 48620 -107380 1 PIX5792_IN
port 5874 n
rlabel metal5 50020 -107480 50120 -107380 1 PIX5793_IN
port 5875 n
rlabel metal5 51520 -107480 51620 -107380 1 PIX5794_IN
port 5876 n
rlabel metal5 53020 -107480 53120 -107380 1 PIX5795_IN
port 5877 n
rlabel metal5 54520 -107480 54620 -107380 1 PIX5796_IN
port 5878 n
rlabel metal5 56020 -107480 56120 -107380 1 PIX5797_IN
port 5879 n
rlabel metal5 57520 -107480 57620 -107380 1 PIX5798_IN
port 5880 n
rlabel metal5 59020 -107480 59120 -107380 1 PIX5799_IN
port 5881 n
rlabel metal5 60520 -107480 60620 -107380 1 PIX5800_IN
port 5882 n
rlabel metal5 62020 -107480 62120 -107380 1 PIX5801_IN
port 5883 n
rlabel metal5 63520 -107480 63620 -107380 1 PIX5802_IN
port 5884 n
rlabel metal5 65020 -107480 65120 -107380 1 PIX5803_IN
port 5885 n
rlabel metal5 66520 -107480 66620 -107380 1 PIX5804_IN
port 5886 n
rlabel metal5 68020 -107480 68120 -107380 1 PIX5805_IN
port 5887 n
rlabel metal5 69520 -107480 69620 -107380 1 PIX5806_IN
port 5888 n
rlabel metal5 71020 -107480 71120 -107380 1 PIX5807_IN
port 5889 n
rlabel metal5 72520 -107480 72620 -107380 1 PIX5808_IN
port 5890 n
rlabel metal5 74020 -107480 74120 -107380 1 PIX5809_IN
port 5891 n
rlabel metal5 75520 -107480 75620 -107380 1 PIX5810_IN
port 5892 n
rlabel metal5 77020 -107480 77120 -107380 1 PIX5811_IN
port 5893 n
rlabel metal5 78520 -107480 78620 -107380 1 PIX5812_IN
port 5894 n
rlabel metal5 80020 -107480 80120 -107380 1 PIX5813_IN
port 5895 n
rlabel metal5 81520 -107480 81620 -107380 1 PIX5814_IN
port 5896 n
rlabel metal5 83020 -107480 83120 -107380 1 PIX5815_IN
port 5897 n
rlabel metal5 84520 -107480 84620 -107380 1 PIX5816_IN
port 5898 n
rlabel metal5 86020 -107480 86120 -107380 1 PIX5817_IN
port 5899 n
rlabel metal5 87520 -107480 87620 -107380 1 PIX5818_IN
port 5900 n
rlabel metal5 89020 -107480 89120 -107380 1 PIX5819_IN
port 5901 n
rlabel metal5 90520 -107480 90620 -107380 1 PIX5820_IN
port 5902 n
rlabel metal5 92020 -107480 92120 -107380 1 PIX5821_IN
port 5903 n
rlabel metal5 93520 -107480 93620 -107380 1 PIX5822_IN
port 5904 n
rlabel metal5 95020 -107480 95120 -107380 1 PIX5823_IN
port 5905 n
rlabel metal5 96520 -107480 96620 -107380 1 PIX5824_IN
port 5906 n
rlabel metal5 98020 -107480 98120 -107380 1 PIX5825_IN
port 5907 n
rlabel metal5 99520 -107480 99620 -107380 1 PIX5826_IN
port 5908 n
rlabel metal5 101020 -107480 101120 -107380 1 PIX5827_IN
port 5909 n
rlabel metal5 102520 -107480 102620 -107380 1 PIX5828_IN
port 5910 n
rlabel metal5 104020 -107480 104120 -107380 1 PIX5829_IN
port 5911 n
rlabel metal5 105520 -107480 105620 -107380 1 PIX5830_IN
port 5912 n
rlabel metal5 107020 -107480 107120 -107380 1 PIX5831_IN
port 5913 n
rlabel metal5 108520 -107480 108620 -107380 1 PIX5832_IN
port 5914 n
rlabel metal5 110020 -107480 110120 -107380 1 PIX5833_IN
port 5915 n
rlabel metal5 111520 -107480 111620 -107380 1 PIX5834_IN
port 5916 n
rlabel metal5 113020 -107480 113120 -107380 1 PIX5835_IN
port 5917 n
rlabel metal5 114520 -107480 114620 -107380 1 PIX5836_IN
port 5918 n
rlabel metal5 116020 -107480 116120 -107380 1 PIX5837_IN
port 5919 n
rlabel metal5 117520 -107480 117620 -107380 1 PIX5838_IN
port 5920 n
rlabel metal5 119020 -107480 119120 -107380 1 PIX5839_IN
port 5921 n
rlabel metal5 520 -108980 620 -108880 1 PIX5840_IN
port 5922 n
rlabel metal2 -1500 -108760 -1500 -108715 3 ROW_SEL73
port 5923 e
rlabel metal5 2020 -108980 2120 -108880 1 PIX5841_IN
port 5924 n
rlabel metal5 3520 -108980 3620 -108880 1 PIX5842_IN
port 5925 n
rlabel metal5 5020 -108980 5120 -108880 1 PIX5843_IN
port 5926 n
rlabel metal5 6520 -108980 6620 -108880 1 PIX5844_IN
port 5927 n
rlabel metal5 8020 -108980 8120 -108880 1 PIX5845_IN
port 5928 n
rlabel metal5 9520 -108980 9620 -108880 1 PIX5846_IN
port 5929 n
rlabel metal5 11020 -108980 11120 -108880 1 PIX5847_IN
port 5930 n
rlabel metal5 12520 -108980 12620 -108880 1 PIX5848_IN
port 5931 n
rlabel metal5 14020 -108980 14120 -108880 1 PIX5849_IN
port 5932 n
rlabel metal5 15520 -108980 15620 -108880 1 PIX5850_IN
port 5933 n
rlabel metal5 17020 -108980 17120 -108880 1 PIX5851_IN
port 5934 n
rlabel metal5 18520 -108980 18620 -108880 1 PIX5852_IN
port 5935 n
rlabel metal5 20020 -108980 20120 -108880 1 PIX5853_IN
port 5936 n
rlabel metal5 21520 -108980 21620 -108880 1 PIX5854_IN
port 5937 n
rlabel metal5 23020 -108980 23120 -108880 1 PIX5855_IN
port 5938 n
rlabel metal5 24520 -108980 24620 -108880 1 PIX5856_IN
port 5939 n
rlabel metal5 26020 -108980 26120 -108880 1 PIX5857_IN
port 5940 n
rlabel metal5 27520 -108980 27620 -108880 1 PIX5858_IN
port 5941 n
rlabel metal5 29020 -108980 29120 -108880 1 PIX5859_IN
port 5942 n
rlabel metal5 30520 -108980 30620 -108880 1 PIX5860_IN
port 5943 n
rlabel metal5 32020 -108980 32120 -108880 1 PIX5861_IN
port 5944 n
rlabel metal5 33520 -108980 33620 -108880 1 PIX5862_IN
port 5945 n
rlabel metal5 35020 -108980 35120 -108880 1 PIX5863_IN
port 5946 n
rlabel metal5 36520 -108980 36620 -108880 1 PIX5864_IN
port 5947 n
rlabel metal5 38020 -108980 38120 -108880 1 PIX5865_IN
port 5948 n
rlabel metal5 39520 -108980 39620 -108880 1 PIX5866_IN
port 5949 n
rlabel metal5 41020 -108980 41120 -108880 1 PIX5867_IN
port 5950 n
rlabel metal5 42520 -108980 42620 -108880 1 PIX5868_IN
port 5951 n
rlabel metal5 44020 -108980 44120 -108880 1 PIX5869_IN
port 5952 n
rlabel metal5 45520 -108980 45620 -108880 1 PIX5870_IN
port 5953 n
rlabel metal5 47020 -108980 47120 -108880 1 PIX5871_IN
port 5954 n
rlabel metal5 48520 -108980 48620 -108880 1 PIX5872_IN
port 5955 n
rlabel metal5 50020 -108980 50120 -108880 1 PIX5873_IN
port 5956 n
rlabel metal5 51520 -108980 51620 -108880 1 PIX5874_IN
port 5957 n
rlabel metal5 53020 -108980 53120 -108880 1 PIX5875_IN
port 5958 n
rlabel metal5 54520 -108980 54620 -108880 1 PIX5876_IN
port 5959 n
rlabel metal5 56020 -108980 56120 -108880 1 PIX5877_IN
port 5960 n
rlabel metal5 57520 -108980 57620 -108880 1 PIX5878_IN
port 5961 n
rlabel metal5 59020 -108980 59120 -108880 1 PIX5879_IN
port 5962 n
rlabel metal5 60520 -108980 60620 -108880 1 PIX5880_IN
port 5963 n
rlabel metal5 62020 -108980 62120 -108880 1 PIX5881_IN
port 5964 n
rlabel metal5 63520 -108980 63620 -108880 1 PIX5882_IN
port 5965 n
rlabel metal5 65020 -108980 65120 -108880 1 PIX5883_IN
port 5966 n
rlabel metal5 66520 -108980 66620 -108880 1 PIX5884_IN
port 5967 n
rlabel metal5 68020 -108980 68120 -108880 1 PIX5885_IN
port 5968 n
rlabel metal5 69520 -108980 69620 -108880 1 PIX5886_IN
port 5969 n
rlabel metal5 71020 -108980 71120 -108880 1 PIX5887_IN
port 5970 n
rlabel metal5 72520 -108980 72620 -108880 1 PIX5888_IN
port 5971 n
rlabel metal5 74020 -108980 74120 -108880 1 PIX5889_IN
port 5972 n
rlabel metal5 75520 -108980 75620 -108880 1 PIX5890_IN
port 5973 n
rlabel metal5 77020 -108980 77120 -108880 1 PIX5891_IN
port 5974 n
rlabel metal5 78520 -108980 78620 -108880 1 PIX5892_IN
port 5975 n
rlabel metal5 80020 -108980 80120 -108880 1 PIX5893_IN
port 5976 n
rlabel metal5 81520 -108980 81620 -108880 1 PIX5894_IN
port 5977 n
rlabel metal5 83020 -108980 83120 -108880 1 PIX5895_IN
port 5978 n
rlabel metal5 84520 -108980 84620 -108880 1 PIX5896_IN
port 5979 n
rlabel metal5 86020 -108980 86120 -108880 1 PIX5897_IN
port 5980 n
rlabel metal5 87520 -108980 87620 -108880 1 PIX5898_IN
port 5981 n
rlabel metal5 89020 -108980 89120 -108880 1 PIX5899_IN
port 5982 n
rlabel metal5 90520 -108980 90620 -108880 1 PIX5900_IN
port 5983 n
rlabel metal5 92020 -108980 92120 -108880 1 PIX5901_IN
port 5984 n
rlabel metal5 93520 -108980 93620 -108880 1 PIX5902_IN
port 5985 n
rlabel metal5 95020 -108980 95120 -108880 1 PIX5903_IN
port 5986 n
rlabel metal5 96520 -108980 96620 -108880 1 PIX5904_IN
port 5987 n
rlabel metal5 98020 -108980 98120 -108880 1 PIX5905_IN
port 5988 n
rlabel metal5 99520 -108980 99620 -108880 1 PIX5906_IN
port 5989 n
rlabel metal5 101020 -108980 101120 -108880 1 PIX5907_IN
port 5990 n
rlabel metal5 102520 -108980 102620 -108880 1 PIX5908_IN
port 5991 n
rlabel metal5 104020 -108980 104120 -108880 1 PIX5909_IN
port 5992 n
rlabel metal5 105520 -108980 105620 -108880 1 PIX5910_IN
port 5993 n
rlabel metal5 107020 -108980 107120 -108880 1 PIX5911_IN
port 5994 n
rlabel metal5 108520 -108980 108620 -108880 1 PIX5912_IN
port 5995 n
rlabel metal5 110020 -108980 110120 -108880 1 PIX5913_IN
port 5996 n
rlabel metal5 111520 -108980 111620 -108880 1 PIX5914_IN
port 5997 n
rlabel metal5 113020 -108980 113120 -108880 1 PIX5915_IN
port 5998 n
rlabel metal5 114520 -108980 114620 -108880 1 PIX5916_IN
port 5999 n
rlabel metal5 116020 -108980 116120 -108880 1 PIX5917_IN
port 6000 n
rlabel metal5 117520 -108980 117620 -108880 1 PIX5918_IN
port 6001 n
rlabel metal5 119020 -108980 119120 -108880 1 PIX5919_IN
port 6002 n
rlabel metal5 520 -110480 620 -110380 1 PIX5920_IN
port 6003 n
rlabel metal2 -1500 -110260 -1500 -110215 3 ROW_SEL74
port 6004 e
rlabel metal5 2020 -110480 2120 -110380 1 PIX5921_IN
port 6005 n
rlabel metal5 3520 -110480 3620 -110380 1 PIX5922_IN
port 6006 n
rlabel metal5 5020 -110480 5120 -110380 1 PIX5923_IN
port 6007 n
rlabel metal5 6520 -110480 6620 -110380 1 PIX5924_IN
port 6008 n
rlabel metal5 8020 -110480 8120 -110380 1 PIX5925_IN
port 6009 n
rlabel metal5 9520 -110480 9620 -110380 1 PIX5926_IN
port 6010 n
rlabel metal5 11020 -110480 11120 -110380 1 PIX5927_IN
port 6011 n
rlabel metal5 12520 -110480 12620 -110380 1 PIX5928_IN
port 6012 n
rlabel metal5 14020 -110480 14120 -110380 1 PIX5929_IN
port 6013 n
rlabel metal5 15520 -110480 15620 -110380 1 PIX5930_IN
port 6014 n
rlabel metal5 17020 -110480 17120 -110380 1 PIX5931_IN
port 6015 n
rlabel metal5 18520 -110480 18620 -110380 1 PIX5932_IN
port 6016 n
rlabel metal5 20020 -110480 20120 -110380 1 PIX5933_IN
port 6017 n
rlabel metal5 21520 -110480 21620 -110380 1 PIX5934_IN
port 6018 n
rlabel metal5 23020 -110480 23120 -110380 1 PIX5935_IN
port 6019 n
rlabel metal5 24520 -110480 24620 -110380 1 PIX5936_IN
port 6020 n
rlabel metal5 26020 -110480 26120 -110380 1 PIX5937_IN
port 6021 n
rlabel metal5 27520 -110480 27620 -110380 1 PIX5938_IN
port 6022 n
rlabel metal5 29020 -110480 29120 -110380 1 PIX5939_IN
port 6023 n
rlabel metal5 30520 -110480 30620 -110380 1 PIX5940_IN
port 6024 n
rlabel metal5 32020 -110480 32120 -110380 1 PIX5941_IN
port 6025 n
rlabel metal5 33520 -110480 33620 -110380 1 PIX5942_IN
port 6026 n
rlabel metal5 35020 -110480 35120 -110380 1 PIX5943_IN
port 6027 n
rlabel metal5 36520 -110480 36620 -110380 1 PIX5944_IN
port 6028 n
rlabel metal5 38020 -110480 38120 -110380 1 PIX5945_IN
port 6029 n
rlabel metal5 39520 -110480 39620 -110380 1 PIX5946_IN
port 6030 n
rlabel metal5 41020 -110480 41120 -110380 1 PIX5947_IN
port 6031 n
rlabel metal5 42520 -110480 42620 -110380 1 PIX5948_IN
port 6032 n
rlabel metal5 44020 -110480 44120 -110380 1 PIX5949_IN
port 6033 n
rlabel metal5 45520 -110480 45620 -110380 1 PIX5950_IN
port 6034 n
rlabel metal5 47020 -110480 47120 -110380 1 PIX5951_IN
port 6035 n
rlabel metal5 48520 -110480 48620 -110380 1 PIX5952_IN
port 6036 n
rlabel metal5 50020 -110480 50120 -110380 1 PIX5953_IN
port 6037 n
rlabel metal5 51520 -110480 51620 -110380 1 PIX5954_IN
port 6038 n
rlabel metal5 53020 -110480 53120 -110380 1 PIX5955_IN
port 6039 n
rlabel metal5 54520 -110480 54620 -110380 1 PIX5956_IN
port 6040 n
rlabel metal5 56020 -110480 56120 -110380 1 PIX5957_IN
port 6041 n
rlabel metal5 57520 -110480 57620 -110380 1 PIX5958_IN
port 6042 n
rlabel metal5 59020 -110480 59120 -110380 1 PIX5959_IN
port 6043 n
rlabel metal5 60520 -110480 60620 -110380 1 PIX5960_IN
port 6044 n
rlabel metal5 62020 -110480 62120 -110380 1 PIX5961_IN
port 6045 n
rlabel metal5 63520 -110480 63620 -110380 1 PIX5962_IN
port 6046 n
rlabel metal5 65020 -110480 65120 -110380 1 PIX5963_IN
port 6047 n
rlabel metal5 66520 -110480 66620 -110380 1 PIX5964_IN
port 6048 n
rlabel metal5 68020 -110480 68120 -110380 1 PIX5965_IN
port 6049 n
rlabel metal5 69520 -110480 69620 -110380 1 PIX5966_IN
port 6050 n
rlabel metal5 71020 -110480 71120 -110380 1 PIX5967_IN
port 6051 n
rlabel metal5 72520 -110480 72620 -110380 1 PIX5968_IN
port 6052 n
rlabel metal5 74020 -110480 74120 -110380 1 PIX5969_IN
port 6053 n
rlabel metal5 75520 -110480 75620 -110380 1 PIX5970_IN
port 6054 n
rlabel metal5 77020 -110480 77120 -110380 1 PIX5971_IN
port 6055 n
rlabel metal5 78520 -110480 78620 -110380 1 PIX5972_IN
port 6056 n
rlabel metal5 80020 -110480 80120 -110380 1 PIX5973_IN
port 6057 n
rlabel metal5 81520 -110480 81620 -110380 1 PIX5974_IN
port 6058 n
rlabel metal5 83020 -110480 83120 -110380 1 PIX5975_IN
port 6059 n
rlabel metal5 84520 -110480 84620 -110380 1 PIX5976_IN
port 6060 n
rlabel metal5 86020 -110480 86120 -110380 1 PIX5977_IN
port 6061 n
rlabel metal5 87520 -110480 87620 -110380 1 PIX5978_IN
port 6062 n
rlabel metal5 89020 -110480 89120 -110380 1 PIX5979_IN
port 6063 n
rlabel metal5 90520 -110480 90620 -110380 1 PIX5980_IN
port 6064 n
rlabel metal5 92020 -110480 92120 -110380 1 PIX5981_IN
port 6065 n
rlabel metal5 93520 -110480 93620 -110380 1 PIX5982_IN
port 6066 n
rlabel metal5 95020 -110480 95120 -110380 1 PIX5983_IN
port 6067 n
rlabel metal5 96520 -110480 96620 -110380 1 PIX5984_IN
port 6068 n
rlabel metal5 98020 -110480 98120 -110380 1 PIX5985_IN
port 6069 n
rlabel metal5 99520 -110480 99620 -110380 1 PIX5986_IN
port 6070 n
rlabel metal5 101020 -110480 101120 -110380 1 PIX5987_IN
port 6071 n
rlabel metal5 102520 -110480 102620 -110380 1 PIX5988_IN
port 6072 n
rlabel metal5 104020 -110480 104120 -110380 1 PIX5989_IN
port 6073 n
rlabel metal5 105520 -110480 105620 -110380 1 PIX5990_IN
port 6074 n
rlabel metal5 107020 -110480 107120 -110380 1 PIX5991_IN
port 6075 n
rlabel metal5 108520 -110480 108620 -110380 1 PIX5992_IN
port 6076 n
rlabel metal5 110020 -110480 110120 -110380 1 PIX5993_IN
port 6077 n
rlabel metal5 111520 -110480 111620 -110380 1 PIX5994_IN
port 6078 n
rlabel metal5 113020 -110480 113120 -110380 1 PIX5995_IN
port 6079 n
rlabel metal5 114520 -110480 114620 -110380 1 PIX5996_IN
port 6080 n
rlabel metal5 116020 -110480 116120 -110380 1 PIX5997_IN
port 6081 n
rlabel metal5 117520 -110480 117620 -110380 1 PIX5998_IN
port 6082 n
rlabel metal5 119020 -110480 119120 -110380 1 PIX5999_IN
port 6083 n
rlabel metal5 520 -111980 620 -111880 1 PIX6000_IN
port 6084 n
rlabel metal2 -1500 -111760 -1500 -111715 3 ROW_SEL75
port 6085 e
rlabel metal5 2020 -111980 2120 -111880 1 PIX6001_IN
port 6086 n
rlabel metal5 3520 -111980 3620 -111880 1 PIX6002_IN
port 6087 n
rlabel metal5 5020 -111980 5120 -111880 1 PIX6003_IN
port 6088 n
rlabel metal5 6520 -111980 6620 -111880 1 PIX6004_IN
port 6089 n
rlabel metal5 8020 -111980 8120 -111880 1 PIX6005_IN
port 6090 n
rlabel metal5 9520 -111980 9620 -111880 1 PIX6006_IN
port 6091 n
rlabel metal5 11020 -111980 11120 -111880 1 PIX6007_IN
port 6092 n
rlabel metal5 12520 -111980 12620 -111880 1 PIX6008_IN
port 6093 n
rlabel metal5 14020 -111980 14120 -111880 1 PIX6009_IN
port 6094 n
rlabel metal5 15520 -111980 15620 -111880 1 PIX6010_IN
port 6095 n
rlabel metal5 17020 -111980 17120 -111880 1 PIX6011_IN
port 6096 n
rlabel metal5 18520 -111980 18620 -111880 1 PIX6012_IN
port 6097 n
rlabel metal5 20020 -111980 20120 -111880 1 PIX6013_IN
port 6098 n
rlabel metal5 21520 -111980 21620 -111880 1 PIX6014_IN
port 6099 n
rlabel metal5 23020 -111980 23120 -111880 1 PIX6015_IN
port 6100 n
rlabel metal5 24520 -111980 24620 -111880 1 PIX6016_IN
port 6101 n
rlabel metal5 26020 -111980 26120 -111880 1 PIX6017_IN
port 6102 n
rlabel metal5 27520 -111980 27620 -111880 1 PIX6018_IN
port 6103 n
rlabel metal5 29020 -111980 29120 -111880 1 PIX6019_IN
port 6104 n
rlabel metal5 30520 -111980 30620 -111880 1 PIX6020_IN
port 6105 n
rlabel metal5 32020 -111980 32120 -111880 1 PIX6021_IN
port 6106 n
rlabel metal5 33520 -111980 33620 -111880 1 PIX6022_IN
port 6107 n
rlabel metal5 35020 -111980 35120 -111880 1 PIX6023_IN
port 6108 n
rlabel metal5 36520 -111980 36620 -111880 1 PIX6024_IN
port 6109 n
rlabel metal5 38020 -111980 38120 -111880 1 PIX6025_IN
port 6110 n
rlabel metal5 39520 -111980 39620 -111880 1 PIX6026_IN
port 6111 n
rlabel metal5 41020 -111980 41120 -111880 1 PIX6027_IN
port 6112 n
rlabel metal5 42520 -111980 42620 -111880 1 PIX6028_IN
port 6113 n
rlabel metal5 44020 -111980 44120 -111880 1 PIX6029_IN
port 6114 n
rlabel metal5 45520 -111980 45620 -111880 1 PIX6030_IN
port 6115 n
rlabel metal5 47020 -111980 47120 -111880 1 PIX6031_IN
port 6116 n
rlabel metal5 48520 -111980 48620 -111880 1 PIX6032_IN
port 6117 n
rlabel metal5 50020 -111980 50120 -111880 1 PIX6033_IN
port 6118 n
rlabel metal5 51520 -111980 51620 -111880 1 PIX6034_IN
port 6119 n
rlabel metal5 53020 -111980 53120 -111880 1 PIX6035_IN
port 6120 n
rlabel metal5 54520 -111980 54620 -111880 1 PIX6036_IN
port 6121 n
rlabel metal5 56020 -111980 56120 -111880 1 PIX6037_IN
port 6122 n
rlabel metal5 57520 -111980 57620 -111880 1 PIX6038_IN
port 6123 n
rlabel metal5 59020 -111980 59120 -111880 1 PIX6039_IN
port 6124 n
rlabel metal5 60520 -111980 60620 -111880 1 PIX6040_IN
port 6125 n
rlabel metal5 62020 -111980 62120 -111880 1 PIX6041_IN
port 6126 n
rlabel metal5 63520 -111980 63620 -111880 1 PIX6042_IN
port 6127 n
rlabel metal5 65020 -111980 65120 -111880 1 PIX6043_IN
port 6128 n
rlabel metal5 66520 -111980 66620 -111880 1 PIX6044_IN
port 6129 n
rlabel metal5 68020 -111980 68120 -111880 1 PIX6045_IN
port 6130 n
rlabel metal5 69520 -111980 69620 -111880 1 PIX6046_IN
port 6131 n
rlabel metal5 71020 -111980 71120 -111880 1 PIX6047_IN
port 6132 n
rlabel metal5 72520 -111980 72620 -111880 1 PIX6048_IN
port 6133 n
rlabel metal5 74020 -111980 74120 -111880 1 PIX6049_IN
port 6134 n
rlabel metal5 75520 -111980 75620 -111880 1 PIX6050_IN
port 6135 n
rlabel metal5 77020 -111980 77120 -111880 1 PIX6051_IN
port 6136 n
rlabel metal5 78520 -111980 78620 -111880 1 PIX6052_IN
port 6137 n
rlabel metal5 80020 -111980 80120 -111880 1 PIX6053_IN
port 6138 n
rlabel metal5 81520 -111980 81620 -111880 1 PIX6054_IN
port 6139 n
rlabel metal5 83020 -111980 83120 -111880 1 PIX6055_IN
port 6140 n
rlabel metal5 84520 -111980 84620 -111880 1 PIX6056_IN
port 6141 n
rlabel metal5 86020 -111980 86120 -111880 1 PIX6057_IN
port 6142 n
rlabel metal5 87520 -111980 87620 -111880 1 PIX6058_IN
port 6143 n
rlabel metal5 89020 -111980 89120 -111880 1 PIX6059_IN
port 6144 n
rlabel metal5 90520 -111980 90620 -111880 1 PIX6060_IN
port 6145 n
rlabel metal5 92020 -111980 92120 -111880 1 PIX6061_IN
port 6146 n
rlabel metal5 93520 -111980 93620 -111880 1 PIX6062_IN
port 6147 n
rlabel metal5 95020 -111980 95120 -111880 1 PIX6063_IN
port 6148 n
rlabel metal5 96520 -111980 96620 -111880 1 PIX6064_IN
port 6149 n
rlabel metal5 98020 -111980 98120 -111880 1 PIX6065_IN
port 6150 n
rlabel metal5 99520 -111980 99620 -111880 1 PIX6066_IN
port 6151 n
rlabel metal5 101020 -111980 101120 -111880 1 PIX6067_IN
port 6152 n
rlabel metal5 102520 -111980 102620 -111880 1 PIX6068_IN
port 6153 n
rlabel metal5 104020 -111980 104120 -111880 1 PIX6069_IN
port 6154 n
rlabel metal5 105520 -111980 105620 -111880 1 PIX6070_IN
port 6155 n
rlabel metal5 107020 -111980 107120 -111880 1 PIX6071_IN
port 6156 n
rlabel metal5 108520 -111980 108620 -111880 1 PIX6072_IN
port 6157 n
rlabel metal5 110020 -111980 110120 -111880 1 PIX6073_IN
port 6158 n
rlabel metal5 111520 -111980 111620 -111880 1 PIX6074_IN
port 6159 n
rlabel metal5 113020 -111980 113120 -111880 1 PIX6075_IN
port 6160 n
rlabel metal5 114520 -111980 114620 -111880 1 PIX6076_IN
port 6161 n
rlabel metal5 116020 -111980 116120 -111880 1 PIX6077_IN
port 6162 n
rlabel metal5 117520 -111980 117620 -111880 1 PIX6078_IN
port 6163 n
rlabel metal5 119020 -111980 119120 -111880 1 PIX6079_IN
port 6164 n
rlabel metal5 520 -113480 620 -113380 1 PIX6080_IN
port 6165 n
rlabel metal2 -1500 -113260 -1500 -113215 3 ROW_SEL76
port 6166 e
rlabel metal5 2020 -113480 2120 -113380 1 PIX6081_IN
port 6167 n
rlabel metal5 3520 -113480 3620 -113380 1 PIX6082_IN
port 6168 n
rlabel metal5 5020 -113480 5120 -113380 1 PIX6083_IN
port 6169 n
rlabel metal5 6520 -113480 6620 -113380 1 PIX6084_IN
port 6170 n
rlabel metal5 8020 -113480 8120 -113380 1 PIX6085_IN
port 6171 n
rlabel metal5 9520 -113480 9620 -113380 1 PIX6086_IN
port 6172 n
rlabel metal5 11020 -113480 11120 -113380 1 PIX6087_IN
port 6173 n
rlabel metal5 12520 -113480 12620 -113380 1 PIX6088_IN
port 6174 n
rlabel metal5 14020 -113480 14120 -113380 1 PIX6089_IN
port 6175 n
rlabel metal5 15520 -113480 15620 -113380 1 PIX6090_IN
port 6176 n
rlabel metal5 17020 -113480 17120 -113380 1 PIX6091_IN
port 6177 n
rlabel metal5 18520 -113480 18620 -113380 1 PIX6092_IN
port 6178 n
rlabel metal5 20020 -113480 20120 -113380 1 PIX6093_IN
port 6179 n
rlabel metal5 21520 -113480 21620 -113380 1 PIX6094_IN
port 6180 n
rlabel metal5 23020 -113480 23120 -113380 1 PIX6095_IN
port 6181 n
rlabel metal5 24520 -113480 24620 -113380 1 PIX6096_IN
port 6182 n
rlabel metal5 26020 -113480 26120 -113380 1 PIX6097_IN
port 6183 n
rlabel metal5 27520 -113480 27620 -113380 1 PIX6098_IN
port 6184 n
rlabel metal5 29020 -113480 29120 -113380 1 PIX6099_IN
port 6185 n
rlabel metal5 30520 -113480 30620 -113380 1 PIX6100_IN
port 6186 n
rlabel metal5 32020 -113480 32120 -113380 1 PIX6101_IN
port 6187 n
rlabel metal5 33520 -113480 33620 -113380 1 PIX6102_IN
port 6188 n
rlabel metal5 35020 -113480 35120 -113380 1 PIX6103_IN
port 6189 n
rlabel metal5 36520 -113480 36620 -113380 1 PIX6104_IN
port 6190 n
rlabel metal5 38020 -113480 38120 -113380 1 PIX6105_IN
port 6191 n
rlabel metal5 39520 -113480 39620 -113380 1 PIX6106_IN
port 6192 n
rlabel metal5 41020 -113480 41120 -113380 1 PIX6107_IN
port 6193 n
rlabel metal5 42520 -113480 42620 -113380 1 PIX6108_IN
port 6194 n
rlabel metal5 44020 -113480 44120 -113380 1 PIX6109_IN
port 6195 n
rlabel metal5 45520 -113480 45620 -113380 1 PIX6110_IN
port 6196 n
rlabel metal5 47020 -113480 47120 -113380 1 PIX6111_IN
port 6197 n
rlabel metal5 48520 -113480 48620 -113380 1 PIX6112_IN
port 6198 n
rlabel metal5 50020 -113480 50120 -113380 1 PIX6113_IN
port 6199 n
rlabel metal5 51520 -113480 51620 -113380 1 PIX6114_IN
port 6200 n
rlabel metal5 53020 -113480 53120 -113380 1 PIX6115_IN
port 6201 n
rlabel metal5 54520 -113480 54620 -113380 1 PIX6116_IN
port 6202 n
rlabel metal5 56020 -113480 56120 -113380 1 PIX6117_IN
port 6203 n
rlabel metal5 57520 -113480 57620 -113380 1 PIX6118_IN
port 6204 n
rlabel metal5 59020 -113480 59120 -113380 1 PIX6119_IN
port 6205 n
rlabel metal5 60520 -113480 60620 -113380 1 PIX6120_IN
port 6206 n
rlabel metal5 62020 -113480 62120 -113380 1 PIX6121_IN
port 6207 n
rlabel metal5 63520 -113480 63620 -113380 1 PIX6122_IN
port 6208 n
rlabel metal5 65020 -113480 65120 -113380 1 PIX6123_IN
port 6209 n
rlabel metal5 66520 -113480 66620 -113380 1 PIX6124_IN
port 6210 n
rlabel metal5 68020 -113480 68120 -113380 1 PIX6125_IN
port 6211 n
rlabel metal5 69520 -113480 69620 -113380 1 PIX6126_IN
port 6212 n
rlabel metal5 71020 -113480 71120 -113380 1 PIX6127_IN
port 6213 n
rlabel metal5 72520 -113480 72620 -113380 1 PIX6128_IN
port 6214 n
rlabel metal5 74020 -113480 74120 -113380 1 PIX6129_IN
port 6215 n
rlabel metal5 75520 -113480 75620 -113380 1 PIX6130_IN
port 6216 n
rlabel metal5 77020 -113480 77120 -113380 1 PIX6131_IN
port 6217 n
rlabel metal5 78520 -113480 78620 -113380 1 PIX6132_IN
port 6218 n
rlabel metal5 80020 -113480 80120 -113380 1 PIX6133_IN
port 6219 n
rlabel metal5 81520 -113480 81620 -113380 1 PIX6134_IN
port 6220 n
rlabel metal5 83020 -113480 83120 -113380 1 PIX6135_IN
port 6221 n
rlabel metal5 84520 -113480 84620 -113380 1 PIX6136_IN
port 6222 n
rlabel metal5 86020 -113480 86120 -113380 1 PIX6137_IN
port 6223 n
rlabel metal5 87520 -113480 87620 -113380 1 PIX6138_IN
port 6224 n
rlabel metal5 89020 -113480 89120 -113380 1 PIX6139_IN
port 6225 n
rlabel metal5 90520 -113480 90620 -113380 1 PIX6140_IN
port 6226 n
rlabel metal5 92020 -113480 92120 -113380 1 PIX6141_IN
port 6227 n
rlabel metal5 93520 -113480 93620 -113380 1 PIX6142_IN
port 6228 n
rlabel metal5 95020 -113480 95120 -113380 1 PIX6143_IN
port 6229 n
rlabel metal5 96520 -113480 96620 -113380 1 PIX6144_IN
port 6230 n
rlabel metal5 98020 -113480 98120 -113380 1 PIX6145_IN
port 6231 n
rlabel metal5 99520 -113480 99620 -113380 1 PIX6146_IN
port 6232 n
rlabel metal5 101020 -113480 101120 -113380 1 PIX6147_IN
port 6233 n
rlabel metal5 102520 -113480 102620 -113380 1 PIX6148_IN
port 6234 n
rlabel metal5 104020 -113480 104120 -113380 1 PIX6149_IN
port 6235 n
rlabel metal5 105520 -113480 105620 -113380 1 PIX6150_IN
port 6236 n
rlabel metal5 107020 -113480 107120 -113380 1 PIX6151_IN
port 6237 n
rlabel metal5 108520 -113480 108620 -113380 1 PIX6152_IN
port 6238 n
rlabel metal5 110020 -113480 110120 -113380 1 PIX6153_IN
port 6239 n
rlabel metal5 111520 -113480 111620 -113380 1 PIX6154_IN
port 6240 n
rlabel metal5 113020 -113480 113120 -113380 1 PIX6155_IN
port 6241 n
rlabel metal5 114520 -113480 114620 -113380 1 PIX6156_IN
port 6242 n
rlabel metal5 116020 -113480 116120 -113380 1 PIX6157_IN
port 6243 n
rlabel metal5 117520 -113480 117620 -113380 1 PIX6158_IN
port 6244 n
rlabel metal5 119020 -113480 119120 -113380 1 PIX6159_IN
port 6245 n
rlabel metal5 520 -114980 620 -114880 1 PIX6160_IN
port 6246 n
rlabel metal2 -1500 -114760 -1500 -114715 3 ROW_SEL77
port 6247 e
rlabel metal5 2020 -114980 2120 -114880 1 PIX6161_IN
port 6248 n
rlabel metal5 3520 -114980 3620 -114880 1 PIX6162_IN
port 6249 n
rlabel metal5 5020 -114980 5120 -114880 1 PIX6163_IN
port 6250 n
rlabel metal5 6520 -114980 6620 -114880 1 PIX6164_IN
port 6251 n
rlabel metal5 8020 -114980 8120 -114880 1 PIX6165_IN
port 6252 n
rlabel metal5 9520 -114980 9620 -114880 1 PIX6166_IN
port 6253 n
rlabel metal5 11020 -114980 11120 -114880 1 PIX6167_IN
port 6254 n
rlabel metal5 12520 -114980 12620 -114880 1 PIX6168_IN
port 6255 n
rlabel metal5 14020 -114980 14120 -114880 1 PIX6169_IN
port 6256 n
rlabel metal5 15520 -114980 15620 -114880 1 PIX6170_IN
port 6257 n
rlabel metal5 17020 -114980 17120 -114880 1 PIX6171_IN
port 6258 n
rlabel metal5 18520 -114980 18620 -114880 1 PIX6172_IN
port 6259 n
rlabel metal5 20020 -114980 20120 -114880 1 PIX6173_IN
port 6260 n
rlabel metal5 21520 -114980 21620 -114880 1 PIX6174_IN
port 6261 n
rlabel metal5 23020 -114980 23120 -114880 1 PIX6175_IN
port 6262 n
rlabel metal5 24520 -114980 24620 -114880 1 PIX6176_IN
port 6263 n
rlabel metal5 26020 -114980 26120 -114880 1 PIX6177_IN
port 6264 n
rlabel metal5 27520 -114980 27620 -114880 1 PIX6178_IN
port 6265 n
rlabel metal5 29020 -114980 29120 -114880 1 PIX6179_IN
port 6266 n
rlabel metal5 30520 -114980 30620 -114880 1 PIX6180_IN
port 6267 n
rlabel metal5 32020 -114980 32120 -114880 1 PIX6181_IN
port 6268 n
rlabel metal5 33520 -114980 33620 -114880 1 PIX6182_IN
port 6269 n
rlabel metal5 35020 -114980 35120 -114880 1 PIX6183_IN
port 6270 n
rlabel metal5 36520 -114980 36620 -114880 1 PIX6184_IN
port 6271 n
rlabel metal5 38020 -114980 38120 -114880 1 PIX6185_IN
port 6272 n
rlabel metal5 39520 -114980 39620 -114880 1 PIX6186_IN
port 6273 n
rlabel metal5 41020 -114980 41120 -114880 1 PIX6187_IN
port 6274 n
rlabel metal5 42520 -114980 42620 -114880 1 PIX6188_IN
port 6275 n
rlabel metal5 44020 -114980 44120 -114880 1 PIX6189_IN
port 6276 n
rlabel metal5 45520 -114980 45620 -114880 1 PIX6190_IN
port 6277 n
rlabel metal5 47020 -114980 47120 -114880 1 PIX6191_IN
port 6278 n
rlabel metal5 48520 -114980 48620 -114880 1 PIX6192_IN
port 6279 n
rlabel metal5 50020 -114980 50120 -114880 1 PIX6193_IN
port 6280 n
rlabel metal5 51520 -114980 51620 -114880 1 PIX6194_IN
port 6281 n
rlabel metal5 53020 -114980 53120 -114880 1 PIX6195_IN
port 6282 n
rlabel metal5 54520 -114980 54620 -114880 1 PIX6196_IN
port 6283 n
rlabel metal5 56020 -114980 56120 -114880 1 PIX6197_IN
port 6284 n
rlabel metal5 57520 -114980 57620 -114880 1 PIX6198_IN
port 6285 n
rlabel metal5 59020 -114980 59120 -114880 1 PIX6199_IN
port 6286 n
rlabel metal5 60520 -114980 60620 -114880 1 PIX6200_IN
port 6287 n
rlabel metal5 62020 -114980 62120 -114880 1 PIX6201_IN
port 6288 n
rlabel metal5 63520 -114980 63620 -114880 1 PIX6202_IN
port 6289 n
rlabel metal5 65020 -114980 65120 -114880 1 PIX6203_IN
port 6290 n
rlabel metal5 66520 -114980 66620 -114880 1 PIX6204_IN
port 6291 n
rlabel metal5 68020 -114980 68120 -114880 1 PIX6205_IN
port 6292 n
rlabel metal5 69520 -114980 69620 -114880 1 PIX6206_IN
port 6293 n
rlabel metal5 71020 -114980 71120 -114880 1 PIX6207_IN
port 6294 n
rlabel metal5 72520 -114980 72620 -114880 1 PIX6208_IN
port 6295 n
rlabel metal5 74020 -114980 74120 -114880 1 PIX6209_IN
port 6296 n
rlabel metal5 75520 -114980 75620 -114880 1 PIX6210_IN
port 6297 n
rlabel metal5 77020 -114980 77120 -114880 1 PIX6211_IN
port 6298 n
rlabel metal5 78520 -114980 78620 -114880 1 PIX6212_IN
port 6299 n
rlabel metal5 80020 -114980 80120 -114880 1 PIX6213_IN
port 6300 n
rlabel metal5 81520 -114980 81620 -114880 1 PIX6214_IN
port 6301 n
rlabel metal5 83020 -114980 83120 -114880 1 PIX6215_IN
port 6302 n
rlabel metal5 84520 -114980 84620 -114880 1 PIX6216_IN
port 6303 n
rlabel metal5 86020 -114980 86120 -114880 1 PIX6217_IN
port 6304 n
rlabel metal5 87520 -114980 87620 -114880 1 PIX6218_IN
port 6305 n
rlabel metal5 89020 -114980 89120 -114880 1 PIX6219_IN
port 6306 n
rlabel metal5 90520 -114980 90620 -114880 1 PIX6220_IN
port 6307 n
rlabel metal5 92020 -114980 92120 -114880 1 PIX6221_IN
port 6308 n
rlabel metal5 93520 -114980 93620 -114880 1 PIX6222_IN
port 6309 n
rlabel metal5 95020 -114980 95120 -114880 1 PIX6223_IN
port 6310 n
rlabel metal5 96520 -114980 96620 -114880 1 PIX6224_IN
port 6311 n
rlabel metal5 98020 -114980 98120 -114880 1 PIX6225_IN
port 6312 n
rlabel metal5 99520 -114980 99620 -114880 1 PIX6226_IN
port 6313 n
rlabel metal5 101020 -114980 101120 -114880 1 PIX6227_IN
port 6314 n
rlabel metal5 102520 -114980 102620 -114880 1 PIX6228_IN
port 6315 n
rlabel metal5 104020 -114980 104120 -114880 1 PIX6229_IN
port 6316 n
rlabel metal5 105520 -114980 105620 -114880 1 PIX6230_IN
port 6317 n
rlabel metal5 107020 -114980 107120 -114880 1 PIX6231_IN
port 6318 n
rlabel metal5 108520 -114980 108620 -114880 1 PIX6232_IN
port 6319 n
rlabel metal5 110020 -114980 110120 -114880 1 PIX6233_IN
port 6320 n
rlabel metal5 111520 -114980 111620 -114880 1 PIX6234_IN
port 6321 n
rlabel metal5 113020 -114980 113120 -114880 1 PIX6235_IN
port 6322 n
rlabel metal5 114520 -114980 114620 -114880 1 PIX6236_IN
port 6323 n
rlabel metal5 116020 -114980 116120 -114880 1 PIX6237_IN
port 6324 n
rlabel metal5 117520 -114980 117620 -114880 1 PIX6238_IN
port 6325 n
rlabel metal5 119020 -114980 119120 -114880 1 PIX6239_IN
port 6326 n
rlabel metal5 520 -116480 620 -116380 1 PIX6240_IN
port 6327 n
rlabel metal2 -1500 -116260 -1500 -116215 3 ROW_SEL78
port 6328 e
rlabel metal5 2020 -116480 2120 -116380 1 PIX6241_IN
port 6329 n
rlabel metal5 3520 -116480 3620 -116380 1 PIX6242_IN
port 6330 n
rlabel metal5 5020 -116480 5120 -116380 1 PIX6243_IN
port 6331 n
rlabel metal5 6520 -116480 6620 -116380 1 PIX6244_IN
port 6332 n
rlabel metal5 8020 -116480 8120 -116380 1 PIX6245_IN
port 6333 n
rlabel metal5 9520 -116480 9620 -116380 1 PIX6246_IN
port 6334 n
rlabel metal5 11020 -116480 11120 -116380 1 PIX6247_IN
port 6335 n
rlabel metal5 12520 -116480 12620 -116380 1 PIX6248_IN
port 6336 n
rlabel metal5 14020 -116480 14120 -116380 1 PIX6249_IN
port 6337 n
rlabel metal5 15520 -116480 15620 -116380 1 PIX6250_IN
port 6338 n
rlabel metal5 17020 -116480 17120 -116380 1 PIX6251_IN
port 6339 n
rlabel metal5 18520 -116480 18620 -116380 1 PIX6252_IN
port 6340 n
rlabel metal5 20020 -116480 20120 -116380 1 PIX6253_IN
port 6341 n
rlabel metal5 21520 -116480 21620 -116380 1 PIX6254_IN
port 6342 n
rlabel metal5 23020 -116480 23120 -116380 1 PIX6255_IN
port 6343 n
rlabel metal5 24520 -116480 24620 -116380 1 PIX6256_IN
port 6344 n
rlabel metal5 26020 -116480 26120 -116380 1 PIX6257_IN
port 6345 n
rlabel metal5 27520 -116480 27620 -116380 1 PIX6258_IN
port 6346 n
rlabel metal5 29020 -116480 29120 -116380 1 PIX6259_IN
port 6347 n
rlabel metal5 30520 -116480 30620 -116380 1 PIX6260_IN
port 6348 n
rlabel metal5 32020 -116480 32120 -116380 1 PIX6261_IN
port 6349 n
rlabel metal5 33520 -116480 33620 -116380 1 PIX6262_IN
port 6350 n
rlabel metal5 35020 -116480 35120 -116380 1 PIX6263_IN
port 6351 n
rlabel metal5 36520 -116480 36620 -116380 1 PIX6264_IN
port 6352 n
rlabel metal5 38020 -116480 38120 -116380 1 PIX6265_IN
port 6353 n
rlabel metal5 39520 -116480 39620 -116380 1 PIX6266_IN
port 6354 n
rlabel metal5 41020 -116480 41120 -116380 1 PIX6267_IN
port 6355 n
rlabel metal5 42520 -116480 42620 -116380 1 PIX6268_IN
port 6356 n
rlabel metal5 44020 -116480 44120 -116380 1 PIX6269_IN
port 6357 n
rlabel metal5 45520 -116480 45620 -116380 1 PIX6270_IN
port 6358 n
rlabel metal5 47020 -116480 47120 -116380 1 PIX6271_IN
port 6359 n
rlabel metal5 48520 -116480 48620 -116380 1 PIX6272_IN
port 6360 n
rlabel metal5 50020 -116480 50120 -116380 1 PIX6273_IN
port 6361 n
rlabel metal5 51520 -116480 51620 -116380 1 PIX6274_IN
port 6362 n
rlabel metal5 53020 -116480 53120 -116380 1 PIX6275_IN
port 6363 n
rlabel metal5 54520 -116480 54620 -116380 1 PIX6276_IN
port 6364 n
rlabel metal5 56020 -116480 56120 -116380 1 PIX6277_IN
port 6365 n
rlabel metal5 57520 -116480 57620 -116380 1 PIX6278_IN
port 6366 n
rlabel metal5 59020 -116480 59120 -116380 1 PIX6279_IN
port 6367 n
rlabel metal5 60520 -116480 60620 -116380 1 PIX6280_IN
port 6368 n
rlabel metal5 62020 -116480 62120 -116380 1 PIX6281_IN
port 6369 n
rlabel metal5 63520 -116480 63620 -116380 1 PIX6282_IN
port 6370 n
rlabel metal5 65020 -116480 65120 -116380 1 PIX6283_IN
port 6371 n
rlabel metal5 66520 -116480 66620 -116380 1 PIX6284_IN
port 6372 n
rlabel metal5 68020 -116480 68120 -116380 1 PIX6285_IN
port 6373 n
rlabel metal5 69520 -116480 69620 -116380 1 PIX6286_IN
port 6374 n
rlabel metal5 71020 -116480 71120 -116380 1 PIX6287_IN
port 6375 n
rlabel metal5 72520 -116480 72620 -116380 1 PIX6288_IN
port 6376 n
rlabel metal5 74020 -116480 74120 -116380 1 PIX6289_IN
port 6377 n
rlabel metal5 75520 -116480 75620 -116380 1 PIX6290_IN
port 6378 n
rlabel metal5 77020 -116480 77120 -116380 1 PIX6291_IN
port 6379 n
rlabel metal5 78520 -116480 78620 -116380 1 PIX6292_IN
port 6380 n
rlabel metal5 80020 -116480 80120 -116380 1 PIX6293_IN
port 6381 n
rlabel metal5 81520 -116480 81620 -116380 1 PIX6294_IN
port 6382 n
rlabel metal5 83020 -116480 83120 -116380 1 PIX6295_IN
port 6383 n
rlabel metal5 84520 -116480 84620 -116380 1 PIX6296_IN
port 6384 n
rlabel metal5 86020 -116480 86120 -116380 1 PIX6297_IN
port 6385 n
rlabel metal5 87520 -116480 87620 -116380 1 PIX6298_IN
port 6386 n
rlabel metal5 89020 -116480 89120 -116380 1 PIX6299_IN
port 6387 n
rlabel metal5 90520 -116480 90620 -116380 1 PIX6300_IN
port 6388 n
rlabel metal5 92020 -116480 92120 -116380 1 PIX6301_IN
port 6389 n
rlabel metal5 93520 -116480 93620 -116380 1 PIX6302_IN
port 6390 n
rlabel metal5 95020 -116480 95120 -116380 1 PIX6303_IN
port 6391 n
rlabel metal5 96520 -116480 96620 -116380 1 PIX6304_IN
port 6392 n
rlabel metal5 98020 -116480 98120 -116380 1 PIX6305_IN
port 6393 n
rlabel metal5 99520 -116480 99620 -116380 1 PIX6306_IN
port 6394 n
rlabel metal5 101020 -116480 101120 -116380 1 PIX6307_IN
port 6395 n
rlabel metal5 102520 -116480 102620 -116380 1 PIX6308_IN
port 6396 n
rlabel metal5 104020 -116480 104120 -116380 1 PIX6309_IN
port 6397 n
rlabel metal5 105520 -116480 105620 -116380 1 PIX6310_IN
port 6398 n
rlabel metal5 107020 -116480 107120 -116380 1 PIX6311_IN
port 6399 n
rlabel metal5 108520 -116480 108620 -116380 1 PIX6312_IN
port 6400 n
rlabel metal5 110020 -116480 110120 -116380 1 PIX6313_IN
port 6401 n
rlabel metal5 111520 -116480 111620 -116380 1 PIX6314_IN
port 6402 n
rlabel metal5 113020 -116480 113120 -116380 1 PIX6315_IN
port 6403 n
rlabel metal5 114520 -116480 114620 -116380 1 PIX6316_IN
port 6404 n
rlabel metal5 116020 -116480 116120 -116380 1 PIX6317_IN
port 6405 n
rlabel metal5 117520 -116480 117620 -116380 1 PIX6318_IN
port 6406 n
rlabel metal5 119020 -116480 119120 -116380 1 PIX6319_IN
port 6407 n
rlabel metal5 520 -117980 620 -117880 1 PIX6320_IN
port 6408 n
rlabel metal4 1315 -118600 1390 -118500 1 PIX_OUT0
port 6409 n
rlabel metal4 110 -119050 220 -118850 1 COL_SEL0
port 6410 n
rlabel metal4 -240 -119300 -240 -119300 1 CSA_VREF
port 6411 n
rlabel metal2 -1500 -117760 -1500 -117715 3 ROW_SEL79
port 6412 e
rlabel metal5 2020 -117980 2120 -117880 1 PIX6321_IN
port 6413 n
rlabel metal4 2815 -118600 2890 -118500 1 PIX_OUT1
port 6414 n
rlabel metal4 1610 -119050 1720 -118850 1 COL_SEL1
port 6415 n
rlabel metal5 3520 -117980 3620 -117880 1 PIX6322_IN
port 6416 n
rlabel metal4 4315 -118600 4390 -118500 1 PIX_OUT2
port 6417 n
rlabel metal4 3110 -119050 3220 -118850 1 COL_SEL2
port 6418 n
rlabel metal5 5020 -117980 5120 -117880 1 PIX6323_IN
port 6419 n
rlabel metal4 5815 -118600 5890 -118500 1 PIX_OUT3
port 6420 n
rlabel metal4 4610 -119050 4720 -118850 1 COL_SEL3
port 6421 n
rlabel metal5 6520 -117980 6620 -117880 1 PIX6324_IN
port 6422 n
rlabel metal4 7315 -118600 7390 -118500 1 PIX_OUT4
port 6423 n
rlabel metal4 6110 -119050 6220 -118850 1 COL_SEL4
port 6424 n
rlabel metal5 8020 -117980 8120 -117880 1 PIX6325_IN
port 6425 n
rlabel metal4 8815 -118600 8890 -118500 1 PIX_OUT5
port 6426 n
rlabel metal4 7610 -119050 7720 -118850 1 COL_SEL5
port 6427 n
rlabel metal5 9520 -117980 9620 -117880 1 PIX6326_IN
port 6428 n
rlabel metal4 10315 -118600 10390 -118500 1 PIX_OUT6
port 6429 n
rlabel metal4 9110 -119050 9220 -118850 1 COL_SEL6
port 6430 n
rlabel metal5 11020 -117980 11120 -117880 1 PIX6327_IN
port 6431 n
rlabel metal4 11815 -118600 11890 -118500 1 PIX_OUT7
port 6432 n
rlabel metal4 10610 -119050 10720 -118850 1 COL_SEL7
port 6433 n
rlabel metal5 12520 -117980 12620 -117880 1 PIX6328_IN
port 6434 n
rlabel metal4 13315 -118600 13390 -118500 1 PIX_OUT8
port 6435 n
rlabel metal4 12110 -119050 12220 -118850 1 COL_SEL8
port 6436 n
rlabel metal5 14020 -117980 14120 -117880 1 PIX6329_IN
port 6437 n
rlabel metal4 14815 -118600 14890 -118500 1 PIX_OUT9
port 6438 n
rlabel metal4 13610 -119050 13720 -118850 1 COL_SEL9
port 6439 n
rlabel metal5 15520 -117980 15620 -117880 1 PIX6330_IN
port 6440 n
rlabel metal4 16315 -118600 16390 -118500 1 PIX_OUT10
port 6441 n
rlabel metal4 15110 -119050 15220 -118850 1 COL_SEL10
port 6442 n
rlabel metal5 17020 -117980 17120 -117880 1 PIX6331_IN
port 6443 n
rlabel metal4 17815 -118600 17890 -118500 1 PIX_OUT11
port 6444 n
rlabel metal4 16610 -119050 16720 -118850 1 COL_SEL11
port 6445 n
rlabel metal5 18520 -117980 18620 -117880 1 PIX6332_IN
port 6446 n
rlabel metal4 19315 -118600 19390 -118500 1 PIX_OUT12
port 6447 n
rlabel metal4 18110 -119050 18220 -118850 1 COL_SEL12
port 6448 n
rlabel metal5 20020 -117980 20120 -117880 1 PIX6333_IN
port 6449 n
rlabel metal4 20815 -118600 20890 -118500 1 PIX_OUT13
port 6450 n
rlabel metal4 19610 -119050 19720 -118850 1 COL_SEL13
port 6451 n
rlabel metal5 21520 -117980 21620 -117880 1 PIX6334_IN
port 6452 n
rlabel metal4 22315 -118600 22390 -118500 1 PIX_OUT14
port 6453 n
rlabel metal4 21110 -119050 21220 -118850 1 COL_SEL14
port 6454 n
rlabel metal5 23020 -117980 23120 -117880 1 PIX6335_IN
port 6455 n
rlabel metal4 23815 -118600 23890 -118500 1 PIX_OUT15
port 6456 n
rlabel metal4 22610 -119050 22720 -118850 1 COL_SEL15
port 6457 n
rlabel metal5 24520 -117980 24620 -117880 1 PIX6336_IN
port 6458 n
rlabel metal4 25315 -118600 25390 -118500 1 PIX_OUT16
port 6459 n
rlabel metal4 24110 -119050 24220 -118850 1 COL_SEL16
port 6460 n
rlabel metal5 26020 -117980 26120 -117880 1 PIX6337_IN
port 6461 n
rlabel metal4 26815 -118600 26890 -118500 1 PIX_OUT17
port 6462 n
rlabel metal4 25610 -119050 25720 -118850 1 COL_SEL17
port 6463 n
rlabel metal5 27520 -117980 27620 -117880 1 PIX6338_IN
port 6464 n
rlabel metal4 28315 -118600 28390 -118500 1 PIX_OUT18
port 6465 n
rlabel metal4 27110 -119050 27220 -118850 1 COL_SEL18
port 6466 n
rlabel metal5 29020 -117980 29120 -117880 1 PIX6339_IN
port 6467 n
rlabel metal4 29815 -118600 29890 -118500 1 PIX_OUT19
port 6468 n
rlabel metal4 28610 -119050 28720 -118850 1 COL_SEL19
port 6469 n
rlabel metal5 30520 -117980 30620 -117880 1 PIX6340_IN
port 6470 n
rlabel metal4 31315 -118600 31390 -118500 1 PIX_OUT20
port 6471 n
rlabel metal4 30110 -119050 30220 -118850 1 COL_SEL20
port 6472 n
rlabel metal5 32020 -117980 32120 -117880 1 PIX6341_IN
port 6473 n
rlabel metal4 32815 -118600 32890 -118500 1 PIX_OUT21
port 6474 n
rlabel metal4 31610 -119050 31720 -118850 1 COL_SEL21
port 6475 n
rlabel metal5 33520 -117980 33620 -117880 1 PIX6342_IN
port 6476 n
rlabel metal4 34315 -118600 34390 -118500 1 PIX_OUT22
port 6477 n
rlabel metal4 33110 -119050 33220 -118850 1 COL_SEL22
port 6478 n
rlabel metal5 35020 -117980 35120 -117880 1 PIX6343_IN
port 6479 n
rlabel metal4 35815 -118600 35890 -118500 1 PIX_OUT23
port 6480 n
rlabel metal4 34610 -119050 34720 -118850 1 COL_SEL23
port 6481 n
rlabel metal5 36520 -117980 36620 -117880 1 PIX6344_IN
port 6482 n
rlabel metal4 37315 -118600 37390 -118500 1 PIX_OUT24
port 6483 n
rlabel metal4 36110 -119050 36220 -118850 1 COL_SEL24
port 6484 n
rlabel metal5 38020 -117980 38120 -117880 1 PIX6345_IN
port 6485 n
rlabel metal4 38815 -118600 38890 -118500 1 PIX_OUT25
port 6486 n
rlabel metal4 37610 -119050 37720 -118850 1 COL_SEL25
port 6487 n
rlabel metal5 39520 -117980 39620 -117880 1 PIX6346_IN
port 6488 n
rlabel metal4 40315 -118600 40390 -118500 1 PIX_OUT26
port 6489 n
rlabel metal4 39110 -119050 39220 -118850 1 COL_SEL26
port 6490 n
rlabel metal5 41020 -117980 41120 -117880 1 PIX6347_IN
port 6491 n
rlabel metal4 41815 -118600 41890 -118500 1 PIX_OUT27
port 6492 n
rlabel metal4 40610 -119050 40720 -118850 1 COL_SEL27
port 6493 n
rlabel metal5 42520 -117980 42620 -117880 1 PIX6348_IN
port 6494 n
rlabel metal4 43315 -118600 43390 -118500 1 PIX_OUT28
port 6495 n
rlabel metal4 42110 -119050 42220 -118850 1 COL_SEL28
port 6496 n
rlabel metal5 44020 -117980 44120 -117880 1 PIX6349_IN
port 6497 n
rlabel metal4 44815 -118600 44890 -118500 1 PIX_OUT29
port 6498 n
rlabel metal4 43610 -119050 43720 -118850 1 COL_SEL29
port 6499 n
rlabel metal5 45520 -117980 45620 -117880 1 PIX6350_IN
port 6500 n
rlabel metal4 46315 -118600 46390 -118500 1 PIX_OUT30
port 6501 n
rlabel metal4 45110 -119050 45220 -118850 1 COL_SEL30
port 6502 n
rlabel metal5 47020 -117980 47120 -117880 1 PIX6351_IN
port 6503 n
rlabel metal4 47815 -118600 47890 -118500 1 PIX_OUT31
port 6504 n
rlabel metal4 46610 -119050 46720 -118850 1 COL_SEL31
port 6505 n
rlabel metal5 48520 -117980 48620 -117880 1 PIX6352_IN
port 6506 n
rlabel metal4 49315 -118600 49390 -118500 1 PIX_OUT32
port 6507 n
rlabel metal4 48110 -119050 48220 -118850 1 COL_SEL32
port 6508 n
rlabel metal5 50020 -117980 50120 -117880 1 PIX6353_IN
port 6509 n
rlabel metal4 50815 -118600 50890 -118500 1 PIX_OUT33
port 6510 n
rlabel metal4 49610 -119050 49720 -118850 1 COL_SEL33
port 6511 n
rlabel metal5 51520 -117980 51620 -117880 1 PIX6354_IN
port 6512 n
rlabel metal4 52315 -118600 52390 -118500 1 PIX_OUT34
port 6513 n
rlabel metal4 51110 -119050 51220 -118850 1 COL_SEL34
port 6514 n
rlabel metal5 53020 -117980 53120 -117880 1 PIX6355_IN
port 6515 n
rlabel metal4 53815 -118600 53890 -118500 1 PIX_OUT35
port 6516 n
rlabel metal4 52610 -119050 52720 -118850 1 COL_SEL35
port 6517 n
rlabel metal5 54520 -117980 54620 -117880 1 PIX6356_IN
port 6518 n
rlabel metal4 55315 -118600 55390 -118500 1 PIX_OUT36
port 6519 n
rlabel metal4 54110 -119050 54220 -118850 1 COL_SEL36
port 6520 n
rlabel metal5 56020 -117980 56120 -117880 1 PIX6357_IN
port 6521 n
rlabel metal4 56815 -118600 56890 -118500 1 PIX_OUT37
port 6522 n
rlabel metal4 55610 -119050 55720 -118850 1 COL_SEL37
port 6523 n
rlabel metal5 57520 -117980 57620 -117880 1 PIX6358_IN
port 6524 n
rlabel metal4 58315 -118600 58390 -118500 1 PIX_OUT38
port 6525 n
rlabel metal4 57110 -119050 57220 -118850 1 COL_SEL38
port 6526 n
rlabel metal5 59020 -117980 59120 -117880 1 PIX6359_IN
port 6527 n
rlabel metal4 59815 -118600 59890 -118500 1 PIX_OUT39
port 6528 n
rlabel metal4 58610 -119050 58720 -118850 1 COL_SEL39
port 6529 n
rlabel metal5 60520 -117980 60620 -117880 1 PIX6360_IN
port 6530 n
rlabel metal4 61315 -118600 61390 -118500 1 PIX_OUT40
port 6531 n
rlabel metal4 60110 -119050 60220 -118850 1 COL_SEL40
port 6532 n
rlabel metal5 62020 -117980 62120 -117880 1 PIX6361_IN
port 6533 n
rlabel metal4 62815 -118600 62890 -118500 1 PIX_OUT41
port 6534 n
rlabel metal4 61610 -119050 61720 -118850 1 COL_SEL41
port 6535 n
rlabel metal5 63520 -117980 63620 -117880 1 PIX6362_IN
port 6536 n
rlabel metal4 64315 -118600 64390 -118500 1 PIX_OUT42
port 6537 n
rlabel metal4 63110 -119050 63220 -118850 1 COL_SEL42
port 6538 n
rlabel metal5 65020 -117980 65120 -117880 1 PIX6363_IN
port 6539 n
rlabel metal4 65815 -118600 65890 -118500 1 PIX_OUT43
port 6540 n
rlabel metal4 64610 -119050 64720 -118850 1 COL_SEL43
port 6541 n
rlabel metal5 66520 -117980 66620 -117880 1 PIX6364_IN
port 6542 n
rlabel metal4 67315 -118600 67390 -118500 1 PIX_OUT44
port 6543 n
rlabel metal4 66110 -119050 66220 -118850 1 COL_SEL44
port 6544 n
rlabel metal5 68020 -117980 68120 -117880 1 PIX6365_IN
port 6545 n
rlabel metal4 68815 -118600 68890 -118500 1 PIX_OUT45
port 6546 n
rlabel metal4 67610 -119050 67720 -118850 1 COL_SEL45
port 6547 n
rlabel metal5 69520 -117980 69620 -117880 1 PIX6366_IN
port 6548 n
rlabel metal4 70315 -118600 70390 -118500 1 PIX_OUT46
port 6549 n
rlabel metal4 69110 -119050 69220 -118850 1 COL_SEL46
port 6550 n
rlabel metal5 71020 -117980 71120 -117880 1 PIX6367_IN
port 6551 n
rlabel metal4 71815 -118600 71890 -118500 1 PIX_OUT47
port 6552 n
rlabel metal4 70610 -119050 70720 -118850 1 COL_SEL47
port 6553 n
rlabel metal5 72520 -117980 72620 -117880 1 PIX6368_IN
port 6554 n
rlabel metal4 73315 -118600 73390 -118500 1 PIX_OUT48
port 6555 n
rlabel metal4 72110 -119050 72220 -118850 1 COL_SEL48
port 6556 n
rlabel metal5 74020 -117980 74120 -117880 1 PIX6369_IN
port 6557 n
rlabel metal4 74815 -118600 74890 -118500 1 PIX_OUT49
port 6558 n
rlabel metal4 73610 -119050 73720 -118850 1 COL_SEL49
port 6559 n
rlabel metal5 75520 -117980 75620 -117880 1 PIX6370_IN
port 6560 n
rlabel metal4 76315 -118600 76390 -118500 1 PIX_OUT50
port 6561 n
rlabel metal4 75110 -119050 75220 -118850 1 COL_SEL50
port 6562 n
rlabel metal5 77020 -117980 77120 -117880 1 PIX6371_IN
port 6563 n
rlabel metal4 77815 -118600 77890 -118500 1 PIX_OUT51
port 6564 n
rlabel metal4 76610 -119050 76720 -118850 1 COL_SEL51
port 6565 n
rlabel metal5 78520 -117980 78620 -117880 1 PIX6372_IN
port 6566 n
rlabel metal4 79315 -118600 79390 -118500 1 PIX_OUT52
port 6567 n
rlabel metal4 78110 -119050 78220 -118850 1 COL_SEL52
port 6568 n
rlabel metal5 80020 -117980 80120 -117880 1 PIX6373_IN
port 6569 n
rlabel metal4 80815 -118600 80890 -118500 1 PIX_OUT53
port 6570 n
rlabel metal4 79610 -119050 79720 -118850 1 COL_SEL53
port 6571 n
rlabel metal5 81520 -117980 81620 -117880 1 PIX6374_IN
port 6572 n
rlabel metal4 82315 -118600 82390 -118500 1 PIX_OUT54
port 6573 n
rlabel metal4 81110 -119050 81220 -118850 1 COL_SEL54
port 6574 n
rlabel metal5 83020 -117980 83120 -117880 1 PIX6375_IN
port 6575 n
rlabel metal4 83815 -118600 83890 -118500 1 PIX_OUT55
port 6576 n
rlabel metal4 82610 -119050 82720 -118850 1 COL_SEL55
port 6577 n
rlabel metal5 84520 -117980 84620 -117880 1 PIX6376_IN
port 6578 n
rlabel metal4 85315 -118600 85390 -118500 1 PIX_OUT56
port 6579 n
rlabel metal4 84110 -119050 84220 -118850 1 COL_SEL56
port 6580 n
rlabel metal5 86020 -117980 86120 -117880 1 PIX6377_IN
port 6581 n
rlabel metal4 86815 -118600 86890 -118500 1 PIX_OUT57
port 6582 n
rlabel metal4 85610 -119050 85720 -118850 1 COL_SEL57
port 6583 n
rlabel metal5 87520 -117980 87620 -117880 1 PIX6378_IN
port 6584 n
rlabel metal4 88315 -118600 88390 -118500 1 PIX_OUT58
port 6585 n
rlabel metal4 87110 -119050 87220 -118850 1 COL_SEL58
port 6586 n
rlabel metal5 89020 -117980 89120 -117880 1 PIX6379_IN
port 6587 n
rlabel metal4 89815 -118600 89890 -118500 1 PIX_OUT59
port 6588 n
rlabel metal4 88610 -119050 88720 -118850 1 COL_SEL59
port 6589 n
rlabel metal5 90520 -117980 90620 -117880 1 PIX6380_IN
port 6590 n
rlabel metal4 91315 -118600 91390 -118500 1 PIX_OUT60
port 6591 n
rlabel metal4 90110 -119050 90220 -118850 1 COL_SEL60
port 6592 n
rlabel metal5 92020 -117980 92120 -117880 1 PIX6381_IN
port 6593 n
rlabel metal4 92815 -118600 92890 -118500 1 PIX_OUT61
port 6594 n
rlabel metal4 91610 -119050 91720 -118850 1 COL_SEL61
port 6595 n
rlabel metal5 93520 -117980 93620 -117880 1 PIX6382_IN
port 6596 n
rlabel metal4 94315 -118600 94390 -118500 1 PIX_OUT62
port 6597 n
rlabel metal4 93110 -119050 93220 -118850 1 COL_SEL62
port 6598 n
rlabel metal5 95020 -117980 95120 -117880 1 PIX6383_IN
port 6599 n
rlabel metal4 95815 -118600 95890 -118500 1 PIX_OUT63
port 6600 n
rlabel metal4 94610 -119050 94720 -118850 1 COL_SEL63
port 6601 n
rlabel metal5 96520 -117980 96620 -117880 1 PIX6384_IN
port 6602 n
rlabel metal4 97315 -118600 97390 -118500 1 PIX_OUT64
port 6603 n
rlabel metal4 96110 -119050 96220 -118850 1 COL_SEL64
port 6604 n
rlabel metal5 98020 -117980 98120 -117880 1 PIX6385_IN
port 6605 n
rlabel metal4 98815 -118600 98890 -118500 1 PIX_OUT65
port 6606 n
rlabel metal4 97610 -119050 97720 -118850 1 COL_SEL65
port 6607 n
rlabel metal5 99520 -117980 99620 -117880 1 PIX6386_IN
port 6608 n
rlabel metal4 100315 -118600 100390 -118500 1 PIX_OUT66
port 6609 n
rlabel metal4 99110 -119050 99220 -118850 1 COL_SEL66
port 6610 n
rlabel metal5 101020 -117980 101120 -117880 1 PIX6387_IN
port 6611 n
rlabel metal4 101815 -118600 101890 -118500 1 PIX_OUT67
port 6612 n
rlabel metal4 100610 -119050 100720 -118850 1 COL_SEL67
port 6613 n
rlabel metal5 102520 -117980 102620 -117880 1 PIX6388_IN
port 6614 n
rlabel metal4 103315 -118600 103390 -118500 1 PIX_OUT68
port 6615 n
rlabel metal4 102110 -119050 102220 -118850 1 COL_SEL68
port 6616 n
rlabel metal5 104020 -117980 104120 -117880 1 PIX6389_IN
port 6617 n
rlabel metal4 104815 -118600 104890 -118500 1 PIX_OUT69
port 6618 n
rlabel metal4 103610 -119050 103720 -118850 1 COL_SEL69
port 6619 n
rlabel metal5 105520 -117980 105620 -117880 1 PIX6390_IN
port 6620 n
rlabel metal4 106315 -118600 106390 -118500 1 PIX_OUT70
port 6621 n
rlabel metal4 105110 -119050 105220 -118850 1 COL_SEL70
port 6622 n
rlabel metal5 107020 -117980 107120 -117880 1 PIX6391_IN
port 6623 n
rlabel metal4 107815 -118600 107890 -118500 1 PIX_OUT71
port 6624 n
rlabel metal4 106610 -119050 106720 -118850 1 COL_SEL71
port 6625 n
rlabel metal5 108520 -117980 108620 -117880 1 PIX6392_IN
port 6626 n
rlabel metal4 109315 -118600 109390 -118500 1 PIX_OUT72
port 6627 n
rlabel metal4 108110 -119050 108220 -118850 1 COL_SEL72
port 6628 n
rlabel metal5 110020 -117980 110120 -117880 1 PIX6393_IN
port 6629 n
rlabel metal4 110815 -118600 110890 -118500 1 PIX_OUT73
port 6630 n
rlabel metal4 109610 -119050 109720 -118850 1 COL_SEL73
port 6631 n
rlabel metal5 111520 -117980 111620 -117880 1 PIX6394_IN
port 6632 n
rlabel metal4 112315 -118600 112390 -118500 1 PIX_OUT74
port 6633 n
rlabel metal4 111110 -119050 111220 -118850 1 COL_SEL74
port 6634 n
rlabel metal5 113020 -117980 113120 -117880 1 PIX6395_IN
port 6635 n
rlabel metal4 113815 -118600 113890 -118500 1 PIX_OUT75
port 6636 n
rlabel metal4 112610 -119050 112720 -118850 1 COL_SEL75
port 6637 n
rlabel metal5 114520 -117980 114620 -117880 1 PIX6396_IN
port 6638 n
rlabel metal4 115315 -118600 115390 -118500 1 PIX_OUT76
port 6639 n
rlabel metal4 114110 -119050 114220 -118850 1 COL_SEL76
port 6640 n
rlabel metal5 116020 -117980 116120 -117880 1 PIX6397_IN
port 6641 n
rlabel metal4 116815 -118600 116890 -118500 1 PIX_OUT77
port 6642 n
rlabel metal4 115610 -119050 115720 -118850 1 COL_SEL77
port 6643 n
rlabel metal5 117520 -117980 117620 -117880 1 PIX6398_IN
port 6644 n
rlabel metal4 118315 -118600 118390 -118500 1 PIX_OUT78
port 6645 n
rlabel metal4 117110 -119050 117220 -118850 1 COL_SEL78
port 6646 n
rlabel metal5 119020 -117980 119120 -117880 1 PIX6399_IN
port 6647 n
rlabel metal4 119815 -118600 119890 -118500 1 PIX_OUT79
port 6648 n
rlabel metal2 119970 -119050 119970 -119050 1 ARRAY_OUT
port 6649 n
rlabel metal4 118610 -119050 118720 -118850 1 COL_SEL79
port 6650 n
<< end >>
