* SPICE3 file created from pixel_array.ext - technology: sky130A

.option scale=5000u

.subckt pixel_array PIX0_IN VBIAS VREF NB2 VDD SF_IB CSA_VREF NB1 ROW_SEL0 PIX1_IN
+ PIX2_IN GND PIX3_IN ROW_SEL1 PIX4_IN PIX5_IN PIX6_IN PIX_OUT0 COL_SEL0 ROW_SEL2
+ PIX7_IN PIX_OUT1 COL_SEL1 PIX8_IN PIX_OUT2 COL_SEL2
X0 PIX_OUT2 COL_SEL2 ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=256000 pd=6280 as=0 ps=0 w=1600 l=400
X1 PIX_OUT1 COL_SEL1 ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=256000 pd=6280 as=0 ps=0 w=1600 l=400
X2 PIX_OUT0 COL_SEL0 ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=142801 pd=3581 as=0 ps=0 w=1600 l=400
C0 VDD pixel_7/test 2.29fF
C1 PIX4_IN VDD 1.18fF
C2 pixel_4/net2 VDD 1.04fF
C3 VDD pixel_4/net1 1.59fF
C4 pixel_4/a_4350_10# VDD 1.49fF
C5 pixel_4/test VDD 2.18fF
C6 PIX_OUT2 CSA_VREF 1.42fF
C7 NB2 VDD 5.20fF
C8 SF_IB CSA_VREF 9.19fF
C9 VDD PIX3_IN 1.18fF
C10 VREF VDD 3.82fF
C11 VDD VBIAS 3.90fF
C12 CSA_VREF PIX5_IN 1.66fF
C13 pixel_3/net1 VDD 1.59fF
C14 VDD pixel_3/net2 1.04fF
C15 pixel_3/test VDD 2.14fF
C16 VDD pixel_3/a_4350_10# 1.48fF
C17 VDD PIX2_IN 1.18fF
C18 pixel_8/gring PIX7_IN 3.31fF
C19 VDD PIX8_IN 1.18fF
C20 NB2 NB1 1.53fF
C21 PIX4_IN CSA_VREF 1.66fF
C22 NB1 VBIAS 1.90fF
C23 pixel_8/gring PIX6_IN 3.31fF
C24 pixel_8/gring VDD 16.04fF
C25 pixel_2/net2 VDD 1.04fF
C26 pixel_2/net1 VDD 1.59fF
C27 VDD pixel_2/a_4350_10# 1.55fF
C28 pixel_2/test VDD 2.28fF
C29 CSA_VREF PIX3_IN 1.66fF
C30 CSA_VREF VREF 1.10fF
C31 PIX_OUT0 VDD 1.06fF
C32 pixel_8/gring NB1 12.68fF
C33 PIX0_IN pixel_8/gring 3.31fF
C34 pixel_7/a_4350_10# VDD 1.51fF
C35 CSA_VREF PIX2_IN 1.66fF
C36 CSA_VREF PIX8_IN 1.66fF
C37 pixel_8/net1 VDD 1.59fF
C38 PIX8_IN pixel_8/net2 1.91fF
C39 VDD PIX1_IN 1.18fF
C40 pixel_1/net2 PIX1_IN 1.91fF
C41 PIX_OUT0 NB1 1.10fF
C42 pixel_8/gring CSA_VREF 1.64fF
C43 PIX5_IN pixel_5/net2 1.91fF
C44 CSA_VREF PIX_OUT0 1.42fF
C45 PIX7_IN VDD 1.18fF
C46 CSA_VREF PIX1_IN 1.66fF
C47 PIX_OUT1 pixel_8/gring 2.82fF
C48 SF_IB VREF 1.94fF
C49 VDD PIX6_IN 1.18fF
C50 VDD pixel_1/net1 1.59fF
C51 VDD pixel_1/net2 1.04fF
C52 PIX4_IN pixel_4/net2 1.91fF
C53 pixel_8/a_4350_10# VDD 1.55fF
C54 pixel_1/a_4350_10# VDD 1.51fF
C55 VDD pixel_1/test 2.29fF
C56 PIX_OUT2 pixel_8/gring 3.78fF
C57 SF_IB pixel_8/gring 2.95fF
C58 PIX0_IN VDD 1.18fF
C59 pixel_8/gring PIX5_IN 3.31fF
C60 PIX7_IN CSA_VREF 1.66fF
C61 VREF VBIAS 4.55fF
C62 CSA_VREF PIX6_IN 1.66fF
C63 CSA_VREF VDD 22.94fF
C64 pixel_3/net2 PIX3_IN 1.91fF
C65 PIX4_IN pixel_8/gring 3.31fF
C66 VDD pixel_8/net2 1.04fF
C67 pixel_8/gring NB2 1.05fF
C68 pixel_8/gring PIX3_IN 3.31fF
C69 PIX0_IN CSA_VREF 1.66fF
C70 pixel_8/gring VBIAS 1.38fF
C71 pixel_8/gring VREF 5.50fF
C72 PIX_OUT1 VDD 1.06fF
C73 pixel_0/test VDD 2.25fF
C74 pixel_8/gring PIX2_IN 3.31fF
C75 pixel_2/net2 PIX2_IN 1.91fF
C76 pixel_8/gring PIX8_IN 3.31fF
C77 pixel_0/net2 VDD 1.04fF
C78 pixel_0/a_4350_10# VDD 1.55fF
C79 VDD pixel_0/net1 1.59fF
C80 pixel_6/net2 PIX6_IN 1.91fF
C81 VDD pixel_6/net1 1.59fF
C82 pixel_6/net2 VDD 1.04fF
C83 PIX_OUT1 NB1 1.10fF
C84 VDD pixel_6/a_4350_10# 1.55fF
C85 pixel_8/test VDD 2.28fF
C86 pixel_6/test VDD 2.25fF
C87 PIX7_IN pixel_7/net2 1.91fF
C88 PIX_OUT2 VDD 1.06fF
C89 SF_IB VDD 32.01fF
C90 pixel_8/gring PIX_OUT0 2.94fF
C91 PIX5_IN VDD 1.18fF
C92 PIX0_IN pixel_0/net2 1.91fF
C93 pixel_7/net2 VDD 1.04fF
C94 PIX_OUT1 CSA_VREF 1.42fF
C95 pixel_5/net1 VDD 1.59fF
C96 pixel_5/net2 VDD 1.04fF
C97 pixel_5/test VDD 2.29fF
C98 pixel_5/a_4350_10# VDD 1.55fF
C99 pixel_7/net1 VDD 1.59fF
C100 pixel_8/gring PIX1_IN 3.31fF
C101 PIX_OUT2 NB1 1.10fF
C102 SF_IB NB1 3.56fF
Xpixel_0 VREF ROW_SEL0 NB1 VBIAS NB2 PIX0_IN SF_IB PIX_OUT0 CSA_VREF pixel
Xpixel_1 VREF ROW_SEL0 NB1 VBIAS NB2 PIX1_IN SF_IB PIX_OUT1 CSA_VREF pixel
Xpixel_2 VREF ROW_SEL0 NB1 VBIAS NB2 PIX2_IN SF_IB PIX_OUT2 CSA_VREF pixel
Xpixel_3 VREF ROW_SEL1 NB1 VBIAS NB2 PIX3_IN SF_IB PIX_OUT0 CSA_VREF pixel
Xpixel_4 VREF ROW_SEL1 NB1 VBIAS NB2 PIX4_IN SF_IB PIX_OUT1 CSA_VREF pixel
Xpixel_5 VREF ROW_SEL1 NB1 VBIAS NB2 PIX5_IN SF_IB PIX_OUT2 CSA_VREF pixel
Xpixel_6 VREF ROW_SEL2 NB1 VBIAS NB2 PIX6_IN SF_IB PIX_OUT0 CSA_VREF pixel
Xpixel_7 VREF ROW_SEL2 NB1 VBIAS NB2 PIX7_IN SF_IB PIX_OUT1 CSA_VREF pixel
Xpixel_8 VREF ROW_SEL2 NB1 VBIAS NB2 PIX8_IN SF_IB PIX_OUT2 CSA_VREF pixel
C103 COL_SEL2 GND 1.30fF
C104 COL_SEL1 GND 1.30fF
C105 COL_SEL0 GND 1.46fF
C106 ARRAY_OUT GND 8.18fF **FLOATING
C107 PIX_OUT2 GND 9.86fF
C108 PIX8_IN GND 6.48fF
C109 pixel_8/gring GND 10.38fF
C110 pixel_8/net2 GND 1.50fF
C111 NB1 GND 31.00fF
C112 PIX_OUT1 GND 10.07fF
C113 ROW_SEL2 GND 8.90fF
C114 PIX7_IN GND 6.50fF
C115 CSA_VREF GND 1.27fF
C116 VDD GND 71.59fF
C117 pixel_7/net2 GND 1.50fF
C118 PIX_OUT0 GND 8.23fF
C119 PIX6_IN GND 6.49fF
C120 pixel_6/net2 GND 1.50fF
C121 PIX5_IN GND 6.49fF
C122 pixel_5/net2 GND 1.50fF
C123 ROW_SEL1 GND 9.12fF
C124 PIX4_IN GND 6.52fF
C125 pixel_4/net2 GND 1.50fF
C126 NB2 GND 12.00fF
C127 VREF GND 10.73fF
C128 VBIAS GND 10.29fF
C129 PIX3_IN GND 6.62fF
C130 pixel_3/net2 GND 1.50fF
C131 PIX2_IN GND 6.49fF
C132 pixel_2/net2 GND 1.50fF
C133 ROW_SEL0 GND 8.91fF
C134 PIX1_IN GND 6.49fF
C135 pixel_1/net2 GND 1.50fF
C136 PIX0_IN GND 6.49fF
C137 pixel_0/net2 GND 1.50fF
.ends
