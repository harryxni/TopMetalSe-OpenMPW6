magic
tech sky130A
magscale 1 2
timestamp 1608354390
<< nwell >>
rect 408 664 1342 1692
<< pwell >>
rect 500 -247 1179 641
<< psubdiff >>
rect 564 -38 1108 46
rect 564 -215 606 -38
rect 1057 -215 1108 -38
rect 564 -221 1108 -215
<< nsubdiff >>
rect 509 1343 1244 1631
<< psubdiffcont >>
rect 606 -215 1057 -38
<< poly >>
rect 716 901 746 941
rect 812 901 842 943
rect 908 901 938 943
rect 1004 901 1034 943
rect 713 891 1052 901
rect 713 854 731 891
rect 1025 854 1052 891
rect 713 844 1052 854
<< polycont >>
rect 731 854 1025 891
<< locali >>
rect 715 854 731 891
rect 1025 854 1041 891
<< viali >>
rect 508 1343 1241 1626
rect 731 854 1025 891
rect 574 -38 1104 44
rect 574 -215 606 -38
rect 606 -215 1057 -38
rect 1057 -215 1104 -38
rect 574 -219 1104 -215
<< metal1 >>
rect 496 1626 1253 1632
rect 496 1343 508 1626
rect 1241 1343 1253 1626
rect 496 1337 1253 1343
rect 631 940 641 1184
rect 695 940 705 1184
rect 753 945 804 1337
rect 835 937 845 1180
rect 904 937 914 1180
rect 946 954 997 1337
rect 1032 939 1042 1182
rect 1101 939 1111 1182
rect 725 891 1037 903
rect 719 854 731 891
rect 1025 854 1037 891
rect 725 848 1037 854
rect 753 734 901 848
rect 408 586 901 734
rect 753 471 901 586
rect 681 188 691 442
rect 749 188 759 442
rect 808 50 862 439
rect 895 185 905 439
rect 983 185 993 439
rect 562 44 1116 50
rect 562 -219 574 44
rect 1104 -219 1116 44
rect 562 -225 1116 -219
<< via1 >>
rect 641 940 695 1184
rect 845 937 904 1180
rect 1042 939 1101 1182
rect 691 188 749 442
rect 905 185 983 439
<< metal2 >>
rect 641 1184 695 1194
rect 845 1180 904 1190
rect 695 940 845 1179
rect 641 939 845 940
rect 641 930 695 939
rect 733 937 845 939
rect 1042 1182 1101 1192
rect 904 939 1042 1179
rect 1101 939 1103 1179
rect 904 937 963 939
rect 733 766 963 937
rect 1042 929 1101 939
rect 733 536 1318 766
rect 733 452 963 536
rect 691 449 963 452
rect 691 442 983 449
rect 749 439 983 442
rect 749 188 905 439
rect 691 186 905 188
rect 691 178 749 186
rect 905 175 983 185
use sky130_fd_pr__pfet_01v8_5UHRWD  sky130_fd_pr__pfet_01v8_5UHRWD_0
timestamp 1608353910
transform 1 0 875 0 1 1091
box -359 -369 359 369
use sky130_fd_pr__nfet_01v8_WRE4LY  sky130_fd_pr__nfet_01v8_WRE4LY_0
timestamp 1608344059
transform 1 0 831 0 1 318
box -263 -330 263 330
<< labels >>
rlabel metal1 408 586 901 734 1 in
rlabel metal2 733 536 1318 766 1 out
rlabel nsubdiff 509 1343 1244 1631 1 vdd
rlabel pwell 574 -219 1104 44 1 vss
<< end >>
