magic
tech sky130A
magscale 1 2
timestamp 1654643737
<< error_p >>
rect -2920 71 -2862 77
rect -2802 71 -2744 77
rect -2684 71 -2626 77
rect -2566 71 -2508 77
rect -2448 71 -2390 77
rect -2330 71 -2272 77
rect -2212 71 -2154 77
rect -2094 71 -2036 77
rect -1976 71 -1918 77
rect -1858 71 -1800 77
rect -1740 71 -1682 77
rect -1622 71 -1564 77
rect -1504 71 -1446 77
rect -1386 71 -1328 77
rect -1268 71 -1210 77
rect -1150 71 -1092 77
rect -1032 71 -974 77
rect -914 71 -856 77
rect -796 71 -738 77
rect -678 71 -620 77
rect -560 71 -502 77
rect -442 71 -384 77
rect -324 71 -266 77
rect -206 71 -148 77
rect -88 71 -30 77
rect 30 71 88 77
rect 148 71 206 77
rect 266 71 324 77
rect 384 71 442 77
rect 502 71 560 77
rect 620 71 678 77
rect 738 71 796 77
rect 856 71 914 77
rect 974 71 1032 77
rect 1092 71 1150 77
rect 1210 71 1268 77
rect 1328 71 1386 77
rect 1446 71 1504 77
rect 1564 71 1622 77
rect 1682 71 1740 77
rect 1800 71 1858 77
rect 1918 71 1976 77
rect 2036 71 2094 77
rect 2154 71 2212 77
rect 2272 71 2330 77
rect 2390 71 2448 77
rect 2508 71 2566 77
rect 2626 71 2684 77
rect 2744 71 2802 77
rect 2862 71 2920 77
rect -2920 37 -2908 71
rect -2802 37 -2790 71
rect -2684 37 -2672 71
rect -2566 37 -2554 71
rect -2448 37 -2436 71
rect -2330 37 -2318 71
rect -2212 37 -2200 71
rect -2094 37 -2082 71
rect -1976 37 -1964 71
rect -1858 37 -1846 71
rect -1740 37 -1728 71
rect -1622 37 -1610 71
rect -1504 37 -1492 71
rect -1386 37 -1374 71
rect -1268 37 -1256 71
rect -1150 37 -1138 71
rect -1032 37 -1020 71
rect -914 37 -902 71
rect -796 37 -784 71
rect -678 37 -666 71
rect -560 37 -548 71
rect -442 37 -430 71
rect -324 37 -312 71
rect -206 37 -194 71
rect -88 37 -76 71
rect 30 37 42 71
rect 148 37 160 71
rect 266 37 278 71
rect 384 37 396 71
rect 502 37 514 71
rect 620 37 632 71
rect 738 37 750 71
rect 856 37 868 71
rect 974 37 986 71
rect 1092 37 1104 71
rect 1210 37 1222 71
rect 1328 37 1340 71
rect 1446 37 1458 71
rect 1564 37 1576 71
rect 1682 37 1694 71
rect 1800 37 1812 71
rect 1918 37 1930 71
rect 2036 37 2048 71
rect 2154 37 2166 71
rect 2272 37 2284 71
rect 2390 37 2402 71
rect 2508 37 2520 71
rect 2626 37 2638 71
rect 2744 37 2756 71
rect 2862 37 2874 71
rect -2920 31 -2862 37
rect -2802 31 -2744 37
rect -2684 31 -2626 37
rect -2566 31 -2508 37
rect -2448 31 -2390 37
rect -2330 31 -2272 37
rect -2212 31 -2154 37
rect -2094 31 -2036 37
rect -1976 31 -1918 37
rect -1858 31 -1800 37
rect -1740 31 -1682 37
rect -1622 31 -1564 37
rect -1504 31 -1446 37
rect -1386 31 -1328 37
rect -1268 31 -1210 37
rect -1150 31 -1092 37
rect -1032 31 -974 37
rect -914 31 -856 37
rect -796 31 -738 37
rect -678 31 -620 37
rect -560 31 -502 37
rect -442 31 -384 37
rect -324 31 -266 37
rect -206 31 -148 37
rect -88 31 -30 37
rect 30 31 88 37
rect 148 31 206 37
rect 266 31 324 37
rect 384 31 442 37
rect 502 31 560 37
rect 620 31 678 37
rect 738 31 796 37
rect 856 31 914 37
rect 974 31 1032 37
rect 1092 31 1150 37
rect 1210 31 1268 37
rect 1328 31 1386 37
rect 1446 31 1504 37
rect 1564 31 1622 37
rect 1682 31 1740 37
rect 1800 31 1858 37
rect 1918 31 1976 37
rect 2036 31 2094 37
rect 2154 31 2212 37
rect 2272 31 2330 37
rect 2390 31 2448 37
rect 2508 31 2566 37
rect 2626 31 2684 37
rect 2744 31 2802 37
rect 2862 31 2920 37
rect -2920 -37 -2862 -31
rect -2802 -37 -2744 -31
rect -2684 -37 -2626 -31
rect -2566 -37 -2508 -31
rect -2448 -37 -2390 -31
rect -2330 -37 -2272 -31
rect -2212 -37 -2154 -31
rect -2094 -37 -2036 -31
rect -1976 -37 -1918 -31
rect -1858 -37 -1800 -31
rect -1740 -37 -1682 -31
rect -1622 -37 -1564 -31
rect -1504 -37 -1446 -31
rect -1386 -37 -1328 -31
rect -1268 -37 -1210 -31
rect -1150 -37 -1092 -31
rect -1032 -37 -974 -31
rect -914 -37 -856 -31
rect -796 -37 -738 -31
rect -678 -37 -620 -31
rect -560 -37 -502 -31
rect -442 -37 -384 -31
rect -324 -37 -266 -31
rect -206 -37 -148 -31
rect -88 -37 -30 -31
rect 30 -37 88 -31
rect 148 -37 206 -31
rect 266 -37 324 -31
rect 384 -37 442 -31
rect 502 -37 560 -31
rect 620 -37 678 -31
rect 738 -37 796 -31
rect 856 -37 914 -31
rect 974 -37 1032 -31
rect 1092 -37 1150 -31
rect 1210 -37 1268 -31
rect 1328 -37 1386 -31
rect 1446 -37 1504 -31
rect 1564 -37 1622 -31
rect 1682 -37 1740 -31
rect 1800 -37 1858 -31
rect 1918 -37 1976 -31
rect 2036 -37 2094 -31
rect 2154 -37 2212 -31
rect 2272 -37 2330 -31
rect 2390 -37 2448 -31
rect 2508 -37 2566 -31
rect 2626 -37 2684 -31
rect 2744 -37 2802 -31
rect 2862 -37 2920 -31
rect -2920 -71 -2908 -37
rect -2802 -71 -2790 -37
rect -2684 -71 -2672 -37
rect -2566 -71 -2554 -37
rect -2448 -71 -2436 -37
rect -2330 -71 -2318 -37
rect -2212 -71 -2200 -37
rect -2094 -71 -2082 -37
rect -1976 -71 -1964 -37
rect -1858 -71 -1846 -37
rect -1740 -71 -1728 -37
rect -1622 -71 -1610 -37
rect -1504 -71 -1492 -37
rect -1386 -71 -1374 -37
rect -1268 -71 -1256 -37
rect -1150 -71 -1138 -37
rect -1032 -71 -1020 -37
rect -914 -71 -902 -37
rect -796 -71 -784 -37
rect -678 -71 -666 -37
rect -560 -71 -548 -37
rect -442 -71 -430 -37
rect -324 -71 -312 -37
rect -206 -71 -194 -37
rect -88 -71 -76 -37
rect 30 -71 42 -37
rect 148 -71 160 -37
rect 266 -71 278 -37
rect 384 -71 396 -37
rect 502 -71 514 -37
rect 620 -71 632 -37
rect 738 -71 750 -37
rect 856 -71 868 -37
rect 974 -71 986 -37
rect 1092 -71 1104 -37
rect 1210 -71 1222 -37
rect 1328 -71 1340 -37
rect 1446 -71 1458 -37
rect 1564 -71 1576 -37
rect 1682 -71 1694 -37
rect 1800 -71 1812 -37
rect 1918 -71 1930 -37
rect 2036 -71 2048 -37
rect 2154 -71 2166 -37
rect 2272 -71 2284 -37
rect 2390 -71 2402 -37
rect 2508 -71 2520 -37
rect 2626 -71 2638 -37
rect 2744 -71 2756 -37
rect 2862 -71 2874 -37
rect -2920 -77 -2862 -71
rect -2802 -77 -2744 -71
rect -2684 -77 -2626 -71
rect -2566 -77 -2508 -71
rect -2448 -77 -2390 -71
rect -2330 -77 -2272 -71
rect -2212 -77 -2154 -71
rect -2094 -77 -2036 -71
rect -1976 -77 -1918 -71
rect -1858 -77 -1800 -71
rect -1740 -77 -1682 -71
rect -1622 -77 -1564 -71
rect -1504 -77 -1446 -71
rect -1386 -77 -1328 -71
rect -1268 -77 -1210 -71
rect -1150 -77 -1092 -71
rect -1032 -77 -974 -71
rect -914 -77 -856 -71
rect -796 -77 -738 -71
rect -678 -77 -620 -71
rect -560 -77 -502 -71
rect -442 -77 -384 -71
rect -324 -77 -266 -71
rect -206 -77 -148 -71
rect -88 -77 -30 -71
rect 30 -77 88 -71
rect 148 -77 206 -71
rect 266 -77 324 -71
rect 384 -77 442 -71
rect 502 -77 560 -71
rect 620 -77 678 -71
rect 738 -77 796 -71
rect 856 -77 914 -71
rect 974 -77 1032 -71
rect 1092 -77 1150 -71
rect 1210 -77 1268 -71
rect 1328 -77 1386 -71
rect 1446 -77 1504 -71
rect 1564 -77 1622 -71
rect 1682 -77 1740 -71
rect 1800 -77 1858 -71
rect 1918 -77 1976 -71
rect 2036 -77 2094 -71
rect 2154 -77 2212 -71
rect 2272 -77 2330 -71
rect 2390 -77 2448 -71
rect 2508 -77 2566 -71
rect 2626 -77 2684 -71
rect 2744 -77 2802 -71
rect 2862 -77 2920 -71
<< nwell >>
rect -3117 -937 3117 937
<< pmos >>
rect -2921 118 -2861 718
rect -2803 118 -2743 718
rect -2685 118 -2625 718
rect -2567 118 -2507 718
rect -2449 118 -2389 718
rect -2331 118 -2271 718
rect -2213 118 -2153 718
rect -2095 118 -2035 718
rect -1977 118 -1917 718
rect -1859 118 -1799 718
rect -1741 118 -1681 718
rect -1623 118 -1563 718
rect -1505 118 -1445 718
rect -1387 118 -1327 718
rect -1269 118 -1209 718
rect -1151 118 -1091 718
rect -1033 118 -973 718
rect -915 118 -855 718
rect -797 118 -737 718
rect -679 118 -619 718
rect -561 118 -501 718
rect -443 118 -383 718
rect -325 118 -265 718
rect -207 118 -147 718
rect -89 118 -29 718
rect 29 118 89 718
rect 147 118 207 718
rect 265 118 325 718
rect 383 118 443 718
rect 501 118 561 718
rect 619 118 679 718
rect 737 118 797 718
rect 855 118 915 718
rect 973 118 1033 718
rect 1091 118 1151 718
rect 1209 118 1269 718
rect 1327 118 1387 718
rect 1445 118 1505 718
rect 1563 118 1623 718
rect 1681 118 1741 718
rect 1799 118 1859 718
rect 1917 118 1977 718
rect 2035 118 2095 718
rect 2153 118 2213 718
rect 2271 118 2331 718
rect 2389 118 2449 718
rect 2507 118 2567 718
rect 2625 118 2685 718
rect 2743 118 2803 718
rect 2861 118 2921 718
rect -2921 -718 -2861 -118
rect -2803 -718 -2743 -118
rect -2685 -718 -2625 -118
rect -2567 -718 -2507 -118
rect -2449 -718 -2389 -118
rect -2331 -718 -2271 -118
rect -2213 -718 -2153 -118
rect -2095 -718 -2035 -118
rect -1977 -718 -1917 -118
rect -1859 -718 -1799 -118
rect -1741 -718 -1681 -118
rect -1623 -718 -1563 -118
rect -1505 -718 -1445 -118
rect -1387 -718 -1327 -118
rect -1269 -718 -1209 -118
rect -1151 -718 -1091 -118
rect -1033 -718 -973 -118
rect -915 -718 -855 -118
rect -797 -718 -737 -118
rect -679 -718 -619 -118
rect -561 -718 -501 -118
rect -443 -718 -383 -118
rect -325 -718 -265 -118
rect -207 -718 -147 -118
rect -89 -718 -29 -118
rect 29 -718 89 -118
rect 147 -718 207 -118
rect 265 -718 325 -118
rect 383 -718 443 -118
rect 501 -718 561 -118
rect 619 -718 679 -118
rect 737 -718 797 -118
rect 855 -718 915 -118
rect 973 -718 1033 -118
rect 1091 -718 1151 -118
rect 1209 -718 1269 -118
rect 1327 -718 1387 -118
rect 1445 -718 1505 -118
rect 1563 -718 1623 -118
rect 1681 -718 1741 -118
rect 1799 -718 1859 -118
rect 1917 -718 1977 -118
rect 2035 -718 2095 -118
rect 2153 -718 2213 -118
rect 2271 -718 2331 -118
rect 2389 -718 2449 -118
rect 2507 -718 2567 -118
rect 2625 -718 2685 -118
rect 2743 -718 2803 -118
rect 2861 -718 2921 -118
<< pdiff >>
rect -2979 673 -2921 718
rect -2979 639 -2967 673
rect -2933 639 -2921 673
rect -2979 605 -2921 639
rect -2979 571 -2967 605
rect -2933 571 -2921 605
rect -2979 537 -2921 571
rect -2979 503 -2967 537
rect -2933 503 -2921 537
rect -2979 469 -2921 503
rect -2979 435 -2967 469
rect -2933 435 -2921 469
rect -2979 401 -2921 435
rect -2979 367 -2967 401
rect -2933 367 -2921 401
rect -2979 333 -2921 367
rect -2979 299 -2967 333
rect -2933 299 -2921 333
rect -2979 265 -2921 299
rect -2979 231 -2967 265
rect -2933 231 -2921 265
rect -2979 197 -2921 231
rect -2979 163 -2967 197
rect -2933 163 -2921 197
rect -2979 118 -2921 163
rect -2861 673 -2803 718
rect -2861 639 -2849 673
rect -2815 639 -2803 673
rect -2861 605 -2803 639
rect -2861 571 -2849 605
rect -2815 571 -2803 605
rect -2861 537 -2803 571
rect -2861 503 -2849 537
rect -2815 503 -2803 537
rect -2861 469 -2803 503
rect -2861 435 -2849 469
rect -2815 435 -2803 469
rect -2861 401 -2803 435
rect -2861 367 -2849 401
rect -2815 367 -2803 401
rect -2861 333 -2803 367
rect -2861 299 -2849 333
rect -2815 299 -2803 333
rect -2861 265 -2803 299
rect -2861 231 -2849 265
rect -2815 231 -2803 265
rect -2861 197 -2803 231
rect -2861 163 -2849 197
rect -2815 163 -2803 197
rect -2861 118 -2803 163
rect -2743 673 -2685 718
rect -2743 639 -2731 673
rect -2697 639 -2685 673
rect -2743 605 -2685 639
rect -2743 571 -2731 605
rect -2697 571 -2685 605
rect -2743 537 -2685 571
rect -2743 503 -2731 537
rect -2697 503 -2685 537
rect -2743 469 -2685 503
rect -2743 435 -2731 469
rect -2697 435 -2685 469
rect -2743 401 -2685 435
rect -2743 367 -2731 401
rect -2697 367 -2685 401
rect -2743 333 -2685 367
rect -2743 299 -2731 333
rect -2697 299 -2685 333
rect -2743 265 -2685 299
rect -2743 231 -2731 265
rect -2697 231 -2685 265
rect -2743 197 -2685 231
rect -2743 163 -2731 197
rect -2697 163 -2685 197
rect -2743 118 -2685 163
rect -2625 673 -2567 718
rect -2625 639 -2613 673
rect -2579 639 -2567 673
rect -2625 605 -2567 639
rect -2625 571 -2613 605
rect -2579 571 -2567 605
rect -2625 537 -2567 571
rect -2625 503 -2613 537
rect -2579 503 -2567 537
rect -2625 469 -2567 503
rect -2625 435 -2613 469
rect -2579 435 -2567 469
rect -2625 401 -2567 435
rect -2625 367 -2613 401
rect -2579 367 -2567 401
rect -2625 333 -2567 367
rect -2625 299 -2613 333
rect -2579 299 -2567 333
rect -2625 265 -2567 299
rect -2625 231 -2613 265
rect -2579 231 -2567 265
rect -2625 197 -2567 231
rect -2625 163 -2613 197
rect -2579 163 -2567 197
rect -2625 118 -2567 163
rect -2507 673 -2449 718
rect -2507 639 -2495 673
rect -2461 639 -2449 673
rect -2507 605 -2449 639
rect -2507 571 -2495 605
rect -2461 571 -2449 605
rect -2507 537 -2449 571
rect -2507 503 -2495 537
rect -2461 503 -2449 537
rect -2507 469 -2449 503
rect -2507 435 -2495 469
rect -2461 435 -2449 469
rect -2507 401 -2449 435
rect -2507 367 -2495 401
rect -2461 367 -2449 401
rect -2507 333 -2449 367
rect -2507 299 -2495 333
rect -2461 299 -2449 333
rect -2507 265 -2449 299
rect -2507 231 -2495 265
rect -2461 231 -2449 265
rect -2507 197 -2449 231
rect -2507 163 -2495 197
rect -2461 163 -2449 197
rect -2507 118 -2449 163
rect -2389 673 -2331 718
rect -2389 639 -2377 673
rect -2343 639 -2331 673
rect -2389 605 -2331 639
rect -2389 571 -2377 605
rect -2343 571 -2331 605
rect -2389 537 -2331 571
rect -2389 503 -2377 537
rect -2343 503 -2331 537
rect -2389 469 -2331 503
rect -2389 435 -2377 469
rect -2343 435 -2331 469
rect -2389 401 -2331 435
rect -2389 367 -2377 401
rect -2343 367 -2331 401
rect -2389 333 -2331 367
rect -2389 299 -2377 333
rect -2343 299 -2331 333
rect -2389 265 -2331 299
rect -2389 231 -2377 265
rect -2343 231 -2331 265
rect -2389 197 -2331 231
rect -2389 163 -2377 197
rect -2343 163 -2331 197
rect -2389 118 -2331 163
rect -2271 673 -2213 718
rect -2271 639 -2259 673
rect -2225 639 -2213 673
rect -2271 605 -2213 639
rect -2271 571 -2259 605
rect -2225 571 -2213 605
rect -2271 537 -2213 571
rect -2271 503 -2259 537
rect -2225 503 -2213 537
rect -2271 469 -2213 503
rect -2271 435 -2259 469
rect -2225 435 -2213 469
rect -2271 401 -2213 435
rect -2271 367 -2259 401
rect -2225 367 -2213 401
rect -2271 333 -2213 367
rect -2271 299 -2259 333
rect -2225 299 -2213 333
rect -2271 265 -2213 299
rect -2271 231 -2259 265
rect -2225 231 -2213 265
rect -2271 197 -2213 231
rect -2271 163 -2259 197
rect -2225 163 -2213 197
rect -2271 118 -2213 163
rect -2153 673 -2095 718
rect -2153 639 -2141 673
rect -2107 639 -2095 673
rect -2153 605 -2095 639
rect -2153 571 -2141 605
rect -2107 571 -2095 605
rect -2153 537 -2095 571
rect -2153 503 -2141 537
rect -2107 503 -2095 537
rect -2153 469 -2095 503
rect -2153 435 -2141 469
rect -2107 435 -2095 469
rect -2153 401 -2095 435
rect -2153 367 -2141 401
rect -2107 367 -2095 401
rect -2153 333 -2095 367
rect -2153 299 -2141 333
rect -2107 299 -2095 333
rect -2153 265 -2095 299
rect -2153 231 -2141 265
rect -2107 231 -2095 265
rect -2153 197 -2095 231
rect -2153 163 -2141 197
rect -2107 163 -2095 197
rect -2153 118 -2095 163
rect -2035 673 -1977 718
rect -2035 639 -2023 673
rect -1989 639 -1977 673
rect -2035 605 -1977 639
rect -2035 571 -2023 605
rect -1989 571 -1977 605
rect -2035 537 -1977 571
rect -2035 503 -2023 537
rect -1989 503 -1977 537
rect -2035 469 -1977 503
rect -2035 435 -2023 469
rect -1989 435 -1977 469
rect -2035 401 -1977 435
rect -2035 367 -2023 401
rect -1989 367 -1977 401
rect -2035 333 -1977 367
rect -2035 299 -2023 333
rect -1989 299 -1977 333
rect -2035 265 -1977 299
rect -2035 231 -2023 265
rect -1989 231 -1977 265
rect -2035 197 -1977 231
rect -2035 163 -2023 197
rect -1989 163 -1977 197
rect -2035 118 -1977 163
rect -1917 673 -1859 718
rect -1917 639 -1905 673
rect -1871 639 -1859 673
rect -1917 605 -1859 639
rect -1917 571 -1905 605
rect -1871 571 -1859 605
rect -1917 537 -1859 571
rect -1917 503 -1905 537
rect -1871 503 -1859 537
rect -1917 469 -1859 503
rect -1917 435 -1905 469
rect -1871 435 -1859 469
rect -1917 401 -1859 435
rect -1917 367 -1905 401
rect -1871 367 -1859 401
rect -1917 333 -1859 367
rect -1917 299 -1905 333
rect -1871 299 -1859 333
rect -1917 265 -1859 299
rect -1917 231 -1905 265
rect -1871 231 -1859 265
rect -1917 197 -1859 231
rect -1917 163 -1905 197
rect -1871 163 -1859 197
rect -1917 118 -1859 163
rect -1799 673 -1741 718
rect -1799 639 -1787 673
rect -1753 639 -1741 673
rect -1799 605 -1741 639
rect -1799 571 -1787 605
rect -1753 571 -1741 605
rect -1799 537 -1741 571
rect -1799 503 -1787 537
rect -1753 503 -1741 537
rect -1799 469 -1741 503
rect -1799 435 -1787 469
rect -1753 435 -1741 469
rect -1799 401 -1741 435
rect -1799 367 -1787 401
rect -1753 367 -1741 401
rect -1799 333 -1741 367
rect -1799 299 -1787 333
rect -1753 299 -1741 333
rect -1799 265 -1741 299
rect -1799 231 -1787 265
rect -1753 231 -1741 265
rect -1799 197 -1741 231
rect -1799 163 -1787 197
rect -1753 163 -1741 197
rect -1799 118 -1741 163
rect -1681 673 -1623 718
rect -1681 639 -1669 673
rect -1635 639 -1623 673
rect -1681 605 -1623 639
rect -1681 571 -1669 605
rect -1635 571 -1623 605
rect -1681 537 -1623 571
rect -1681 503 -1669 537
rect -1635 503 -1623 537
rect -1681 469 -1623 503
rect -1681 435 -1669 469
rect -1635 435 -1623 469
rect -1681 401 -1623 435
rect -1681 367 -1669 401
rect -1635 367 -1623 401
rect -1681 333 -1623 367
rect -1681 299 -1669 333
rect -1635 299 -1623 333
rect -1681 265 -1623 299
rect -1681 231 -1669 265
rect -1635 231 -1623 265
rect -1681 197 -1623 231
rect -1681 163 -1669 197
rect -1635 163 -1623 197
rect -1681 118 -1623 163
rect -1563 673 -1505 718
rect -1563 639 -1551 673
rect -1517 639 -1505 673
rect -1563 605 -1505 639
rect -1563 571 -1551 605
rect -1517 571 -1505 605
rect -1563 537 -1505 571
rect -1563 503 -1551 537
rect -1517 503 -1505 537
rect -1563 469 -1505 503
rect -1563 435 -1551 469
rect -1517 435 -1505 469
rect -1563 401 -1505 435
rect -1563 367 -1551 401
rect -1517 367 -1505 401
rect -1563 333 -1505 367
rect -1563 299 -1551 333
rect -1517 299 -1505 333
rect -1563 265 -1505 299
rect -1563 231 -1551 265
rect -1517 231 -1505 265
rect -1563 197 -1505 231
rect -1563 163 -1551 197
rect -1517 163 -1505 197
rect -1563 118 -1505 163
rect -1445 673 -1387 718
rect -1445 639 -1433 673
rect -1399 639 -1387 673
rect -1445 605 -1387 639
rect -1445 571 -1433 605
rect -1399 571 -1387 605
rect -1445 537 -1387 571
rect -1445 503 -1433 537
rect -1399 503 -1387 537
rect -1445 469 -1387 503
rect -1445 435 -1433 469
rect -1399 435 -1387 469
rect -1445 401 -1387 435
rect -1445 367 -1433 401
rect -1399 367 -1387 401
rect -1445 333 -1387 367
rect -1445 299 -1433 333
rect -1399 299 -1387 333
rect -1445 265 -1387 299
rect -1445 231 -1433 265
rect -1399 231 -1387 265
rect -1445 197 -1387 231
rect -1445 163 -1433 197
rect -1399 163 -1387 197
rect -1445 118 -1387 163
rect -1327 673 -1269 718
rect -1327 639 -1315 673
rect -1281 639 -1269 673
rect -1327 605 -1269 639
rect -1327 571 -1315 605
rect -1281 571 -1269 605
rect -1327 537 -1269 571
rect -1327 503 -1315 537
rect -1281 503 -1269 537
rect -1327 469 -1269 503
rect -1327 435 -1315 469
rect -1281 435 -1269 469
rect -1327 401 -1269 435
rect -1327 367 -1315 401
rect -1281 367 -1269 401
rect -1327 333 -1269 367
rect -1327 299 -1315 333
rect -1281 299 -1269 333
rect -1327 265 -1269 299
rect -1327 231 -1315 265
rect -1281 231 -1269 265
rect -1327 197 -1269 231
rect -1327 163 -1315 197
rect -1281 163 -1269 197
rect -1327 118 -1269 163
rect -1209 673 -1151 718
rect -1209 639 -1197 673
rect -1163 639 -1151 673
rect -1209 605 -1151 639
rect -1209 571 -1197 605
rect -1163 571 -1151 605
rect -1209 537 -1151 571
rect -1209 503 -1197 537
rect -1163 503 -1151 537
rect -1209 469 -1151 503
rect -1209 435 -1197 469
rect -1163 435 -1151 469
rect -1209 401 -1151 435
rect -1209 367 -1197 401
rect -1163 367 -1151 401
rect -1209 333 -1151 367
rect -1209 299 -1197 333
rect -1163 299 -1151 333
rect -1209 265 -1151 299
rect -1209 231 -1197 265
rect -1163 231 -1151 265
rect -1209 197 -1151 231
rect -1209 163 -1197 197
rect -1163 163 -1151 197
rect -1209 118 -1151 163
rect -1091 673 -1033 718
rect -1091 639 -1079 673
rect -1045 639 -1033 673
rect -1091 605 -1033 639
rect -1091 571 -1079 605
rect -1045 571 -1033 605
rect -1091 537 -1033 571
rect -1091 503 -1079 537
rect -1045 503 -1033 537
rect -1091 469 -1033 503
rect -1091 435 -1079 469
rect -1045 435 -1033 469
rect -1091 401 -1033 435
rect -1091 367 -1079 401
rect -1045 367 -1033 401
rect -1091 333 -1033 367
rect -1091 299 -1079 333
rect -1045 299 -1033 333
rect -1091 265 -1033 299
rect -1091 231 -1079 265
rect -1045 231 -1033 265
rect -1091 197 -1033 231
rect -1091 163 -1079 197
rect -1045 163 -1033 197
rect -1091 118 -1033 163
rect -973 673 -915 718
rect -973 639 -961 673
rect -927 639 -915 673
rect -973 605 -915 639
rect -973 571 -961 605
rect -927 571 -915 605
rect -973 537 -915 571
rect -973 503 -961 537
rect -927 503 -915 537
rect -973 469 -915 503
rect -973 435 -961 469
rect -927 435 -915 469
rect -973 401 -915 435
rect -973 367 -961 401
rect -927 367 -915 401
rect -973 333 -915 367
rect -973 299 -961 333
rect -927 299 -915 333
rect -973 265 -915 299
rect -973 231 -961 265
rect -927 231 -915 265
rect -973 197 -915 231
rect -973 163 -961 197
rect -927 163 -915 197
rect -973 118 -915 163
rect -855 673 -797 718
rect -855 639 -843 673
rect -809 639 -797 673
rect -855 605 -797 639
rect -855 571 -843 605
rect -809 571 -797 605
rect -855 537 -797 571
rect -855 503 -843 537
rect -809 503 -797 537
rect -855 469 -797 503
rect -855 435 -843 469
rect -809 435 -797 469
rect -855 401 -797 435
rect -855 367 -843 401
rect -809 367 -797 401
rect -855 333 -797 367
rect -855 299 -843 333
rect -809 299 -797 333
rect -855 265 -797 299
rect -855 231 -843 265
rect -809 231 -797 265
rect -855 197 -797 231
rect -855 163 -843 197
rect -809 163 -797 197
rect -855 118 -797 163
rect -737 673 -679 718
rect -737 639 -725 673
rect -691 639 -679 673
rect -737 605 -679 639
rect -737 571 -725 605
rect -691 571 -679 605
rect -737 537 -679 571
rect -737 503 -725 537
rect -691 503 -679 537
rect -737 469 -679 503
rect -737 435 -725 469
rect -691 435 -679 469
rect -737 401 -679 435
rect -737 367 -725 401
rect -691 367 -679 401
rect -737 333 -679 367
rect -737 299 -725 333
rect -691 299 -679 333
rect -737 265 -679 299
rect -737 231 -725 265
rect -691 231 -679 265
rect -737 197 -679 231
rect -737 163 -725 197
rect -691 163 -679 197
rect -737 118 -679 163
rect -619 673 -561 718
rect -619 639 -607 673
rect -573 639 -561 673
rect -619 605 -561 639
rect -619 571 -607 605
rect -573 571 -561 605
rect -619 537 -561 571
rect -619 503 -607 537
rect -573 503 -561 537
rect -619 469 -561 503
rect -619 435 -607 469
rect -573 435 -561 469
rect -619 401 -561 435
rect -619 367 -607 401
rect -573 367 -561 401
rect -619 333 -561 367
rect -619 299 -607 333
rect -573 299 -561 333
rect -619 265 -561 299
rect -619 231 -607 265
rect -573 231 -561 265
rect -619 197 -561 231
rect -619 163 -607 197
rect -573 163 -561 197
rect -619 118 -561 163
rect -501 673 -443 718
rect -501 639 -489 673
rect -455 639 -443 673
rect -501 605 -443 639
rect -501 571 -489 605
rect -455 571 -443 605
rect -501 537 -443 571
rect -501 503 -489 537
rect -455 503 -443 537
rect -501 469 -443 503
rect -501 435 -489 469
rect -455 435 -443 469
rect -501 401 -443 435
rect -501 367 -489 401
rect -455 367 -443 401
rect -501 333 -443 367
rect -501 299 -489 333
rect -455 299 -443 333
rect -501 265 -443 299
rect -501 231 -489 265
rect -455 231 -443 265
rect -501 197 -443 231
rect -501 163 -489 197
rect -455 163 -443 197
rect -501 118 -443 163
rect -383 673 -325 718
rect -383 639 -371 673
rect -337 639 -325 673
rect -383 605 -325 639
rect -383 571 -371 605
rect -337 571 -325 605
rect -383 537 -325 571
rect -383 503 -371 537
rect -337 503 -325 537
rect -383 469 -325 503
rect -383 435 -371 469
rect -337 435 -325 469
rect -383 401 -325 435
rect -383 367 -371 401
rect -337 367 -325 401
rect -383 333 -325 367
rect -383 299 -371 333
rect -337 299 -325 333
rect -383 265 -325 299
rect -383 231 -371 265
rect -337 231 -325 265
rect -383 197 -325 231
rect -383 163 -371 197
rect -337 163 -325 197
rect -383 118 -325 163
rect -265 673 -207 718
rect -265 639 -253 673
rect -219 639 -207 673
rect -265 605 -207 639
rect -265 571 -253 605
rect -219 571 -207 605
rect -265 537 -207 571
rect -265 503 -253 537
rect -219 503 -207 537
rect -265 469 -207 503
rect -265 435 -253 469
rect -219 435 -207 469
rect -265 401 -207 435
rect -265 367 -253 401
rect -219 367 -207 401
rect -265 333 -207 367
rect -265 299 -253 333
rect -219 299 -207 333
rect -265 265 -207 299
rect -265 231 -253 265
rect -219 231 -207 265
rect -265 197 -207 231
rect -265 163 -253 197
rect -219 163 -207 197
rect -265 118 -207 163
rect -147 673 -89 718
rect -147 639 -135 673
rect -101 639 -89 673
rect -147 605 -89 639
rect -147 571 -135 605
rect -101 571 -89 605
rect -147 537 -89 571
rect -147 503 -135 537
rect -101 503 -89 537
rect -147 469 -89 503
rect -147 435 -135 469
rect -101 435 -89 469
rect -147 401 -89 435
rect -147 367 -135 401
rect -101 367 -89 401
rect -147 333 -89 367
rect -147 299 -135 333
rect -101 299 -89 333
rect -147 265 -89 299
rect -147 231 -135 265
rect -101 231 -89 265
rect -147 197 -89 231
rect -147 163 -135 197
rect -101 163 -89 197
rect -147 118 -89 163
rect -29 673 29 718
rect -29 639 -17 673
rect 17 639 29 673
rect -29 605 29 639
rect -29 571 -17 605
rect 17 571 29 605
rect -29 537 29 571
rect -29 503 -17 537
rect 17 503 29 537
rect -29 469 29 503
rect -29 435 -17 469
rect 17 435 29 469
rect -29 401 29 435
rect -29 367 -17 401
rect 17 367 29 401
rect -29 333 29 367
rect -29 299 -17 333
rect 17 299 29 333
rect -29 265 29 299
rect -29 231 -17 265
rect 17 231 29 265
rect -29 197 29 231
rect -29 163 -17 197
rect 17 163 29 197
rect -29 118 29 163
rect 89 673 147 718
rect 89 639 101 673
rect 135 639 147 673
rect 89 605 147 639
rect 89 571 101 605
rect 135 571 147 605
rect 89 537 147 571
rect 89 503 101 537
rect 135 503 147 537
rect 89 469 147 503
rect 89 435 101 469
rect 135 435 147 469
rect 89 401 147 435
rect 89 367 101 401
rect 135 367 147 401
rect 89 333 147 367
rect 89 299 101 333
rect 135 299 147 333
rect 89 265 147 299
rect 89 231 101 265
rect 135 231 147 265
rect 89 197 147 231
rect 89 163 101 197
rect 135 163 147 197
rect 89 118 147 163
rect 207 673 265 718
rect 207 639 219 673
rect 253 639 265 673
rect 207 605 265 639
rect 207 571 219 605
rect 253 571 265 605
rect 207 537 265 571
rect 207 503 219 537
rect 253 503 265 537
rect 207 469 265 503
rect 207 435 219 469
rect 253 435 265 469
rect 207 401 265 435
rect 207 367 219 401
rect 253 367 265 401
rect 207 333 265 367
rect 207 299 219 333
rect 253 299 265 333
rect 207 265 265 299
rect 207 231 219 265
rect 253 231 265 265
rect 207 197 265 231
rect 207 163 219 197
rect 253 163 265 197
rect 207 118 265 163
rect 325 673 383 718
rect 325 639 337 673
rect 371 639 383 673
rect 325 605 383 639
rect 325 571 337 605
rect 371 571 383 605
rect 325 537 383 571
rect 325 503 337 537
rect 371 503 383 537
rect 325 469 383 503
rect 325 435 337 469
rect 371 435 383 469
rect 325 401 383 435
rect 325 367 337 401
rect 371 367 383 401
rect 325 333 383 367
rect 325 299 337 333
rect 371 299 383 333
rect 325 265 383 299
rect 325 231 337 265
rect 371 231 383 265
rect 325 197 383 231
rect 325 163 337 197
rect 371 163 383 197
rect 325 118 383 163
rect 443 673 501 718
rect 443 639 455 673
rect 489 639 501 673
rect 443 605 501 639
rect 443 571 455 605
rect 489 571 501 605
rect 443 537 501 571
rect 443 503 455 537
rect 489 503 501 537
rect 443 469 501 503
rect 443 435 455 469
rect 489 435 501 469
rect 443 401 501 435
rect 443 367 455 401
rect 489 367 501 401
rect 443 333 501 367
rect 443 299 455 333
rect 489 299 501 333
rect 443 265 501 299
rect 443 231 455 265
rect 489 231 501 265
rect 443 197 501 231
rect 443 163 455 197
rect 489 163 501 197
rect 443 118 501 163
rect 561 673 619 718
rect 561 639 573 673
rect 607 639 619 673
rect 561 605 619 639
rect 561 571 573 605
rect 607 571 619 605
rect 561 537 619 571
rect 561 503 573 537
rect 607 503 619 537
rect 561 469 619 503
rect 561 435 573 469
rect 607 435 619 469
rect 561 401 619 435
rect 561 367 573 401
rect 607 367 619 401
rect 561 333 619 367
rect 561 299 573 333
rect 607 299 619 333
rect 561 265 619 299
rect 561 231 573 265
rect 607 231 619 265
rect 561 197 619 231
rect 561 163 573 197
rect 607 163 619 197
rect 561 118 619 163
rect 679 673 737 718
rect 679 639 691 673
rect 725 639 737 673
rect 679 605 737 639
rect 679 571 691 605
rect 725 571 737 605
rect 679 537 737 571
rect 679 503 691 537
rect 725 503 737 537
rect 679 469 737 503
rect 679 435 691 469
rect 725 435 737 469
rect 679 401 737 435
rect 679 367 691 401
rect 725 367 737 401
rect 679 333 737 367
rect 679 299 691 333
rect 725 299 737 333
rect 679 265 737 299
rect 679 231 691 265
rect 725 231 737 265
rect 679 197 737 231
rect 679 163 691 197
rect 725 163 737 197
rect 679 118 737 163
rect 797 673 855 718
rect 797 639 809 673
rect 843 639 855 673
rect 797 605 855 639
rect 797 571 809 605
rect 843 571 855 605
rect 797 537 855 571
rect 797 503 809 537
rect 843 503 855 537
rect 797 469 855 503
rect 797 435 809 469
rect 843 435 855 469
rect 797 401 855 435
rect 797 367 809 401
rect 843 367 855 401
rect 797 333 855 367
rect 797 299 809 333
rect 843 299 855 333
rect 797 265 855 299
rect 797 231 809 265
rect 843 231 855 265
rect 797 197 855 231
rect 797 163 809 197
rect 843 163 855 197
rect 797 118 855 163
rect 915 673 973 718
rect 915 639 927 673
rect 961 639 973 673
rect 915 605 973 639
rect 915 571 927 605
rect 961 571 973 605
rect 915 537 973 571
rect 915 503 927 537
rect 961 503 973 537
rect 915 469 973 503
rect 915 435 927 469
rect 961 435 973 469
rect 915 401 973 435
rect 915 367 927 401
rect 961 367 973 401
rect 915 333 973 367
rect 915 299 927 333
rect 961 299 973 333
rect 915 265 973 299
rect 915 231 927 265
rect 961 231 973 265
rect 915 197 973 231
rect 915 163 927 197
rect 961 163 973 197
rect 915 118 973 163
rect 1033 673 1091 718
rect 1033 639 1045 673
rect 1079 639 1091 673
rect 1033 605 1091 639
rect 1033 571 1045 605
rect 1079 571 1091 605
rect 1033 537 1091 571
rect 1033 503 1045 537
rect 1079 503 1091 537
rect 1033 469 1091 503
rect 1033 435 1045 469
rect 1079 435 1091 469
rect 1033 401 1091 435
rect 1033 367 1045 401
rect 1079 367 1091 401
rect 1033 333 1091 367
rect 1033 299 1045 333
rect 1079 299 1091 333
rect 1033 265 1091 299
rect 1033 231 1045 265
rect 1079 231 1091 265
rect 1033 197 1091 231
rect 1033 163 1045 197
rect 1079 163 1091 197
rect 1033 118 1091 163
rect 1151 673 1209 718
rect 1151 639 1163 673
rect 1197 639 1209 673
rect 1151 605 1209 639
rect 1151 571 1163 605
rect 1197 571 1209 605
rect 1151 537 1209 571
rect 1151 503 1163 537
rect 1197 503 1209 537
rect 1151 469 1209 503
rect 1151 435 1163 469
rect 1197 435 1209 469
rect 1151 401 1209 435
rect 1151 367 1163 401
rect 1197 367 1209 401
rect 1151 333 1209 367
rect 1151 299 1163 333
rect 1197 299 1209 333
rect 1151 265 1209 299
rect 1151 231 1163 265
rect 1197 231 1209 265
rect 1151 197 1209 231
rect 1151 163 1163 197
rect 1197 163 1209 197
rect 1151 118 1209 163
rect 1269 673 1327 718
rect 1269 639 1281 673
rect 1315 639 1327 673
rect 1269 605 1327 639
rect 1269 571 1281 605
rect 1315 571 1327 605
rect 1269 537 1327 571
rect 1269 503 1281 537
rect 1315 503 1327 537
rect 1269 469 1327 503
rect 1269 435 1281 469
rect 1315 435 1327 469
rect 1269 401 1327 435
rect 1269 367 1281 401
rect 1315 367 1327 401
rect 1269 333 1327 367
rect 1269 299 1281 333
rect 1315 299 1327 333
rect 1269 265 1327 299
rect 1269 231 1281 265
rect 1315 231 1327 265
rect 1269 197 1327 231
rect 1269 163 1281 197
rect 1315 163 1327 197
rect 1269 118 1327 163
rect 1387 673 1445 718
rect 1387 639 1399 673
rect 1433 639 1445 673
rect 1387 605 1445 639
rect 1387 571 1399 605
rect 1433 571 1445 605
rect 1387 537 1445 571
rect 1387 503 1399 537
rect 1433 503 1445 537
rect 1387 469 1445 503
rect 1387 435 1399 469
rect 1433 435 1445 469
rect 1387 401 1445 435
rect 1387 367 1399 401
rect 1433 367 1445 401
rect 1387 333 1445 367
rect 1387 299 1399 333
rect 1433 299 1445 333
rect 1387 265 1445 299
rect 1387 231 1399 265
rect 1433 231 1445 265
rect 1387 197 1445 231
rect 1387 163 1399 197
rect 1433 163 1445 197
rect 1387 118 1445 163
rect 1505 673 1563 718
rect 1505 639 1517 673
rect 1551 639 1563 673
rect 1505 605 1563 639
rect 1505 571 1517 605
rect 1551 571 1563 605
rect 1505 537 1563 571
rect 1505 503 1517 537
rect 1551 503 1563 537
rect 1505 469 1563 503
rect 1505 435 1517 469
rect 1551 435 1563 469
rect 1505 401 1563 435
rect 1505 367 1517 401
rect 1551 367 1563 401
rect 1505 333 1563 367
rect 1505 299 1517 333
rect 1551 299 1563 333
rect 1505 265 1563 299
rect 1505 231 1517 265
rect 1551 231 1563 265
rect 1505 197 1563 231
rect 1505 163 1517 197
rect 1551 163 1563 197
rect 1505 118 1563 163
rect 1623 673 1681 718
rect 1623 639 1635 673
rect 1669 639 1681 673
rect 1623 605 1681 639
rect 1623 571 1635 605
rect 1669 571 1681 605
rect 1623 537 1681 571
rect 1623 503 1635 537
rect 1669 503 1681 537
rect 1623 469 1681 503
rect 1623 435 1635 469
rect 1669 435 1681 469
rect 1623 401 1681 435
rect 1623 367 1635 401
rect 1669 367 1681 401
rect 1623 333 1681 367
rect 1623 299 1635 333
rect 1669 299 1681 333
rect 1623 265 1681 299
rect 1623 231 1635 265
rect 1669 231 1681 265
rect 1623 197 1681 231
rect 1623 163 1635 197
rect 1669 163 1681 197
rect 1623 118 1681 163
rect 1741 673 1799 718
rect 1741 639 1753 673
rect 1787 639 1799 673
rect 1741 605 1799 639
rect 1741 571 1753 605
rect 1787 571 1799 605
rect 1741 537 1799 571
rect 1741 503 1753 537
rect 1787 503 1799 537
rect 1741 469 1799 503
rect 1741 435 1753 469
rect 1787 435 1799 469
rect 1741 401 1799 435
rect 1741 367 1753 401
rect 1787 367 1799 401
rect 1741 333 1799 367
rect 1741 299 1753 333
rect 1787 299 1799 333
rect 1741 265 1799 299
rect 1741 231 1753 265
rect 1787 231 1799 265
rect 1741 197 1799 231
rect 1741 163 1753 197
rect 1787 163 1799 197
rect 1741 118 1799 163
rect 1859 673 1917 718
rect 1859 639 1871 673
rect 1905 639 1917 673
rect 1859 605 1917 639
rect 1859 571 1871 605
rect 1905 571 1917 605
rect 1859 537 1917 571
rect 1859 503 1871 537
rect 1905 503 1917 537
rect 1859 469 1917 503
rect 1859 435 1871 469
rect 1905 435 1917 469
rect 1859 401 1917 435
rect 1859 367 1871 401
rect 1905 367 1917 401
rect 1859 333 1917 367
rect 1859 299 1871 333
rect 1905 299 1917 333
rect 1859 265 1917 299
rect 1859 231 1871 265
rect 1905 231 1917 265
rect 1859 197 1917 231
rect 1859 163 1871 197
rect 1905 163 1917 197
rect 1859 118 1917 163
rect 1977 673 2035 718
rect 1977 639 1989 673
rect 2023 639 2035 673
rect 1977 605 2035 639
rect 1977 571 1989 605
rect 2023 571 2035 605
rect 1977 537 2035 571
rect 1977 503 1989 537
rect 2023 503 2035 537
rect 1977 469 2035 503
rect 1977 435 1989 469
rect 2023 435 2035 469
rect 1977 401 2035 435
rect 1977 367 1989 401
rect 2023 367 2035 401
rect 1977 333 2035 367
rect 1977 299 1989 333
rect 2023 299 2035 333
rect 1977 265 2035 299
rect 1977 231 1989 265
rect 2023 231 2035 265
rect 1977 197 2035 231
rect 1977 163 1989 197
rect 2023 163 2035 197
rect 1977 118 2035 163
rect 2095 673 2153 718
rect 2095 639 2107 673
rect 2141 639 2153 673
rect 2095 605 2153 639
rect 2095 571 2107 605
rect 2141 571 2153 605
rect 2095 537 2153 571
rect 2095 503 2107 537
rect 2141 503 2153 537
rect 2095 469 2153 503
rect 2095 435 2107 469
rect 2141 435 2153 469
rect 2095 401 2153 435
rect 2095 367 2107 401
rect 2141 367 2153 401
rect 2095 333 2153 367
rect 2095 299 2107 333
rect 2141 299 2153 333
rect 2095 265 2153 299
rect 2095 231 2107 265
rect 2141 231 2153 265
rect 2095 197 2153 231
rect 2095 163 2107 197
rect 2141 163 2153 197
rect 2095 118 2153 163
rect 2213 673 2271 718
rect 2213 639 2225 673
rect 2259 639 2271 673
rect 2213 605 2271 639
rect 2213 571 2225 605
rect 2259 571 2271 605
rect 2213 537 2271 571
rect 2213 503 2225 537
rect 2259 503 2271 537
rect 2213 469 2271 503
rect 2213 435 2225 469
rect 2259 435 2271 469
rect 2213 401 2271 435
rect 2213 367 2225 401
rect 2259 367 2271 401
rect 2213 333 2271 367
rect 2213 299 2225 333
rect 2259 299 2271 333
rect 2213 265 2271 299
rect 2213 231 2225 265
rect 2259 231 2271 265
rect 2213 197 2271 231
rect 2213 163 2225 197
rect 2259 163 2271 197
rect 2213 118 2271 163
rect 2331 673 2389 718
rect 2331 639 2343 673
rect 2377 639 2389 673
rect 2331 605 2389 639
rect 2331 571 2343 605
rect 2377 571 2389 605
rect 2331 537 2389 571
rect 2331 503 2343 537
rect 2377 503 2389 537
rect 2331 469 2389 503
rect 2331 435 2343 469
rect 2377 435 2389 469
rect 2331 401 2389 435
rect 2331 367 2343 401
rect 2377 367 2389 401
rect 2331 333 2389 367
rect 2331 299 2343 333
rect 2377 299 2389 333
rect 2331 265 2389 299
rect 2331 231 2343 265
rect 2377 231 2389 265
rect 2331 197 2389 231
rect 2331 163 2343 197
rect 2377 163 2389 197
rect 2331 118 2389 163
rect 2449 673 2507 718
rect 2449 639 2461 673
rect 2495 639 2507 673
rect 2449 605 2507 639
rect 2449 571 2461 605
rect 2495 571 2507 605
rect 2449 537 2507 571
rect 2449 503 2461 537
rect 2495 503 2507 537
rect 2449 469 2507 503
rect 2449 435 2461 469
rect 2495 435 2507 469
rect 2449 401 2507 435
rect 2449 367 2461 401
rect 2495 367 2507 401
rect 2449 333 2507 367
rect 2449 299 2461 333
rect 2495 299 2507 333
rect 2449 265 2507 299
rect 2449 231 2461 265
rect 2495 231 2507 265
rect 2449 197 2507 231
rect 2449 163 2461 197
rect 2495 163 2507 197
rect 2449 118 2507 163
rect 2567 673 2625 718
rect 2567 639 2579 673
rect 2613 639 2625 673
rect 2567 605 2625 639
rect 2567 571 2579 605
rect 2613 571 2625 605
rect 2567 537 2625 571
rect 2567 503 2579 537
rect 2613 503 2625 537
rect 2567 469 2625 503
rect 2567 435 2579 469
rect 2613 435 2625 469
rect 2567 401 2625 435
rect 2567 367 2579 401
rect 2613 367 2625 401
rect 2567 333 2625 367
rect 2567 299 2579 333
rect 2613 299 2625 333
rect 2567 265 2625 299
rect 2567 231 2579 265
rect 2613 231 2625 265
rect 2567 197 2625 231
rect 2567 163 2579 197
rect 2613 163 2625 197
rect 2567 118 2625 163
rect 2685 673 2743 718
rect 2685 639 2697 673
rect 2731 639 2743 673
rect 2685 605 2743 639
rect 2685 571 2697 605
rect 2731 571 2743 605
rect 2685 537 2743 571
rect 2685 503 2697 537
rect 2731 503 2743 537
rect 2685 469 2743 503
rect 2685 435 2697 469
rect 2731 435 2743 469
rect 2685 401 2743 435
rect 2685 367 2697 401
rect 2731 367 2743 401
rect 2685 333 2743 367
rect 2685 299 2697 333
rect 2731 299 2743 333
rect 2685 265 2743 299
rect 2685 231 2697 265
rect 2731 231 2743 265
rect 2685 197 2743 231
rect 2685 163 2697 197
rect 2731 163 2743 197
rect 2685 118 2743 163
rect 2803 673 2861 718
rect 2803 639 2815 673
rect 2849 639 2861 673
rect 2803 605 2861 639
rect 2803 571 2815 605
rect 2849 571 2861 605
rect 2803 537 2861 571
rect 2803 503 2815 537
rect 2849 503 2861 537
rect 2803 469 2861 503
rect 2803 435 2815 469
rect 2849 435 2861 469
rect 2803 401 2861 435
rect 2803 367 2815 401
rect 2849 367 2861 401
rect 2803 333 2861 367
rect 2803 299 2815 333
rect 2849 299 2861 333
rect 2803 265 2861 299
rect 2803 231 2815 265
rect 2849 231 2861 265
rect 2803 197 2861 231
rect 2803 163 2815 197
rect 2849 163 2861 197
rect 2803 118 2861 163
rect 2921 673 2979 718
rect 2921 639 2933 673
rect 2967 639 2979 673
rect 2921 605 2979 639
rect 2921 571 2933 605
rect 2967 571 2979 605
rect 2921 537 2979 571
rect 2921 503 2933 537
rect 2967 503 2979 537
rect 2921 469 2979 503
rect 2921 435 2933 469
rect 2967 435 2979 469
rect 2921 401 2979 435
rect 2921 367 2933 401
rect 2967 367 2979 401
rect 2921 333 2979 367
rect 2921 299 2933 333
rect 2967 299 2979 333
rect 2921 265 2979 299
rect 2921 231 2933 265
rect 2967 231 2979 265
rect 2921 197 2979 231
rect 2921 163 2933 197
rect 2967 163 2979 197
rect 2921 118 2979 163
rect -2979 -163 -2921 -118
rect -2979 -197 -2967 -163
rect -2933 -197 -2921 -163
rect -2979 -231 -2921 -197
rect -2979 -265 -2967 -231
rect -2933 -265 -2921 -231
rect -2979 -299 -2921 -265
rect -2979 -333 -2967 -299
rect -2933 -333 -2921 -299
rect -2979 -367 -2921 -333
rect -2979 -401 -2967 -367
rect -2933 -401 -2921 -367
rect -2979 -435 -2921 -401
rect -2979 -469 -2967 -435
rect -2933 -469 -2921 -435
rect -2979 -503 -2921 -469
rect -2979 -537 -2967 -503
rect -2933 -537 -2921 -503
rect -2979 -571 -2921 -537
rect -2979 -605 -2967 -571
rect -2933 -605 -2921 -571
rect -2979 -639 -2921 -605
rect -2979 -673 -2967 -639
rect -2933 -673 -2921 -639
rect -2979 -718 -2921 -673
rect -2861 -163 -2803 -118
rect -2861 -197 -2849 -163
rect -2815 -197 -2803 -163
rect -2861 -231 -2803 -197
rect -2861 -265 -2849 -231
rect -2815 -265 -2803 -231
rect -2861 -299 -2803 -265
rect -2861 -333 -2849 -299
rect -2815 -333 -2803 -299
rect -2861 -367 -2803 -333
rect -2861 -401 -2849 -367
rect -2815 -401 -2803 -367
rect -2861 -435 -2803 -401
rect -2861 -469 -2849 -435
rect -2815 -469 -2803 -435
rect -2861 -503 -2803 -469
rect -2861 -537 -2849 -503
rect -2815 -537 -2803 -503
rect -2861 -571 -2803 -537
rect -2861 -605 -2849 -571
rect -2815 -605 -2803 -571
rect -2861 -639 -2803 -605
rect -2861 -673 -2849 -639
rect -2815 -673 -2803 -639
rect -2861 -718 -2803 -673
rect -2743 -163 -2685 -118
rect -2743 -197 -2731 -163
rect -2697 -197 -2685 -163
rect -2743 -231 -2685 -197
rect -2743 -265 -2731 -231
rect -2697 -265 -2685 -231
rect -2743 -299 -2685 -265
rect -2743 -333 -2731 -299
rect -2697 -333 -2685 -299
rect -2743 -367 -2685 -333
rect -2743 -401 -2731 -367
rect -2697 -401 -2685 -367
rect -2743 -435 -2685 -401
rect -2743 -469 -2731 -435
rect -2697 -469 -2685 -435
rect -2743 -503 -2685 -469
rect -2743 -537 -2731 -503
rect -2697 -537 -2685 -503
rect -2743 -571 -2685 -537
rect -2743 -605 -2731 -571
rect -2697 -605 -2685 -571
rect -2743 -639 -2685 -605
rect -2743 -673 -2731 -639
rect -2697 -673 -2685 -639
rect -2743 -718 -2685 -673
rect -2625 -163 -2567 -118
rect -2625 -197 -2613 -163
rect -2579 -197 -2567 -163
rect -2625 -231 -2567 -197
rect -2625 -265 -2613 -231
rect -2579 -265 -2567 -231
rect -2625 -299 -2567 -265
rect -2625 -333 -2613 -299
rect -2579 -333 -2567 -299
rect -2625 -367 -2567 -333
rect -2625 -401 -2613 -367
rect -2579 -401 -2567 -367
rect -2625 -435 -2567 -401
rect -2625 -469 -2613 -435
rect -2579 -469 -2567 -435
rect -2625 -503 -2567 -469
rect -2625 -537 -2613 -503
rect -2579 -537 -2567 -503
rect -2625 -571 -2567 -537
rect -2625 -605 -2613 -571
rect -2579 -605 -2567 -571
rect -2625 -639 -2567 -605
rect -2625 -673 -2613 -639
rect -2579 -673 -2567 -639
rect -2625 -718 -2567 -673
rect -2507 -163 -2449 -118
rect -2507 -197 -2495 -163
rect -2461 -197 -2449 -163
rect -2507 -231 -2449 -197
rect -2507 -265 -2495 -231
rect -2461 -265 -2449 -231
rect -2507 -299 -2449 -265
rect -2507 -333 -2495 -299
rect -2461 -333 -2449 -299
rect -2507 -367 -2449 -333
rect -2507 -401 -2495 -367
rect -2461 -401 -2449 -367
rect -2507 -435 -2449 -401
rect -2507 -469 -2495 -435
rect -2461 -469 -2449 -435
rect -2507 -503 -2449 -469
rect -2507 -537 -2495 -503
rect -2461 -537 -2449 -503
rect -2507 -571 -2449 -537
rect -2507 -605 -2495 -571
rect -2461 -605 -2449 -571
rect -2507 -639 -2449 -605
rect -2507 -673 -2495 -639
rect -2461 -673 -2449 -639
rect -2507 -718 -2449 -673
rect -2389 -163 -2331 -118
rect -2389 -197 -2377 -163
rect -2343 -197 -2331 -163
rect -2389 -231 -2331 -197
rect -2389 -265 -2377 -231
rect -2343 -265 -2331 -231
rect -2389 -299 -2331 -265
rect -2389 -333 -2377 -299
rect -2343 -333 -2331 -299
rect -2389 -367 -2331 -333
rect -2389 -401 -2377 -367
rect -2343 -401 -2331 -367
rect -2389 -435 -2331 -401
rect -2389 -469 -2377 -435
rect -2343 -469 -2331 -435
rect -2389 -503 -2331 -469
rect -2389 -537 -2377 -503
rect -2343 -537 -2331 -503
rect -2389 -571 -2331 -537
rect -2389 -605 -2377 -571
rect -2343 -605 -2331 -571
rect -2389 -639 -2331 -605
rect -2389 -673 -2377 -639
rect -2343 -673 -2331 -639
rect -2389 -718 -2331 -673
rect -2271 -163 -2213 -118
rect -2271 -197 -2259 -163
rect -2225 -197 -2213 -163
rect -2271 -231 -2213 -197
rect -2271 -265 -2259 -231
rect -2225 -265 -2213 -231
rect -2271 -299 -2213 -265
rect -2271 -333 -2259 -299
rect -2225 -333 -2213 -299
rect -2271 -367 -2213 -333
rect -2271 -401 -2259 -367
rect -2225 -401 -2213 -367
rect -2271 -435 -2213 -401
rect -2271 -469 -2259 -435
rect -2225 -469 -2213 -435
rect -2271 -503 -2213 -469
rect -2271 -537 -2259 -503
rect -2225 -537 -2213 -503
rect -2271 -571 -2213 -537
rect -2271 -605 -2259 -571
rect -2225 -605 -2213 -571
rect -2271 -639 -2213 -605
rect -2271 -673 -2259 -639
rect -2225 -673 -2213 -639
rect -2271 -718 -2213 -673
rect -2153 -163 -2095 -118
rect -2153 -197 -2141 -163
rect -2107 -197 -2095 -163
rect -2153 -231 -2095 -197
rect -2153 -265 -2141 -231
rect -2107 -265 -2095 -231
rect -2153 -299 -2095 -265
rect -2153 -333 -2141 -299
rect -2107 -333 -2095 -299
rect -2153 -367 -2095 -333
rect -2153 -401 -2141 -367
rect -2107 -401 -2095 -367
rect -2153 -435 -2095 -401
rect -2153 -469 -2141 -435
rect -2107 -469 -2095 -435
rect -2153 -503 -2095 -469
rect -2153 -537 -2141 -503
rect -2107 -537 -2095 -503
rect -2153 -571 -2095 -537
rect -2153 -605 -2141 -571
rect -2107 -605 -2095 -571
rect -2153 -639 -2095 -605
rect -2153 -673 -2141 -639
rect -2107 -673 -2095 -639
rect -2153 -718 -2095 -673
rect -2035 -163 -1977 -118
rect -2035 -197 -2023 -163
rect -1989 -197 -1977 -163
rect -2035 -231 -1977 -197
rect -2035 -265 -2023 -231
rect -1989 -265 -1977 -231
rect -2035 -299 -1977 -265
rect -2035 -333 -2023 -299
rect -1989 -333 -1977 -299
rect -2035 -367 -1977 -333
rect -2035 -401 -2023 -367
rect -1989 -401 -1977 -367
rect -2035 -435 -1977 -401
rect -2035 -469 -2023 -435
rect -1989 -469 -1977 -435
rect -2035 -503 -1977 -469
rect -2035 -537 -2023 -503
rect -1989 -537 -1977 -503
rect -2035 -571 -1977 -537
rect -2035 -605 -2023 -571
rect -1989 -605 -1977 -571
rect -2035 -639 -1977 -605
rect -2035 -673 -2023 -639
rect -1989 -673 -1977 -639
rect -2035 -718 -1977 -673
rect -1917 -163 -1859 -118
rect -1917 -197 -1905 -163
rect -1871 -197 -1859 -163
rect -1917 -231 -1859 -197
rect -1917 -265 -1905 -231
rect -1871 -265 -1859 -231
rect -1917 -299 -1859 -265
rect -1917 -333 -1905 -299
rect -1871 -333 -1859 -299
rect -1917 -367 -1859 -333
rect -1917 -401 -1905 -367
rect -1871 -401 -1859 -367
rect -1917 -435 -1859 -401
rect -1917 -469 -1905 -435
rect -1871 -469 -1859 -435
rect -1917 -503 -1859 -469
rect -1917 -537 -1905 -503
rect -1871 -537 -1859 -503
rect -1917 -571 -1859 -537
rect -1917 -605 -1905 -571
rect -1871 -605 -1859 -571
rect -1917 -639 -1859 -605
rect -1917 -673 -1905 -639
rect -1871 -673 -1859 -639
rect -1917 -718 -1859 -673
rect -1799 -163 -1741 -118
rect -1799 -197 -1787 -163
rect -1753 -197 -1741 -163
rect -1799 -231 -1741 -197
rect -1799 -265 -1787 -231
rect -1753 -265 -1741 -231
rect -1799 -299 -1741 -265
rect -1799 -333 -1787 -299
rect -1753 -333 -1741 -299
rect -1799 -367 -1741 -333
rect -1799 -401 -1787 -367
rect -1753 -401 -1741 -367
rect -1799 -435 -1741 -401
rect -1799 -469 -1787 -435
rect -1753 -469 -1741 -435
rect -1799 -503 -1741 -469
rect -1799 -537 -1787 -503
rect -1753 -537 -1741 -503
rect -1799 -571 -1741 -537
rect -1799 -605 -1787 -571
rect -1753 -605 -1741 -571
rect -1799 -639 -1741 -605
rect -1799 -673 -1787 -639
rect -1753 -673 -1741 -639
rect -1799 -718 -1741 -673
rect -1681 -163 -1623 -118
rect -1681 -197 -1669 -163
rect -1635 -197 -1623 -163
rect -1681 -231 -1623 -197
rect -1681 -265 -1669 -231
rect -1635 -265 -1623 -231
rect -1681 -299 -1623 -265
rect -1681 -333 -1669 -299
rect -1635 -333 -1623 -299
rect -1681 -367 -1623 -333
rect -1681 -401 -1669 -367
rect -1635 -401 -1623 -367
rect -1681 -435 -1623 -401
rect -1681 -469 -1669 -435
rect -1635 -469 -1623 -435
rect -1681 -503 -1623 -469
rect -1681 -537 -1669 -503
rect -1635 -537 -1623 -503
rect -1681 -571 -1623 -537
rect -1681 -605 -1669 -571
rect -1635 -605 -1623 -571
rect -1681 -639 -1623 -605
rect -1681 -673 -1669 -639
rect -1635 -673 -1623 -639
rect -1681 -718 -1623 -673
rect -1563 -163 -1505 -118
rect -1563 -197 -1551 -163
rect -1517 -197 -1505 -163
rect -1563 -231 -1505 -197
rect -1563 -265 -1551 -231
rect -1517 -265 -1505 -231
rect -1563 -299 -1505 -265
rect -1563 -333 -1551 -299
rect -1517 -333 -1505 -299
rect -1563 -367 -1505 -333
rect -1563 -401 -1551 -367
rect -1517 -401 -1505 -367
rect -1563 -435 -1505 -401
rect -1563 -469 -1551 -435
rect -1517 -469 -1505 -435
rect -1563 -503 -1505 -469
rect -1563 -537 -1551 -503
rect -1517 -537 -1505 -503
rect -1563 -571 -1505 -537
rect -1563 -605 -1551 -571
rect -1517 -605 -1505 -571
rect -1563 -639 -1505 -605
rect -1563 -673 -1551 -639
rect -1517 -673 -1505 -639
rect -1563 -718 -1505 -673
rect -1445 -163 -1387 -118
rect -1445 -197 -1433 -163
rect -1399 -197 -1387 -163
rect -1445 -231 -1387 -197
rect -1445 -265 -1433 -231
rect -1399 -265 -1387 -231
rect -1445 -299 -1387 -265
rect -1445 -333 -1433 -299
rect -1399 -333 -1387 -299
rect -1445 -367 -1387 -333
rect -1445 -401 -1433 -367
rect -1399 -401 -1387 -367
rect -1445 -435 -1387 -401
rect -1445 -469 -1433 -435
rect -1399 -469 -1387 -435
rect -1445 -503 -1387 -469
rect -1445 -537 -1433 -503
rect -1399 -537 -1387 -503
rect -1445 -571 -1387 -537
rect -1445 -605 -1433 -571
rect -1399 -605 -1387 -571
rect -1445 -639 -1387 -605
rect -1445 -673 -1433 -639
rect -1399 -673 -1387 -639
rect -1445 -718 -1387 -673
rect -1327 -163 -1269 -118
rect -1327 -197 -1315 -163
rect -1281 -197 -1269 -163
rect -1327 -231 -1269 -197
rect -1327 -265 -1315 -231
rect -1281 -265 -1269 -231
rect -1327 -299 -1269 -265
rect -1327 -333 -1315 -299
rect -1281 -333 -1269 -299
rect -1327 -367 -1269 -333
rect -1327 -401 -1315 -367
rect -1281 -401 -1269 -367
rect -1327 -435 -1269 -401
rect -1327 -469 -1315 -435
rect -1281 -469 -1269 -435
rect -1327 -503 -1269 -469
rect -1327 -537 -1315 -503
rect -1281 -537 -1269 -503
rect -1327 -571 -1269 -537
rect -1327 -605 -1315 -571
rect -1281 -605 -1269 -571
rect -1327 -639 -1269 -605
rect -1327 -673 -1315 -639
rect -1281 -673 -1269 -639
rect -1327 -718 -1269 -673
rect -1209 -163 -1151 -118
rect -1209 -197 -1197 -163
rect -1163 -197 -1151 -163
rect -1209 -231 -1151 -197
rect -1209 -265 -1197 -231
rect -1163 -265 -1151 -231
rect -1209 -299 -1151 -265
rect -1209 -333 -1197 -299
rect -1163 -333 -1151 -299
rect -1209 -367 -1151 -333
rect -1209 -401 -1197 -367
rect -1163 -401 -1151 -367
rect -1209 -435 -1151 -401
rect -1209 -469 -1197 -435
rect -1163 -469 -1151 -435
rect -1209 -503 -1151 -469
rect -1209 -537 -1197 -503
rect -1163 -537 -1151 -503
rect -1209 -571 -1151 -537
rect -1209 -605 -1197 -571
rect -1163 -605 -1151 -571
rect -1209 -639 -1151 -605
rect -1209 -673 -1197 -639
rect -1163 -673 -1151 -639
rect -1209 -718 -1151 -673
rect -1091 -163 -1033 -118
rect -1091 -197 -1079 -163
rect -1045 -197 -1033 -163
rect -1091 -231 -1033 -197
rect -1091 -265 -1079 -231
rect -1045 -265 -1033 -231
rect -1091 -299 -1033 -265
rect -1091 -333 -1079 -299
rect -1045 -333 -1033 -299
rect -1091 -367 -1033 -333
rect -1091 -401 -1079 -367
rect -1045 -401 -1033 -367
rect -1091 -435 -1033 -401
rect -1091 -469 -1079 -435
rect -1045 -469 -1033 -435
rect -1091 -503 -1033 -469
rect -1091 -537 -1079 -503
rect -1045 -537 -1033 -503
rect -1091 -571 -1033 -537
rect -1091 -605 -1079 -571
rect -1045 -605 -1033 -571
rect -1091 -639 -1033 -605
rect -1091 -673 -1079 -639
rect -1045 -673 -1033 -639
rect -1091 -718 -1033 -673
rect -973 -163 -915 -118
rect -973 -197 -961 -163
rect -927 -197 -915 -163
rect -973 -231 -915 -197
rect -973 -265 -961 -231
rect -927 -265 -915 -231
rect -973 -299 -915 -265
rect -973 -333 -961 -299
rect -927 -333 -915 -299
rect -973 -367 -915 -333
rect -973 -401 -961 -367
rect -927 -401 -915 -367
rect -973 -435 -915 -401
rect -973 -469 -961 -435
rect -927 -469 -915 -435
rect -973 -503 -915 -469
rect -973 -537 -961 -503
rect -927 -537 -915 -503
rect -973 -571 -915 -537
rect -973 -605 -961 -571
rect -927 -605 -915 -571
rect -973 -639 -915 -605
rect -973 -673 -961 -639
rect -927 -673 -915 -639
rect -973 -718 -915 -673
rect -855 -163 -797 -118
rect -855 -197 -843 -163
rect -809 -197 -797 -163
rect -855 -231 -797 -197
rect -855 -265 -843 -231
rect -809 -265 -797 -231
rect -855 -299 -797 -265
rect -855 -333 -843 -299
rect -809 -333 -797 -299
rect -855 -367 -797 -333
rect -855 -401 -843 -367
rect -809 -401 -797 -367
rect -855 -435 -797 -401
rect -855 -469 -843 -435
rect -809 -469 -797 -435
rect -855 -503 -797 -469
rect -855 -537 -843 -503
rect -809 -537 -797 -503
rect -855 -571 -797 -537
rect -855 -605 -843 -571
rect -809 -605 -797 -571
rect -855 -639 -797 -605
rect -855 -673 -843 -639
rect -809 -673 -797 -639
rect -855 -718 -797 -673
rect -737 -163 -679 -118
rect -737 -197 -725 -163
rect -691 -197 -679 -163
rect -737 -231 -679 -197
rect -737 -265 -725 -231
rect -691 -265 -679 -231
rect -737 -299 -679 -265
rect -737 -333 -725 -299
rect -691 -333 -679 -299
rect -737 -367 -679 -333
rect -737 -401 -725 -367
rect -691 -401 -679 -367
rect -737 -435 -679 -401
rect -737 -469 -725 -435
rect -691 -469 -679 -435
rect -737 -503 -679 -469
rect -737 -537 -725 -503
rect -691 -537 -679 -503
rect -737 -571 -679 -537
rect -737 -605 -725 -571
rect -691 -605 -679 -571
rect -737 -639 -679 -605
rect -737 -673 -725 -639
rect -691 -673 -679 -639
rect -737 -718 -679 -673
rect -619 -163 -561 -118
rect -619 -197 -607 -163
rect -573 -197 -561 -163
rect -619 -231 -561 -197
rect -619 -265 -607 -231
rect -573 -265 -561 -231
rect -619 -299 -561 -265
rect -619 -333 -607 -299
rect -573 -333 -561 -299
rect -619 -367 -561 -333
rect -619 -401 -607 -367
rect -573 -401 -561 -367
rect -619 -435 -561 -401
rect -619 -469 -607 -435
rect -573 -469 -561 -435
rect -619 -503 -561 -469
rect -619 -537 -607 -503
rect -573 -537 -561 -503
rect -619 -571 -561 -537
rect -619 -605 -607 -571
rect -573 -605 -561 -571
rect -619 -639 -561 -605
rect -619 -673 -607 -639
rect -573 -673 -561 -639
rect -619 -718 -561 -673
rect -501 -163 -443 -118
rect -501 -197 -489 -163
rect -455 -197 -443 -163
rect -501 -231 -443 -197
rect -501 -265 -489 -231
rect -455 -265 -443 -231
rect -501 -299 -443 -265
rect -501 -333 -489 -299
rect -455 -333 -443 -299
rect -501 -367 -443 -333
rect -501 -401 -489 -367
rect -455 -401 -443 -367
rect -501 -435 -443 -401
rect -501 -469 -489 -435
rect -455 -469 -443 -435
rect -501 -503 -443 -469
rect -501 -537 -489 -503
rect -455 -537 -443 -503
rect -501 -571 -443 -537
rect -501 -605 -489 -571
rect -455 -605 -443 -571
rect -501 -639 -443 -605
rect -501 -673 -489 -639
rect -455 -673 -443 -639
rect -501 -718 -443 -673
rect -383 -163 -325 -118
rect -383 -197 -371 -163
rect -337 -197 -325 -163
rect -383 -231 -325 -197
rect -383 -265 -371 -231
rect -337 -265 -325 -231
rect -383 -299 -325 -265
rect -383 -333 -371 -299
rect -337 -333 -325 -299
rect -383 -367 -325 -333
rect -383 -401 -371 -367
rect -337 -401 -325 -367
rect -383 -435 -325 -401
rect -383 -469 -371 -435
rect -337 -469 -325 -435
rect -383 -503 -325 -469
rect -383 -537 -371 -503
rect -337 -537 -325 -503
rect -383 -571 -325 -537
rect -383 -605 -371 -571
rect -337 -605 -325 -571
rect -383 -639 -325 -605
rect -383 -673 -371 -639
rect -337 -673 -325 -639
rect -383 -718 -325 -673
rect -265 -163 -207 -118
rect -265 -197 -253 -163
rect -219 -197 -207 -163
rect -265 -231 -207 -197
rect -265 -265 -253 -231
rect -219 -265 -207 -231
rect -265 -299 -207 -265
rect -265 -333 -253 -299
rect -219 -333 -207 -299
rect -265 -367 -207 -333
rect -265 -401 -253 -367
rect -219 -401 -207 -367
rect -265 -435 -207 -401
rect -265 -469 -253 -435
rect -219 -469 -207 -435
rect -265 -503 -207 -469
rect -265 -537 -253 -503
rect -219 -537 -207 -503
rect -265 -571 -207 -537
rect -265 -605 -253 -571
rect -219 -605 -207 -571
rect -265 -639 -207 -605
rect -265 -673 -253 -639
rect -219 -673 -207 -639
rect -265 -718 -207 -673
rect -147 -163 -89 -118
rect -147 -197 -135 -163
rect -101 -197 -89 -163
rect -147 -231 -89 -197
rect -147 -265 -135 -231
rect -101 -265 -89 -231
rect -147 -299 -89 -265
rect -147 -333 -135 -299
rect -101 -333 -89 -299
rect -147 -367 -89 -333
rect -147 -401 -135 -367
rect -101 -401 -89 -367
rect -147 -435 -89 -401
rect -147 -469 -135 -435
rect -101 -469 -89 -435
rect -147 -503 -89 -469
rect -147 -537 -135 -503
rect -101 -537 -89 -503
rect -147 -571 -89 -537
rect -147 -605 -135 -571
rect -101 -605 -89 -571
rect -147 -639 -89 -605
rect -147 -673 -135 -639
rect -101 -673 -89 -639
rect -147 -718 -89 -673
rect -29 -163 29 -118
rect -29 -197 -17 -163
rect 17 -197 29 -163
rect -29 -231 29 -197
rect -29 -265 -17 -231
rect 17 -265 29 -231
rect -29 -299 29 -265
rect -29 -333 -17 -299
rect 17 -333 29 -299
rect -29 -367 29 -333
rect -29 -401 -17 -367
rect 17 -401 29 -367
rect -29 -435 29 -401
rect -29 -469 -17 -435
rect 17 -469 29 -435
rect -29 -503 29 -469
rect -29 -537 -17 -503
rect 17 -537 29 -503
rect -29 -571 29 -537
rect -29 -605 -17 -571
rect 17 -605 29 -571
rect -29 -639 29 -605
rect -29 -673 -17 -639
rect 17 -673 29 -639
rect -29 -718 29 -673
rect 89 -163 147 -118
rect 89 -197 101 -163
rect 135 -197 147 -163
rect 89 -231 147 -197
rect 89 -265 101 -231
rect 135 -265 147 -231
rect 89 -299 147 -265
rect 89 -333 101 -299
rect 135 -333 147 -299
rect 89 -367 147 -333
rect 89 -401 101 -367
rect 135 -401 147 -367
rect 89 -435 147 -401
rect 89 -469 101 -435
rect 135 -469 147 -435
rect 89 -503 147 -469
rect 89 -537 101 -503
rect 135 -537 147 -503
rect 89 -571 147 -537
rect 89 -605 101 -571
rect 135 -605 147 -571
rect 89 -639 147 -605
rect 89 -673 101 -639
rect 135 -673 147 -639
rect 89 -718 147 -673
rect 207 -163 265 -118
rect 207 -197 219 -163
rect 253 -197 265 -163
rect 207 -231 265 -197
rect 207 -265 219 -231
rect 253 -265 265 -231
rect 207 -299 265 -265
rect 207 -333 219 -299
rect 253 -333 265 -299
rect 207 -367 265 -333
rect 207 -401 219 -367
rect 253 -401 265 -367
rect 207 -435 265 -401
rect 207 -469 219 -435
rect 253 -469 265 -435
rect 207 -503 265 -469
rect 207 -537 219 -503
rect 253 -537 265 -503
rect 207 -571 265 -537
rect 207 -605 219 -571
rect 253 -605 265 -571
rect 207 -639 265 -605
rect 207 -673 219 -639
rect 253 -673 265 -639
rect 207 -718 265 -673
rect 325 -163 383 -118
rect 325 -197 337 -163
rect 371 -197 383 -163
rect 325 -231 383 -197
rect 325 -265 337 -231
rect 371 -265 383 -231
rect 325 -299 383 -265
rect 325 -333 337 -299
rect 371 -333 383 -299
rect 325 -367 383 -333
rect 325 -401 337 -367
rect 371 -401 383 -367
rect 325 -435 383 -401
rect 325 -469 337 -435
rect 371 -469 383 -435
rect 325 -503 383 -469
rect 325 -537 337 -503
rect 371 -537 383 -503
rect 325 -571 383 -537
rect 325 -605 337 -571
rect 371 -605 383 -571
rect 325 -639 383 -605
rect 325 -673 337 -639
rect 371 -673 383 -639
rect 325 -718 383 -673
rect 443 -163 501 -118
rect 443 -197 455 -163
rect 489 -197 501 -163
rect 443 -231 501 -197
rect 443 -265 455 -231
rect 489 -265 501 -231
rect 443 -299 501 -265
rect 443 -333 455 -299
rect 489 -333 501 -299
rect 443 -367 501 -333
rect 443 -401 455 -367
rect 489 -401 501 -367
rect 443 -435 501 -401
rect 443 -469 455 -435
rect 489 -469 501 -435
rect 443 -503 501 -469
rect 443 -537 455 -503
rect 489 -537 501 -503
rect 443 -571 501 -537
rect 443 -605 455 -571
rect 489 -605 501 -571
rect 443 -639 501 -605
rect 443 -673 455 -639
rect 489 -673 501 -639
rect 443 -718 501 -673
rect 561 -163 619 -118
rect 561 -197 573 -163
rect 607 -197 619 -163
rect 561 -231 619 -197
rect 561 -265 573 -231
rect 607 -265 619 -231
rect 561 -299 619 -265
rect 561 -333 573 -299
rect 607 -333 619 -299
rect 561 -367 619 -333
rect 561 -401 573 -367
rect 607 -401 619 -367
rect 561 -435 619 -401
rect 561 -469 573 -435
rect 607 -469 619 -435
rect 561 -503 619 -469
rect 561 -537 573 -503
rect 607 -537 619 -503
rect 561 -571 619 -537
rect 561 -605 573 -571
rect 607 -605 619 -571
rect 561 -639 619 -605
rect 561 -673 573 -639
rect 607 -673 619 -639
rect 561 -718 619 -673
rect 679 -163 737 -118
rect 679 -197 691 -163
rect 725 -197 737 -163
rect 679 -231 737 -197
rect 679 -265 691 -231
rect 725 -265 737 -231
rect 679 -299 737 -265
rect 679 -333 691 -299
rect 725 -333 737 -299
rect 679 -367 737 -333
rect 679 -401 691 -367
rect 725 -401 737 -367
rect 679 -435 737 -401
rect 679 -469 691 -435
rect 725 -469 737 -435
rect 679 -503 737 -469
rect 679 -537 691 -503
rect 725 -537 737 -503
rect 679 -571 737 -537
rect 679 -605 691 -571
rect 725 -605 737 -571
rect 679 -639 737 -605
rect 679 -673 691 -639
rect 725 -673 737 -639
rect 679 -718 737 -673
rect 797 -163 855 -118
rect 797 -197 809 -163
rect 843 -197 855 -163
rect 797 -231 855 -197
rect 797 -265 809 -231
rect 843 -265 855 -231
rect 797 -299 855 -265
rect 797 -333 809 -299
rect 843 -333 855 -299
rect 797 -367 855 -333
rect 797 -401 809 -367
rect 843 -401 855 -367
rect 797 -435 855 -401
rect 797 -469 809 -435
rect 843 -469 855 -435
rect 797 -503 855 -469
rect 797 -537 809 -503
rect 843 -537 855 -503
rect 797 -571 855 -537
rect 797 -605 809 -571
rect 843 -605 855 -571
rect 797 -639 855 -605
rect 797 -673 809 -639
rect 843 -673 855 -639
rect 797 -718 855 -673
rect 915 -163 973 -118
rect 915 -197 927 -163
rect 961 -197 973 -163
rect 915 -231 973 -197
rect 915 -265 927 -231
rect 961 -265 973 -231
rect 915 -299 973 -265
rect 915 -333 927 -299
rect 961 -333 973 -299
rect 915 -367 973 -333
rect 915 -401 927 -367
rect 961 -401 973 -367
rect 915 -435 973 -401
rect 915 -469 927 -435
rect 961 -469 973 -435
rect 915 -503 973 -469
rect 915 -537 927 -503
rect 961 -537 973 -503
rect 915 -571 973 -537
rect 915 -605 927 -571
rect 961 -605 973 -571
rect 915 -639 973 -605
rect 915 -673 927 -639
rect 961 -673 973 -639
rect 915 -718 973 -673
rect 1033 -163 1091 -118
rect 1033 -197 1045 -163
rect 1079 -197 1091 -163
rect 1033 -231 1091 -197
rect 1033 -265 1045 -231
rect 1079 -265 1091 -231
rect 1033 -299 1091 -265
rect 1033 -333 1045 -299
rect 1079 -333 1091 -299
rect 1033 -367 1091 -333
rect 1033 -401 1045 -367
rect 1079 -401 1091 -367
rect 1033 -435 1091 -401
rect 1033 -469 1045 -435
rect 1079 -469 1091 -435
rect 1033 -503 1091 -469
rect 1033 -537 1045 -503
rect 1079 -537 1091 -503
rect 1033 -571 1091 -537
rect 1033 -605 1045 -571
rect 1079 -605 1091 -571
rect 1033 -639 1091 -605
rect 1033 -673 1045 -639
rect 1079 -673 1091 -639
rect 1033 -718 1091 -673
rect 1151 -163 1209 -118
rect 1151 -197 1163 -163
rect 1197 -197 1209 -163
rect 1151 -231 1209 -197
rect 1151 -265 1163 -231
rect 1197 -265 1209 -231
rect 1151 -299 1209 -265
rect 1151 -333 1163 -299
rect 1197 -333 1209 -299
rect 1151 -367 1209 -333
rect 1151 -401 1163 -367
rect 1197 -401 1209 -367
rect 1151 -435 1209 -401
rect 1151 -469 1163 -435
rect 1197 -469 1209 -435
rect 1151 -503 1209 -469
rect 1151 -537 1163 -503
rect 1197 -537 1209 -503
rect 1151 -571 1209 -537
rect 1151 -605 1163 -571
rect 1197 -605 1209 -571
rect 1151 -639 1209 -605
rect 1151 -673 1163 -639
rect 1197 -673 1209 -639
rect 1151 -718 1209 -673
rect 1269 -163 1327 -118
rect 1269 -197 1281 -163
rect 1315 -197 1327 -163
rect 1269 -231 1327 -197
rect 1269 -265 1281 -231
rect 1315 -265 1327 -231
rect 1269 -299 1327 -265
rect 1269 -333 1281 -299
rect 1315 -333 1327 -299
rect 1269 -367 1327 -333
rect 1269 -401 1281 -367
rect 1315 -401 1327 -367
rect 1269 -435 1327 -401
rect 1269 -469 1281 -435
rect 1315 -469 1327 -435
rect 1269 -503 1327 -469
rect 1269 -537 1281 -503
rect 1315 -537 1327 -503
rect 1269 -571 1327 -537
rect 1269 -605 1281 -571
rect 1315 -605 1327 -571
rect 1269 -639 1327 -605
rect 1269 -673 1281 -639
rect 1315 -673 1327 -639
rect 1269 -718 1327 -673
rect 1387 -163 1445 -118
rect 1387 -197 1399 -163
rect 1433 -197 1445 -163
rect 1387 -231 1445 -197
rect 1387 -265 1399 -231
rect 1433 -265 1445 -231
rect 1387 -299 1445 -265
rect 1387 -333 1399 -299
rect 1433 -333 1445 -299
rect 1387 -367 1445 -333
rect 1387 -401 1399 -367
rect 1433 -401 1445 -367
rect 1387 -435 1445 -401
rect 1387 -469 1399 -435
rect 1433 -469 1445 -435
rect 1387 -503 1445 -469
rect 1387 -537 1399 -503
rect 1433 -537 1445 -503
rect 1387 -571 1445 -537
rect 1387 -605 1399 -571
rect 1433 -605 1445 -571
rect 1387 -639 1445 -605
rect 1387 -673 1399 -639
rect 1433 -673 1445 -639
rect 1387 -718 1445 -673
rect 1505 -163 1563 -118
rect 1505 -197 1517 -163
rect 1551 -197 1563 -163
rect 1505 -231 1563 -197
rect 1505 -265 1517 -231
rect 1551 -265 1563 -231
rect 1505 -299 1563 -265
rect 1505 -333 1517 -299
rect 1551 -333 1563 -299
rect 1505 -367 1563 -333
rect 1505 -401 1517 -367
rect 1551 -401 1563 -367
rect 1505 -435 1563 -401
rect 1505 -469 1517 -435
rect 1551 -469 1563 -435
rect 1505 -503 1563 -469
rect 1505 -537 1517 -503
rect 1551 -537 1563 -503
rect 1505 -571 1563 -537
rect 1505 -605 1517 -571
rect 1551 -605 1563 -571
rect 1505 -639 1563 -605
rect 1505 -673 1517 -639
rect 1551 -673 1563 -639
rect 1505 -718 1563 -673
rect 1623 -163 1681 -118
rect 1623 -197 1635 -163
rect 1669 -197 1681 -163
rect 1623 -231 1681 -197
rect 1623 -265 1635 -231
rect 1669 -265 1681 -231
rect 1623 -299 1681 -265
rect 1623 -333 1635 -299
rect 1669 -333 1681 -299
rect 1623 -367 1681 -333
rect 1623 -401 1635 -367
rect 1669 -401 1681 -367
rect 1623 -435 1681 -401
rect 1623 -469 1635 -435
rect 1669 -469 1681 -435
rect 1623 -503 1681 -469
rect 1623 -537 1635 -503
rect 1669 -537 1681 -503
rect 1623 -571 1681 -537
rect 1623 -605 1635 -571
rect 1669 -605 1681 -571
rect 1623 -639 1681 -605
rect 1623 -673 1635 -639
rect 1669 -673 1681 -639
rect 1623 -718 1681 -673
rect 1741 -163 1799 -118
rect 1741 -197 1753 -163
rect 1787 -197 1799 -163
rect 1741 -231 1799 -197
rect 1741 -265 1753 -231
rect 1787 -265 1799 -231
rect 1741 -299 1799 -265
rect 1741 -333 1753 -299
rect 1787 -333 1799 -299
rect 1741 -367 1799 -333
rect 1741 -401 1753 -367
rect 1787 -401 1799 -367
rect 1741 -435 1799 -401
rect 1741 -469 1753 -435
rect 1787 -469 1799 -435
rect 1741 -503 1799 -469
rect 1741 -537 1753 -503
rect 1787 -537 1799 -503
rect 1741 -571 1799 -537
rect 1741 -605 1753 -571
rect 1787 -605 1799 -571
rect 1741 -639 1799 -605
rect 1741 -673 1753 -639
rect 1787 -673 1799 -639
rect 1741 -718 1799 -673
rect 1859 -163 1917 -118
rect 1859 -197 1871 -163
rect 1905 -197 1917 -163
rect 1859 -231 1917 -197
rect 1859 -265 1871 -231
rect 1905 -265 1917 -231
rect 1859 -299 1917 -265
rect 1859 -333 1871 -299
rect 1905 -333 1917 -299
rect 1859 -367 1917 -333
rect 1859 -401 1871 -367
rect 1905 -401 1917 -367
rect 1859 -435 1917 -401
rect 1859 -469 1871 -435
rect 1905 -469 1917 -435
rect 1859 -503 1917 -469
rect 1859 -537 1871 -503
rect 1905 -537 1917 -503
rect 1859 -571 1917 -537
rect 1859 -605 1871 -571
rect 1905 -605 1917 -571
rect 1859 -639 1917 -605
rect 1859 -673 1871 -639
rect 1905 -673 1917 -639
rect 1859 -718 1917 -673
rect 1977 -163 2035 -118
rect 1977 -197 1989 -163
rect 2023 -197 2035 -163
rect 1977 -231 2035 -197
rect 1977 -265 1989 -231
rect 2023 -265 2035 -231
rect 1977 -299 2035 -265
rect 1977 -333 1989 -299
rect 2023 -333 2035 -299
rect 1977 -367 2035 -333
rect 1977 -401 1989 -367
rect 2023 -401 2035 -367
rect 1977 -435 2035 -401
rect 1977 -469 1989 -435
rect 2023 -469 2035 -435
rect 1977 -503 2035 -469
rect 1977 -537 1989 -503
rect 2023 -537 2035 -503
rect 1977 -571 2035 -537
rect 1977 -605 1989 -571
rect 2023 -605 2035 -571
rect 1977 -639 2035 -605
rect 1977 -673 1989 -639
rect 2023 -673 2035 -639
rect 1977 -718 2035 -673
rect 2095 -163 2153 -118
rect 2095 -197 2107 -163
rect 2141 -197 2153 -163
rect 2095 -231 2153 -197
rect 2095 -265 2107 -231
rect 2141 -265 2153 -231
rect 2095 -299 2153 -265
rect 2095 -333 2107 -299
rect 2141 -333 2153 -299
rect 2095 -367 2153 -333
rect 2095 -401 2107 -367
rect 2141 -401 2153 -367
rect 2095 -435 2153 -401
rect 2095 -469 2107 -435
rect 2141 -469 2153 -435
rect 2095 -503 2153 -469
rect 2095 -537 2107 -503
rect 2141 -537 2153 -503
rect 2095 -571 2153 -537
rect 2095 -605 2107 -571
rect 2141 -605 2153 -571
rect 2095 -639 2153 -605
rect 2095 -673 2107 -639
rect 2141 -673 2153 -639
rect 2095 -718 2153 -673
rect 2213 -163 2271 -118
rect 2213 -197 2225 -163
rect 2259 -197 2271 -163
rect 2213 -231 2271 -197
rect 2213 -265 2225 -231
rect 2259 -265 2271 -231
rect 2213 -299 2271 -265
rect 2213 -333 2225 -299
rect 2259 -333 2271 -299
rect 2213 -367 2271 -333
rect 2213 -401 2225 -367
rect 2259 -401 2271 -367
rect 2213 -435 2271 -401
rect 2213 -469 2225 -435
rect 2259 -469 2271 -435
rect 2213 -503 2271 -469
rect 2213 -537 2225 -503
rect 2259 -537 2271 -503
rect 2213 -571 2271 -537
rect 2213 -605 2225 -571
rect 2259 -605 2271 -571
rect 2213 -639 2271 -605
rect 2213 -673 2225 -639
rect 2259 -673 2271 -639
rect 2213 -718 2271 -673
rect 2331 -163 2389 -118
rect 2331 -197 2343 -163
rect 2377 -197 2389 -163
rect 2331 -231 2389 -197
rect 2331 -265 2343 -231
rect 2377 -265 2389 -231
rect 2331 -299 2389 -265
rect 2331 -333 2343 -299
rect 2377 -333 2389 -299
rect 2331 -367 2389 -333
rect 2331 -401 2343 -367
rect 2377 -401 2389 -367
rect 2331 -435 2389 -401
rect 2331 -469 2343 -435
rect 2377 -469 2389 -435
rect 2331 -503 2389 -469
rect 2331 -537 2343 -503
rect 2377 -537 2389 -503
rect 2331 -571 2389 -537
rect 2331 -605 2343 -571
rect 2377 -605 2389 -571
rect 2331 -639 2389 -605
rect 2331 -673 2343 -639
rect 2377 -673 2389 -639
rect 2331 -718 2389 -673
rect 2449 -163 2507 -118
rect 2449 -197 2461 -163
rect 2495 -197 2507 -163
rect 2449 -231 2507 -197
rect 2449 -265 2461 -231
rect 2495 -265 2507 -231
rect 2449 -299 2507 -265
rect 2449 -333 2461 -299
rect 2495 -333 2507 -299
rect 2449 -367 2507 -333
rect 2449 -401 2461 -367
rect 2495 -401 2507 -367
rect 2449 -435 2507 -401
rect 2449 -469 2461 -435
rect 2495 -469 2507 -435
rect 2449 -503 2507 -469
rect 2449 -537 2461 -503
rect 2495 -537 2507 -503
rect 2449 -571 2507 -537
rect 2449 -605 2461 -571
rect 2495 -605 2507 -571
rect 2449 -639 2507 -605
rect 2449 -673 2461 -639
rect 2495 -673 2507 -639
rect 2449 -718 2507 -673
rect 2567 -163 2625 -118
rect 2567 -197 2579 -163
rect 2613 -197 2625 -163
rect 2567 -231 2625 -197
rect 2567 -265 2579 -231
rect 2613 -265 2625 -231
rect 2567 -299 2625 -265
rect 2567 -333 2579 -299
rect 2613 -333 2625 -299
rect 2567 -367 2625 -333
rect 2567 -401 2579 -367
rect 2613 -401 2625 -367
rect 2567 -435 2625 -401
rect 2567 -469 2579 -435
rect 2613 -469 2625 -435
rect 2567 -503 2625 -469
rect 2567 -537 2579 -503
rect 2613 -537 2625 -503
rect 2567 -571 2625 -537
rect 2567 -605 2579 -571
rect 2613 -605 2625 -571
rect 2567 -639 2625 -605
rect 2567 -673 2579 -639
rect 2613 -673 2625 -639
rect 2567 -718 2625 -673
rect 2685 -163 2743 -118
rect 2685 -197 2697 -163
rect 2731 -197 2743 -163
rect 2685 -231 2743 -197
rect 2685 -265 2697 -231
rect 2731 -265 2743 -231
rect 2685 -299 2743 -265
rect 2685 -333 2697 -299
rect 2731 -333 2743 -299
rect 2685 -367 2743 -333
rect 2685 -401 2697 -367
rect 2731 -401 2743 -367
rect 2685 -435 2743 -401
rect 2685 -469 2697 -435
rect 2731 -469 2743 -435
rect 2685 -503 2743 -469
rect 2685 -537 2697 -503
rect 2731 -537 2743 -503
rect 2685 -571 2743 -537
rect 2685 -605 2697 -571
rect 2731 -605 2743 -571
rect 2685 -639 2743 -605
rect 2685 -673 2697 -639
rect 2731 -673 2743 -639
rect 2685 -718 2743 -673
rect 2803 -163 2861 -118
rect 2803 -197 2815 -163
rect 2849 -197 2861 -163
rect 2803 -231 2861 -197
rect 2803 -265 2815 -231
rect 2849 -265 2861 -231
rect 2803 -299 2861 -265
rect 2803 -333 2815 -299
rect 2849 -333 2861 -299
rect 2803 -367 2861 -333
rect 2803 -401 2815 -367
rect 2849 -401 2861 -367
rect 2803 -435 2861 -401
rect 2803 -469 2815 -435
rect 2849 -469 2861 -435
rect 2803 -503 2861 -469
rect 2803 -537 2815 -503
rect 2849 -537 2861 -503
rect 2803 -571 2861 -537
rect 2803 -605 2815 -571
rect 2849 -605 2861 -571
rect 2803 -639 2861 -605
rect 2803 -673 2815 -639
rect 2849 -673 2861 -639
rect 2803 -718 2861 -673
rect 2921 -163 2979 -118
rect 2921 -197 2933 -163
rect 2967 -197 2979 -163
rect 2921 -231 2979 -197
rect 2921 -265 2933 -231
rect 2967 -265 2979 -231
rect 2921 -299 2979 -265
rect 2921 -333 2933 -299
rect 2967 -333 2979 -299
rect 2921 -367 2979 -333
rect 2921 -401 2933 -367
rect 2967 -401 2979 -367
rect 2921 -435 2979 -401
rect 2921 -469 2933 -435
rect 2967 -469 2979 -435
rect 2921 -503 2979 -469
rect 2921 -537 2933 -503
rect 2967 -537 2979 -503
rect 2921 -571 2979 -537
rect 2921 -605 2933 -571
rect 2967 -605 2979 -571
rect 2921 -639 2979 -605
rect 2921 -673 2933 -639
rect 2967 -673 2979 -639
rect 2921 -718 2979 -673
<< pdiffc >>
rect -2967 639 -2933 673
rect -2967 571 -2933 605
rect -2967 503 -2933 537
rect -2967 435 -2933 469
rect -2967 367 -2933 401
rect -2967 299 -2933 333
rect -2967 231 -2933 265
rect -2967 163 -2933 197
rect -2849 639 -2815 673
rect -2849 571 -2815 605
rect -2849 503 -2815 537
rect -2849 435 -2815 469
rect -2849 367 -2815 401
rect -2849 299 -2815 333
rect -2849 231 -2815 265
rect -2849 163 -2815 197
rect -2731 639 -2697 673
rect -2731 571 -2697 605
rect -2731 503 -2697 537
rect -2731 435 -2697 469
rect -2731 367 -2697 401
rect -2731 299 -2697 333
rect -2731 231 -2697 265
rect -2731 163 -2697 197
rect -2613 639 -2579 673
rect -2613 571 -2579 605
rect -2613 503 -2579 537
rect -2613 435 -2579 469
rect -2613 367 -2579 401
rect -2613 299 -2579 333
rect -2613 231 -2579 265
rect -2613 163 -2579 197
rect -2495 639 -2461 673
rect -2495 571 -2461 605
rect -2495 503 -2461 537
rect -2495 435 -2461 469
rect -2495 367 -2461 401
rect -2495 299 -2461 333
rect -2495 231 -2461 265
rect -2495 163 -2461 197
rect -2377 639 -2343 673
rect -2377 571 -2343 605
rect -2377 503 -2343 537
rect -2377 435 -2343 469
rect -2377 367 -2343 401
rect -2377 299 -2343 333
rect -2377 231 -2343 265
rect -2377 163 -2343 197
rect -2259 639 -2225 673
rect -2259 571 -2225 605
rect -2259 503 -2225 537
rect -2259 435 -2225 469
rect -2259 367 -2225 401
rect -2259 299 -2225 333
rect -2259 231 -2225 265
rect -2259 163 -2225 197
rect -2141 639 -2107 673
rect -2141 571 -2107 605
rect -2141 503 -2107 537
rect -2141 435 -2107 469
rect -2141 367 -2107 401
rect -2141 299 -2107 333
rect -2141 231 -2107 265
rect -2141 163 -2107 197
rect -2023 639 -1989 673
rect -2023 571 -1989 605
rect -2023 503 -1989 537
rect -2023 435 -1989 469
rect -2023 367 -1989 401
rect -2023 299 -1989 333
rect -2023 231 -1989 265
rect -2023 163 -1989 197
rect -1905 639 -1871 673
rect -1905 571 -1871 605
rect -1905 503 -1871 537
rect -1905 435 -1871 469
rect -1905 367 -1871 401
rect -1905 299 -1871 333
rect -1905 231 -1871 265
rect -1905 163 -1871 197
rect -1787 639 -1753 673
rect -1787 571 -1753 605
rect -1787 503 -1753 537
rect -1787 435 -1753 469
rect -1787 367 -1753 401
rect -1787 299 -1753 333
rect -1787 231 -1753 265
rect -1787 163 -1753 197
rect -1669 639 -1635 673
rect -1669 571 -1635 605
rect -1669 503 -1635 537
rect -1669 435 -1635 469
rect -1669 367 -1635 401
rect -1669 299 -1635 333
rect -1669 231 -1635 265
rect -1669 163 -1635 197
rect -1551 639 -1517 673
rect -1551 571 -1517 605
rect -1551 503 -1517 537
rect -1551 435 -1517 469
rect -1551 367 -1517 401
rect -1551 299 -1517 333
rect -1551 231 -1517 265
rect -1551 163 -1517 197
rect -1433 639 -1399 673
rect -1433 571 -1399 605
rect -1433 503 -1399 537
rect -1433 435 -1399 469
rect -1433 367 -1399 401
rect -1433 299 -1399 333
rect -1433 231 -1399 265
rect -1433 163 -1399 197
rect -1315 639 -1281 673
rect -1315 571 -1281 605
rect -1315 503 -1281 537
rect -1315 435 -1281 469
rect -1315 367 -1281 401
rect -1315 299 -1281 333
rect -1315 231 -1281 265
rect -1315 163 -1281 197
rect -1197 639 -1163 673
rect -1197 571 -1163 605
rect -1197 503 -1163 537
rect -1197 435 -1163 469
rect -1197 367 -1163 401
rect -1197 299 -1163 333
rect -1197 231 -1163 265
rect -1197 163 -1163 197
rect -1079 639 -1045 673
rect -1079 571 -1045 605
rect -1079 503 -1045 537
rect -1079 435 -1045 469
rect -1079 367 -1045 401
rect -1079 299 -1045 333
rect -1079 231 -1045 265
rect -1079 163 -1045 197
rect -961 639 -927 673
rect -961 571 -927 605
rect -961 503 -927 537
rect -961 435 -927 469
rect -961 367 -927 401
rect -961 299 -927 333
rect -961 231 -927 265
rect -961 163 -927 197
rect -843 639 -809 673
rect -843 571 -809 605
rect -843 503 -809 537
rect -843 435 -809 469
rect -843 367 -809 401
rect -843 299 -809 333
rect -843 231 -809 265
rect -843 163 -809 197
rect -725 639 -691 673
rect -725 571 -691 605
rect -725 503 -691 537
rect -725 435 -691 469
rect -725 367 -691 401
rect -725 299 -691 333
rect -725 231 -691 265
rect -725 163 -691 197
rect -607 639 -573 673
rect -607 571 -573 605
rect -607 503 -573 537
rect -607 435 -573 469
rect -607 367 -573 401
rect -607 299 -573 333
rect -607 231 -573 265
rect -607 163 -573 197
rect -489 639 -455 673
rect -489 571 -455 605
rect -489 503 -455 537
rect -489 435 -455 469
rect -489 367 -455 401
rect -489 299 -455 333
rect -489 231 -455 265
rect -489 163 -455 197
rect -371 639 -337 673
rect -371 571 -337 605
rect -371 503 -337 537
rect -371 435 -337 469
rect -371 367 -337 401
rect -371 299 -337 333
rect -371 231 -337 265
rect -371 163 -337 197
rect -253 639 -219 673
rect -253 571 -219 605
rect -253 503 -219 537
rect -253 435 -219 469
rect -253 367 -219 401
rect -253 299 -219 333
rect -253 231 -219 265
rect -253 163 -219 197
rect -135 639 -101 673
rect -135 571 -101 605
rect -135 503 -101 537
rect -135 435 -101 469
rect -135 367 -101 401
rect -135 299 -101 333
rect -135 231 -101 265
rect -135 163 -101 197
rect -17 639 17 673
rect -17 571 17 605
rect -17 503 17 537
rect -17 435 17 469
rect -17 367 17 401
rect -17 299 17 333
rect -17 231 17 265
rect -17 163 17 197
rect 101 639 135 673
rect 101 571 135 605
rect 101 503 135 537
rect 101 435 135 469
rect 101 367 135 401
rect 101 299 135 333
rect 101 231 135 265
rect 101 163 135 197
rect 219 639 253 673
rect 219 571 253 605
rect 219 503 253 537
rect 219 435 253 469
rect 219 367 253 401
rect 219 299 253 333
rect 219 231 253 265
rect 219 163 253 197
rect 337 639 371 673
rect 337 571 371 605
rect 337 503 371 537
rect 337 435 371 469
rect 337 367 371 401
rect 337 299 371 333
rect 337 231 371 265
rect 337 163 371 197
rect 455 639 489 673
rect 455 571 489 605
rect 455 503 489 537
rect 455 435 489 469
rect 455 367 489 401
rect 455 299 489 333
rect 455 231 489 265
rect 455 163 489 197
rect 573 639 607 673
rect 573 571 607 605
rect 573 503 607 537
rect 573 435 607 469
rect 573 367 607 401
rect 573 299 607 333
rect 573 231 607 265
rect 573 163 607 197
rect 691 639 725 673
rect 691 571 725 605
rect 691 503 725 537
rect 691 435 725 469
rect 691 367 725 401
rect 691 299 725 333
rect 691 231 725 265
rect 691 163 725 197
rect 809 639 843 673
rect 809 571 843 605
rect 809 503 843 537
rect 809 435 843 469
rect 809 367 843 401
rect 809 299 843 333
rect 809 231 843 265
rect 809 163 843 197
rect 927 639 961 673
rect 927 571 961 605
rect 927 503 961 537
rect 927 435 961 469
rect 927 367 961 401
rect 927 299 961 333
rect 927 231 961 265
rect 927 163 961 197
rect 1045 639 1079 673
rect 1045 571 1079 605
rect 1045 503 1079 537
rect 1045 435 1079 469
rect 1045 367 1079 401
rect 1045 299 1079 333
rect 1045 231 1079 265
rect 1045 163 1079 197
rect 1163 639 1197 673
rect 1163 571 1197 605
rect 1163 503 1197 537
rect 1163 435 1197 469
rect 1163 367 1197 401
rect 1163 299 1197 333
rect 1163 231 1197 265
rect 1163 163 1197 197
rect 1281 639 1315 673
rect 1281 571 1315 605
rect 1281 503 1315 537
rect 1281 435 1315 469
rect 1281 367 1315 401
rect 1281 299 1315 333
rect 1281 231 1315 265
rect 1281 163 1315 197
rect 1399 639 1433 673
rect 1399 571 1433 605
rect 1399 503 1433 537
rect 1399 435 1433 469
rect 1399 367 1433 401
rect 1399 299 1433 333
rect 1399 231 1433 265
rect 1399 163 1433 197
rect 1517 639 1551 673
rect 1517 571 1551 605
rect 1517 503 1551 537
rect 1517 435 1551 469
rect 1517 367 1551 401
rect 1517 299 1551 333
rect 1517 231 1551 265
rect 1517 163 1551 197
rect 1635 639 1669 673
rect 1635 571 1669 605
rect 1635 503 1669 537
rect 1635 435 1669 469
rect 1635 367 1669 401
rect 1635 299 1669 333
rect 1635 231 1669 265
rect 1635 163 1669 197
rect 1753 639 1787 673
rect 1753 571 1787 605
rect 1753 503 1787 537
rect 1753 435 1787 469
rect 1753 367 1787 401
rect 1753 299 1787 333
rect 1753 231 1787 265
rect 1753 163 1787 197
rect 1871 639 1905 673
rect 1871 571 1905 605
rect 1871 503 1905 537
rect 1871 435 1905 469
rect 1871 367 1905 401
rect 1871 299 1905 333
rect 1871 231 1905 265
rect 1871 163 1905 197
rect 1989 639 2023 673
rect 1989 571 2023 605
rect 1989 503 2023 537
rect 1989 435 2023 469
rect 1989 367 2023 401
rect 1989 299 2023 333
rect 1989 231 2023 265
rect 1989 163 2023 197
rect 2107 639 2141 673
rect 2107 571 2141 605
rect 2107 503 2141 537
rect 2107 435 2141 469
rect 2107 367 2141 401
rect 2107 299 2141 333
rect 2107 231 2141 265
rect 2107 163 2141 197
rect 2225 639 2259 673
rect 2225 571 2259 605
rect 2225 503 2259 537
rect 2225 435 2259 469
rect 2225 367 2259 401
rect 2225 299 2259 333
rect 2225 231 2259 265
rect 2225 163 2259 197
rect 2343 639 2377 673
rect 2343 571 2377 605
rect 2343 503 2377 537
rect 2343 435 2377 469
rect 2343 367 2377 401
rect 2343 299 2377 333
rect 2343 231 2377 265
rect 2343 163 2377 197
rect 2461 639 2495 673
rect 2461 571 2495 605
rect 2461 503 2495 537
rect 2461 435 2495 469
rect 2461 367 2495 401
rect 2461 299 2495 333
rect 2461 231 2495 265
rect 2461 163 2495 197
rect 2579 639 2613 673
rect 2579 571 2613 605
rect 2579 503 2613 537
rect 2579 435 2613 469
rect 2579 367 2613 401
rect 2579 299 2613 333
rect 2579 231 2613 265
rect 2579 163 2613 197
rect 2697 639 2731 673
rect 2697 571 2731 605
rect 2697 503 2731 537
rect 2697 435 2731 469
rect 2697 367 2731 401
rect 2697 299 2731 333
rect 2697 231 2731 265
rect 2697 163 2731 197
rect 2815 639 2849 673
rect 2815 571 2849 605
rect 2815 503 2849 537
rect 2815 435 2849 469
rect 2815 367 2849 401
rect 2815 299 2849 333
rect 2815 231 2849 265
rect 2815 163 2849 197
rect 2933 639 2967 673
rect 2933 571 2967 605
rect 2933 503 2967 537
rect 2933 435 2967 469
rect 2933 367 2967 401
rect 2933 299 2967 333
rect 2933 231 2967 265
rect 2933 163 2967 197
rect -2967 -197 -2933 -163
rect -2967 -265 -2933 -231
rect -2967 -333 -2933 -299
rect -2967 -401 -2933 -367
rect -2967 -469 -2933 -435
rect -2967 -537 -2933 -503
rect -2967 -605 -2933 -571
rect -2967 -673 -2933 -639
rect -2849 -197 -2815 -163
rect -2849 -265 -2815 -231
rect -2849 -333 -2815 -299
rect -2849 -401 -2815 -367
rect -2849 -469 -2815 -435
rect -2849 -537 -2815 -503
rect -2849 -605 -2815 -571
rect -2849 -673 -2815 -639
rect -2731 -197 -2697 -163
rect -2731 -265 -2697 -231
rect -2731 -333 -2697 -299
rect -2731 -401 -2697 -367
rect -2731 -469 -2697 -435
rect -2731 -537 -2697 -503
rect -2731 -605 -2697 -571
rect -2731 -673 -2697 -639
rect -2613 -197 -2579 -163
rect -2613 -265 -2579 -231
rect -2613 -333 -2579 -299
rect -2613 -401 -2579 -367
rect -2613 -469 -2579 -435
rect -2613 -537 -2579 -503
rect -2613 -605 -2579 -571
rect -2613 -673 -2579 -639
rect -2495 -197 -2461 -163
rect -2495 -265 -2461 -231
rect -2495 -333 -2461 -299
rect -2495 -401 -2461 -367
rect -2495 -469 -2461 -435
rect -2495 -537 -2461 -503
rect -2495 -605 -2461 -571
rect -2495 -673 -2461 -639
rect -2377 -197 -2343 -163
rect -2377 -265 -2343 -231
rect -2377 -333 -2343 -299
rect -2377 -401 -2343 -367
rect -2377 -469 -2343 -435
rect -2377 -537 -2343 -503
rect -2377 -605 -2343 -571
rect -2377 -673 -2343 -639
rect -2259 -197 -2225 -163
rect -2259 -265 -2225 -231
rect -2259 -333 -2225 -299
rect -2259 -401 -2225 -367
rect -2259 -469 -2225 -435
rect -2259 -537 -2225 -503
rect -2259 -605 -2225 -571
rect -2259 -673 -2225 -639
rect -2141 -197 -2107 -163
rect -2141 -265 -2107 -231
rect -2141 -333 -2107 -299
rect -2141 -401 -2107 -367
rect -2141 -469 -2107 -435
rect -2141 -537 -2107 -503
rect -2141 -605 -2107 -571
rect -2141 -673 -2107 -639
rect -2023 -197 -1989 -163
rect -2023 -265 -1989 -231
rect -2023 -333 -1989 -299
rect -2023 -401 -1989 -367
rect -2023 -469 -1989 -435
rect -2023 -537 -1989 -503
rect -2023 -605 -1989 -571
rect -2023 -673 -1989 -639
rect -1905 -197 -1871 -163
rect -1905 -265 -1871 -231
rect -1905 -333 -1871 -299
rect -1905 -401 -1871 -367
rect -1905 -469 -1871 -435
rect -1905 -537 -1871 -503
rect -1905 -605 -1871 -571
rect -1905 -673 -1871 -639
rect -1787 -197 -1753 -163
rect -1787 -265 -1753 -231
rect -1787 -333 -1753 -299
rect -1787 -401 -1753 -367
rect -1787 -469 -1753 -435
rect -1787 -537 -1753 -503
rect -1787 -605 -1753 -571
rect -1787 -673 -1753 -639
rect -1669 -197 -1635 -163
rect -1669 -265 -1635 -231
rect -1669 -333 -1635 -299
rect -1669 -401 -1635 -367
rect -1669 -469 -1635 -435
rect -1669 -537 -1635 -503
rect -1669 -605 -1635 -571
rect -1669 -673 -1635 -639
rect -1551 -197 -1517 -163
rect -1551 -265 -1517 -231
rect -1551 -333 -1517 -299
rect -1551 -401 -1517 -367
rect -1551 -469 -1517 -435
rect -1551 -537 -1517 -503
rect -1551 -605 -1517 -571
rect -1551 -673 -1517 -639
rect -1433 -197 -1399 -163
rect -1433 -265 -1399 -231
rect -1433 -333 -1399 -299
rect -1433 -401 -1399 -367
rect -1433 -469 -1399 -435
rect -1433 -537 -1399 -503
rect -1433 -605 -1399 -571
rect -1433 -673 -1399 -639
rect -1315 -197 -1281 -163
rect -1315 -265 -1281 -231
rect -1315 -333 -1281 -299
rect -1315 -401 -1281 -367
rect -1315 -469 -1281 -435
rect -1315 -537 -1281 -503
rect -1315 -605 -1281 -571
rect -1315 -673 -1281 -639
rect -1197 -197 -1163 -163
rect -1197 -265 -1163 -231
rect -1197 -333 -1163 -299
rect -1197 -401 -1163 -367
rect -1197 -469 -1163 -435
rect -1197 -537 -1163 -503
rect -1197 -605 -1163 -571
rect -1197 -673 -1163 -639
rect -1079 -197 -1045 -163
rect -1079 -265 -1045 -231
rect -1079 -333 -1045 -299
rect -1079 -401 -1045 -367
rect -1079 -469 -1045 -435
rect -1079 -537 -1045 -503
rect -1079 -605 -1045 -571
rect -1079 -673 -1045 -639
rect -961 -197 -927 -163
rect -961 -265 -927 -231
rect -961 -333 -927 -299
rect -961 -401 -927 -367
rect -961 -469 -927 -435
rect -961 -537 -927 -503
rect -961 -605 -927 -571
rect -961 -673 -927 -639
rect -843 -197 -809 -163
rect -843 -265 -809 -231
rect -843 -333 -809 -299
rect -843 -401 -809 -367
rect -843 -469 -809 -435
rect -843 -537 -809 -503
rect -843 -605 -809 -571
rect -843 -673 -809 -639
rect -725 -197 -691 -163
rect -725 -265 -691 -231
rect -725 -333 -691 -299
rect -725 -401 -691 -367
rect -725 -469 -691 -435
rect -725 -537 -691 -503
rect -725 -605 -691 -571
rect -725 -673 -691 -639
rect -607 -197 -573 -163
rect -607 -265 -573 -231
rect -607 -333 -573 -299
rect -607 -401 -573 -367
rect -607 -469 -573 -435
rect -607 -537 -573 -503
rect -607 -605 -573 -571
rect -607 -673 -573 -639
rect -489 -197 -455 -163
rect -489 -265 -455 -231
rect -489 -333 -455 -299
rect -489 -401 -455 -367
rect -489 -469 -455 -435
rect -489 -537 -455 -503
rect -489 -605 -455 -571
rect -489 -673 -455 -639
rect -371 -197 -337 -163
rect -371 -265 -337 -231
rect -371 -333 -337 -299
rect -371 -401 -337 -367
rect -371 -469 -337 -435
rect -371 -537 -337 -503
rect -371 -605 -337 -571
rect -371 -673 -337 -639
rect -253 -197 -219 -163
rect -253 -265 -219 -231
rect -253 -333 -219 -299
rect -253 -401 -219 -367
rect -253 -469 -219 -435
rect -253 -537 -219 -503
rect -253 -605 -219 -571
rect -253 -673 -219 -639
rect -135 -197 -101 -163
rect -135 -265 -101 -231
rect -135 -333 -101 -299
rect -135 -401 -101 -367
rect -135 -469 -101 -435
rect -135 -537 -101 -503
rect -135 -605 -101 -571
rect -135 -673 -101 -639
rect -17 -197 17 -163
rect -17 -265 17 -231
rect -17 -333 17 -299
rect -17 -401 17 -367
rect -17 -469 17 -435
rect -17 -537 17 -503
rect -17 -605 17 -571
rect -17 -673 17 -639
rect 101 -197 135 -163
rect 101 -265 135 -231
rect 101 -333 135 -299
rect 101 -401 135 -367
rect 101 -469 135 -435
rect 101 -537 135 -503
rect 101 -605 135 -571
rect 101 -673 135 -639
rect 219 -197 253 -163
rect 219 -265 253 -231
rect 219 -333 253 -299
rect 219 -401 253 -367
rect 219 -469 253 -435
rect 219 -537 253 -503
rect 219 -605 253 -571
rect 219 -673 253 -639
rect 337 -197 371 -163
rect 337 -265 371 -231
rect 337 -333 371 -299
rect 337 -401 371 -367
rect 337 -469 371 -435
rect 337 -537 371 -503
rect 337 -605 371 -571
rect 337 -673 371 -639
rect 455 -197 489 -163
rect 455 -265 489 -231
rect 455 -333 489 -299
rect 455 -401 489 -367
rect 455 -469 489 -435
rect 455 -537 489 -503
rect 455 -605 489 -571
rect 455 -673 489 -639
rect 573 -197 607 -163
rect 573 -265 607 -231
rect 573 -333 607 -299
rect 573 -401 607 -367
rect 573 -469 607 -435
rect 573 -537 607 -503
rect 573 -605 607 -571
rect 573 -673 607 -639
rect 691 -197 725 -163
rect 691 -265 725 -231
rect 691 -333 725 -299
rect 691 -401 725 -367
rect 691 -469 725 -435
rect 691 -537 725 -503
rect 691 -605 725 -571
rect 691 -673 725 -639
rect 809 -197 843 -163
rect 809 -265 843 -231
rect 809 -333 843 -299
rect 809 -401 843 -367
rect 809 -469 843 -435
rect 809 -537 843 -503
rect 809 -605 843 -571
rect 809 -673 843 -639
rect 927 -197 961 -163
rect 927 -265 961 -231
rect 927 -333 961 -299
rect 927 -401 961 -367
rect 927 -469 961 -435
rect 927 -537 961 -503
rect 927 -605 961 -571
rect 927 -673 961 -639
rect 1045 -197 1079 -163
rect 1045 -265 1079 -231
rect 1045 -333 1079 -299
rect 1045 -401 1079 -367
rect 1045 -469 1079 -435
rect 1045 -537 1079 -503
rect 1045 -605 1079 -571
rect 1045 -673 1079 -639
rect 1163 -197 1197 -163
rect 1163 -265 1197 -231
rect 1163 -333 1197 -299
rect 1163 -401 1197 -367
rect 1163 -469 1197 -435
rect 1163 -537 1197 -503
rect 1163 -605 1197 -571
rect 1163 -673 1197 -639
rect 1281 -197 1315 -163
rect 1281 -265 1315 -231
rect 1281 -333 1315 -299
rect 1281 -401 1315 -367
rect 1281 -469 1315 -435
rect 1281 -537 1315 -503
rect 1281 -605 1315 -571
rect 1281 -673 1315 -639
rect 1399 -197 1433 -163
rect 1399 -265 1433 -231
rect 1399 -333 1433 -299
rect 1399 -401 1433 -367
rect 1399 -469 1433 -435
rect 1399 -537 1433 -503
rect 1399 -605 1433 -571
rect 1399 -673 1433 -639
rect 1517 -197 1551 -163
rect 1517 -265 1551 -231
rect 1517 -333 1551 -299
rect 1517 -401 1551 -367
rect 1517 -469 1551 -435
rect 1517 -537 1551 -503
rect 1517 -605 1551 -571
rect 1517 -673 1551 -639
rect 1635 -197 1669 -163
rect 1635 -265 1669 -231
rect 1635 -333 1669 -299
rect 1635 -401 1669 -367
rect 1635 -469 1669 -435
rect 1635 -537 1669 -503
rect 1635 -605 1669 -571
rect 1635 -673 1669 -639
rect 1753 -197 1787 -163
rect 1753 -265 1787 -231
rect 1753 -333 1787 -299
rect 1753 -401 1787 -367
rect 1753 -469 1787 -435
rect 1753 -537 1787 -503
rect 1753 -605 1787 -571
rect 1753 -673 1787 -639
rect 1871 -197 1905 -163
rect 1871 -265 1905 -231
rect 1871 -333 1905 -299
rect 1871 -401 1905 -367
rect 1871 -469 1905 -435
rect 1871 -537 1905 -503
rect 1871 -605 1905 -571
rect 1871 -673 1905 -639
rect 1989 -197 2023 -163
rect 1989 -265 2023 -231
rect 1989 -333 2023 -299
rect 1989 -401 2023 -367
rect 1989 -469 2023 -435
rect 1989 -537 2023 -503
rect 1989 -605 2023 -571
rect 1989 -673 2023 -639
rect 2107 -197 2141 -163
rect 2107 -265 2141 -231
rect 2107 -333 2141 -299
rect 2107 -401 2141 -367
rect 2107 -469 2141 -435
rect 2107 -537 2141 -503
rect 2107 -605 2141 -571
rect 2107 -673 2141 -639
rect 2225 -197 2259 -163
rect 2225 -265 2259 -231
rect 2225 -333 2259 -299
rect 2225 -401 2259 -367
rect 2225 -469 2259 -435
rect 2225 -537 2259 -503
rect 2225 -605 2259 -571
rect 2225 -673 2259 -639
rect 2343 -197 2377 -163
rect 2343 -265 2377 -231
rect 2343 -333 2377 -299
rect 2343 -401 2377 -367
rect 2343 -469 2377 -435
rect 2343 -537 2377 -503
rect 2343 -605 2377 -571
rect 2343 -673 2377 -639
rect 2461 -197 2495 -163
rect 2461 -265 2495 -231
rect 2461 -333 2495 -299
rect 2461 -401 2495 -367
rect 2461 -469 2495 -435
rect 2461 -537 2495 -503
rect 2461 -605 2495 -571
rect 2461 -673 2495 -639
rect 2579 -197 2613 -163
rect 2579 -265 2613 -231
rect 2579 -333 2613 -299
rect 2579 -401 2613 -367
rect 2579 -469 2613 -435
rect 2579 -537 2613 -503
rect 2579 -605 2613 -571
rect 2579 -673 2613 -639
rect 2697 -197 2731 -163
rect 2697 -265 2731 -231
rect 2697 -333 2731 -299
rect 2697 -401 2731 -367
rect 2697 -469 2731 -435
rect 2697 -537 2731 -503
rect 2697 -605 2731 -571
rect 2697 -673 2731 -639
rect 2815 -197 2849 -163
rect 2815 -265 2849 -231
rect 2815 -333 2849 -299
rect 2815 -401 2849 -367
rect 2815 -469 2849 -435
rect 2815 -537 2849 -503
rect 2815 -605 2849 -571
rect 2815 -673 2849 -639
rect 2933 -197 2967 -163
rect 2933 -265 2967 -231
rect 2933 -333 2967 -299
rect 2933 -401 2967 -367
rect 2933 -469 2967 -435
rect 2933 -537 2967 -503
rect 2933 -605 2967 -571
rect 2933 -673 2967 -639
<< nsubdiff >>
rect -3081 867 -2975 901
rect -2941 867 -2907 901
rect -2873 867 -2839 901
rect -2805 867 -2771 901
rect -2737 867 -2703 901
rect -2669 867 -2635 901
rect -2601 867 -2567 901
rect -2533 867 -2499 901
rect -2465 867 -2431 901
rect -2397 867 -2363 901
rect -2329 867 -2295 901
rect -2261 867 -2227 901
rect -2193 867 -2159 901
rect -2125 867 -2091 901
rect -2057 867 -2023 901
rect -1989 867 -1955 901
rect -1921 867 -1887 901
rect -1853 867 -1819 901
rect -1785 867 -1751 901
rect -1717 867 -1683 901
rect -1649 867 -1615 901
rect -1581 867 -1547 901
rect -1513 867 -1479 901
rect -1445 867 -1411 901
rect -1377 867 -1343 901
rect -1309 867 -1275 901
rect -1241 867 -1207 901
rect -1173 867 -1139 901
rect -1105 867 -1071 901
rect -1037 867 -1003 901
rect -969 867 -935 901
rect -901 867 -867 901
rect -833 867 -799 901
rect -765 867 -731 901
rect -697 867 -663 901
rect -629 867 -595 901
rect -561 867 -527 901
rect -493 867 -459 901
rect -425 867 -391 901
rect -357 867 -323 901
rect -289 867 -255 901
rect -221 867 -187 901
rect -153 867 -119 901
rect -85 867 -51 901
rect -17 867 17 901
rect 51 867 85 901
rect 119 867 153 901
rect 187 867 221 901
rect 255 867 289 901
rect 323 867 357 901
rect 391 867 425 901
rect 459 867 493 901
rect 527 867 561 901
rect 595 867 629 901
rect 663 867 697 901
rect 731 867 765 901
rect 799 867 833 901
rect 867 867 901 901
rect 935 867 969 901
rect 1003 867 1037 901
rect 1071 867 1105 901
rect 1139 867 1173 901
rect 1207 867 1241 901
rect 1275 867 1309 901
rect 1343 867 1377 901
rect 1411 867 1445 901
rect 1479 867 1513 901
rect 1547 867 1581 901
rect 1615 867 1649 901
rect 1683 867 1717 901
rect 1751 867 1785 901
rect 1819 867 1853 901
rect 1887 867 1921 901
rect 1955 867 1989 901
rect 2023 867 2057 901
rect 2091 867 2125 901
rect 2159 867 2193 901
rect 2227 867 2261 901
rect 2295 867 2329 901
rect 2363 867 2397 901
rect 2431 867 2465 901
rect 2499 867 2533 901
rect 2567 867 2601 901
rect 2635 867 2669 901
rect 2703 867 2737 901
rect 2771 867 2805 901
rect 2839 867 2873 901
rect 2907 867 2941 901
rect 2975 867 3081 901
rect -3081 799 -3047 867
rect -3081 731 -3047 765
rect 3047 799 3081 867
rect 3047 731 3081 765
rect -3081 663 -3047 697
rect -3081 595 -3047 629
rect -3081 527 -3047 561
rect -3081 459 -3047 493
rect -3081 391 -3047 425
rect -3081 323 -3047 357
rect -3081 255 -3047 289
rect -3081 187 -3047 221
rect -3081 119 -3047 153
rect 3047 663 3081 697
rect 3047 595 3081 629
rect 3047 527 3081 561
rect 3047 459 3081 493
rect 3047 391 3081 425
rect 3047 323 3081 357
rect 3047 255 3081 289
rect 3047 187 3081 221
rect 3047 119 3081 153
rect -3081 51 -3047 85
rect 3047 51 3081 85
rect -3081 -17 -3047 17
rect 3047 -17 3081 17
rect -3081 -85 -3047 -51
rect 3047 -85 3081 -51
rect -3081 -153 -3047 -119
rect -3081 -221 -3047 -187
rect -3081 -289 -3047 -255
rect -3081 -357 -3047 -323
rect -3081 -425 -3047 -391
rect -3081 -493 -3047 -459
rect -3081 -561 -3047 -527
rect -3081 -629 -3047 -595
rect -3081 -697 -3047 -663
rect 3047 -153 3081 -119
rect 3047 -221 3081 -187
rect 3047 -289 3081 -255
rect 3047 -357 3081 -323
rect 3047 -425 3081 -391
rect 3047 -493 3081 -459
rect 3047 -561 3081 -527
rect 3047 -629 3081 -595
rect 3047 -697 3081 -663
rect -3081 -765 -3047 -731
rect -3081 -867 -3047 -799
rect 3047 -765 3081 -731
rect 3047 -867 3081 -799
rect -3081 -901 -2975 -867
rect -2941 -901 -2907 -867
rect -2873 -901 -2839 -867
rect -2805 -901 -2771 -867
rect -2737 -901 -2703 -867
rect -2669 -901 -2635 -867
rect -2601 -901 -2567 -867
rect -2533 -901 -2499 -867
rect -2465 -901 -2431 -867
rect -2397 -901 -2363 -867
rect -2329 -901 -2295 -867
rect -2261 -901 -2227 -867
rect -2193 -901 -2159 -867
rect -2125 -901 -2091 -867
rect -2057 -901 -2023 -867
rect -1989 -901 -1955 -867
rect -1921 -901 -1887 -867
rect -1853 -901 -1819 -867
rect -1785 -901 -1751 -867
rect -1717 -901 -1683 -867
rect -1649 -901 -1615 -867
rect -1581 -901 -1547 -867
rect -1513 -901 -1479 -867
rect -1445 -901 -1411 -867
rect -1377 -901 -1343 -867
rect -1309 -901 -1275 -867
rect -1241 -901 -1207 -867
rect -1173 -901 -1139 -867
rect -1105 -901 -1071 -867
rect -1037 -901 -1003 -867
rect -969 -901 -935 -867
rect -901 -901 -867 -867
rect -833 -901 -799 -867
rect -765 -901 -731 -867
rect -697 -901 -663 -867
rect -629 -901 -595 -867
rect -561 -901 -527 -867
rect -493 -901 -459 -867
rect -425 -901 -391 -867
rect -357 -901 -323 -867
rect -289 -901 -255 -867
rect -221 -901 -187 -867
rect -153 -901 -119 -867
rect -85 -901 -51 -867
rect -17 -901 17 -867
rect 51 -901 85 -867
rect 119 -901 153 -867
rect 187 -901 221 -867
rect 255 -901 289 -867
rect 323 -901 357 -867
rect 391 -901 425 -867
rect 459 -901 493 -867
rect 527 -901 561 -867
rect 595 -901 629 -867
rect 663 -901 697 -867
rect 731 -901 765 -867
rect 799 -901 833 -867
rect 867 -901 901 -867
rect 935 -901 969 -867
rect 1003 -901 1037 -867
rect 1071 -901 1105 -867
rect 1139 -901 1173 -867
rect 1207 -901 1241 -867
rect 1275 -901 1309 -867
rect 1343 -901 1377 -867
rect 1411 -901 1445 -867
rect 1479 -901 1513 -867
rect 1547 -901 1581 -867
rect 1615 -901 1649 -867
rect 1683 -901 1717 -867
rect 1751 -901 1785 -867
rect 1819 -901 1853 -867
rect 1887 -901 1921 -867
rect 1955 -901 1989 -867
rect 2023 -901 2057 -867
rect 2091 -901 2125 -867
rect 2159 -901 2193 -867
rect 2227 -901 2261 -867
rect 2295 -901 2329 -867
rect 2363 -901 2397 -867
rect 2431 -901 2465 -867
rect 2499 -901 2533 -867
rect 2567 -901 2601 -867
rect 2635 -901 2669 -867
rect 2703 -901 2737 -867
rect 2771 -901 2805 -867
rect 2839 -901 2873 -867
rect 2907 -901 2941 -867
rect 2975 -901 3081 -867
<< nsubdiffcont >>
rect -2975 867 -2941 901
rect -2907 867 -2873 901
rect -2839 867 -2805 901
rect -2771 867 -2737 901
rect -2703 867 -2669 901
rect -2635 867 -2601 901
rect -2567 867 -2533 901
rect -2499 867 -2465 901
rect -2431 867 -2397 901
rect -2363 867 -2329 901
rect -2295 867 -2261 901
rect -2227 867 -2193 901
rect -2159 867 -2125 901
rect -2091 867 -2057 901
rect -2023 867 -1989 901
rect -1955 867 -1921 901
rect -1887 867 -1853 901
rect -1819 867 -1785 901
rect -1751 867 -1717 901
rect -1683 867 -1649 901
rect -1615 867 -1581 901
rect -1547 867 -1513 901
rect -1479 867 -1445 901
rect -1411 867 -1377 901
rect -1343 867 -1309 901
rect -1275 867 -1241 901
rect -1207 867 -1173 901
rect -1139 867 -1105 901
rect -1071 867 -1037 901
rect -1003 867 -969 901
rect -935 867 -901 901
rect -867 867 -833 901
rect -799 867 -765 901
rect -731 867 -697 901
rect -663 867 -629 901
rect -595 867 -561 901
rect -527 867 -493 901
rect -459 867 -425 901
rect -391 867 -357 901
rect -323 867 -289 901
rect -255 867 -221 901
rect -187 867 -153 901
rect -119 867 -85 901
rect -51 867 -17 901
rect 17 867 51 901
rect 85 867 119 901
rect 153 867 187 901
rect 221 867 255 901
rect 289 867 323 901
rect 357 867 391 901
rect 425 867 459 901
rect 493 867 527 901
rect 561 867 595 901
rect 629 867 663 901
rect 697 867 731 901
rect 765 867 799 901
rect 833 867 867 901
rect 901 867 935 901
rect 969 867 1003 901
rect 1037 867 1071 901
rect 1105 867 1139 901
rect 1173 867 1207 901
rect 1241 867 1275 901
rect 1309 867 1343 901
rect 1377 867 1411 901
rect 1445 867 1479 901
rect 1513 867 1547 901
rect 1581 867 1615 901
rect 1649 867 1683 901
rect 1717 867 1751 901
rect 1785 867 1819 901
rect 1853 867 1887 901
rect 1921 867 1955 901
rect 1989 867 2023 901
rect 2057 867 2091 901
rect 2125 867 2159 901
rect 2193 867 2227 901
rect 2261 867 2295 901
rect 2329 867 2363 901
rect 2397 867 2431 901
rect 2465 867 2499 901
rect 2533 867 2567 901
rect 2601 867 2635 901
rect 2669 867 2703 901
rect 2737 867 2771 901
rect 2805 867 2839 901
rect 2873 867 2907 901
rect 2941 867 2975 901
rect -3081 765 -3047 799
rect 3047 765 3081 799
rect -3081 697 -3047 731
rect -3081 629 -3047 663
rect -3081 561 -3047 595
rect -3081 493 -3047 527
rect -3081 425 -3047 459
rect -3081 357 -3047 391
rect -3081 289 -3047 323
rect -3081 221 -3047 255
rect -3081 153 -3047 187
rect -3081 85 -3047 119
rect 3047 697 3081 731
rect 3047 629 3081 663
rect 3047 561 3081 595
rect 3047 493 3081 527
rect 3047 425 3081 459
rect 3047 357 3081 391
rect 3047 289 3081 323
rect 3047 221 3081 255
rect 3047 153 3081 187
rect -3081 17 -3047 51
rect 3047 85 3081 119
rect -3081 -51 -3047 -17
rect 3047 17 3081 51
rect -3081 -119 -3047 -85
rect 3047 -51 3081 -17
rect -3081 -187 -3047 -153
rect -3081 -255 -3047 -221
rect -3081 -323 -3047 -289
rect -3081 -391 -3047 -357
rect -3081 -459 -3047 -425
rect -3081 -527 -3047 -493
rect -3081 -595 -3047 -561
rect -3081 -663 -3047 -629
rect -3081 -731 -3047 -697
rect 3047 -119 3081 -85
rect 3047 -187 3081 -153
rect 3047 -255 3081 -221
rect 3047 -323 3081 -289
rect 3047 -391 3081 -357
rect 3047 -459 3081 -425
rect 3047 -527 3081 -493
rect 3047 -595 3081 -561
rect 3047 -663 3081 -629
rect 3047 -731 3081 -697
rect -3081 -799 -3047 -765
rect 3047 -799 3081 -765
rect -2975 -901 -2941 -867
rect -2907 -901 -2873 -867
rect -2839 -901 -2805 -867
rect -2771 -901 -2737 -867
rect -2703 -901 -2669 -867
rect -2635 -901 -2601 -867
rect -2567 -901 -2533 -867
rect -2499 -901 -2465 -867
rect -2431 -901 -2397 -867
rect -2363 -901 -2329 -867
rect -2295 -901 -2261 -867
rect -2227 -901 -2193 -867
rect -2159 -901 -2125 -867
rect -2091 -901 -2057 -867
rect -2023 -901 -1989 -867
rect -1955 -901 -1921 -867
rect -1887 -901 -1853 -867
rect -1819 -901 -1785 -867
rect -1751 -901 -1717 -867
rect -1683 -901 -1649 -867
rect -1615 -901 -1581 -867
rect -1547 -901 -1513 -867
rect -1479 -901 -1445 -867
rect -1411 -901 -1377 -867
rect -1343 -901 -1309 -867
rect -1275 -901 -1241 -867
rect -1207 -901 -1173 -867
rect -1139 -901 -1105 -867
rect -1071 -901 -1037 -867
rect -1003 -901 -969 -867
rect -935 -901 -901 -867
rect -867 -901 -833 -867
rect -799 -901 -765 -867
rect -731 -901 -697 -867
rect -663 -901 -629 -867
rect -595 -901 -561 -867
rect -527 -901 -493 -867
rect -459 -901 -425 -867
rect -391 -901 -357 -867
rect -323 -901 -289 -867
rect -255 -901 -221 -867
rect -187 -901 -153 -867
rect -119 -901 -85 -867
rect -51 -901 -17 -867
rect 17 -901 51 -867
rect 85 -901 119 -867
rect 153 -901 187 -867
rect 221 -901 255 -867
rect 289 -901 323 -867
rect 357 -901 391 -867
rect 425 -901 459 -867
rect 493 -901 527 -867
rect 561 -901 595 -867
rect 629 -901 663 -867
rect 697 -901 731 -867
rect 765 -901 799 -867
rect 833 -901 867 -867
rect 901 -901 935 -867
rect 969 -901 1003 -867
rect 1037 -901 1071 -867
rect 1105 -901 1139 -867
rect 1173 -901 1207 -867
rect 1241 -901 1275 -867
rect 1309 -901 1343 -867
rect 1377 -901 1411 -867
rect 1445 -901 1479 -867
rect 1513 -901 1547 -867
rect 1581 -901 1615 -867
rect 1649 -901 1683 -867
rect 1717 -901 1751 -867
rect 1785 -901 1819 -867
rect 1853 -901 1887 -867
rect 1921 -901 1955 -867
rect 1989 -901 2023 -867
rect 2057 -901 2091 -867
rect 2125 -901 2159 -867
rect 2193 -901 2227 -867
rect 2261 -901 2295 -867
rect 2329 -901 2363 -867
rect 2397 -901 2431 -867
rect 2465 -901 2499 -867
rect 2533 -901 2567 -867
rect 2601 -901 2635 -867
rect 2669 -901 2703 -867
rect 2737 -901 2771 -867
rect 2805 -901 2839 -867
rect 2873 -901 2907 -867
rect 2941 -901 2975 -867
<< poly >>
rect -2924 749 -2858 815
rect -2806 749 -2740 815
rect -2688 749 -2622 815
rect -2570 749 -2504 815
rect -2452 749 -2386 815
rect -2334 749 -2268 815
rect -2216 749 -2150 815
rect -2098 749 -2032 815
rect -1980 749 -1914 815
rect -1862 749 -1796 815
rect -1744 749 -1678 815
rect -1626 749 -1560 815
rect -1508 749 -1442 815
rect -1390 749 -1324 815
rect -1272 749 -1206 815
rect -1154 749 -1088 815
rect -1036 749 -970 815
rect -918 749 -852 815
rect -800 749 -734 815
rect -682 749 -616 815
rect -564 749 -498 815
rect -446 749 -380 815
rect -328 749 -262 815
rect -210 749 -144 815
rect -92 749 -26 815
rect 26 749 92 815
rect 144 749 210 815
rect 262 749 328 815
rect 380 749 446 815
rect 498 749 564 815
rect 616 749 682 815
rect 734 749 800 815
rect 852 749 918 815
rect 970 749 1036 815
rect 1088 749 1154 815
rect 1206 749 1272 815
rect 1324 749 1390 815
rect 1442 749 1508 815
rect 1560 749 1626 815
rect 1678 749 1744 815
rect 1796 749 1862 815
rect 1914 749 1980 815
rect 2032 749 2098 815
rect 2150 749 2216 815
rect 2268 749 2334 815
rect 2386 749 2452 815
rect 2504 749 2570 815
rect 2622 749 2688 815
rect 2740 749 2806 815
rect 2858 749 2924 815
rect -2921 718 -2861 749
rect -2803 718 -2743 749
rect -2685 718 -2625 749
rect -2567 718 -2507 749
rect -2449 718 -2389 749
rect -2331 718 -2271 749
rect -2213 718 -2153 749
rect -2095 718 -2035 749
rect -1977 718 -1917 749
rect -1859 718 -1799 749
rect -1741 718 -1681 749
rect -1623 718 -1563 749
rect -1505 718 -1445 749
rect -1387 718 -1327 749
rect -1269 718 -1209 749
rect -1151 718 -1091 749
rect -1033 718 -973 749
rect -915 718 -855 749
rect -797 718 -737 749
rect -679 718 -619 749
rect -561 718 -501 749
rect -443 718 -383 749
rect -325 718 -265 749
rect -207 718 -147 749
rect -89 718 -29 749
rect 29 718 89 749
rect 147 718 207 749
rect 265 718 325 749
rect 383 718 443 749
rect 501 718 561 749
rect 619 718 679 749
rect 737 718 797 749
rect 855 718 915 749
rect 973 718 1033 749
rect 1091 718 1151 749
rect 1209 718 1269 749
rect 1327 718 1387 749
rect 1445 718 1505 749
rect 1563 718 1623 749
rect 1681 718 1741 749
rect 1799 718 1859 749
rect 1917 718 1977 749
rect 2035 718 2095 749
rect 2153 718 2213 749
rect 2271 718 2331 749
rect 2389 718 2449 749
rect 2507 718 2567 749
rect 2625 718 2685 749
rect 2743 718 2803 749
rect 2861 718 2921 749
rect -2921 87 -2861 118
rect -2803 87 -2743 118
rect -2685 87 -2625 118
rect -2567 87 -2507 118
rect -2449 87 -2389 118
rect -2331 87 -2271 118
rect -2213 87 -2153 118
rect -2095 87 -2035 118
rect -1977 87 -1917 118
rect -1859 87 -1799 118
rect -1741 87 -1681 118
rect -1623 87 -1563 118
rect -1505 87 -1445 118
rect -1387 87 -1327 118
rect -1269 87 -1209 118
rect -1151 87 -1091 118
rect -1033 87 -973 118
rect -915 87 -855 118
rect -797 87 -737 118
rect -679 87 -619 118
rect -561 87 -501 118
rect -443 87 -383 118
rect -325 87 -265 118
rect -207 87 -147 118
rect -89 87 -29 118
rect 29 87 89 118
rect 147 87 207 118
rect 265 87 325 118
rect 383 87 443 118
rect 501 87 561 118
rect 619 87 679 118
rect 737 87 797 118
rect 855 87 915 118
rect 973 87 1033 118
rect 1091 87 1151 118
rect 1209 87 1269 118
rect 1327 87 1387 118
rect 1445 87 1505 118
rect 1563 87 1623 118
rect 1681 87 1741 118
rect 1799 87 1859 118
rect 1917 87 1977 118
rect 2035 87 2095 118
rect 2153 87 2213 118
rect 2271 87 2331 118
rect 2389 87 2449 118
rect 2507 87 2567 118
rect 2625 87 2685 118
rect 2743 87 2803 118
rect 2861 87 2921 118
rect -2924 71 -2858 87
rect -2924 37 -2908 71
rect -2874 37 -2858 71
rect -2924 21 -2858 37
rect -2806 71 -2740 87
rect -2806 37 -2790 71
rect -2756 37 -2740 71
rect -2806 21 -2740 37
rect -2688 71 -2622 87
rect -2688 37 -2672 71
rect -2638 37 -2622 71
rect -2688 21 -2622 37
rect -2570 71 -2504 87
rect -2570 37 -2554 71
rect -2520 37 -2504 71
rect -2570 21 -2504 37
rect -2452 71 -2386 87
rect -2452 37 -2436 71
rect -2402 37 -2386 71
rect -2452 21 -2386 37
rect -2334 71 -2268 87
rect -2334 37 -2318 71
rect -2284 37 -2268 71
rect -2334 21 -2268 37
rect -2216 71 -2150 87
rect -2216 37 -2200 71
rect -2166 37 -2150 71
rect -2216 21 -2150 37
rect -2098 71 -2032 87
rect -2098 37 -2082 71
rect -2048 37 -2032 71
rect -2098 21 -2032 37
rect -1980 71 -1914 87
rect -1980 37 -1964 71
rect -1930 37 -1914 71
rect -1980 21 -1914 37
rect -1862 71 -1796 87
rect -1862 37 -1846 71
rect -1812 37 -1796 71
rect -1862 21 -1796 37
rect -1744 71 -1678 87
rect -1744 37 -1728 71
rect -1694 37 -1678 71
rect -1744 21 -1678 37
rect -1626 71 -1560 87
rect -1626 37 -1610 71
rect -1576 37 -1560 71
rect -1626 21 -1560 37
rect -1508 71 -1442 87
rect -1508 37 -1492 71
rect -1458 37 -1442 71
rect -1508 21 -1442 37
rect -1390 71 -1324 87
rect -1390 37 -1374 71
rect -1340 37 -1324 71
rect -1390 21 -1324 37
rect -1272 71 -1206 87
rect -1272 37 -1256 71
rect -1222 37 -1206 71
rect -1272 21 -1206 37
rect -1154 71 -1088 87
rect -1154 37 -1138 71
rect -1104 37 -1088 71
rect -1154 21 -1088 37
rect -1036 71 -970 87
rect -1036 37 -1020 71
rect -986 37 -970 71
rect -1036 21 -970 37
rect -918 71 -852 87
rect -918 37 -902 71
rect -868 37 -852 71
rect -918 21 -852 37
rect -800 71 -734 87
rect -800 37 -784 71
rect -750 37 -734 71
rect -800 21 -734 37
rect -682 71 -616 87
rect -682 37 -666 71
rect -632 37 -616 71
rect -682 21 -616 37
rect -564 71 -498 87
rect -564 37 -548 71
rect -514 37 -498 71
rect -564 21 -498 37
rect -446 71 -380 87
rect -446 37 -430 71
rect -396 37 -380 71
rect -446 21 -380 37
rect -328 71 -262 87
rect -328 37 -312 71
rect -278 37 -262 71
rect -328 21 -262 37
rect -210 71 -144 87
rect -210 37 -194 71
rect -160 37 -144 71
rect -210 21 -144 37
rect -92 71 -26 87
rect -92 37 -76 71
rect -42 37 -26 71
rect -92 21 -26 37
rect 26 71 92 87
rect 26 37 42 71
rect 76 37 92 71
rect 26 21 92 37
rect 144 71 210 87
rect 144 37 160 71
rect 194 37 210 71
rect 144 21 210 37
rect 262 71 328 87
rect 262 37 278 71
rect 312 37 328 71
rect 262 21 328 37
rect 380 71 446 87
rect 380 37 396 71
rect 430 37 446 71
rect 380 21 446 37
rect 498 71 564 87
rect 498 37 514 71
rect 548 37 564 71
rect 498 21 564 37
rect 616 71 682 87
rect 616 37 632 71
rect 666 37 682 71
rect 616 21 682 37
rect 734 71 800 87
rect 734 37 750 71
rect 784 37 800 71
rect 734 21 800 37
rect 852 71 918 87
rect 852 37 868 71
rect 902 37 918 71
rect 852 21 918 37
rect 970 71 1036 87
rect 970 37 986 71
rect 1020 37 1036 71
rect 970 21 1036 37
rect 1088 71 1154 87
rect 1088 37 1104 71
rect 1138 37 1154 71
rect 1088 21 1154 37
rect 1206 71 1272 87
rect 1206 37 1222 71
rect 1256 37 1272 71
rect 1206 21 1272 37
rect 1324 71 1390 87
rect 1324 37 1340 71
rect 1374 37 1390 71
rect 1324 21 1390 37
rect 1442 71 1508 87
rect 1442 37 1458 71
rect 1492 37 1508 71
rect 1442 21 1508 37
rect 1560 71 1626 87
rect 1560 37 1576 71
rect 1610 37 1626 71
rect 1560 21 1626 37
rect 1678 71 1744 87
rect 1678 37 1694 71
rect 1728 37 1744 71
rect 1678 21 1744 37
rect 1796 71 1862 87
rect 1796 37 1812 71
rect 1846 37 1862 71
rect 1796 21 1862 37
rect 1914 71 1980 87
rect 1914 37 1930 71
rect 1964 37 1980 71
rect 1914 21 1980 37
rect 2032 71 2098 87
rect 2032 37 2048 71
rect 2082 37 2098 71
rect 2032 21 2098 37
rect 2150 71 2216 87
rect 2150 37 2166 71
rect 2200 37 2216 71
rect 2150 21 2216 37
rect 2268 71 2334 87
rect 2268 37 2284 71
rect 2318 37 2334 71
rect 2268 21 2334 37
rect 2386 71 2452 87
rect 2386 37 2402 71
rect 2436 37 2452 71
rect 2386 21 2452 37
rect 2504 71 2570 87
rect 2504 37 2520 71
rect 2554 37 2570 71
rect 2504 21 2570 37
rect 2622 71 2688 87
rect 2622 37 2638 71
rect 2672 37 2688 71
rect 2622 21 2688 37
rect 2740 71 2806 87
rect 2740 37 2756 71
rect 2790 37 2806 71
rect 2740 21 2806 37
rect 2858 71 2924 87
rect 2858 37 2874 71
rect 2908 37 2924 71
rect 2858 21 2924 37
rect -2924 -37 -2858 -21
rect -2924 -71 -2908 -37
rect -2874 -71 -2858 -37
rect -2924 -87 -2858 -71
rect -2806 -37 -2740 -21
rect -2806 -71 -2790 -37
rect -2756 -71 -2740 -37
rect -2806 -87 -2740 -71
rect -2688 -37 -2622 -21
rect -2688 -71 -2672 -37
rect -2638 -71 -2622 -37
rect -2688 -87 -2622 -71
rect -2570 -37 -2504 -21
rect -2570 -71 -2554 -37
rect -2520 -71 -2504 -37
rect -2570 -87 -2504 -71
rect -2452 -37 -2386 -21
rect -2452 -71 -2436 -37
rect -2402 -71 -2386 -37
rect -2452 -87 -2386 -71
rect -2334 -37 -2268 -21
rect -2334 -71 -2318 -37
rect -2284 -71 -2268 -37
rect -2334 -87 -2268 -71
rect -2216 -37 -2150 -21
rect -2216 -71 -2200 -37
rect -2166 -71 -2150 -37
rect -2216 -87 -2150 -71
rect -2098 -37 -2032 -21
rect -2098 -71 -2082 -37
rect -2048 -71 -2032 -37
rect -2098 -87 -2032 -71
rect -1980 -37 -1914 -21
rect -1980 -71 -1964 -37
rect -1930 -71 -1914 -37
rect -1980 -87 -1914 -71
rect -1862 -37 -1796 -21
rect -1862 -71 -1846 -37
rect -1812 -71 -1796 -37
rect -1862 -87 -1796 -71
rect -1744 -37 -1678 -21
rect -1744 -71 -1728 -37
rect -1694 -71 -1678 -37
rect -1744 -87 -1678 -71
rect -1626 -37 -1560 -21
rect -1626 -71 -1610 -37
rect -1576 -71 -1560 -37
rect -1626 -87 -1560 -71
rect -1508 -37 -1442 -21
rect -1508 -71 -1492 -37
rect -1458 -71 -1442 -37
rect -1508 -87 -1442 -71
rect -1390 -37 -1324 -21
rect -1390 -71 -1374 -37
rect -1340 -71 -1324 -37
rect -1390 -87 -1324 -71
rect -1272 -37 -1206 -21
rect -1272 -71 -1256 -37
rect -1222 -71 -1206 -37
rect -1272 -87 -1206 -71
rect -1154 -37 -1088 -21
rect -1154 -71 -1138 -37
rect -1104 -71 -1088 -37
rect -1154 -87 -1088 -71
rect -1036 -37 -970 -21
rect -1036 -71 -1020 -37
rect -986 -71 -970 -37
rect -1036 -87 -970 -71
rect -918 -37 -852 -21
rect -918 -71 -902 -37
rect -868 -71 -852 -37
rect -918 -87 -852 -71
rect -800 -37 -734 -21
rect -800 -71 -784 -37
rect -750 -71 -734 -37
rect -800 -87 -734 -71
rect -682 -37 -616 -21
rect -682 -71 -666 -37
rect -632 -71 -616 -37
rect -682 -87 -616 -71
rect -564 -37 -498 -21
rect -564 -71 -548 -37
rect -514 -71 -498 -37
rect -564 -87 -498 -71
rect -446 -37 -380 -21
rect -446 -71 -430 -37
rect -396 -71 -380 -37
rect -446 -87 -380 -71
rect -328 -37 -262 -21
rect -328 -71 -312 -37
rect -278 -71 -262 -37
rect -328 -87 -262 -71
rect -210 -37 -144 -21
rect -210 -71 -194 -37
rect -160 -71 -144 -37
rect -210 -87 -144 -71
rect -92 -37 -26 -21
rect -92 -71 -76 -37
rect -42 -71 -26 -37
rect -92 -87 -26 -71
rect 26 -37 92 -21
rect 26 -71 42 -37
rect 76 -71 92 -37
rect 26 -87 92 -71
rect 144 -37 210 -21
rect 144 -71 160 -37
rect 194 -71 210 -37
rect 144 -87 210 -71
rect 262 -37 328 -21
rect 262 -71 278 -37
rect 312 -71 328 -37
rect 262 -87 328 -71
rect 380 -37 446 -21
rect 380 -71 396 -37
rect 430 -71 446 -37
rect 380 -87 446 -71
rect 498 -37 564 -21
rect 498 -71 514 -37
rect 548 -71 564 -37
rect 498 -87 564 -71
rect 616 -37 682 -21
rect 616 -71 632 -37
rect 666 -71 682 -37
rect 616 -87 682 -71
rect 734 -37 800 -21
rect 734 -71 750 -37
rect 784 -71 800 -37
rect 734 -87 800 -71
rect 852 -37 918 -21
rect 852 -71 868 -37
rect 902 -71 918 -37
rect 852 -87 918 -71
rect 970 -37 1036 -21
rect 970 -71 986 -37
rect 1020 -71 1036 -37
rect 970 -87 1036 -71
rect 1088 -37 1154 -21
rect 1088 -71 1104 -37
rect 1138 -71 1154 -37
rect 1088 -87 1154 -71
rect 1206 -37 1272 -21
rect 1206 -71 1222 -37
rect 1256 -71 1272 -37
rect 1206 -87 1272 -71
rect 1324 -37 1390 -21
rect 1324 -71 1340 -37
rect 1374 -71 1390 -37
rect 1324 -87 1390 -71
rect 1442 -37 1508 -21
rect 1442 -71 1458 -37
rect 1492 -71 1508 -37
rect 1442 -87 1508 -71
rect 1560 -37 1626 -21
rect 1560 -71 1576 -37
rect 1610 -71 1626 -37
rect 1560 -87 1626 -71
rect 1678 -37 1744 -21
rect 1678 -71 1694 -37
rect 1728 -71 1744 -37
rect 1678 -87 1744 -71
rect 1796 -37 1862 -21
rect 1796 -71 1812 -37
rect 1846 -71 1862 -37
rect 1796 -87 1862 -71
rect 1914 -37 1980 -21
rect 1914 -71 1930 -37
rect 1964 -71 1980 -37
rect 1914 -87 1980 -71
rect 2032 -37 2098 -21
rect 2032 -71 2048 -37
rect 2082 -71 2098 -37
rect 2032 -87 2098 -71
rect 2150 -37 2216 -21
rect 2150 -71 2166 -37
rect 2200 -71 2216 -37
rect 2150 -87 2216 -71
rect 2268 -37 2334 -21
rect 2268 -71 2284 -37
rect 2318 -71 2334 -37
rect 2268 -87 2334 -71
rect 2386 -37 2452 -21
rect 2386 -71 2402 -37
rect 2436 -71 2452 -37
rect 2386 -87 2452 -71
rect 2504 -37 2570 -21
rect 2504 -71 2520 -37
rect 2554 -71 2570 -37
rect 2504 -87 2570 -71
rect 2622 -37 2688 -21
rect 2622 -71 2638 -37
rect 2672 -71 2688 -37
rect 2622 -87 2688 -71
rect 2740 -37 2806 -21
rect 2740 -71 2756 -37
rect 2790 -71 2806 -37
rect 2740 -87 2806 -71
rect 2858 -37 2924 -21
rect 2858 -71 2874 -37
rect 2908 -71 2924 -37
rect 2858 -87 2924 -71
rect -2921 -118 -2861 -87
rect -2803 -118 -2743 -87
rect -2685 -118 -2625 -87
rect -2567 -118 -2507 -87
rect -2449 -118 -2389 -87
rect -2331 -118 -2271 -87
rect -2213 -118 -2153 -87
rect -2095 -118 -2035 -87
rect -1977 -118 -1917 -87
rect -1859 -118 -1799 -87
rect -1741 -118 -1681 -87
rect -1623 -118 -1563 -87
rect -1505 -118 -1445 -87
rect -1387 -118 -1327 -87
rect -1269 -118 -1209 -87
rect -1151 -118 -1091 -87
rect -1033 -118 -973 -87
rect -915 -118 -855 -87
rect -797 -118 -737 -87
rect -679 -118 -619 -87
rect -561 -118 -501 -87
rect -443 -118 -383 -87
rect -325 -118 -265 -87
rect -207 -118 -147 -87
rect -89 -118 -29 -87
rect 29 -118 89 -87
rect 147 -118 207 -87
rect 265 -118 325 -87
rect 383 -118 443 -87
rect 501 -118 561 -87
rect 619 -118 679 -87
rect 737 -118 797 -87
rect 855 -118 915 -87
rect 973 -118 1033 -87
rect 1091 -118 1151 -87
rect 1209 -118 1269 -87
rect 1327 -118 1387 -87
rect 1445 -118 1505 -87
rect 1563 -118 1623 -87
rect 1681 -118 1741 -87
rect 1799 -118 1859 -87
rect 1917 -118 1977 -87
rect 2035 -118 2095 -87
rect 2153 -118 2213 -87
rect 2271 -118 2331 -87
rect 2389 -118 2449 -87
rect 2507 -118 2567 -87
rect 2625 -118 2685 -87
rect 2743 -118 2803 -87
rect 2861 -118 2921 -87
rect -2921 -749 -2861 -718
rect -2803 -749 -2743 -718
rect -2685 -749 -2625 -718
rect -2567 -749 -2507 -718
rect -2449 -749 -2389 -718
rect -2331 -749 -2271 -718
rect -2213 -749 -2153 -718
rect -2095 -749 -2035 -718
rect -1977 -749 -1917 -718
rect -1859 -749 -1799 -718
rect -1741 -749 -1681 -718
rect -1623 -749 -1563 -718
rect -1505 -749 -1445 -718
rect -1387 -749 -1327 -718
rect -1269 -749 -1209 -718
rect -1151 -749 -1091 -718
rect -1033 -749 -973 -718
rect -915 -749 -855 -718
rect -797 -749 -737 -718
rect -679 -749 -619 -718
rect -561 -749 -501 -718
rect -443 -749 -383 -718
rect -325 -749 -265 -718
rect -207 -749 -147 -718
rect -89 -749 -29 -718
rect 29 -749 89 -718
rect 147 -749 207 -718
rect 265 -749 325 -718
rect 383 -749 443 -718
rect 501 -749 561 -718
rect 619 -749 679 -718
rect 737 -749 797 -718
rect 855 -749 915 -718
rect 973 -749 1033 -718
rect 1091 -749 1151 -718
rect 1209 -749 1269 -718
rect 1327 -749 1387 -718
rect 1445 -749 1505 -718
rect 1563 -749 1623 -718
rect 1681 -749 1741 -718
rect 1799 -749 1859 -718
rect 1917 -749 1977 -718
rect 2035 -749 2095 -718
rect 2153 -749 2213 -718
rect 2271 -749 2331 -718
rect 2389 -749 2449 -718
rect 2507 -749 2567 -718
rect 2625 -749 2685 -718
rect 2743 -749 2803 -718
rect 2861 -749 2921 -718
rect -2924 -815 -2858 -749
rect -2806 -815 -2740 -749
rect -2688 -815 -2622 -749
rect -2570 -815 -2504 -749
rect -2452 -815 -2386 -749
rect -2334 -815 -2268 -749
rect -2216 -815 -2150 -749
rect -2098 -815 -2032 -749
rect -1980 -815 -1914 -749
rect -1862 -815 -1796 -749
rect -1744 -815 -1678 -749
rect -1626 -815 -1560 -749
rect -1508 -815 -1442 -749
rect -1390 -815 -1324 -749
rect -1272 -815 -1206 -749
rect -1154 -815 -1088 -749
rect -1036 -815 -970 -749
rect -918 -815 -852 -749
rect -800 -815 -734 -749
rect -682 -815 -616 -749
rect -564 -815 -498 -749
rect -446 -815 -380 -749
rect -328 -815 -262 -749
rect -210 -815 -144 -749
rect -92 -815 -26 -749
rect 26 -815 92 -749
rect 144 -815 210 -749
rect 262 -815 328 -749
rect 380 -815 446 -749
rect 498 -815 564 -749
rect 616 -815 682 -749
rect 734 -815 800 -749
rect 852 -815 918 -749
rect 970 -815 1036 -749
rect 1088 -815 1154 -749
rect 1206 -815 1272 -749
rect 1324 -815 1390 -749
rect 1442 -815 1508 -749
rect 1560 -815 1626 -749
rect 1678 -815 1744 -749
rect 1796 -815 1862 -749
rect 1914 -815 1980 -749
rect 2032 -815 2098 -749
rect 2150 -815 2216 -749
rect 2268 -815 2334 -749
rect 2386 -815 2452 -749
rect 2504 -815 2570 -749
rect 2622 -815 2688 -749
rect 2740 -815 2806 -749
rect 2858 -815 2924 -749
<< polycont >>
rect -2908 37 -2874 71
rect -2790 37 -2756 71
rect -2672 37 -2638 71
rect -2554 37 -2520 71
rect -2436 37 -2402 71
rect -2318 37 -2284 71
rect -2200 37 -2166 71
rect -2082 37 -2048 71
rect -1964 37 -1930 71
rect -1846 37 -1812 71
rect -1728 37 -1694 71
rect -1610 37 -1576 71
rect -1492 37 -1458 71
rect -1374 37 -1340 71
rect -1256 37 -1222 71
rect -1138 37 -1104 71
rect -1020 37 -986 71
rect -902 37 -868 71
rect -784 37 -750 71
rect -666 37 -632 71
rect -548 37 -514 71
rect -430 37 -396 71
rect -312 37 -278 71
rect -194 37 -160 71
rect -76 37 -42 71
rect 42 37 76 71
rect 160 37 194 71
rect 278 37 312 71
rect 396 37 430 71
rect 514 37 548 71
rect 632 37 666 71
rect 750 37 784 71
rect 868 37 902 71
rect 986 37 1020 71
rect 1104 37 1138 71
rect 1222 37 1256 71
rect 1340 37 1374 71
rect 1458 37 1492 71
rect 1576 37 1610 71
rect 1694 37 1728 71
rect 1812 37 1846 71
rect 1930 37 1964 71
rect 2048 37 2082 71
rect 2166 37 2200 71
rect 2284 37 2318 71
rect 2402 37 2436 71
rect 2520 37 2554 71
rect 2638 37 2672 71
rect 2756 37 2790 71
rect 2874 37 2908 71
rect -2908 -71 -2874 -37
rect -2790 -71 -2756 -37
rect -2672 -71 -2638 -37
rect -2554 -71 -2520 -37
rect -2436 -71 -2402 -37
rect -2318 -71 -2284 -37
rect -2200 -71 -2166 -37
rect -2082 -71 -2048 -37
rect -1964 -71 -1930 -37
rect -1846 -71 -1812 -37
rect -1728 -71 -1694 -37
rect -1610 -71 -1576 -37
rect -1492 -71 -1458 -37
rect -1374 -71 -1340 -37
rect -1256 -71 -1222 -37
rect -1138 -71 -1104 -37
rect -1020 -71 -986 -37
rect -902 -71 -868 -37
rect -784 -71 -750 -37
rect -666 -71 -632 -37
rect -548 -71 -514 -37
rect -430 -71 -396 -37
rect -312 -71 -278 -37
rect -194 -71 -160 -37
rect -76 -71 -42 -37
rect 42 -71 76 -37
rect 160 -71 194 -37
rect 278 -71 312 -37
rect 396 -71 430 -37
rect 514 -71 548 -37
rect 632 -71 666 -37
rect 750 -71 784 -37
rect 868 -71 902 -37
rect 986 -71 1020 -37
rect 1104 -71 1138 -37
rect 1222 -71 1256 -37
rect 1340 -71 1374 -37
rect 1458 -71 1492 -37
rect 1576 -71 1610 -37
rect 1694 -71 1728 -37
rect 1812 -71 1846 -37
rect 1930 -71 1964 -37
rect 2048 -71 2082 -37
rect 2166 -71 2200 -37
rect 2284 -71 2318 -37
rect 2402 -71 2436 -37
rect 2520 -71 2554 -37
rect 2638 -71 2672 -37
rect 2756 -71 2790 -37
rect 2874 -71 2908 -37
<< locali >>
rect -3081 867 -2975 901
rect -2941 867 -2907 901
rect -2873 867 -2839 901
rect -2805 867 -2771 901
rect -2737 867 -2703 901
rect -2669 867 -2635 901
rect -2601 867 -2567 901
rect -2533 867 -2499 901
rect -2465 867 -2431 901
rect -2397 867 -2363 901
rect -2329 867 -2295 901
rect -2261 867 -2227 901
rect -2193 867 -2159 901
rect -2125 867 -2091 901
rect -2057 867 -2023 901
rect -1989 867 -1955 901
rect -1921 867 -1887 901
rect -1853 867 -1819 901
rect -1785 867 -1751 901
rect -1717 867 -1683 901
rect -1649 867 -1615 901
rect -1581 867 -1547 901
rect -1513 867 -1479 901
rect -1445 867 -1411 901
rect -1377 867 -1343 901
rect -1309 867 -1275 901
rect -1241 867 -1207 901
rect -1173 867 -1139 901
rect -1105 867 -1071 901
rect -1037 867 -1003 901
rect -969 867 -935 901
rect -901 867 -867 901
rect -833 867 -799 901
rect -765 867 -731 901
rect -697 867 -663 901
rect -629 867 -595 901
rect -561 867 -527 901
rect -493 867 -459 901
rect -425 867 -391 901
rect -357 867 -323 901
rect -289 867 -255 901
rect -221 867 -187 901
rect -153 867 -119 901
rect -85 867 -51 901
rect -17 867 17 901
rect 51 867 85 901
rect 119 867 153 901
rect 187 867 221 901
rect 255 867 289 901
rect 323 867 357 901
rect 391 867 425 901
rect 459 867 493 901
rect 527 867 561 901
rect 595 867 629 901
rect 663 867 697 901
rect 731 867 765 901
rect 799 867 833 901
rect 867 867 901 901
rect 935 867 969 901
rect 1003 867 1037 901
rect 1071 867 1105 901
rect 1139 867 1173 901
rect 1207 867 1241 901
rect 1275 867 1309 901
rect 1343 867 1377 901
rect 1411 867 1445 901
rect 1479 867 1513 901
rect 1547 867 1581 901
rect 1615 867 1649 901
rect 1683 867 1717 901
rect 1751 867 1785 901
rect 1819 867 1853 901
rect 1887 867 1921 901
rect 1955 867 1989 901
rect 2023 867 2057 901
rect 2091 867 2125 901
rect 2159 867 2193 901
rect 2227 867 2261 901
rect 2295 867 2329 901
rect 2363 867 2397 901
rect 2431 867 2465 901
rect 2499 867 2533 901
rect 2567 867 2601 901
rect 2635 867 2669 901
rect 2703 867 2737 901
rect 2771 867 2805 901
rect 2839 867 2873 901
rect 2907 867 2941 901
rect 2975 867 3081 901
rect -3081 799 -3047 867
rect -3081 731 -3047 765
rect 3047 799 3081 867
rect 3047 731 3081 765
rect -3081 663 -3047 697
rect -3081 595 -3047 629
rect -3081 527 -3047 561
rect -3081 459 -3047 493
rect -3081 391 -3047 425
rect -3081 323 -3047 357
rect -3081 255 -3047 289
rect -3081 187 -3047 221
rect -3081 119 -3047 153
rect -2967 687 -2933 722
rect -2967 615 -2933 639
rect -2967 543 -2933 571
rect -2967 471 -2933 503
rect -2967 401 -2933 435
rect -2967 333 -2933 365
rect -2967 265 -2933 293
rect -2967 197 -2933 221
rect -2967 114 -2933 149
rect -2849 687 -2815 722
rect -2849 615 -2815 639
rect -2849 543 -2815 571
rect -2849 471 -2815 503
rect -2849 401 -2815 435
rect -2849 333 -2815 365
rect -2849 265 -2815 293
rect -2849 197 -2815 221
rect -2849 114 -2815 149
rect -2731 687 -2697 722
rect -2731 615 -2697 639
rect -2731 543 -2697 571
rect -2731 471 -2697 503
rect -2731 401 -2697 435
rect -2731 333 -2697 365
rect -2731 265 -2697 293
rect -2731 197 -2697 221
rect -2731 114 -2697 149
rect -2613 687 -2579 722
rect -2613 615 -2579 639
rect -2613 543 -2579 571
rect -2613 471 -2579 503
rect -2613 401 -2579 435
rect -2613 333 -2579 365
rect -2613 265 -2579 293
rect -2613 197 -2579 221
rect -2613 114 -2579 149
rect -2495 687 -2461 722
rect -2495 615 -2461 639
rect -2495 543 -2461 571
rect -2495 471 -2461 503
rect -2495 401 -2461 435
rect -2495 333 -2461 365
rect -2495 265 -2461 293
rect -2495 197 -2461 221
rect -2495 114 -2461 149
rect -2377 687 -2343 722
rect -2377 615 -2343 639
rect -2377 543 -2343 571
rect -2377 471 -2343 503
rect -2377 401 -2343 435
rect -2377 333 -2343 365
rect -2377 265 -2343 293
rect -2377 197 -2343 221
rect -2377 114 -2343 149
rect -2259 687 -2225 722
rect -2259 615 -2225 639
rect -2259 543 -2225 571
rect -2259 471 -2225 503
rect -2259 401 -2225 435
rect -2259 333 -2225 365
rect -2259 265 -2225 293
rect -2259 197 -2225 221
rect -2259 114 -2225 149
rect -2141 687 -2107 722
rect -2141 615 -2107 639
rect -2141 543 -2107 571
rect -2141 471 -2107 503
rect -2141 401 -2107 435
rect -2141 333 -2107 365
rect -2141 265 -2107 293
rect -2141 197 -2107 221
rect -2141 114 -2107 149
rect -2023 687 -1989 722
rect -2023 615 -1989 639
rect -2023 543 -1989 571
rect -2023 471 -1989 503
rect -2023 401 -1989 435
rect -2023 333 -1989 365
rect -2023 265 -1989 293
rect -2023 197 -1989 221
rect -2023 114 -1989 149
rect -1905 687 -1871 722
rect -1905 615 -1871 639
rect -1905 543 -1871 571
rect -1905 471 -1871 503
rect -1905 401 -1871 435
rect -1905 333 -1871 365
rect -1905 265 -1871 293
rect -1905 197 -1871 221
rect -1905 114 -1871 149
rect -1787 687 -1753 722
rect -1787 615 -1753 639
rect -1787 543 -1753 571
rect -1787 471 -1753 503
rect -1787 401 -1753 435
rect -1787 333 -1753 365
rect -1787 265 -1753 293
rect -1787 197 -1753 221
rect -1787 114 -1753 149
rect -1669 687 -1635 722
rect -1669 615 -1635 639
rect -1669 543 -1635 571
rect -1669 471 -1635 503
rect -1669 401 -1635 435
rect -1669 333 -1635 365
rect -1669 265 -1635 293
rect -1669 197 -1635 221
rect -1669 114 -1635 149
rect -1551 687 -1517 722
rect -1551 615 -1517 639
rect -1551 543 -1517 571
rect -1551 471 -1517 503
rect -1551 401 -1517 435
rect -1551 333 -1517 365
rect -1551 265 -1517 293
rect -1551 197 -1517 221
rect -1551 114 -1517 149
rect -1433 687 -1399 722
rect -1433 615 -1399 639
rect -1433 543 -1399 571
rect -1433 471 -1399 503
rect -1433 401 -1399 435
rect -1433 333 -1399 365
rect -1433 265 -1399 293
rect -1433 197 -1399 221
rect -1433 114 -1399 149
rect -1315 687 -1281 722
rect -1315 615 -1281 639
rect -1315 543 -1281 571
rect -1315 471 -1281 503
rect -1315 401 -1281 435
rect -1315 333 -1281 365
rect -1315 265 -1281 293
rect -1315 197 -1281 221
rect -1315 114 -1281 149
rect -1197 687 -1163 722
rect -1197 615 -1163 639
rect -1197 543 -1163 571
rect -1197 471 -1163 503
rect -1197 401 -1163 435
rect -1197 333 -1163 365
rect -1197 265 -1163 293
rect -1197 197 -1163 221
rect -1197 114 -1163 149
rect -1079 687 -1045 722
rect -1079 615 -1045 639
rect -1079 543 -1045 571
rect -1079 471 -1045 503
rect -1079 401 -1045 435
rect -1079 333 -1045 365
rect -1079 265 -1045 293
rect -1079 197 -1045 221
rect -1079 114 -1045 149
rect -961 687 -927 722
rect -961 615 -927 639
rect -961 543 -927 571
rect -961 471 -927 503
rect -961 401 -927 435
rect -961 333 -927 365
rect -961 265 -927 293
rect -961 197 -927 221
rect -961 114 -927 149
rect -843 687 -809 722
rect -843 615 -809 639
rect -843 543 -809 571
rect -843 471 -809 503
rect -843 401 -809 435
rect -843 333 -809 365
rect -843 265 -809 293
rect -843 197 -809 221
rect -843 114 -809 149
rect -725 687 -691 722
rect -725 615 -691 639
rect -725 543 -691 571
rect -725 471 -691 503
rect -725 401 -691 435
rect -725 333 -691 365
rect -725 265 -691 293
rect -725 197 -691 221
rect -725 114 -691 149
rect -607 687 -573 722
rect -607 615 -573 639
rect -607 543 -573 571
rect -607 471 -573 503
rect -607 401 -573 435
rect -607 333 -573 365
rect -607 265 -573 293
rect -607 197 -573 221
rect -607 114 -573 149
rect -489 687 -455 722
rect -489 615 -455 639
rect -489 543 -455 571
rect -489 471 -455 503
rect -489 401 -455 435
rect -489 333 -455 365
rect -489 265 -455 293
rect -489 197 -455 221
rect -489 114 -455 149
rect -371 687 -337 722
rect -371 615 -337 639
rect -371 543 -337 571
rect -371 471 -337 503
rect -371 401 -337 435
rect -371 333 -337 365
rect -371 265 -337 293
rect -371 197 -337 221
rect -371 114 -337 149
rect -253 687 -219 722
rect -253 615 -219 639
rect -253 543 -219 571
rect -253 471 -219 503
rect -253 401 -219 435
rect -253 333 -219 365
rect -253 265 -219 293
rect -253 197 -219 221
rect -253 114 -219 149
rect -135 687 -101 722
rect -135 615 -101 639
rect -135 543 -101 571
rect -135 471 -101 503
rect -135 401 -101 435
rect -135 333 -101 365
rect -135 265 -101 293
rect -135 197 -101 221
rect -135 114 -101 149
rect -17 687 17 722
rect -17 615 17 639
rect -17 543 17 571
rect -17 471 17 503
rect -17 401 17 435
rect -17 333 17 365
rect -17 265 17 293
rect -17 197 17 221
rect -17 114 17 149
rect 101 687 135 722
rect 101 615 135 639
rect 101 543 135 571
rect 101 471 135 503
rect 101 401 135 435
rect 101 333 135 365
rect 101 265 135 293
rect 101 197 135 221
rect 101 114 135 149
rect 219 687 253 722
rect 219 615 253 639
rect 219 543 253 571
rect 219 471 253 503
rect 219 401 253 435
rect 219 333 253 365
rect 219 265 253 293
rect 219 197 253 221
rect 219 114 253 149
rect 337 687 371 722
rect 337 615 371 639
rect 337 543 371 571
rect 337 471 371 503
rect 337 401 371 435
rect 337 333 371 365
rect 337 265 371 293
rect 337 197 371 221
rect 337 114 371 149
rect 455 687 489 722
rect 455 615 489 639
rect 455 543 489 571
rect 455 471 489 503
rect 455 401 489 435
rect 455 333 489 365
rect 455 265 489 293
rect 455 197 489 221
rect 455 114 489 149
rect 573 687 607 722
rect 573 615 607 639
rect 573 543 607 571
rect 573 471 607 503
rect 573 401 607 435
rect 573 333 607 365
rect 573 265 607 293
rect 573 197 607 221
rect 573 114 607 149
rect 691 687 725 722
rect 691 615 725 639
rect 691 543 725 571
rect 691 471 725 503
rect 691 401 725 435
rect 691 333 725 365
rect 691 265 725 293
rect 691 197 725 221
rect 691 114 725 149
rect 809 687 843 722
rect 809 615 843 639
rect 809 543 843 571
rect 809 471 843 503
rect 809 401 843 435
rect 809 333 843 365
rect 809 265 843 293
rect 809 197 843 221
rect 809 114 843 149
rect 927 687 961 722
rect 927 615 961 639
rect 927 543 961 571
rect 927 471 961 503
rect 927 401 961 435
rect 927 333 961 365
rect 927 265 961 293
rect 927 197 961 221
rect 927 114 961 149
rect 1045 687 1079 722
rect 1045 615 1079 639
rect 1045 543 1079 571
rect 1045 471 1079 503
rect 1045 401 1079 435
rect 1045 333 1079 365
rect 1045 265 1079 293
rect 1045 197 1079 221
rect 1045 114 1079 149
rect 1163 687 1197 722
rect 1163 615 1197 639
rect 1163 543 1197 571
rect 1163 471 1197 503
rect 1163 401 1197 435
rect 1163 333 1197 365
rect 1163 265 1197 293
rect 1163 197 1197 221
rect 1163 114 1197 149
rect 1281 687 1315 722
rect 1281 615 1315 639
rect 1281 543 1315 571
rect 1281 471 1315 503
rect 1281 401 1315 435
rect 1281 333 1315 365
rect 1281 265 1315 293
rect 1281 197 1315 221
rect 1281 114 1315 149
rect 1399 687 1433 722
rect 1399 615 1433 639
rect 1399 543 1433 571
rect 1399 471 1433 503
rect 1399 401 1433 435
rect 1399 333 1433 365
rect 1399 265 1433 293
rect 1399 197 1433 221
rect 1399 114 1433 149
rect 1517 687 1551 722
rect 1517 615 1551 639
rect 1517 543 1551 571
rect 1517 471 1551 503
rect 1517 401 1551 435
rect 1517 333 1551 365
rect 1517 265 1551 293
rect 1517 197 1551 221
rect 1517 114 1551 149
rect 1635 687 1669 722
rect 1635 615 1669 639
rect 1635 543 1669 571
rect 1635 471 1669 503
rect 1635 401 1669 435
rect 1635 333 1669 365
rect 1635 265 1669 293
rect 1635 197 1669 221
rect 1635 114 1669 149
rect 1753 687 1787 722
rect 1753 615 1787 639
rect 1753 543 1787 571
rect 1753 471 1787 503
rect 1753 401 1787 435
rect 1753 333 1787 365
rect 1753 265 1787 293
rect 1753 197 1787 221
rect 1753 114 1787 149
rect 1871 687 1905 722
rect 1871 615 1905 639
rect 1871 543 1905 571
rect 1871 471 1905 503
rect 1871 401 1905 435
rect 1871 333 1905 365
rect 1871 265 1905 293
rect 1871 197 1905 221
rect 1871 114 1905 149
rect 1989 687 2023 722
rect 1989 615 2023 639
rect 1989 543 2023 571
rect 1989 471 2023 503
rect 1989 401 2023 435
rect 1989 333 2023 365
rect 1989 265 2023 293
rect 1989 197 2023 221
rect 1989 114 2023 149
rect 2107 687 2141 722
rect 2107 615 2141 639
rect 2107 543 2141 571
rect 2107 471 2141 503
rect 2107 401 2141 435
rect 2107 333 2141 365
rect 2107 265 2141 293
rect 2107 197 2141 221
rect 2107 114 2141 149
rect 2225 687 2259 722
rect 2225 615 2259 639
rect 2225 543 2259 571
rect 2225 471 2259 503
rect 2225 401 2259 435
rect 2225 333 2259 365
rect 2225 265 2259 293
rect 2225 197 2259 221
rect 2225 114 2259 149
rect 2343 687 2377 722
rect 2343 615 2377 639
rect 2343 543 2377 571
rect 2343 471 2377 503
rect 2343 401 2377 435
rect 2343 333 2377 365
rect 2343 265 2377 293
rect 2343 197 2377 221
rect 2343 114 2377 149
rect 2461 687 2495 722
rect 2461 615 2495 639
rect 2461 543 2495 571
rect 2461 471 2495 503
rect 2461 401 2495 435
rect 2461 333 2495 365
rect 2461 265 2495 293
rect 2461 197 2495 221
rect 2461 114 2495 149
rect 2579 687 2613 722
rect 2579 615 2613 639
rect 2579 543 2613 571
rect 2579 471 2613 503
rect 2579 401 2613 435
rect 2579 333 2613 365
rect 2579 265 2613 293
rect 2579 197 2613 221
rect 2579 114 2613 149
rect 2697 687 2731 722
rect 2697 615 2731 639
rect 2697 543 2731 571
rect 2697 471 2731 503
rect 2697 401 2731 435
rect 2697 333 2731 365
rect 2697 265 2731 293
rect 2697 197 2731 221
rect 2697 114 2731 149
rect 2815 687 2849 722
rect 2815 615 2849 639
rect 2815 543 2849 571
rect 2815 471 2849 503
rect 2815 401 2849 435
rect 2815 333 2849 365
rect 2815 265 2849 293
rect 2815 197 2849 221
rect 2815 114 2849 149
rect 2933 687 2967 722
rect 2933 615 2967 639
rect 2933 543 2967 571
rect 2933 471 2967 503
rect 2933 401 2967 435
rect 2933 333 2967 365
rect 2933 265 2967 293
rect 2933 197 2967 221
rect 2933 114 2967 149
rect 3047 663 3081 697
rect 3047 595 3081 629
rect 3047 527 3081 561
rect 3047 459 3081 493
rect 3047 391 3081 425
rect 3047 323 3081 357
rect 3047 255 3081 289
rect 3047 187 3081 221
rect 3047 119 3081 153
rect -3081 51 -3047 85
rect -2924 37 -2908 71
rect -2874 37 -2858 71
rect -2806 37 -2790 71
rect -2756 37 -2740 71
rect -2688 37 -2672 71
rect -2638 37 -2622 71
rect -2570 37 -2554 71
rect -2520 37 -2504 71
rect -2452 37 -2436 71
rect -2402 37 -2386 71
rect -2334 37 -2318 71
rect -2284 37 -2268 71
rect -2216 37 -2200 71
rect -2166 37 -2150 71
rect -2098 37 -2082 71
rect -2048 37 -2032 71
rect -1980 37 -1964 71
rect -1930 37 -1914 71
rect -1862 37 -1846 71
rect -1812 37 -1796 71
rect -1744 37 -1728 71
rect -1694 37 -1678 71
rect -1626 37 -1610 71
rect -1576 37 -1560 71
rect -1508 37 -1492 71
rect -1458 37 -1442 71
rect -1390 37 -1374 71
rect -1340 37 -1324 71
rect -1272 37 -1256 71
rect -1222 37 -1206 71
rect -1154 37 -1138 71
rect -1104 37 -1088 71
rect -1036 37 -1020 71
rect -986 37 -970 71
rect -918 37 -902 71
rect -868 37 -852 71
rect -800 37 -784 71
rect -750 37 -734 71
rect -682 37 -666 71
rect -632 37 -616 71
rect -564 37 -548 71
rect -514 37 -498 71
rect -446 37 -430 71
rect -396 37 -380 71
rect -328 37 -312 71
rect -278 37 -262 71
rect -210 37 -194 71
rect -160 37 -144 71
rect -92 37 -76 71
rect -42 37 -26 71
rect 26 37 42 71
rect 76 37 92 71
rect 144 37 160 71
rect 194 37 210 71
rect 262 37 278 71
rect 312 37 328 71
rect 380 37 396 71
rect 430 37 446 71
rect 498 37 514 71
rect 548 37 564 71
rect 616 37 632 71
rect 666 37 682 71
rect 734 37 750 71
rect 784 37 800 71
rect 852 37 868 71
rect 902 37 918 71
rect 970 37 986 71
rect 1020 37 1036 71
rect 1088 37 1104 71
rect 1138 37 1154 71
rect 1206 37 1222 71
rect 1256 37 1272 71
rect 1324 37 1340 71
rect 1374 37 1390 71
rect 1442 37 1458 71
rect 1492 37 1508 71
rect 1560 37 1576 71
rect 1610 37 1626 71
rect 1678 37 1694 71
rect 1728 37 1744 71
rect 1796 37 1812 71
rect 1846 37 1862 71
rect 1914 37 1930 71
rect 1964 37 1980 71
rect 2032 37 2048 71
rect 2082 37 2098 71
rect 2150 37 2166 71
rect 2200 37 2216 71
rect 2268 37 2284 71
rect 2318 37 2334 71
rect 2386 37 2402 71
rect 2436 37 2452 71
rect 2504 37 2520 71
rect 2554 37 2570 71
rect 2622 37 2638 71
rect 2672 37 2688 71
rect 2740 37 2756 71
rect 2790 37 2806 71
rect 2858 37 2874 71
rect 2908 37 2924 71
rect 3047 51 3081 85
rect -3081 -17 -3047 17
rect 3047 -17 3081 17
rect -3081 -85 -3047 -51
rect -2924 -71 -2908 -37
rect -2874 -71 -2858 -37
rect -2806 -71 -2790 -37
rect -2756 -71 -2740 -37
rect -2688 -71 -2672 -37
rect -2638 -71 -2622 -37
rect -2570 -71 -2554 -37
rect -2520 -71 -2504 -37
rect -2452 -71 -2436 -37
rect -2402 -71 -2386 -37
rect -2334 -71 -2318 -37
rect -2284 -71 -2268 -37
rect -2216 -71 -2200 -37
rect -2166 -71 -2150 -37
rect -2098 -71 -2082 -37
rect -2048 -71 -2032 -37
rect -1980 -71 -1964 -37
rect -1930 -71 -1914 -37
rect -1862 -71 -1846 -37
rect -1812 -71 -1796 -37
rect -1744 -71 -1728 -37
rect -1694 -71 -1678 -37
rect -1626 -71 -1610 -37
rect -1576 -71 -1560 -37
rect -1508 -71 -1492 -37
rect -1458 -71 -1442 -37
rect -1390 -71 -1374 -37
rect -1340 -71 -1324 -37
rect -1272 -71 -1256 -37
rect -1222 -71 -1206 -37
rect -1154 -71 -1138 -37
rect -1104 -71 -1088 -37
rect -1036 -71 -1020 -37
rect -986 -71 -970 -37
rect -918 -71 -902 -37
rect -868 -71 -852 -37
rect -800 -71 -784 -37
rect -750 -71 -734 -37
rect -682 -71 -666 -37
rect -632 -71 -616 -37
rect -564 -71 -548 -37
rect -514 -71 -498 -37
rect -446 -71 -430 -37
rect -396 -71 -380 -37
rect -328 -71 -312 -37
rect -278 -71 -262 -37
rect -210 -71 -194 -37
rect -160 -71 -144 -37
rect -92 -71 -76 -37
rect -42 -71 -26 -37
rect 26 -71 42 -37
rect 76 -71 92 -37
rect 144 -71 160 -37
rect 194 -71 210 -37
rect 262 -71 278 -37
rect 312 -71 328 -37
rect 380 -71 396 -37
rect 430 -71 446 -37
rect 498 -71 514 -37
rect 548 -71 564 -37
rect 616 -71 632 -37
rect 666 -71 682 -37
rect 734 -71 750 -37
rect 784 -71 800 -37
rect 852 -71 868 -37
rect 902 -71 918 -37
rect 970 -71 986 -37
rect 1020 -71 1036 -37
rect 1088 -71 1104 -37
rect 1138 -71 1154 -37
rect 1206 -71 1222 -37
rect 1256 -71 1272 -37
rect 1324 -71 1340 -37
rect 1374 -71 1390 -37
rect 1442 -71 1458 -37
rect 1492 -71 1508 -37
rect 1560 -71 1576 -37
rect 1610 -71 1626 -37
rect 1678 -71 1694 -37
rect 1728 -71 1744 -37
rect 1796 -71 1812 -37
rect 1846 -71 1862 -37
rect 1914 -71 1930 -37
rect 1964 -71 1980 -37
rect 2032 -71 2048 -37
rect 2082 -71 2098 -37
rect 2150 -71 2166 -37
rect 2200 -71 2216 -37
rect 2268 -71 2284 -37
rect 2318 -71 2334 -37
rect 2386 -71 2402 -37
rect 2436 -71 2452 -37
rect 2504 -71 2520 -37
rect 2554 -71 2570 -37
rect 2622 -71 2638 -37
rect 2672 -71 2688 -37
rect 2740 -71 2756 -37
rect 2790 -71 2806 -37
rect 2858 -71 2874 -37
rect 2908 -71 2924 -37
rect 3047 -85 3081 -51
rect -3081 -153 -3047 -119
rect -3081 -221 -3047 -187
rect -3081 -289 -3047 -255
rect -3081 -357 -3047 -323
rect -3081 -425 -3047 -391
rect -3081 -493 -3047 -459
rect -3081 -561 -3047 -527
rect -3081 -629 -3047 -595
rect -3081 -697 -3047 -663
rect -2967 -149 -2933 -114
rect -2967 -221 -2933 -197
rect -2967 -293 -2933 -265
rect -2967 -365 -2933 -333
rect -2967 -435 -2933 -401
rect -2967 -503 -2933 -471
rect -2967 -571 -2933 -543
rect -2967 -639 -2933 -615
rect -2967 -722 -2933 -687
rect -2849 -149 -2815 -114
rect -2849 -221 -2815 -197
rect -2849 -293 -2815 -265
rect -2849 -365 -2815 -333
rect -2849 -435 -2815 -401
rect -2849 -503 -2815 -471
rect -2849 -571 -2815 -543
rect -2849 -639 -2815 -615
rect -2849 -722 -2815 -687
rect -2731 -149 -2697 -114
rect -2731 -221 -2697 -197
rect -2731 -293 -2697 -265
rect -2731 -365 -2697 -333
rect -2731 -435 -2697 -401
rect -2731 -503 -2697 -471
rect -2731 -571 -2697 -543
rect -2731 -639 -2697 -615
rect -2731 -722 -2697 -687
rect -2613 -149 -2579 -114
rect -2613 -221 -2579 -197
rect -2613 -293 -2579 -265
rect -2613 -365 -2579 -333
rect -2613 -435 -2579 -401
rect -2613 -503 -2579 -471
rect -2613 -571 -2579 -543
rect -2613 -639 -2579 -615
rect -2613 -722 -2579 -687
rect -2495 -149 -2461 -114
rect -2495 -221 -2461 -197
rect -2495 -293 -2461 -265
rect -2495 -365 -2461 -333
rect -2495 -435 -2461 -401
rect -2495 -503 -2461 -471
rect -2495 -571 -2461 -543
rect -2495 -639 -2461 -615
rect -2495 -722 -2461 -687
rect -2377 -149 -2343 -114
rect -2377 -221 -2343 -197
rect -2377 -293 -2343 -265
rect -2377 -365 -2343 -333
rect -2377 -435 -2343 -401
rect -2377 -503 -2343 -471
rect -2377 -571 -2343 -543
rect -2377 -639 -2343 -615
rect -2377 -722 -2343 -687
rect -2259 -149 -2225 -114
rect -2259 -221 -2225 -197
rect -2259 -293 -2225 -265
rect -2259 -365 -2225 -333
rect -2259 -435 -2225 -401
rect -2259 -503 -2225 -471
rect -2259 -571 -2225 -543
rect -2259 -639 -2225 -615
rect -2259 -722 -2225 -687
rect -2141 -149 -2107 -114
rect -2141 -221 -2107 -197
rect -2141 -293 -2107 -265
rect -2141 -365 -2107 -333
rect -2141 -435 -2107 -401
rect -2141 -503 -2107 -471
rect -2141 -571 -2107 -543
rect -2141 -639 -2107 -615
rect -2141 -722 -2107 -687
rect -2023 -149 -1989 -114
rect -2023 -221 -1989 -197
rect -2023 -293 -1989 -265
rect -2023 -365 -1989 -333
rect -2023 -435 -1989 -401
rect -2023 -503 -1989 -471
rect -2023 -571 -1989 -543
rect -2023 -639 -1989 -615
rect -2023 -722 -1989 -687
rect -1905 -149 -1871 -114
rect -1905 -221 -1871 -197
rect -1905 -293 -1871 -265
rect -1905 -365 -1871 -333
rect -1905 -435 -1871 -401
rect -1905 -503 -1871 -471
rect -1905 -571 -1871 -543
rect -1905 -639 -1871 -615
rect -1905 -722 -1871 -687
rect -1787 -149 -1753 -114
rect -1787 -221 -1753 -197
rect -1787 -293 -1753 -265
rect -1787 -365 -1753 -333
rect -1787 -435 -1753 -401
rect -1787 -503 -1753 -471
rect -1787 -571 -1753 -543
rect -1787 -639 -1753 -615
rect -1787 -722 -1753 -687
rect -1669 -149 -1635 -114
rect -1669 -221 -1635 -197
rect -1669 -293 -1635 -265
rect -1669 -365 -1635 -333
rect -1669 -435 -1635 -401
rect -1669 -503 -1635 -471
rect -1669 -571 -1635 -543
rect -1669 -639 -1635 -615
rect -1669 -722 -1635 -687
rect -1551 -149 -1517 -114
rect -1551 -221 -1517 -197
rect -1551 -293 -1517 -265
rect -1551 -365 -1517 -333
rect -1551 -435 -1517 -401
rect -1551 -503 -1517 -471
rect -1551 -571 -1517 -543
rect -1551 -639 -1517 -615
rect -1551 -722 -1517 -687
rect -1433 -149 -1399 -114
rect -1433 -221 -1399 -197
rect -1433 -293 -1399 -265
rect -1433 -365 -1399 -333
rect -1433 -435 -1399 -401
rect -1433 -503 -1399 -471
rect -1433 -571 -1399 -543
rect -1433 -639 -1399 -615
rect -1433 -722 -1399 -687
rect -1315 -149 -1281 -114
rect -1315 -221 -1281 -197
rect -1315 -293 -1281 -265
rect -1315 -365 -1281 -333
rect -1315 -435 -1281 -401
rect -1315 -503 -1281 -471
rect -1315 -571 -1281 -543
rect -1315 -639 -1281 -615
rect -1315 -722 -1281 -687
rect -1197 -149 -1163 -114
rect -1197 -221 -1163 -197
rect -1197 -293 -1163 -265
rect -1197 -365 -1163 -333
rect -1197 -435 -1163 -401
rect -1197 -503 -1163 -471
rect -1197 -571 -1163 -543
rect -1197 -639 -1163 -615
rect -1197 -722 -1163 -687
rect -1079 -149 -1045 -114
rect -1079 -221 -1045 -197
rect -1079 -293 -1045 -265
rect -1079 -365 -1045 -333
rect -1079 -435 -1045 -401
rect -1079 -503 -1045 -471
rect -1079 -571 -1045 -543
rect -1079 -639 -1045 -615
rect -1079 -722 -1045 -687
rect -961 -149 -927 -114
rect -961 -221 -927 -197
rect -961 -293 -927 -265
rect -961 -365 -927 -333
rect -961 -435 -927 -401
rect -961 -503 -927 -471
rect -961 -571 -927 -543
rect -961 -639 -927 -615
rect -961 -722 -927 -687
rect -843 -149 -809 -114
rect -843 -221 -809 -197
rect -843 -293 -809 -265
rect -843 -365 -809 -333
rect -843 -435 -809 -401
rect -843 -503 -809 -471
rect -843 -571 -809 -543
rect -843 -639 -809 -615
rect -843 -722 -809 -687
rect -725 -149 -691 -114
rect -725 -221 -691 -197
rect -725 -293 -691 -265
rect -725 -365 -691 -333
rect -725 -435 -691 -401
rect -725 -503 -691 -471
rect -725 -571 -691 -543
rect -725 -639 -691 -615
rect -725 -722 -691 -687
rect -607 -149 -573 -114
rect -607 -221 -573 -197
rect -607 -293 -573 -265
rect -607 -365 -573 -333
rect -607 -435 -573 -401
rect -607 -503 -573 -471
rect -607 -571 -573 -543
rect -607 -639 -573 -615
rect -607 -722 -573 -687
rect -489 -149 -455 -114
rect -489 -221 -455 -197
rect -489 -293 -455 -265
rect -489 -365 -455 -333
rect -489 -435 -455 -401
rect -489 -503 -455 -471
rect -489 -571 -455 -543
rect -489 -639 -455 -615
rect -489 -722 -455 -687
rect -371 -149 -337 -114
rect -371 -221 -337 -197
rect -371 -293 -337 -265
rect -371 -365 -337 -333
rect -371 -435 -337 -401
rect -371 -503 -337 -471
rect -371 -571 -337 -543
rect -371 -639 -337 -615
rect -371 -722 -337 -687
rect -253 -149 -219 -114
rect -253 -221 -219 -197
rect -253 -293 -219 -265
rect -253 -365 -219 -333
rect -253 -435 -219 -401
rect -253 -503 -219 -471
rect -253 -571 -219 -543
rect -253 -639 -219 -615
rect -253 -722 -219 -687
rect -135 -149 -101 -114
rect -135 -221 -101 -197
rect -135 -293 -101 -265
rect -135 -365 -101 -333
rect -135 -435 -101 -401
rect -135 -503 -101 -471
rect -135 -571 -101 -543
rect -135 -639 -101 -615
rect -135 -722 -101 -687
rect -17 -149 17 -114
rect -17 -221 17 -197
rect -17 -293 17 -265
rect -17 -365 17 -333
rect -17 -435 17 -401
rect -17 -503 17 -471
rect -17 -571 17 -543
rect -17 -639 17 -615
rect -17 -722 17 -687
rect 101 -149 135 -114
rect 101 -221 135 -197
rect 101 -293 135 -265
rect 101 -365 135 -333
rect 101 -435 135 -401
rect 101 -503 135 -471
rect 101 -571 135 -543
rect 101 -639 135 -615
rect 101 -722 135 -687
rect 219 -149 253 -114
rect 219 -221 253 -197
rect 219 -293 253 -265
rect 219 -365 253 -333
rect 219 -435 253 -401
rect 219 -503 253 -471
rect 219 -571 253 -543
rect 219 -639 253 -615
rect 219 -722 253 -687
rect 337 -149 371 -114
rect 337 -221 371 -197
rect 337 -293 371 -265
rect 337 -365 371 -333
rect 337 -435 371 -401
rect 337 -503 371 -471
rect 337 -571 371 -543
rect 337 -639 371 -615
rect 337 -722 371 -687
rect 455 -149 489 -114
rect 455 -221 489 -197
rect 455 -293 489 -265
rect 455 -365 489 -333
rect 455 -435 489 -401
rect 455 -503 489 -471
rect 455 -571 489 -543
rect 455 -639 489 -615
rect 455 -722 489 -687
rect 573 -149 607 -114
rect 573 -221 607 -197
rect 573 -293 607 -265
rect 573 -365 607 -333
rect 573 -435 607 -401
rect 573 -503 607 -471
rect 573 -571 607 -543
rect 573 -639 607 -615
rect 573 -722 607 -687
rect 691 -149 725 -114
rect 691 -221 725 -197
rect 691 -293 725 -265
rect 691 -365 725 -333
rect 691 -435 725 -401
rect 691 -503 725 -471
rect 691 -571 725 -543
rect 691 -639 725 -615
rect 691 -722 725 -687
rect 809 -149 843 -114
rect 809 -221 843 -197
rect 809 -293 843 -265
rect 809 -365 843 -333
rect 809 -435 843 -401
rect 809 -503 843 -471
rect 809 -571 843 -543
rect 809 -639 843 -615
rect 809 -722 843 -687
rect 927 -149 961 -114
rect 927 -221 961 -197
rect 927 -293 961 -265
rect 927 -365 961 -333
rect 927 -435 961 -401
rect 927 -503 961 -471
rect 927 -571 961 -543
rect 927 -639 961 -615
rect 927 -722 961 -687
rect 1045 -149 1079 -114
rect 1045 -221 1079 -197
rect 1045 -293 1079 -265
rect 1045 -365 1079 -333
rect 1045 -435 1079 -401
rect 1045 -503 1079 -471
rect 1045 -571 1079 -543
rect 1045 -639 1079 -615
rect 1045 -722 1079 -687
rect 1163 -149 1197 -114
rect 1163 -221 1197 -197
rect 1163 -293 1197 -265
rect 1163 -365 1197 -333
rect 1163 -435 1197 -401
rect 1163 -503 1197 -471
rect 1163 -571 1197 -543
rect 1163 -639 1197 -615
rect 1163 -722 1197 -687
rect 1281 -149 1315 -114
rect 1281 -221 1315 -197
rect 1281 -293 1315 -265
rect 1281 -365 1315 -333
rect 1281 -435 1315 -401
rect 1281 -503 1315 -471
rect 1281 -571 1315 -543
rect 1281 -639 1315 -615
rect 1281 -722 1315 -687
rect 1399 -149 1433 -114
rect 1399 -221 1433 -197
rect 1399 -293 1433 -265
rect 1399 -365 1433 -333
rect 1399 -435 1433 -401
rect 1399 -503 1433 -471
rect 1399 -571 1433 -543
rect 1399 -639 1433 -615
rect 1399 -722 1433 -687
rect 1517 -149 1551 -114
rect 1517 -221 1551 -197
rect 1517 -293 1551 -265
rect 1517 -365 1551 -333
rect 1517 -435 1551 -401
rect 1517 -503 1551 -471
rect 1517 -571 1551 -543
rect 1517 -639 1551 -615
rect 1517 -722 1551 -687
rect 1635 -149 1669 -114
rect 1635 -221 1669 -197
rect 1635 -293 1669 -265
rect 1635 -365 1669 -333
rect 1635 -435 1669 -401
rect 1635 -503 1669 -471
rect 1635 -571 1669 -543
rect 1635 -639 1669 -615
rect 1635 -722 1669 -687
rect 1753 -149 1787 -114
rect 1753 -221 1787 -197
rect 1753 -293 1787 -265
rect 1753 -365 1787 -333
rect 1753 -435 1787 -401
rect 1753 -503 1787 -471
rect 1753 -571 1787 -543
rect 1753 -639 1787 -615
rect 1753 -722 1787 -687
rect 1871 -149 1905 -114
rect 1871 -221 1905 -197
rect 1871 -293 1905 -265
rect 1871 -365 1905 -333
rect 1871 -435 1905 -401
rect 1871 -503 1905 -471
rect 1871 -571 1905 -543
rect 1871 -639 1905 -615
rect 1871 -722 1905 -687
rect 1989 -149 2023 -114
rect 1989 -221 2023 -197
rect 1989 -293 2023 -265
rect 1989 -365 2023 -333
rect 1989 -435 2023 -401
rect 1989 -503 2023 -471
rect 1989 -571 2023 -543
rect 1989 -639 2023 -615
rect 1989 -722 2023 -687
rect 2107 -149 2141 -114
rect 2107 -221 2141 -197
rect 2107 -293 2141 -265
rect 2107 -365 2141 -333
rect 2107 -435 2141 -401
rect 2107 -503 2141 -471
rect 2107 -571 2141 -543
rect 2107 -639 2141 -615
rect 2107 -722 2141 -687
rect 2225 -149 2259 -114
rect 2225 -221 2259 -197
rect 2225 -293 2259 -265
rect 2225 -365 2259 -333
rect 2225 -435 2259 -401
rect 2225 -503 2259 -471
rect 2225 -571 2259 -543
rect 2225 -639 2259 -615
rect 2225 -722 2259 -687
rect 2343 -149 2377 -114
rect 2343 -221 2377 -197
rect 2343 -293 2377 -265
rect 2343 -365 2377 -333
rect 2343 -435 2377 -401
rect 2343 -503 2377 -471
rect 2343 -571 2377 -543
rect 2343 -639 2377 -615
rect 2343 -722 2377 -687
rect 2461 -149 2495 -114
rect 2461 -221 2495 -197
rect 2461 -293 2495 -265
rect 2461 -365 2495 -333
rect 2461 -435 2495 -401
rect 2461 -503 2495 -471
rect 2461 -571 2495 -543
rect 2461 -639 2495 -615
rect 2461 -722 2495 -687
rect 2579 -149 2613 -114
rect 2579 -221 2613 -197
rect 2579 -293 2613 -265
rect 2579 -365 2613 -333
rect 2579 -435 2613 -401
rect 2579 -503 2613 -471
rect 2579 -571 2613 -543
rect 2579 -639 2613 -615
rect 2579 -722 2613 -687
rect 2697 -149 2731 -114
rect 2697 -221 2731 -197
rect 2697 -293 2731 -265
rect 2697 -365 2731 -333
rect 2697 -435 2731 -401
rect 2697 -503 2731 -471
rect 2697 -571 2731 -543
rect 2697 -639 2731 -615
rect 2697 -722 2731 -687
rect 2815 -149 2849 -114
rect 2815 -221 2849 -197
rect 2815 -293 2849 -265
rect 2815 -365 2849 -333
rect 2815 -435 2849 -401
rect 2815 -503 2849 -471
rect 2815 -571 2849 -543
rect 2815 -639 2849 -615
rect 2815 -722 2849 -687
rect 2933 -149 2967 -114
rect 2933 -221 2967 -197
rect 2933 -293 2967 -265
rect 2933 -365 2967 -333
rect 2933 -435 2967 -401
rect 2933 -503 2967 -471
rect 2933 -571 2967 -543
rect 2933 -639 2967 -615
rect 2933 -722 2967 -687
rect 3047 -153 3081 -119
rect 3047 -221 3081 -187
rect 3047 -289 3081 -255
rect 3047 -357 3081 -323
rect 3047 -425 3081 -391
rect 3047 -493 3081 -459
rect 3047 -561 3081 -527
rect 3047 -629 3081 -595
rect 3047 -697 3081 -663
rect -3081 -765 -3047 -731
rect -3081 -867 -3047 -799
rect 3047 -765 3081 -731
rect 3047 -867 3081 -799
rect -3081 -901 -2975 -867
rect -2941 -901 -2907 -867
rect -2873 -901 -2839 -867
rect -2805 -901 -2771 -867
rect -2737 -901 -2703 -867
rect -2669 -901 -2635 -867
rect -2601 -901 -2567 -867
rect -2533 -901 -2499 -867
rect -2465 -901 -2431 -867
rect -2397 -901 -2363 -867
rect -2329 -901 -2295 -867
rect -2261 -901 -2227 -867
rect -2193 -901 -2159 -867
rect -2125 -901 -2091 -867
rect -2057 -901 -2023 -867
rect -1989 -901 -1955 -867
rect -1921 -901 -1887 -867
rect -1853 -901 -1819 -867
rect -1785 -901 -1751 -867
rect -1717 -901 -1683 -867
rect -1649 -901 -1615 -867
rect -1581 -901 -1547 -867
rect -1513 -901 -1479 -867
rect -1445 -901 -1411 -867
rect -1377 -901 -1343 -867
rect -1309 -901 -1275 -867
rect -1241 -901 -1207 -867
rect -1173 -901 -1139 -867
rect -1105 -901 -1071 -867
rect -1037 -901 -1003 -867
rect -969 -901 -935 -867
rect -901 -901 -867 -867
rect -833 -901 -799 -867
rect -765 -901 -731 -867
rect -697 -901 -663 -867
rect -629 -901 -595 -867
rect -561 -901 -527 -867
rect -493 -901 -459 -867
rect -425 -901 -391 -867
rect -357 -901 -323 -867
rect -289 -901 -255 -867
rect -221 -901 -187 -867
rect -153 -901 -119 -867
rect -85 -901 -51 -867
rect -17 -901 17 -867
rect 51 -901 85 -867
rect 119 -901 153 -867
rect 187 -901 221 -867
rect 255 -901 289 -867
rect 323 -901 357 -867
rect 391 -901 425 -867
rect 459 -901 493 -867
rect 527 -901 561 -867
rect 595 -901 629 -867
rect 663 -901 697 -867
rect 731 -901 765 -867
rect 799 -901 833 -867
rect 867 -901 901 -867
rect 935 -901 969 -867
rect 1003 -901 1037 -867
rect 1071 -901 1105 -867
rect 1139 -901 1173 -867
rect 1207 -901 1241 -867
rect 1275 -901 1309 -867
rect 1343 -901 1377 -867
rect 1411 -901 1445 -867
rect 1479 -901 1513 -867
rect 1547 -901 1581 -867
rect 1615 -901 1649 -867
rect 1683 -901 1717 -867
rect 1751 -901 1785 -867
rect 1819 -901 1853 -867
rect 1887 -901 1921 -867
rect 1955 -901 1989 -867
rect 2023 -901 2057 -867
rect 2091 -901 2125 -867
rect 2159 -901 2193 -867
rect 2227 -901 2261 -867
rect 2295 -901 2329 -867
rect 2363 -901 2397 -867
rect 2431 -901 2465 -867
rect 2499 -901 2533 -867
rect 2567 -901 2601 -867
rect 2635 -901 2669 -867
rect 2703 -901 2737 -867
rect 2771 -901 2805 -867
rect 2839 -901 2873 -867
rect 2907 -901 2941 -867
rect 2975 -901 3081 -867
<< viali >>
rect -2967 673 -2933 687
rect -2967 653 -2933 673
rect -2967 605 -2933 615
rect -2967 581 -2933 605
rect -2967 537 -2933 543
rect -2967 509 -2933 537
rect -2967 469 -2933 471
rect -2967 437 -2933 469
rect -2967 367 -2933 399
rect -2967 365 -2933 367
rect -2967 299 -2933 327
rect -2967 293 -2933 299
rect -2967 231 -2933 255
rect -2967 221 -2933 231
rect -2967 163 -2933 183
rect -2967 149 -2933 163
rect -2849 673 -2815 687
rect -2849 653 -2815 673
rect -2849 605 -2815 615
rect -2849 581 -2815 605
rect -2849 537 -2815 543
rect -2849 509 -2815 537
rect -2849 469 -2815 471
rect -2849 437 -2815 469
rect -2849 367 -2815 399
rect -2849 365 -2815 367
rect -2849 299 -2815 327
rect -2849 293 -2815 299
rect -2849 231 -2815 255
rect -2849 221 -2815 231
rect -2849 163 -2815 183
rect -2849 149 -2815 163
rect -2731 673 -2697 687
rect -2731 653 -2697 673
rect -2731 605 -2697 615
rect -2731 581 -2697 605
rect -2731 537 -2697 543
rect -2731 509 -2697 537
rect -2731 469 -2697 471
rect -2731 437 -2697 469
rect -2731 367 -2697 399
rect -2731 365 -2697 367
rect -2731 299 -2697 327
rect -2731 293 -2697 299
rect -2731 231 -2697 255
rect -2731 221 -2697 231
rect -2731 163 -2697 183
rect -2731 149 -2697 163
rect -2613 673 -2579 687
rect -2613 653 -2579 673
rect -2613 605 -2579 615
rect -2613 581 -2579 605
rect -2613 537 -2579 543
rect -2613 509 -2579 537
rect -2613 469 -2579 471
rect -2613 437 -2579 469
rect -2613 367 -2579 399
rect -2613 365 -2579 367
rect -2613 299 -2579 327
rect -2613 293 -2579 299
rect -2613 231 -2579 255
rect -2613 221 -2579 231
rect -2613 163 -2579 183
rect -2613 149 -2579 163
rect -2495 673 -2461 687
rect -2495 653 -2461 673
rect -2495 605 -2461 615
rect -2495 581 -2461 605
rect -2495 537 -2461 543
rect -2495 509 -2461 537
rect -2495 469 -2461 471
rect -2495 437 -2461 469
rect -2495 367 -2461 399
rect -2495 365 -2461 367
rect -2495 299 -2461 327
rect -2495 293 -2461 299
rect -2495 231 -2461 255
rect -2495 221 -2461 231
rect -2495 163 -2461 183
rect -2495 149 -2461 163
rect -2377 673 -2343 687
rect -2377 653 -2343 673
rect -2377 605 -2343 615
rect -2377 581 -2343 605
rect -2377 537 -2343 543
rect -2377 509 -2343 537
rect -2377 469 -2343 471
rect -2377 437 -2343 469
rect -2377 367 -2343 399
rect -2377 365 -2343 367
rect -2377 299 -2343 327
rect -2377 293 -2343 299
rect -2377 231 -2343 255
rect -2377 221 -2343 231
rect -2377 163 -2343 183
rect -2377 149 -2343 163
rect -2259 673 -2225 687
rect -2259 653 -2225 673
rect -2259 605 -2225 615
rect -2259 581 -2225 605
rect -2259 537 -2225 543
rect -2259 509 -2225 537
rect -2259 469 -2225 471
rect -2259 437 -2225 469
rect -2259 367 -2225 399
rect -2259 365 -2225 367
rect -2259 299 -2225 327
rect -2259 293 -2225 299
rect -2259 231 -2225 255
rect -2259 221 -2225 231
rect -2259 163 -2225 183
rect -2259 149 -2225 163
rect -2141 673 -2107 687
rect -2141 653 -2107 673
rect -2141 605 -2107 615
rect -2141 581 -2107 605
rect -2141 537 -2107 543
rect -2141 509 -2107 537
rect -2141 469 -2107 471
rect -2141 437 -2107 469
rect -2141 367 -2107 399
rect -2141 365 -2107 367
rect -2141 299 -2107 327
rect -2141 293 -2107 299
rect -2141 231 -2107 255
rect -2141 221 -2107 231
rect -2141 163 -2107 183
rect -2141 149 -2107 163
rect -2023 673 -1989 687
rect -2023 653 -1989 673
rect -2023 605 -1989 615
rect -2023 581 -1989 605
rect -2023 537 -1989 543
rect -2023 509 -1989 537
rect -2023 469 -1989 471
rect -2023 437 -1989 469
rect -2023 367 -1989 399
rect -2023 365 -1989 367
rect -2023 299 -1989 327
rect -2023 293 -1989 299
rect -2023 231 -1989 255
rect -2023 221 -1989 231
rect -2023 163 -1989 183
rect -2023 149 -1989 163
rect -1905 673 -1871 687
rect -1905 653 -1871 673
rect -1905 605 -1871 615
rect -1905 581 -1871 605
rect -1905 537 -1871 543
rect -1905 509 -1871 537
rect -1905 469 -1871 471
rect -1905 437 -1871 469
rect -1905 367 -1871 399
rect -1905 365 -1871 367
rect -1905 299 -1871 327
rect -1905 293 -1871 299
rect -1905 231 -1871 255
rect -1905 221 -1871 231
rect -1905 163 -1871 183
rect -1905 149 -1871 163
rect -1787 673 -1753 687
rect -1787 653 -1753 673
rect -1787 605 -1753 615
rect -1787 581 -1753 605
rect -1787 537 -1753 543
rect -1787 509 -1753 537
rect -1787 469 -1753 471
rect -1787 437 -1753 469
rect -1787 367 -1753 399
rect -1787 365 -1753 367
rect -1787 299 -1753 327
rect -1787 293 -1753 299
rect -1787 231 -1753 255
rect -1787 221 -1753 231
rect -1787 163 -1753 183
rect -1787 149 -1753 163
rect -1669 673 -1635 687
rect -1669 653 -1635 673
rect -1669 605 -1635 615
rect -1669 581 -1635 605
rect -1669 537 -1635 543
rect -1669 509 -1635 537
rect -1669 469 -1635 471
rect -1669 437 -1635 469
rect -1669 367 -1635 399
rect -1669 365 -1635 367
rect -1669 299 -1635 327
rect -1669 293 -1635 299
rect -1669 231 -1635 255
rect -1669 221 -1635 231
rect -1669 163 -1635 183
rect -1669 149 -1635 163
rect -1551 673 -1517 687
rect -1551 653 -1517 673
rect -1551 605 -1517 615
rect -1551 581 -1517 605
rect -1551 537 -1517 543
rect -1551 509 -1517 537
rect -1551 469 -1517 471
rect -1551 437 -1517 469
rect -1551 367 -1517 399
rect -1551 365 -1517 367
rect -1551 299 -1517 327
rect -1551 293 -1517 299
rect -1551 231 -1517 255
rect -1551 221 -1517 231
rect -1551 163 -1517 183
rect -1551 149 -1517 163
rect -1433 673 -1399 687
rect -1433 653 -1399 673
rect -1433 605 -1399 615
rect -1433 581 -1399 605
rect -1433 537 -1399 543
rect -1433 509 -1399 537
rect -1433 469 -1399 471
rect -1433 437 -1399 469
rect -1433 367 -1399 399
rect -1433 365 -1399 367
rect -1433 299 -1399 327
rect -1433 293 -1399 299
rect -1433 231 -1399 255
rect -1433 221 -1399 231
rect -1433 163 -1399 183
rect -1433 149 -1399 163
rect -1315 673 -1281 687
rect -1315 653 -1281 673
rect -1315 605 -1281 615
rect -1315 581 -1281 605
rect -1315 537 -1281 543
rect -1315 509 -1281 537
rect -1315 469 -1281 471
rect -1315 437 -1281 469
rect -1315 367 -1281 399
rect -1315 365 -1281 367
rect -1315 299 -1281 327
rect -1315 293 -1281 299
rect -1315 231 -1281 255
rect -1315 221 -1281 231
rect -1315 163 -1281 183
rect -1315 149 -1281 163
rect -1197 673 -1163 687
rect -1197 653 -1163 673
rect -1197 605 -1163 615
rect -1197 581 -1163 605
rect -1197 537 -1163 543
rect -1197 509 -1163 537
rect -1197 469 -1163 471
rect -1197 437 -1163 469
rect -1197 367 -1163 399
rect -1197 365 -1163 367
rect -1197 299 -1163 327
rect -1197 293 -1163 299
rect -1197 231 -1163 255
rect -1197 221 -1163 231
rect -1197 163 -1163 183
rect -1197 149 -1163 163
rect -1079 673 -1045 687
rect -1079 653 -1045 673
rect -1079 605 -1045 615
rect -1079 581 -1045 605
rect -1079 537 -1045 543
rect -1079 509 -1045 537
rect -1079 469 -1045 471
rect -1079 437 -1045 469
rect -1079 367 -1045 399
rect -1079 365 -1045 367
rect -1079 299 -1045 327
rect -1079 293 -1045 299
rect -1079 231 -1045 255
rect -1079 221 -1045 231
rect -1079 163 -1045 183
rect -1079 149 -1045 163
rect -961 673 -927 687
rect -961 653 -927 673
rect -961 605 -927 615
rect -961 581 -927 605
rect -961 537 -927 543
rect -961 509 -927 537
rect -961 469 -927 471
rect -961 437 -927 469
rect -961 367 -927 399
rect -961 365 -927 367
rect -961 299 -927 327
rect -961 293 -927 299
rect -961 231 -927 255
rect -961 221 -927 231
rect -961 163 -927 183
rect -961 149 -927 163
rect -843 673 -809 687
rect -843 653 -809 673
rect -843 605 -809 615
rect -843 581 -809 605
rect -843 537 -809 543
rect -843 509 -809 537
rect -843 469 -809 471
rect -843 437 -809 469
rect -843 367 -809 399
rect -843 365 -809 367
rect -843 299 -809 327
rect -843 293 -809 299
rect -843 231 -809 255
rect -843 221 -809 231
rect -843 163 -809 183
rect -843 149 -809 163
rect -725 673 -691 687
rect -725 653 -691 673
rect -725 605 -691 615
rect -725 581 -691 605
rect -725 537 -691 543
rect -725 509 -691 537
rect -725 469 -691 471
rect -725 437 -691 469
rect -725 367 -691 399
rect -725 365 -691 367
rect -725 299 -691 327
rect -725 293 -691 299
rect -725 231 -691 255
rect -725 221 -691 231
rect -725 163 -691 183
rect -725 149 -691 163
rect -607 673 -573 687
rect -607 653 -573 673
rect -607 605 -573 615
rect -607 581 -573 605
rect -607 537 -573 543
rect -607 509 -573 537
rect -607 469 -573 471
rect -607 437 -573 469
rect -607 367 -573 399
rect -607 365 -573 367
rect -607 299 -573 327
rect -607 293 -573 299
rect -607 231 -573 255
rect -607 221 -573 231
rect -607 163 -573 183
rect -607 149 -573 163
rect -489 673 -455 687
rect -489 653 -455 673
rect -489 605 -455 615
rect -489 581 -455 605
rect -489 537 -455 543
rect -489 509 -455 537
rect -489 469 -455 471
rect -489 437 -455 469
rect -489 367 -455 399
rect -489 365 -455 367
rect -489 299 -455 327
rect -489 293 -455 299
rect -489 231 -455 255
rect -489 221 -455 231
rect -489 163 -455 183
rect -489 149 -455 163
rect -371 673 -337 687
rect -371 653 -337 673
rect -371 605 -337 615
rect -371 581 -337 605
rect -371 537 -337 543
rect -371 509 -337 537
rect -371 469 -337 471
rect -371 437 -337 469
rect -371 367 -337 399
rect -371 365 -337 367
rect -371 299 -337 327
rect -371 293 -337 299
rect -371 231 -337 255
rect -371 221 -337 231
rect -371 163 -337 183
rect -371 149 -337 163
rect -253 673 -219 687
rect -253 653 -219 673
rect -253 605 -219 615
rect -253 581 -219 605
rect -253 537 -219 543
rect -253 509 -219 537
rect -253 469 -219 471
rect -253 437 -219 469
rect -253 367 -219 399
rect -253 365 -219 367
rect -253 299 -219 327
rect -253 293 -219 299
rect -253 231 -219 255
rect -253 221 -219 231
rect -253 163 -219 183
rect -253 149 -219 163
rect -135 673 -101 687
rect -135 653 -101 673
rect -135 605 -101 615
rect -135 581 -101 605
rect -135 537 -101 543
rect -135 509 -101 537
rect -135 469 -101 471
rect -135 437 -101 469
rect -135 367 -101 399
rect -135 365 -101 367
rect -135 299 -101 327
rect -135 293 -101 299
rect -135 231 -101 255
rect -135 221 -101 231
rect -135 163 -101 183
rect -135 149 -101 163
rect -17 673 17 687
rect -17 653 17 673
rect -17 605 17 615
rect -17 581 17 605
rect -17 537 17 543
rect -17 509 17 537
rect -17 469 17 471
rect -17 437 17 469
rect -17 367 17 399
rect -17 365 17 367
rect -17 299 17 327
rect -17 293 17 299
rect -17 231 17 255
rect -17 221 17 231
rect -17 163 17 183
rect -17 149 17 163
rect 101 673 135 687
rect 101 653 135 673
rect 101 605 135 615
rect 101 581 135 605
rect 101 537 135 543
rect 101 509 135 537
rect 101 469 135 471
rect 101 437 135 469
rect 101 367 135 399
rect 101 365 135 367
rect 101 299 135 327
rect 101 293 135 299
rect 101 231 135 255
rect 101 221 135 231
rect 101 163 135 183
rect 101 149 135 163
rect 219 673 253 687
rect 219 653 253 673
rect 219 605 253 615
rect 219 581 253 605
rect 219 537 253 543
rect 219 509 253 537
rect 219 469 253 471
rect 219 437 253 469
rect 219 367 253 399
rect 219 365 253 367
rect 219 299 253 327
rect 219 293 253 299
rect 219 231 253 255
rect 219 221 253 231
rect 219 163 253 183
rect 219 149 253 163
rect 337 673 371 687
rect 337 653 371 673
rect 337 605 371 615
rect 337 581 371 605
rect 337 537 371 543
rect 337 509 371 537
rect 337 469 371 471
rect 337 437 371 469
rect 337 367 371 399
rect 337 365 371 367
rect 337 299 371 327
rect 337 293 371 299
rect 337 231 371 255
rect 337 221 371 231
rect 337 163 371 183
rect 337 149 371 163
rect 455 673 489 687
rect 455 653 489 673
rect 455 605 489 615
rect 455 581 489 605
rect 455 537 489 543
rect 455 509 489 537
rect 455 469 489 471
rect 455 437 489 469
rect 455 367 489 399
rect 455 365 489 367
rect 455 299 489 327
rect 455 293 489 299
rect 455 231 489 255
rect 455 221 489 231
rect 455 163 489 183
rect 455 149 489 163
rect 573 673 607 687
rect 573 653 607 673
rect 573 605 607 615
rect 573 581 607 605
rect 573 537 607 543
rect 573 509 607 537
rect 573 469 607 471
rect 573 437 607 469
rect 573 367 607 399
rect 573 365 607 367
rect 573 299 607 327
rect 573 293 607 299
rect 573 231 607 255
rect 573 221 607 231
rect 573 163 607 183
rect 573 149 607 163
rect 691 673 725 687
rect 691 653 725 673
rect 691 605 725 615
rect 691 581 725 605
rect 691 537 725 543
rect 691 509 725 537
rect 691 469 725 471
rect 691 437 725 469
rect 691 367 725 399
rect 691 365 725 367
rect 691 299 725 327
rect 691 293 725 299
rect 691 231 725 255
rect 691 221 725 231
rect 691 163 725 183
rect 691 149 725 163
rect 809 673 843 687
rect 809 653 843 673
rect 809 605 843 615
rect 809 581 843 605
rect 809 537 843 543
rect 809 509 843 537
rect 809 469 843 471
rect 809 437 843 469
rect 809 367 843 399
rect 809 365 843 367
rect 809 299 843 327
rect 809 293 843 299
rect 809 231 843 255
rect 809 221 843 231
rect 809 163 843 183
rect 809 149 843 163
rect 927 673 961 687
rect 927 653 961 673
rect 927 605 961 615
rect 927 581 961 605
rect 927 537 961 543
rect 927 509 961 537
rect 927 469 961 471
rect 927 437 961 469
rect 927 367 961 399
rect 927 365 961 367
rect 927 299 961 327
rect 927 293 961 299
rect 927 231 961 255
rect 927 221 961 231
rect 927 163 961 183
rect 927 149 961 163
rect 1045 673 1079 687
rect 1045 653 1079 673
rect 1045 605 1079 615
rect 1045 581 1079 605
rect 1045 537 1079 543
rect 1045 509 1079 537
rect 1045 469 1079 471
rect 1045 437 1079 469
rect 1045 367 1079 399
rect 1045 365 1079 367
rect 1045 299 1079 327
rect 1045 293 1079 299
rect 1045 231 1079 255
rect 1045 221 1079 231
rect 1045 163 1079 183
rect 1045 149 1079 163
rect 1163 673 1197 687
rect 1163 653 1197 673
rect 1163 605 1197 615
rect 1163 581 1197 605
rect 1163 537 1197 543
rect 1163 509 1197 537
rect 1163 469 1197 471
rect 1163 437 1197 469
rect 1163 367 1197 399
rect 1163 365 1197 367
rect 1163 299 1197 327
rect 1163 293 1197 299
rect 1163 231 1197 255
rect 1163 221 1197 231
rect 1163 163 1197 183
rect 1163 149 1197 163
rect 1281 673 1315 687
rect 1281 653 1315 673
rect 1281 605 1315 615
rect 1281 581 1315 605
rect 1281 537 1315 543
rect 1281 509 1315 537
rect 1281 469 1315 471
rect 1281 437 1315 469
rect 1281 367 1315 399
rect 1281 365 1315 367
rect 1281 299 1315 327
rect 1281 293 1315 299
rect 1281 231 1315 255
rect 1281 221 1315 231
rect 1281 163 1315 183
rect 1281 149 1315 163
rect 1399 673 1433 687
rect 1399 653 1433 673
rect 1399 605 1433 615
rect 1399 581 1433 605
rect 1399 537 1433 543
rect 1399 509 1433 537
rect 1399 469 1433 471
rect 1399 437 1433 469
rect 1399 367 1433 399
rect 1399 365 1433 367
rect 1399 299 1433 327
rect 1399 293 1433 299
rect 1399 231 1433 255
rect 1399 221 1433 231
rect 1399 163 1433 183
rect 1399 149 1433 163
rect 1517 673 1551 687
rect 1517 653 1551 673
rect 1517 605 1551 615
rect 1517 581 1551 605
rect 1517 537 1551 543
rect 1517 509 1551 537
rect 1517 469 1551 471
rect 1517 437 1551 469
rect 1517 367 1551 399
rect 1517 365 1551 367
rect 1517 299 1551 327
rect 1517 293 1551 299
rect 1517 231 1551 255
rect 1517 221 1551 231
rect 1517 163 1551 183
rect 1517 149 1551 163
rect 1635 673 1669 687
rect 1635 653 1669 673
rect 1635 605 1669 615
rect 1635 581 1669 605
rect 1635 537 1669 543
rect 1635 509 1669 537
rect 1635 469 1669 471
rect 1635 437 1669 469
rect 1635 367 1669 399
rect 1635 365 1669 367
rect 1635 299 1669 327
rect 1635 293 1669 299
rect 1635 231 1669 255
rect 1635 221 1669 231
rect 1635 163 1669 183
rect 1635 149 1669 163
rect 1753 673 1787 687
rect 1753 653 1787 673
rect 1753 605 1787 615
rect 1753 581 1787 605
rect 1753 537 1787 543
rect 1753 509 1787 537
rect 1753 469 1787 471
rect 1753 437 1787 469
rect 1753 367 1787 399
rect 1753 365 1787 367
rect 1753 299 1787 327
rect 1753 293 1787 299
rect 1753 231 1787 255
rect 1753 221 1787 231
rect 1753 163 1787 183
rect 1753 149 1787 163
rect 1871 673 1905 687
rect 1871 653 1905 673
rect 1871 605 1905 615
rect 1871 581 1905 605
rect 1871 537 1905 543
rect 1871 509 1905 537
rect 1871 469 1905 471
rect 1871 437 1905 469
rect 1871 367 1905 399
rect 1871 365 1905 367
rect 1871 299 1905 327
rect 1871 293 1905 299
rect 1871 231 1905 255
rect 1871 221 1905 231
rect 1871 163 1905 183
rect 1871 149 1905 163
rect 1989 673 2023 687
rect 1989 653 2023 673
rect 1989 605 2023 615
rect 1989 581 2023 605
rect 1989 537 2023 543
rect 1989 509 2023 537
rect 1989 469 2023 471
rect 1989 437 2023 469
rect 1989 367 2023 399
rect 1989 365 2023 367
rect 1989 299 2023 327
rect 1989 293 2023 299
rect 1989 231 2023 255
rect 1989 221 2023 231
rect 1989 163 2023 183
rect 1989 149 2023 163
rect 2107 673 2141 687
rect 2107 653 2141 673
rect 2107 605 2141 615
rect 2107 581 2141 605
rect 2107 537 2141 543
rect 2107 509 2141 537
rect 2107 469 2141 471
rect 2107 437 2141 469
rect 2107 367 2141 399
rect 2107 365 2141 367
rect 2107 299 2141 327
rect 2107 293 2141 299
rect 2107 231 2141 255
rect 2107 221 2141 231
rect 2107 163 2141 183
rect 2107 149 2141 163
rect 2225 673 2259 687
rect 2225 653 2259 673
rect 2225 605 2259 615
rect 2225 581 2259 605
rect 2225 537 2259 543
rect 2225 509 2259 537
rect 2225 469 2259 471
rect 2225 437 2259 469
rect 2225 367 2259 399
rect 2225 365 2259 367
rect 2225 299 2259 327
rect 2225 293 2259 299
rect 2225 231 2259 255
rect 2225 221 2259 231
rect 2225 163 2259 183
rect 2225 149 2259 163
rect 2343 673 2377 687
rect 2343 653 2377 673
rect 2343 605 2377 615
rect 2343 581 2377 605
rect 2343 537 2377 543
rect 2343 509 2377 537
rect 2343 469 2377 471
rect 2343 437 2377 469
rect 2343 367 2377 399
rect 2343 365 2377 367
rect 2343 299 2377 327
rect 2343 293 2377 299
rect 2343 231 2377 255
rect 2343 221 2377 231
rect 2343 163 2377 183
rect 2343 149 2377 163
rect 2461 673 2495 687
rect 2461 653 2495 673
rect 2461 605 2495 615
rect 2461 581 2495 605
rect 2461 537 2495 543
rect 2461 509 2495 537
rect 2461 469 2495 471
rect 2461 437 2495 469
rect 2461 367 2495 399
rect 2461 365 2495 367
rect 2461 299 2495 327
rect 2461 293 2495 299
rect 2461 231 2495 255
rect 2461 221 2495 231
rect 2461 163 2495 183
rect 2461 149 2495 163
rect 2579 673 2613 687
rect 2579 653 2613 673
rect 2579 605 2613 615
rect 2579 581 2613 605
rect 2579 537 2613 543
rect 2579 509 2613 537
rect 2579 469 2613 471
rect 2579 437 2613 469
rect 2579 367 2613 399
rect 2579 365 2613 367
rect 2579 299 2613 327
rect 2579 293 2613 299
rect 2579 231 2613 255
rect 2579 221 2613 231
rect 2579 163 2613 183
rect 2579 149 2613 163
rect 2697 673 2731 687
rect 2697 653 2731 673
rect 2697 605 2731 615
rect 2697 581 2731 605
rect 2697 537 2731 543
rect 2697 509 2731 537
rect 2697 469 2731 471
rect 2697 437 2731 469
rect 2697 367 2731 399
rect 2697 365 2731 367
rect 2697 299 2731 327
rect 2697 293 2731 299
rect 2697 231 2731 255
rect 2697 221 2731 231
rect 2697 163 2731 183
rect 2697 149 2731 163
rect 2815 673 2849 687
rect 2815 653 2849 673
rect 2815 605 2849 615
rect 2815 581 2849 605
rect 2815 537 2849 543
rect 2815 509 2849 537
rect 2815 469 2849 471
rect 2815 437 2849 469
rect 2815 367 2849 399
rect 2815 365 2849 367
rect 2815 299 2849 327
rect 2815 293 2849 299
rect 2815 231 2849 255
rect 2815 221 2849 231
rect 2815 163 2849 183
rect 2815 149 2849 163
rect 2933 673 2967 687
rect 2933 653 2967 673
rect 2933 605 2967 615
rect 2933 581 2967 605
rect 2933 537 2967 543
rect 2933 509 2967 537
rect 2933 469 2967 471
rect 2933 437 2967 469
rect 2933 367 2967 399
rect 2933 365 2967 367
rect 2933 299 2967 327
rect 2933 293 2967 299
rect 2933 231 2967 255
rect 2933 221 2967 231
rect 2933 163 2967 183
rect 2933 149 2967 163
rect -2908 37 -2874 71
rect -2790 37 -2756 71
rect -2672 37 -2638 71
rect -2554 37 -2520 71
rect -2436 37 -2402 71
rect -2318 37 -2284 71
rect -2200 37 -2166 71
rect -2082 37 -2048 71
rect -1964 37 -1930 71
rect -1846 37 -1812 71
rect -1728 37 -1694 71
rect -1610 37 -1576 71
rect -1492 37 -1458 71
rect -1374 37 -1340 71
rect -1256 37 -1222 71
rect -1138 37 -1104 71
rect -1020 37 -986 71
rect -902 37 -868 71
rect -784 37 -750 71
rect -666 37 -632 71
rect -548 37 -514 71
rect -430 37 -396 71
rect -312 37 -278 71
rect -194 37 -160 71
rect -76 37 -42 71
rect 42 37 76 71
rect 160 37 194 71
rect 278 37 312 71
rect 396 37 430 71
rect 514 37 548 71
rect 632 37 666 71
rect 750 37 784 71
rect 868 37 902 71
rect 986 37 1020 71
rect 1104 37 1138 71
rect 1222 37 1256 71
rect 1340 37 1374 71
rect 1458 37 1492 71
rect 1576 37 1610 71
rect 1694 37 1728 71
rect 1812 37 1846 71
rect 1930 37 1964 71
rect 2048 37 2082 71
rect 2166 37 2200 71
rect 2284 37 2318 71
rect 2402 37 2436 71
rect 2520 37 2554 71
rect 2638 37 2672 71
rect 2756 37 2790 71
rect 2874 37 2908 71
rect -2908 -71 -2874 -37
rect -2790 -71 -2756 -37
rect -2672 -71 -2638 -37
rect -2554 -71 -2520 -37
rect -2436 -71 -2402 -37
rect -2318 -71 -2284 -37
rect -2200 -71 -2166 -37
rect -2082 -71 -2048 -37
rect -1964 -71 -1930 -37
rect -1846 -71 -1812 -37
rect -1728 -71 -1694 -37
rect -1610 -71 -1576 -37
rect -1492 -71 -1458 -37
rect -1374 -71 -1340 -37
rect -1256 -71 -1222 -37
rect -1138 -71 -1104 -37
rect -1020 -71 -986 -37
rect -902 -71 -868 -37
rect -784 -71 -750 -37
rect -666 -71 -632 -37
rect -548 -71 -514 -37
rect -430 -71 -396 -37
rect -312 -71 -278 -37
rect -194 -71 -160 -37
rect -76 -71 -42 -37
rect 42 -71 76 -37
rect 160 -71 194 -37
rect 278 -71 312 -37
rect 396 -71 430 -37
rect 514 -71 548 -37
rect 632 -71 666 -37
rect 750 -71 784 -37
rect 868 -71 902 -37
rect 986 -71 1020 -37
rect 1104 -71 1138 -37
rect 1222 -71 1256 -37
rect 1340 -71 1374 -37
rect 1458 -71 1492 -37
rect 1576 -71 1610 -37
rect 1694 -71 1728 -37
rect 1812 -71 1846 -37
rect 1930 -71 1964 -37
rect 2048 -71 2082 -37
rect 2166 -71 2200 -37
rect 2284 -71 2318 -37
rect 2402 -71 2436 -37
rect 2520 -71 2554 -37
rect 2638 -71 2672 -37
rect 2756 -71 2790 -37
rect 2874 -71 2908 -37
rect -2967 -163 -2933 -149
rect -2967 -183 -2933 -163
rect -2967 -231 -2933 -221
rect -2967 -255 -2933 -231
rect -2967 -299 -2933 -293
rect -2967 -327 -2933 -299
rect -2967 -367 -2933 -365
rect -2967 -399 -2933 -367
rect -2967 -469 -2933 -437
rect -2967 -471 -2933 -469
rect -2967 -537 -2933 -509
rect -2967 -543 -2933 -537
rect -2967 -605 -2933 -581
rect -2967 -615 -2933 -605
rect -2967 -673 -2933 -653
rect -2967 -687 -2933 -673
rect -2849 -163 -2815 -149
rect -2849 -183 -2815 -163
rect -2849 -231 -2815 -221
rect -2849 -255 -2815 -231
rect -2849 -299 -2815 -293
rect -2849 -327 -2815 -299
rect -2849 -367 -2815 -365
rect -2849 -399 -2815 -367
rect -2849 -469 -2815 -437
rect -2849 -471 -2815 -469
rect -2849 -537 -2815 -509
rect -2849 -543 -2815 -537
rect -2849 -605 -2815 -581
rect -2849 -615 -2815 -605
rect -2849 -673 -2815 -653
rect -2849 -687 -2815 -673
rect -2731 -163 -2697 -149
rect -2731 -183 -2697 -163
rect -2731 -231 -2697 -221
rect -2731 -255 -2697 -231
rect -2731 -299 -2697 -293
rect -2731 -327 -2697 -299
rect -2731 -367 -2697 -365
rect -2731 -399 -2697 -367
rect -2731 -469 -2697 -437
rect -2731 -471 -2697 -469
rect -2731 -537 -2697 -509
rect -2731 -543 -2697 -537
rect -2731 -605 -2697 -581
rect -2731 -615 -2697 -605
rect -2731 -673 -2697 -653
rect -2731 -687 -2697 -673
rect -2613 -163 -2579 -149
rect -2613 -183 -2579 -163
rect -2613 -231 -2579 -221
rect -2613 -255 -2579 -231
rect -2613 -299 -2579 -293
rect -2613 -327 -2579 -299
rect -2613 -367 -2579 -365
rect -2613 -399 -2579 -367
rect -2613 -469 -2579 -437
rect -2613 -471 -2579 -469
rect -2613 -537 -2579 -509
rect -2613 -543 -2579 -537
rect -2613 -605 -2579 -581
rect -2613 -615 -2579 -605
rect -2613 -673 -2579 -653
rect -2613 -687 -2579 -673
rect -2495 -163 -2461 -149
rect -2495 -183 -2461 -163
rect -2495 -231 -2461 -221
rect -2495 -255 -2461 -231
rect -2495 -299 -2461 -293
rect -2495 -327 -2461 -299
rect -2495 -367 -2461 -365
rect -2495 -399 -2461 -367
rect -2495 -469 -2461 -437
rect -2495 -471 -2461 -469
rect -2495 -537 -2461 -509
rect -2495 -543 -2461 -537
rect -2495 -605 -2461 -581
rect -2495 -615 -2461 -605
rect -2495 -673 -2461 -653
rect -2495 -687 -2461 -673
rect -2377 -163 -2343 -149
rect -2377 -183 -2343 -163
rect -2377 -231 -2343 -221
rect -2377 -255 -2343 -231
rect -2377 -299 -2343 -293
rect -2377 -327 -2343 -299
rect -2377 -367 -2343 -365
rect -2377 -399 -2343 -367
rect -2377 -469 -2343 -437
rect -2377 -471 -2343 -469
rect -2377 -537 -2343 -509
rect -2377 -543 -2343 -537
rect -2377 -605 -2343 -581
rect -2377 -615 -2343 -605
rect -2377 -673 -2343 -653
rect -2377 -687 -2343 -673
rect -2259 -163 -2225 -149
rect -2259 -183 -2225 -163
rect -2259 -231 -2225 -221
rect -2259 -255 -2225 -231
rect -2259 -299 -2225 -293
rect -2259 -327 -2225 -299
rect -2259 -367 -2225 -365
rect -2259 -399 -2225 -367
rect -2259 -469 -2225 -437
rect -2259 -471 -2225 -469
rect -2259 -537 -2225 -509
rect -2259 -543 -2225 -537
rect -2259 -605 -2225 -581
rect -2259 -615 -2225 -605
rect -2259 -673 -2225 -653
rect -2259 -687 -2225 -673
rect -2141 -163 -2107 -149
rect -2141 -183 -2107 -163
rect -2141 -231 -2107 -221
rect -2141 -255 -2107 -231
rect -2141 -299 -2107 -293
rect -2141 -327 -2107 -299
rect -2141 -367 -2107 -365
rect -2141 -399 -2107 -367
rect -2141 -469 -2107 -437
rect -2141 -471 -2107 -469
rect -2141 -537 -2107 -509
rect -2141 -543 -2107 -537
rect -2141 -605 -2107 -581
rect -2141 -615 -2107 -605
rect -2141 -673 -2107 -653
rect -2141 -687 -2107 -673
rect -2023 -163 -1989 -149
rect -2023 -183 -1989 -163
rect -2023 -231 -1989 -221
rect -2023 -255 -1989 -231
rect -2023 -299 -1989 -293
rect -2023 -327 -1989 -299
rect -2023 -367 -1989 -365
rect -2023 -399 -1989 -367
rect -2023 -469 -1989 -437
rect -2023 -471 -1989 -469
rect -2023 -537 -1989 -509
rect -2023 -543 -1989 -537
rect -2023 -605 -1989 -581
rect -2023 -615 -1989 -605
rect -2023 -673 -1989 -653
rect -2023 -687 -1989 -673
rect -1905 -163 -1871 -149
rect -1905 -183 -1871 -163
rect -1905 -231 -1871 -221
rect -1905 -255 -1871 -231
rect -1905 -299 -1871 -293
rect -1905 -327 -1871 -299
rect -1905 -367 -1871 -365
rect -1905 -399 -1871 -367
rect -1905 -469 -1871 -437
rect -1905 -471 -1871 -469
rect -1905 -537 -1871 -509
rect -1905 -543 -1871 -537
rect -1905 -605 -1871 -581
rect -1905 -615 -1871 -605
rect -1905 -673 -1871 -653
rect -1905 -687 -1871 -673
rect -1787 -163 -1753 -149
rect -1787 -183 -1753 -163
rect -1787 -231 -1753 -221
rect -1787 -255 -1753 -231
rect -1787 -299 -1753 -293
rect -1787 -327 -1753 -299
rect -1787 -367 -1753 -365
rect -1787 -399 -1753 -367
rect -1787 -469 -1753 -437
rect -1787 -471 -1753 -469
rect -1787 -537 -1753 -509
rect -1787 -543 -1753 -537
rect -1787 -605 -1753 -581
rect -1787 -615 -1753 -605
rect -1787 -673 -1753 -653
rect -1787 -687 -1753 -673
rect -1669 -163 -1635 -149
rect -1669 -183 -1635 -163
rect -1669 -231 -1635 -221
rect -1669 -255 -1635 -231
rect -1669 -299 -1635 -293
rect -1669 -327 -1635 -299
rect -1669 -367 -1635 -365
rect -1669 -399 -1635 -367
rect -1669 -469 -1635 -437
rect -1669 -471 -1635 -469
rect -1669 -537 -1635 -509
rect -1669 -543 -1635 -537
rect -1669 -605 -1635 -581
rect -1669 -615 -1635 -605
rect -1669 -673 -1635 -653
rect -1669 -687 -1635 -673
rect -1551 -163 -1517 -149
rect -1551 -183 -1517 -163
rect -1551 -231 -1517 -221
rect -1551 -255 -1517 -231
rect -1551 -299 -1517 -293
rect -1551 -327 -1517 -299
rect -1551 -367 -1517 -365
rect -1551 -399 -1517 -367
rect -1551 -469 -1517 -437
rect -1551 -471 -1517 -469
rect -1551 -537 -1517 -509
rect -1551 -543 -1517 -537
rect -1551 -605 -1517 -581
rect -1551 -615 -1517 -605
rect -1551 -673 -1517 -653
rect -1551 -687 -1517 -673
rect -1433 -163 -1399 -149
rect -1433 -183 -1399 -163
rect -1433 -231 -1399 -221
rect -1433 -255 -1399 -231
rect -1433 -299 -1399 -293
rect -1433 -327 -1399 -299
rect -1433 -367 -1399 -365
rect -1433 -399 -1399 -367
rect -1433 -469 -1399 -437
rect -1433 -471 -1399 -469
rect -1433 -537 -1399 -509
rect -1433 -543 -1399 -537
rect -1433 -605 -1399 -581
rect -1433 -615 -1399 -605
rect -1433 -673 -1399 -653
rect -1433 -687 -1399 -673
rect -1315 -163 -1281 -149
rect -1315 -183 -1281 -163
rect -1315 -231 -1281 -221
rect -1315 -255 -1281 -231
rect -1315 -299 -1281 -293
rect -1315 -327 -1281 -299
rect -1315 -367 -1281 -365
rect -1315 -399 -1281 -367
rect -1315 -469 -1281 -437
rect -1315 -471 -1281 -469
rect -1315 -537 -1281 -509
rect -1315 -543 -1281 -537
rect -1315 -605 -1281 -581
rect -1315 -615 -1281 -605
rect -1315 -673 -1281 -653
rect -1315 -687 -1281 -673
rect -1197 -163 -1163 -149
rect -1197 -183 -1163 -163
rect -1197 -231 -1163 -221
rect -1197 -255 -1163 -231
rect -1197 -299 -1163 -293
rect -1197 -327 -1163 -299
rect -1197 -367 -1163 -365
rect -1197 -399 -1163 -367
rect -1197 -469 -1163 -437
rect -1197 -471 -1163 -469
rect -1197 -537 -1163 -509
rect -1197 -543 -1163 -537
rect -1197 -605 -1163 -581
rect -1197 -615 -1163 -605
rect -1197 -673 -1163 -653
rect -1197 -687 -1163 -673
rect -1079 -163 -1045 -149
rect -1079 -183 -1045 -163
rect -1079 -231 -1045 -221
rect -1079 -255 -1045 -231
rect -1079 -299 -1045 -293
rect -1079 -327 -1045 -299
rect -1079 -367 -1045 -365
rect -1079 -399 -1045 -367
rect -1079 -469 -1045 -437
rect -1079 -471 -1045 -469
rect -1079 -537 -1045 -509
rect -1079 -543 -1045 -537
rect -1079 -605 -1045 -581
rect -1079 -615 -1045 -605
rect -1079 -673 -1045 -653
rect -1079 -687 -1045 -673
rect -961 -163 -927 -149
rect -961 -183 -927 -163
rect -961 -231 -927 -221
rect -961 -255 -927 -231
rect -961 -299 -927 -293
rect -961 -327 -927 -299
rect -961 -367 -927 -365
rect -961 -399 -927 -367
rect -961 -469 -927 -437
rect -961 -471 -927 -469
rect -961 -537 -927 -509
rect -961 -543 -927 -537
rect -961 -605 -927 -581
rect -961 -615 -927 -605
rect -961 -673 -927 -653
rect -961 -687 -927 -673
rect -843 -163 -809 -149
rect -843 -183 -809 -163
rect -843 -231 -809 -221
rect -843 -255 -809 -231
rect -843 -299 -809 -293
rect -843 -327 -809 -299
rect -843 -367 -809 -365
rect -843 -399 -809 -367
rect -843 -469 -809 -437
rect -843 -471 -809 -469
rect -843 -537 -809 -509
rect -843 -543 -809 -537
rect -843 -605 -809 -581
rect -843 -615 -809 -605
rect -843 -673 -809 -653
rect -843 -687 -809 -673
rect -725 -163 -691 -149
rect -725 -183 -691 -163
rect -725 -231 -691 -221
rect -725 -255 -691 -231
rect -725 -299 -691 -293
rect -725 -327 -691 -299
rect -725 -367 -691 -365
rect -725 -399 -691 -367
rect -725 -469 -691 -437
rect -725 -471 -691 -469
rect -725 -537 -691 -509
rect -725 -543 -691 -537
rect -725 -605 -691 -581
rect -725 -615 -691 -605
rect -725 -673 -691 -653
rect -725 -687 -691 -673
rect -607 -163 -573 -149
rect -607 -183 -573 -163
rect -607 -231 -573 -221
rect -607 -255 -573 -231
rect -607 -299 -573 -293
rect -607 -327 -573 -299
rect -607 -367 -573 -365
rect -607 -399 -573 -367
rect -607 -469 -573 -437
rect -607 -471 -573 -469
rect -607 -537 -573 -509
rect -607 -543 -573 -537
rect -607 -605 -573 -581
rect -607 -615 -573 -605
rect -607 -673 -573 -653
rect -607 -687 -573 -673
rect -489 -163 -455 -149
rect -489 -183 -455 -163
rect -489 -231 -455 -221
rect -489 -255 -455 -231
rect -489 -299 -455 -293
rect -489 -327 -455 -299
rect -489 -367 -455 -365
rect -489 -399 -455 -367
rect -489 -469 -455 -437
rect -489 -471 -455 -469
rect -489 -537 -455 -509
rect -489 -543 -455 -537
rect -489 -605 -455 -581
rect -489 -615 -455 -605
rect -489 -673 -455 -653
rect -489 -687 -455 -673
rect -371 -163 -337 -149
rect -371 -183 -337 -163
rect -371 -231 -337 -221
rect -371 -255 -337 -231
rect -371 -299 -337 -293
rect -371 -327 -337 -299
rect -371 -367 -337 -365
rect -371 -399 -337 -367
rect -371 -469 -337 -437
rect -371 -471 -337 -469
rect -371 -537 -337 -509
rect -371 -543 -337 -537
rect -371 -605 -337 -581
rect -371 -615 -337 -605
rect -371 -673 -337 -653
rect -371 -687 -337 -673
rect -253 -163 -219 -149
rect -253 -183 -219 -163
rect -253 -231 -219 -221
rect -253 -255 -219 -231
rect -253 -299 -219 -293
rect -253 -327 -219 -299
rect -253 -367 -219 -365
rect -253 -399 -219 -367
rect -253 -469 -219 -437
rect -253 -471 -219 -469
rect -253 -537 -219 -509
rect -253 -543 -219 -537
rect -253 -605 -219 -581
rect -253 -615 -219 -605
rect -253 -673 -219 -653
rect -253 -687 -219 -673
rect -135 -163 -101 -149
rect -135 -183 -101 -163
rect -135 -231 -101 -221
rect -135 -255 -101 -231
rect -135 -299 -101 -293
rect -135 -327 -101 -299
rect -135 -367 -101 -365
rect -135 -399 -101 -367
rect -135 -469 -101 -437
rect -135 -471 -101 -469
rect -135 -537 -101 -509
rect -135 -543 -101 -537
rect -135 -605 -101 -581
rect -135 -615 -101 -605
rect -135 -673 -101 -653
rect -135 -687 -101 -673
rect -17 -163 17 -149
rect -17 -183 17 -163
rect -17 -231 17 -221
rect -17 -255 17 -231
rect -17 -299 17 -293
rect -17 -327 17 -299
rect -17 -367 17 -365
rect -17 -399 17 -367
rect -17 -469 17 -437
rect -17 -471 17 -469
rect -17 -537 17 -509
rect -17 -543 17 -537
rect -17 -605 17 -581
rect -17 -615 17 -605
rect -17 -673 17 -653
rect -17 -687 17 -673
rect 101 -163 135 -149
rect 101 -183 135 -163
rect 101 -231 135 -221
rect 101 -255 135 -231
rect 101 -299 135 -293
rect 101 -327 135 -299
rect 101 -367 135 -365
rect 101 -399 135 -367
rect 101 -469 135 -437
rect 101 -471 135 -469
rect 101 -537 135 -509
rect 101 -543 135 -537
rect 101 -605 135 -581
rect 101 -615 135 -605
rect 101 -673 135 -653
rect 101 -687 135 -673
rect 219 -163 253 -149
rect 219 -183 253 -163
rect 219 -231 253 -221
rect 219 -255 253 -231
rect 219 -299 253 -293
rect 219 -327 253 -299
rect 219 -367 253 -365
rect 219 -399 253 -367
rect 219 -469 253 -437
rect 219 -471 253 -469
rect 219 -537 253 -509
rect 219 -543 253 -537
rect 219 -605 253 -581
rect 219 -615 253 -605
rect 219 -673 253 -653
rect 219 -687 253 -673
rect 337 -163 371 -149
rect 337 -183 371 -163
rect 337 -231 371 -221
rect 337 -255 371 -231
rect 337 -299 371 -293
rect 337 -327 371 -299
rect 337 -367 371 -365
rect 337 -399 371 -367
rect 337 -469 371 -437
rect 337 -471 371 -469
rect 337 -537 371 -509
rect 337 -543 371 -537
rect 337 -605 371 -581
rect 337 -615 371 -605
rect 337 -673 371 -653
rect 337 -687 371 -673
rect 455 -163 489 -149
rect 455 -183 489 -163
rect 455 -231 489 -221
rect 455 -255 489 -231
rect 455 -299 489 -293
rect 455 -327 489 -299
rect 455 -367 489 -365
rect 455 -399 489 -367
rect 455 -469 489 -437
rect 455 -471 489 -469
rect 455 -537 489 -509
rect 455 -543 489 -537
rect 455 -605 489 -581
rect 455 -615 489 -605
rect 455 -673 489 -653
rect 455 -687 489 -673
rect 573 -163 607 -149
rect 573 -183 607 -163
rect 573 -231 607 -221
rect 573 -255 607 -231
rect 573 -299 607 -293
rect 573 -327 607 -299
rect 573 -367 607 -365
rect 573 -399 607 -367
rect 573 -469 607 -437
rect 573 -471 607 -469
rect 573 -537 607 -509
rect 573 -543 607 -537
rect 573 -605 607 -581
rect 573 -615 607 -605
rect 573 -673 607 -653
rect 573 -687 607 -673
rect 691 -163 725 -149
rect 691 -183 725 -163
rect 691 -231 725 -221
rect 691 -255 725 -231
rect 691 -299 725 -293
rect 691 -327 725 -299
rect 691 -367 725 -365
rect 691 -399 725 -367
rect 691 -469 725 -437
rect 691 -471 725 -469
rect 691 -537 725 -509
rect 691 -543 725 -537
rect 691 -605 725 -581
rect 691 -615 725 -605
rect 691 -673 725 -653
rect 691 -687 725 -673
rect 809 -163 843 -149
rect 809 -183 843 -163
rect 809 -231 843 -221
rect 809 -255 843 -231
rect 809 -299 843 -293
rect 809 -327 843 -299
rect 809 -367 843 -365
rect 809 -399 843 -367
rect 809 -469 843 -437
rect 809 -471 843 -469
rect 809 -537 843 -509
rect 809 -543 843 -537
rect 809 -605 843 -581
rect 809 -615 843 -605
rect 809 -673 843 -653
rect 809 -687 843 -673
rect 927 -163 961 -149
rect 927 -183 961 -163
rect 927 -231 961 -221
rect 927 -255 961 -231
rect 927 -299 961 -293
rect 927 -327 961 -299
rect 927 -367 961 -365
rect 927 -399 961 -367
rect 927 -469 961 -437
rect 927 -471 961 -469
rect 927 -537 961 -509
rect 927 -543 961 -537
rect 927 -605 961 -581
rect 927 -615 961 -605
rect 927 -673 961 -653
rect 927 -687 961 -673
rect 1045 -163 1079 -149
rect 1045 -183 1079 -163
rect 1045 -231 1079 -221
rect 1045 -255 1079 -231
rect 1045 -299 1079 -293
rect 1045 -327 1079 -299
rect 1045 -367 1079 -365
rect 1045 -399 1079 -367
rect 1045 -469 1079 -437
rect 1045 -471 1079 -469
rect 1045 -537 1079 -509
rect 1045 -543 1079 -537
rect 1045 -605 1079 -581
rect 1045 -615 1079 -605
rect 1045 -673 1079 -653
rect 1045 -687 1079 -673
rect 1163 -163 1197 -149
rect 1163 -183 1197 -163
rect 1163 -231 1197 -221
rect 1163 -255 1197 -231
rect 1163 -299 1197 -293
rect 1163 -327 1197 -299
rect 1163 -367 1197 -365
rect 1163 -399 1197 -367
rect 1163 -469 1197 -437
rect 1163 -471 1197 -469
rect 1163 -537 1197 -509
rect 1163 -543 1197 -537
rect 1163 -605 1197 -581
rect 1163 -615 1197 -605
rect 1163 -673 1197 -653
rect 1163 -687 1197 -673
rect 1281 -163 1315 -149
rect 1281 -183 1315 -163
rect 1281 -231 1315 -221
rect 1281 -255 1315 -231
rect 1281 -299 1315 -293
rect 1281 -327 1315 -299
rect 1281 -367 1315 -365
rect 1281 -399 1315 -367
rect 1281 -469 1315 -437
rect 1281 -471 1315 -469
rect 1281 -537 1315 -509
rect 1281 -543 1315 -537
rect 1281 -605 1315 -581
rect 1281 -615 1315 -605
rect 1281 -673 1315 -653
rect 1281 -687 1315 -673
rect 1399 -163 1433 -149
rect 1399 -183 1433 -163
rect 1399 -231 1433 -221
rect 1399 -255 1433 -231
rect 1399 -299 1433 -293
rect 1399 -327 1433 -299
rect 1399 -367 1433 -365
rect 1399 -399 1433 -367
rect 1399 -469 1433 -437
rect 1399 -471 1433 -469
rect 1399 -537 1433 -509
rect 1399 -543 1433 -537
rect 1399 -605 1433 -581
rect 1399 -615 1433 -605
rect 1399 -673 1433 -653
rect 1399 -687 1433 -673
rect 1517 -163 1551 -149
rect 1517 -183 1551 -163
rect 1517 -231 1551 -221
rect 1517 -255 1551 -231
rect 1517 -299 1551 -293
rect 1517 -327 1551 -299
rect 1517 -367 1551 -365
rect 1517 -399 1551 -367
rect 1517 -469 1551 -437
rect 1517 -471 1551 -469
rect 1517 -537 1551 -509
rect 1517 -543 1551 -537
rect 1517 -605 1551 -581
rect 1517 -615 1551 -605
rect 1517 -673 1551 -653
rect 1517 -687 1551 -673
rect 1635 -163 1669 -149
rect 1635 -183 1669 -163
rect 1635 -231 1669 -221
rect 1635 -255 1669 -231
rect 1635 -299 1669 -293
rect 1635 -327 1669 -299
rect 1635 -367 1669 -365
rect 1635 -399 1669 -367
rect 1635 -469 1669 -437
rect 1635 -471 1669 -469
rect 1635 -537 1669 -509
rect 1635 -543 1669 -537
rect 1635 -605 1669 -581
rect 1635 -615 1669 -605
rect 1635 -673 1669 -653
rect 1635 -687 1669 -673
rect 1753 -163 1787 -149
rect 1753 -183 1787 -163
rect 1753 -231 1787 -221
rect 1753 -255 1787 -231
rect 1753 -299 1787 -293
rect 1753 -327 1787 -299
rect 1753 -367 1787 -365
rect 1753 -399 1787 -367
rect 1753 -469 1787 -437
rect 1753 -471 1787 -469
rect 1753 -537 1787 -509
rect 1753 -543 1787 -537
rect 1753 -605 1787 -581
rect 1753 -615 1787 -605
rect 1753 -673 1787 -653
rect 1753 -687 1787 -673
rect 1871 -163 1905 -149
rect 1871 -183 1905 -163
rect 1871 -231 1905 -221
rect 1871 -255 1905 -231
rect 1871 -299 1905 -293
rect 1871 -327 1905 -299
rect 1871 -367 1905 -365
rect 1871 -399 1905 -367
rect 1871 -469 1905 -437
rect 1871 -471 1905 -469
rect 1871 -537 1905 -509
rect 1871 -543 1905 -537
rect 1871 -605 1905 -581
rect 1871 -615 1905 -605
rect 1871 -673 1905 -653
rect 1871 -687 1905 -673
rect 1989 -163 2023 -149
rect 1989 -183 2023 -163
rect 1989 -231 2023 -221
rect 1989 -255 2023 -231
rect 1989 -299 2023 -293
rect 1989 -327 2023 -299
rect 1989 -367 2023 -365
rect 1989 -399 2023 -367
rect 1989 -469 2023 -437
rect 1989 -471 2023 -469
rect 1989 -537 2023 -509
rect 1989 -543 2023 -537
rect 1989 -605 2023 -581
rect 1989 -615 2023 -605
rect 1989 -673 2023 -653
rect 1989 -687 2023 -673
rect 2107 -163 2141 -149
rect 2107 -183 2141 -163
rect 2107 -231 2141 -221
rect 2107 -255 2141 -231
rect 2107 -299 2141 -293
rect 2107 -327 2141 -299
rect 2107 -367 2141 -365
rect 2107 -399 2141 -367
rect 2107 -469 2141 -437
rect 2107 -471 2141 -469
rect 2107 -537 2141 -509
rect 2107 -543 2141 -537
rect 2107 -605 2141 -581
rect 2107 -615 2141 -605
rect 2107 -673 2141 -653
rect 2107 -687 2141 -673
rect 2225 -163 2259 -149
rect 2225 -183 2259 -163
rect 2225 -231 2259 -221
rect 2225 -255 2259 -231
rect 2225 -299 2259 -293
rect 2225 -327 2259 -299
rect 2225 -367 2259 -365
rect 2225 -399 2259 -367
rect 2225 -469 2259 -437
rect 2225 -471 2259 -469
rect 2225 -537 2259 -509
rect 2225 -543 2259 -537
rect 2225 -605 2259 -581
rect 2225 -615 2259 -605
rect 2225 -673 2259 -653
rect 2225 -687 2259 -673
rect 2343 -163 2377 -149
rect 2343 -183 2377 -163
rect 2343 -231 2377 -221
rect 2343 -255 2377 -231
rect 2343 -299 2377 -293
rect 2343 -327 2377 -299
rect 2343 -367 2377 -365
rect 2343 -399 2377 -367
rect 2343 -469 2377 -437
rect 2343 -471 2377 -469
rect 2343 -537 2377 -509
rect 2343 -543 2377 -537
rect 2343 -605 2377 -581
rect 2343 -615 2377 -605
rect 2343 -673 2377 -653
rect 2343 -687 2377 -673
rect 2461 -163 2495 -149
rect 2461 -183 2495 -163
rect 2461 -231 2495 -221
rect 2461 -255 2495 -231
rect 2461 -299 2495 -293
rect 2461 -327 2495 -299
rect 2461 -367 2495 -365
rect 2461 -399 2495 -367
rect 2461 -469 2495 -437
rect 2461 -471 2495 -469
rect 2461 -537 2495 -509
rect 2461 -543 2495 -537
rect 2461 -605 2495 -581
rect 2461 -615 2495 -605
rect 2461 -673 2495 -653
rect 2461 -687 2495 -673
rect 2579 -163 2613 -149
rect 2579 -183 2613 -163
rect 2579 -231 2613 -221
rect 2579 -255 2613 -231
rect 2579 -299 2613 -293
rect 2579 -327 2613 -299
rect 2579 -367 2613 -365
rect 2579 -399 2613 -367
rect 2579 -469 2613 -437
rect 2579 -471 2613 -469
rect 2579 -537 2613 -509
rect 2579 -543 2613 -537
rect 2579 -605 2613 -581
rect 2579 -615 2613 -605
rect 2579 -673 2613 -653
rect 2579 -687 2613 -673
rect 2697 -163 2731 -149
rect 2697 -183 2731 -163
rect 2697 -231 2731 -221
rect 2697 -255 2731 -231
rect 2697 -299 2731 -293
rect 2697 -327 2731 -299
rect 2697 -367 2731 -365
rect 2697 -399 2731 -367
rect 2697 -469 2731 -437
rect 2697 -471 2731 -469
rect 2697 -537 2731 -509
rect 2697 -543 2731 -537
rect 2697 -605 2731 -581
rect 2697 -615 2731 -605
rect 2697 -673 2731 -653
rect 2697 -687 2731 -673
rect 2815 -163 2849 -149
rect 2815 -183 2849 -163
rect 2815 -231 2849 -221
rect 2815 -255 2849 -231
rect 2815 -299 2849 -293
rect 2815 -327 2849 -299
rect 2815 -367 2849 -365
rect 2815 -399 2849 -367
rect 2815 -469 2849 -437
rect 2815 -471 2849 -469
rect 2815 -537 2849 -509
rect 2815 -543 2849 -537
rect 2815 -605 2849 -581
rect 2815 -615 2849 -605
rect 2815 -673 2849 -653
rect 2815 -687 2849 -673
rect 2933 -163 2967 -149
rect 2933 -183 2967 -163
rect 2933 -231 2967 -221
rect 2933 -255 2967 -231
rect 2933 -299 2967 -293
rect 2933 -327 2967 -299
rect 2933 -367 2967 -365
rect 2933 -399 2967 -367
rect 2933 -469 2967 -437
rect 2933 -471 2967 -469
rect 2933 -537 2967 -509
rect 2933 -543 2967 -537
rect 2933 -605 2967 -581
rect 2933 -615 2967 -605
rect 2933 -673 2967 -653
rect 2933 -687 2967 -673
<< metal1 >>
rect -2973 687 -2927 718
rect -2973 653 -2967 687
rect -2933 653 -2927 687
rect -2973 615 -2927 653
rect -2973 581 -2967 615
rect -2933 581 -2927 615
rect -2973 543 -2927 581
rect -2973 509 -2967 543
rect -2933 509 -2927 543
rect -2973 471 -2927 509
rect -2973 437 -2967 471
rect -2933 437 -2927 471
rect -2973 399 -2927 437
rect -2973 365 -2967 399
rect -2933 365 -2927 399
rect -2973 327 -2927 365
rect -2973 293 -2967 327
rect -2933 293 -2927 327
rect -2973 255 -2927 293
rect -2973 221 -2967 255
rect -2933 221 -2927 255
rect -2973 183 -2927 221
rect -2973 149 -2967 183
rect -2933 149 -2927 183
rect -2973 118 -2927 149
rect -2855 687 -2809 718
rect -2855 653 -2849 687
rect -2815 653 -2809 687
rect -2855 615 -2809 653
rect -2855 581 -2849 615
rect -2815 581 -2809 615
rect -2855 543 -2809 581
rect -2855 509 -2849 543
rect -2815 509 -2809 543
rect -2855 471 -2809 509
rect -2855 437 -2849 471
rect -2815 437 -2809 471
rect -2855 399 -2809 437
rect -2855 365 -2849 399
rect -2815 365 -2809 399
rect -2855 327 -2809 365
rect -2855 293 -2849 327
rect -2815 293 -2809 327
rect -2855 255 -2809 293
rect -2855 221 -2849 255
rect -2815 221 -2809 255
rect -2855 183 -2809 221
rect -2855 149 -2849 183
rect -2815 149 -2809 183
rect -2855 118 -2809 149
rect -2737 687 -2691 718
rect -2737 653 -2731 687
rect -2697 653 -2691 687
rect -2737 615 -2691 653
rect -2737 581 -2731 615
rect -2697 581 -2691 615
rect -2737 543 -2691 581
rect -2737 509 -2731 543
rect -2697 509 -2691 543
rect -2737 471 -2691 509
rect -2737 437 -2731 471
rect -2697 437 -2691 471
rect -2737 399 -2691 437
rect -2737 365 -2731 399
rect -2697 365 -2691 399
rect -2737 327 -2691 365
rect -2737 293 -2731 327
rect -2697 293 -2691 327
rect -2737 255 -2691 293
rect -2737 221 -2731 255
rect -2697 221 -2691 255
rect -2737 183 -2691 221
rect -2737 149 -2731 183
rect -2697 149 -2691 183
rect -2737 118 -2691 149
rect -2619 687 -2573 718
rect -2619 653 -2613 687
rect -2579 653 -2573 687
rect -2619 615 -2573 653
rect -2619 581 -2613 615
rect -2579 581 -2573 615
rect -2619 543 -2573 581
rect -2619 509 -2613 543
rect -2579 509 -2573 543
rect -2619 471 -2573 509
rect -2619 437 -2613 471
rect -2579 437 -2573 471
rect -2619 399 -2573 437
rect -2619 365 -2613 399
rect -2579 365 -2573 399
rect -2619 327 -2573 365
rect -2619 293 -2613 327
rect -2579 293 -2573 327
rect -2619 255 -2573 293
rect -2619 221 -2613 255
rect -2579 221 -2573 255
rect -2619 183 -2573 221
rect -2619 149 -2613 183
rect -2579 149 -2573 183
rect -2619 118 -2573 149
rect -2501 687 -2455 718
rect -2501 653 -2495 687
rect -2461 653 -2455 687
rect -2501 615 -2455 653
rect -2501 581 -2495 615
rect -2461 581 -2455 615
rect -2501 543 -2455 581
rect -2501 509 -2495 543
rect -2461 509 -2455 543
rect -2501 471 -2455 509
rect -2501 437 -2495 471
rect -2461 437 -2455 471
rect -2501 399 -2455 437
rect -2501 365 -2495 399
rect -2461 365 -2455 399
rect -2501 327 -2455 365
rect -2501 293 -2495 327
rect -2461 293 -2455 327
rect -2501 255 -2455 293
rect -2501 221 -2495 255
rect -2461 221 -2455 255
rect -2501 183 -2455 221
rect -2501 149 -2495 183
rect -2461 149 -2455 183
rect -2501 118 -2455 149
rect -2383 687 -2337 718
rect -2383 653 -2377 687
rect -2343 653 -2337 687
rect -2383 615 -2337 653
rect -2383 581 -2377 615
rect -2343 581 -2337 615
rect -2383 543 -2337 581
rect -2383 509 -2377 543
rect -2343 509 -2337 543
rect -2383 471 -2337 509
rect -2383 437 -2377 471
rect -2343 437 -2337 471
rect -2383 399 -2337 437
rect -2383 365 -2377 399
rect -2343 365 -2337 399
rect -2383 327 -2337 365
rect -2383 293 -2377 327
rect -2343 293 -2337 327
rect -2383 255 -2337 293
rect -2383 221 -2377 255
rect -2343 221 -2337 255
rect -2383 183 -2337 221
rect -2383 149 -2377 183
rect -2343 149 -2337 183
rect -2383 118 -2337 149
rect -2265 687 -2219 718
rect -2265 653 -2259 687
rect -2225 653 -2219 687
rect -2265 615 -2219 653
rect -2265 581 -2259 615
rect -2225 581 -2219 615
rect -2265 543 -2219 581
rect -2265 509 -2259 543
rect -2225 509 -2219 543
rect -2265 471 -2219 509
rect -2265 437 -2259 471
rect -2225 437 -2219 471
rect -2265 399 -2219 437
rect -2265 365 -2259 399
rect -2225 365 -2219 399
rect -2265 327 -2219 365
rect -2265 293 -2259 327
rect -2225 293 -2219 327
rect -2265 255 -2219 293
rect -2265 221 -2259 255
rect -2225 221 -2219 255
rect -2265 183 -2219 221
rect -2265 149 -2259 183
rect -2225 149 -2219 183
rect -2265 118 -2219 149
rect -2147 687 -2101 718
rect -2147 653 -2141 687
rect -2107 653 -2101 687
rect -2147 615 -2101 653
rect -2147 581 -2141 615
rect -2107 581 -2101 615
rect -2147 543 -2101 581
rect -2147 509 -2141 543
rect -2107 509 -2101 543
rect -2147 471 -2101 509
rect -2147 437 -2141 471
rect -2107 437 -2101 471
rect -2147 399 -2101 437
rect -2147 365 -2141 399
rect -2107 365 -2101 399
rect -2147 327 -2101 365
rect -2147 293 -2141 327
rect -2107 293 -2101 327
rect -2147 255 -2101 293
rect -2147 221 -2141 255
rect -2107 221 -2101 255
rect -2147 183 -2101 221
rect -2147 149 -2141 183
rect -2107 149 -2101 183
rect -2147 118 -2101 149
rect -2029 687 -1983 718
rect -2029 653 -2023 687
rect -1989 653 -1983 687
rect -2029 615 -1983 653
rect -2029 581 -2023 615
rect -1989 581 -1983 615
rect -2029 543 -1983 581
rect -2029 509 -2023 543
rect -1989 509 -1983 543
rect -2029 471 -1983 509
rect -2029 437 -2023 471
rect -1989 437 -1983 471
rect -2029 399 -1983 437
rect -2029 365 -2023 399
rect -1989 365 -1983 399
rect -2029 327 -1983 365
rect -2029 293 -2023 327
rect -1989 293 -1983 327
rect -2029 255 -1983 293
rect -2029 221 -2023 255
rect -1989 221 -1983 255
rect -2029 183 -1983 221
rect -2029 149 -2023 183
rect -1989 149 -1983 183
rect -2029 118 -1983 149
rect -1911 687 -1865 718
rect -1911 653 -1905 687
rect -1871 653 -1865 687
rect -1911 615 -1865 653
rect -1911 581 -1905 615
rect -1871 581 -1865 615
rect -1911 543 -1865 581
rect -1911 509 -1905 543
rect -1871 509 -1865 543
rect -1911 471 -1865 509
rect -1911 437 -1905 471
rect -1871 437 -1865 471
rect -1911 399 -1865 437
rect -1911 365 -1905 399
rect -1871 365 -1865 399
rect -1911 327 -1865 365
rect -1911 293 -1905 327
rect -1871 293 -1865 327
rect -1911 255 -1865 293
rect -1911 221 -1905 255
rect -1871 221 -1865 255
rect -1911 183 -1865 221
rect -1911 149 -1905 183
rect -1871 149 -1865 183
rect -1911 118 -1865 149
rect -1793 687 -1747 718
rect -1793 653 -1787 687
rect -1753 653 -1747 687
rect -1793 615 -1747 653
rect -1793 581 -1787 615
rect -1753 581 -1747 615
rect -1793 543 -1747 581
rect -1793 509 -1787 543
rect -1753 509 -1747 543
rect -1793 471 -1747 509
rect -1793 437 -1787 471
rect -1753 437 -1747 471
rect -1793 399 -1747 437
rect -1793 365 -1787 399
rect -1753 365 -1747 399
rect -1793 327 -1747 365
rect -1793 293 -1787 327
rect -1753 293 -1747 327
rect -1793 255 -1747 293
rect -1793 221 -1787 255
rect -1753 221 -1747 255
rect -1793 183 -1747 221
rect -1793 149 -1787 183
rect -1753 149 -1747 183
rect -1793 118 -1747 149
rect -1675 687 -1629 718
rect -1675 653 -1669 687
rect -1635 653 -1629 687
rect -1675 615 -1629 653
rect -1675 581 -1669 615
rect -1635 581 -1629 615
rect -1675 543 -1629 581
rect -1675 509 -1669 543
rect -1635 509 -1629 543
rect -1675 471 -1629 509
rect -1675 437 -1669 471
rect -1635 437 -1629 471
rect -1675 399 -1629 437
rect -1675 365 -1669 399
rect -1635 365 -1629 399
rect -1675 327 -1629 365
rect -1675 293 -1669 327
rect -1635 293 -1629 327
rect -1675 255 -1629 293
rect -1675 221 -1669 255
rect -1635 221 -1629 255
rect -1675 183 -1629 221
rect -1675 149 -1669 183
rect -1635 149 -1629 183
rect -1675 118 -1629 149
rect -1557 687 -1511 718
rect -1557 653 -1551 687
rect -1517 653 -1511 687
rect -1557 615 -1511 653
rect -1557 581 -1551 615
rect -1517 581 -1511 615
rect -1557 543 -1511 581
rect -1557 509 -1551 543
rect -1517 509 -1511 543
rect -1557 471 -1511 509
rect -1557 437 -1551 471
rect -1517 437 -1511 471
rect -1557 399 -1511 437
rect -1557 365 -1551 399
rect -1517 365 -1511 399
rect -1557 327 -1511 365
rect -1557 293 -1551 327
rect -1517 293 -1511 327
rect -1557 255 -1511 293
rect -1557 221 -1551 255
rect -1517 221 -1511 255
rect -1557 183 -1511 221
rect -1557 149 -1551 183
rect -1517 149 -1511 183
rect -1557 118 -1511 149
rect -1439 687 -1393 718
rect -1439 653 -1433 687
rect -1399 653 -1393 687
rect -1439 615 -1393 653
rect -1439 581 -1433 615
rect -1399 581 -1393 615
rect -1439 543 -1393 581
rect -1439 509 -1433 543
rect -1399 509 -1393 543
rect -1439 471 -1393 509
rect -1439 437 -1433 471
rect -1399 437 -1393 471
rect -1439 399 -1393 437
rect -1439 365 -1433 399
rect -1399 365 -1393 399
rect -1439 327 -1393 365
rect -1439 293 -1433 327
rect -1399 293 -1393 327
rect -1439 255 -1393 293
rect -1439 221 -1433 255
rect -1399 221 -1393 255
rect -1439 183 -1393 221
rect -1439 149 -1433 183
rect -1399 149 -1393 183
rect -1439 118 -1393 149
rect -1321 687 -1275 718
rect -1321 653 -1315 687
rect -1281 653 -1275 687
rect -1321 615 -1275 653
rect -1321 581 -1315 615
rect -1281 581 -1275 615
rect -1321 543 -1275 581
rect -1321 509 -1315 543
rect -1281 509 -1275 543
rect -1321 471 -1275 509
rect -1321 437 -1315 471
rect -1281 437 -1275 471
rect -1321 399 -1275 437
rect -1321 365 -1315 399
rect -1281 365 -1275 399
rect -1321 327 -1275 365
rect -1321 293 -1315 327
rect -1281 293 -1275 327
rect -1321 255 -1275 293
rect -1321 221 -1315 255
rect -1281 221 -1275 255
rect -1321 183 -1275 221
rect -1321 149 -1315 183
rect -1281 149 -1275 183
rect -1321 118 -1275 149
rect -1203 687 -1157 718
rect -1203 653 -1197 687
rect -1163 653 -1157 687
rect -1203 615 -1157 653
rect -1203 581 -1197 615
rect -1163 581 -1157 615
rect -1203 543 -1157 581
rect -1203 509 -1197 543
rect -1163 509 -1157 543
rect -1203 471 -1157 509
rect -1203 437 -1197 471
rect -1163 437 -1157 471
rect -1203 399 -1157 437
rect -1203 365 -1197 399
rect -1163 365 -1157 399
rect -1203 327 -1157 365
rect -1203 293 -1197 327
rect -1163 293 -1157 327
rect -1203 255 -1157 293
rect -1203 221 -1197 255
rect -1163 221 -1157 255
rect -1203 183 -1157 221
rect -1203 149 -1197 183
rect -1163 149 -1157 183
rect -1203 118 -1157 149
rect -1085 687 -1039 718
rect -1085 653 -1079 687
rect -1045 653 -1039 687
rect -1085 615 -1039 653
rect -1085 581 -1079 615
rect -1045 581 -1039 615
rect -1085 543 -1039 581
rect -1085 509 -1079 543
rect -1045 509 -1039 543
rect -1085 471 -1039 509
rect -1085 437 -1079 471
rect -1045 437 -1039 471
rect -1085 399 -1039 437
rect -1085 365 -1079 399
rect -1045 365 -1039 399
rect -1085 327 -1039 365
rect -1085 293 -1079 327
rect -1045 293 -1039 327
rect -1085 255 -1039 293
rect -1085 221 -1079 255
rect -1045 221 -1039 255
rect -1085 183 -1039 221
rect -1085 149 -1079 183
rect -1045 149 -1039 183
rect -1085 118 -1039 149
rect -967 687 -921 718
rect -967 653 -961 687
rect -927 653 -921 687
rect -967 615 -921 653
rect -967 581 -961 615
rect -927 581 -921 615
rect -967 543 -921 581
rect -967 509 -961 543
rect -927 509 -921 543
rect -967 471 -921 509
rect -967 437 -961 471
rect -927 437 -921 471
rect -967 399 -921 437
rect -967 365 -961 399
rect -927 365 -921 399
rect -967 327 -921 365
rect -967 293 -961 327
rect -927 293 -921 327
rect -967 255 -921 293
rect -967 221 -961 255
rect -927 221 -921 255
rect -967 183 -921 221
rect -967 149 -961 183
rect -927 149 -921 183
rect -967 118 -921 149
rect -849 687 -803 718
rect -849 653 -843 687
rect -809 653 -803 687
rect -849 615 -803 653
rect -849 581 -843 615
rect -809 581 -803 615
rect -849 543 -803 581
rect -849 509 -843 543
rect -809 509 -803 543
rect -849 471 -803 509
rect -849 437 -843 471
rect -809 437 -803 471
rect -849 399 -803 437
rect -849 365 -843 399
rect -809 365 -803 399
rect -849 327 -803 365
rect -849 293 -843 327
rect -809 293 -803 327
rect -849 255 -803 293
rect -849 221 -843 255
rect -809 221 -803 255
rect -849 183 -803 221
rect -849 149 -843 183
rect -809 149 -803 183
rect -849 118 -803 149
rect -731 687 -685 718
rect -731 653 -725 687
rect -691 653 -685 687
rect -731 615 -685 653
rect -731 581 -725 615
rect -691 581 -685 615
rect -731 543 -685 581
rect -731 509 -725 543
rect -691 509 -685 543
rect -731 471 -685 509
rect -731 437 -725 471
rect -691 437 -685 471
rect -731 399 -685 437
rect -731 365 -725 399
rect -691 365 -685 399
rect -731 327 -685 365
rect -731 293 -725 327
rect -691 293 -685 327
rect -731 255 -685 293
rect -731 221 -725 255
rect -691 221 -685 255
rect -731 183 -685 221
rect -731 149 -725 183
rect -691 149 -685 183
rect -731 118 -685 149
rect -613 687 -567 718
rect -613 653 -607 687
rect -573 653 -567 687
rect -613 615 -567 653
rect -613 581 -607 615
rect -573 581 -567 615
rect -613 543 -567 581
rect -613 509 -607 543
rect -573 509 -567 543
rect -613 471 -567 509
rect -613 437 -607 471
rect -573 437 -567 471
rect -613 399 -567 437
rect -613 365 -607 399
rect -573 365 -567 399
rect -613 327 -567 365
rect -613 293 -607 327
rect -573 293 -567 327
rect -613 255 -567 293
rect -613 221 -607 255
rect -573 221 -567 255
rect -613 183 -567 221
rect -613 149 -607 183
rect -573 149 -567 183
rect -613 118 -567 149
rect -495 687 -449 718
rect -495 653 -489 687
rect -455 653 -449 687
rect -495 615 -449 653
rect -495 581 -489 615
rect -455 581 -449 615
rect -495 543 -449 581
rect -495 509 -489 543
rect -455 509 -449 543
rect -495 471 -449 509
rect -495 437 -489 471
rect -455 437 -449 471
rect -495 399 -449 437
rect -495 365 -489 399
rect -455 365 -449 399
rect -495 327 -449 365
rect -495 293 -489 327
rect -455 293 -449 327
rect -495 255 -449 293
rect -495 221 -489 255
rect -455 221 -449 255
rect -495 183 -449 221
rect -495 149 -489 183
rect -455 149 -449 183
rect -495 118 -449 149
rect -377 687 -331 718
rect -377 653 -371 687
rect -337 653 -331 687
rect -377 615 -331 653
rect -377 581 -371 615
rect -337 581 -331 615
rect -377 543 -331 581
rect -377 509 -371 543
rect -337 509 -331 543
rect -377 471 -331 509
rect -377 437 -371 471
rect -337 437 -331 471
rect -377 399 -331 437
rect -377 365 -371 399
rect -337 365 -331 399
rect -377 327 -331 365
rect -377 293 -371 327
rect -337 293 -331 327
rect -377 255 -331 293
rect -377 221 -371 255
rect -337 221 -331 255
rect -377 183 -331 221
rect -377 149 -371 183
rect -337 149 -331 183
rect -377 118 -331 149
rect -259 687 -213 718
rect -259 653 -253 687
rect -219 653 -213 687
rect -259 615 -213 653
rect -259 581 -253 615
rect -219 581 -213 615
rect -259 543 -213 581
rect -259 509 -253 543
rect -219 509 -213 543
rect -259 471 -213 509
rect -259 437 -253 471
rect -219 437 -213 471
rect -259 399 -213 437
rect -259 365 -253 399
rect -219 365 -213 399
rect -259 327 -213 365
rect -259 293 -253 327
rect -219 293 -213 327
rect -259 255 -213 293
rect -259 221 -253 255
rect -219 221 -213 255
rect -259 183 -213 221
rect -259 149 -253 183
rect -219 149 -213 183
rect -259 118 -213 149
rect -141 687 -95 718
rect -141 653 -135 687
rect -101 653 -95 687
rect -141 615 -95 653
rect -141 581 -135 615
rect -101 581 -95 615
rect -141 543 -95 581
rect -141 509 -135 543
rect -101 509 -95 543
rect -141 471 -95 509
rect -141 437 -135 471
rect -101 437 -95 471
rect -141 399 -95 437
rect -141 365 -135 399
rect -101 365 -95 399
rect -141 327 -95 365
rect -141 293 -135 327
rect -101 293 -95 327
rect -141 255 -95 293
rect -141 221 -135 255
rect -101 221 -95 255
rect -141 183 -95 221
rect -141 149 -135 183
rect -101 149 -95 183
rect -141 118 -95 149
rect -23 687 23 718
rect -23 653 -17 687
rect 17 653 23 687
rect -23 615 23 653
rect -23 581 -17 615
rect 17 581 23 615
rect -23 543 23 581
rect -23 509 -17 543
rect 17 509 23 543
rect -23 471 23 509
rect -23 437 -17 471
rect 17 437 23 471
rect -23 399 23 437
rect -23 365 -17 399
rect 17 365 23 399
rect -23 327 23 365
rect -23 293 -17 327
rect 17 293 23 327
rect -23 255 23 293
rect -23 221 -17 255
rect 17 221 23 255
rect -23 183 23 221
rect -23 149 -17 183
rect 17 149 23 183
rect -23 118 23 149
rect 95 687 141 718
rect 95 653 101 687
rect 135 653 141 687
rect 95 615 141 653
rect 95 581 101 615
rect 135 581 141 615
rect 95 543 141 581
rect 95 509 101 543
rect 135 509 141 543
rect 95 471 141 509
rect 95 437 101 471
rect 135 437 141 471
rect 95 399 141 437
rect 95 365 101 399
rect 135 365 141 399
rect 95 327 141 365
rect 95 293 101 327
rect 135 293 141 327
rect 95 255 141 293
rect 95 221 101 255
rect 135 221 141 255
rect 95 183 141 221
rect 95 149 101 183
rect 135 149 141 183
rect 95 118 141 149
rect 213 687 259 718
rect 213 653 219 687
rect 253 653 259 687
rect 213 615 259 653
rect 213 581 219 615
rect 253 581 259 615
rect 213 543 259 581
rect 213 509 219 543
rect 253 509 259 543
rect 213 471 259 509
rect 213 437 219 471
rect 253 437 259 471
rect 213 399 259 437
rect 213 365 219 399
rect 253 365 259 399
rect 213 327 259 365
rect 213 293 219 327
rect 253 293 259 327
rect 213 255 259 293
rect 213 221 219 255
rect 253 221 259 255
rect 213 183 259 221
rect 213 149 219 183
rect 253 149 259 183
rect 213 118 259 149
rect 331 687 377 718
rect 331 653 337 687
rect 371 653 377 687
rect 331 615 377 653
rect 331 581 337 615
rect 371 581 377 615
rect 331 543 377 581
rect 331 509 337 543
rect 371 509 377 543
rect 331 471 377 509
rect 331 437 337 471
rect 371 437 377 471
rect 331 399 377 437
rect 331 365 337 399
rect 371 365 377 399
rect 331 327 377 365
rect 331 293 337 327
rect 371 293 377 327
rect 331 255 377 293
rect 331 221 337 255
rect 371 221 377 255
rect 331 183 377 221
rect 331 149 337 183
rect 371 149 377 183
rect 331 118 377 149
rect 449 687 495 718
rect 449 653 455 687
rect 489 653 495 687
rect 449 615 495 653
rect 449 581 455 615
rect 489 581 495 615
rect 449 543 495 581
rect 449 509 455 543
rect 489 509 495 543
rect 449 471 495 509
rect 449 437 455 471
rect 489 437 495 471
rect 449 399 495 437
rect 449 365 455 399
rect 489 365 495 399
rect 449 327 495 365
rect 449 293 455 327
rect 489 293 495 327
rect 449 255 495 293
rect 449 221 455 255
rect 489 221 495 255
rect 449 183 495 221
rect 449 149 455 183
rect 489 149 495 183
rect 449 118 495 149
rect 567 687 613 718
rect 567 653 573 687
rect 607 653 613 687
rect 567 615 613 653
rect 567 581 573 615
rect 607 581 613 615
rect 567 543 613 581
rect 567 509 573 543
rect 607 509 613 543
rect 567 471 613 509
rect 567 437 573 471
rect 607 437 613 471
rect 567 399 613 437
rect 567 365 573 399
rect 607 365 613 399
rect 567 327 613 365
rect 567 293 573 327
rect 607 293 613 327
rect 567 255 613 293
rect 567 221 573 255
rect 607 221 613 255
rect 567 183 613 221
rect 567 149 573 183
rect 607 149 613 183
rect 567 118 613 149
rect 685 687 731 718
rect 685 653 691 687
rect 725 653 731 687
rect 685 615 731 653
rect 685 581 691 615
rect 725 581 731 615
rect 685 543 731 581
rect 685 509 691 543
rect 725 509 731 543
rect 685 471 731 509
rect 685 437 691 471
rect 725 437 731 471
rect 685 399 731 437
rect 685 365 691 399
rect 725 365 731 399
rect 685 327 731 365
rect 685 293 691 327
rect 725 293 731 327
rect 685 255 731 293
rect 685 221 691 255
rect 725 221 731 255
rect 685 183 731 221
rect 685 149 691 183
rect 725 149 731 183
rect 685 118 731 149
rect 803 687 849 718
rect 803 653 809 687
rect 843 653 849 687
rect 803 615 849 653
rect 803 581 809 615
rect 843 581 849 615
rect 803 543 849 581
rect 803 509 809 543
rect 843 509 849 543
rect 803 471 849 509
rect 803 437 809 471
rect 843 437 849 471
rect 803 399 849 437
rect 803 365 809 399
rect 843 365 849 399
rect 803 327 849 365
rect 803 293 809 327
rect 843 293 849 327
rect 803 255 849 293
rect 803 221 809 255
rect 843 221 849 255
rect 803 183 849 221
rect 803 149 809 183
rect 843 149 849 183
rect 803 118 849 149
rect 921 687 967 718
rect 921 653 927 687
rect 961 653 967 687
rect 921 615 967 653
rect 921 581 927 615
rect 961 581 967 615
rect 921 543 967 581
rect 921 509 927 543
rect 961 509 967 543
rect 921 471 967 509
rect 921 437 927 471
rect 961 437 967 471
rect 921 399 967 437
rect 921 365 927 399
rect 961 365 967 399
rect 921 327 967 365
rect 921 293 927 327
rect 961 293 967 327
rect 921 255 967 293
rect 921 221 927 255
rect 961 221 967 255
rect 921 183 967 221
rect 921 149 927 183
rect 961 149 967 183
rect 921 118 967 149
rect 1039 687 1085 718
rect 1039 653 1045 687
rect 1079 653 1085 687
rect 1039 615 1085 653
rect 1039 581 1045 615
rect 1079 581 1085 615
rect 1039 543 1085 581
rect 1039 509 1045 543
rect 1079 509 1085 543
rect 1039 471 1085 509
rect 1039 437 1045 471
rect 1079 437 1085 471
rect 1039 399 1085 437
rect 1039 365 1045 399
rect 1079 365 1085 399
rect 1039 327 1085 365
rect 1039 293 1045 327
rect 1079 293 1085 327
rect 1039 255 1085 293
rect 1039 221 1045 255
rect 1079 221 1085 255
rect 1039 183 1085 221
rect 1039 149 1045 183
rect 1079 149 1085 183
rect 1039 118 1085 149
rect 1157 687 1203 718
rect 1157 653 1163 687
rect 1197 653 1203 687
rect 1157 615 1203 653
rect 1157 581 1163 615
rect 1197 581 1203 615
rect 1157 543 1203 581
rect 1157 509 1163 543
rect 1197 509 1203 543
rect 1157 471 1203 509
rect 1157 437 1163 471
rect 1197 437 1203 471
rect 1157 399 1203 437
rect 1157 365 1163 399
rect 1197 365 1203 399
rect 1157 327 1203 365
rect 1157 293 1163 327
rect 1197 293 1203 327
rect 1157 255 1203 293
rect 1157 221 1163 255
rect 1197 221 1203 255
rect 1157 183 1203 221
rect 1157 149 1163 183
rect 1197 149 1203 183
rect 1157 118 1203 149
rect 1275 687 1321 718
rect 1275 653 1281 687
rect 1315 653 1321 687
rect 1275 615 1321 653
rect 1275 581 1281 615
rect 1315 581 1321 615
rect 1275 543 1321 581
rect 1275 509 1281 543
rect 1315 509 1321 543
rect 1275 471 1321 509
rect 1275 437 1281 471
rect 1315 437 1321 471
rect 1275 399 1321 437
rect 1275 365 1281 399
rect 1315 365 1321 399
rect 1275 327 1321 365
rect 1275 293 1281 327
rect 1315 293 1321 327
rect 1275 255 1321 293
rect 1275 221 1281 255
rect 1315 221 1321 255
rect 1275 183 1321 221
rect 1275 149 1281 183
rect 1315 149 1321 183
rect 1275 118 1321 149
rect 1393 687 1439 718
rect 1393 653 1399 687
rect 1433 653 1439 687
rect 1393 615 1439 653
rect 1393 581 1399 615
rect 1433 581 1439 615
rect 1393 543 1439 581
rect 1393 509 1399 543
rect 1433 509 1439 543
rect 1393 471 1439 509
rect 1393 437 1399 471
rect 1433 437 1439 471
rect 1393 399 1439 437
rect 1393 365 1399 399
rect 1433 365 1439 399
rect 1393 327 1439 365
rect 1393 293 1399 327
rect 1433 293 1439 327
rect 1393 255 1439 293
rect 1393 221 1399 255
rect 1433 221 1439 255
rect 1393 183 1439 221
rect 1393 149 1399 183
rect 1433 149 1439 183
rect 1393 118 1439 149
rect 1511 687 1557 718
rect 1511 653 1517 687
rect 1551 653 1557 687
rect 1511 615 1557 653
rect 1511 581 1517 615
rect 1551 581 1557 615
rect 1511 543 1557 581
rect 1511 509 1517 543
rect 1551 509 1557 543
rect 1511 471 1557 509
rect 1511 437 1517 471
rect 1551 437 1557 471
rect 1511 399 1557 437
rect 1511 365 1517 399
rect 1551 365 1557 399
rect 1511 327 1557 365
rect 1511 293 1517 327
rect 1551 293 1557 327
rect 1511 255 1557 293
rect 1511 221 1517 255
rect 1551 221 1557 255
rect 1511 183 1557 221
rect 1511 149 1517 183
rect 1551 149 1557 183
rect 1511 118 1557 149
rect 1629 687 1675 718
rect 1629 653 1635 687
rect 1669 653 1675 687
rect 1629 615 1675 653
rect 1629 581 1635 615
rect 1669 581 1675 615
rect 1629 543 1675 581
rect 1629 509 1635 543
rect 1669 509 1675 543
rect 1629 471 1675 509
rect 1629 437 1635 471
rect 1669 437 1675 471
rect 1629 399 1675 437
rect 1629 365 1635 399
rect 1669 365 1675 399
rect 1629 327 1675 365
rect 1629 293 1635 327
rect 1669 293 1675 327
rect 1629 255 1675 293
rect 1629 221 1635 255
rect 1669 221 1675 255
rect 1629 183 1675 221
rect 1629 149 1635 183
rect 1669 149 1675 183
rect 1629 118 1675 149
rect 1747 687 1793 718
rect 1747 653 1753 687
rect 1787 653 1793 687
rect 1747 615 1793 653
rect 1747 581 1753 615
rect 1787 581 1793 615
rect 1747 543 1793 581
rect 1747 509 1753 543
rect 1787 509 1793 543
rect 1747 471 1793 509
rect 1747 437 1753 471
rect 1787 437 1793 471
rect 1747 399 1793 437
rect 1747 365 1753 399
rect 1787 365 1793 399
rect 1747 327 1793 365
rect 1747 293 1753 327
rect 1787 293 1793 327
rect 1747 255 1793 293
rect 1747 221 1753 255
rect 1787 221 1793 255
rect 1747 183 1793 221
rect 1747 149 1753 183
rect 1787 149 1793 183
rect 1747 118 1793 149
rect 1865 687 1911 718
rect 1865 653 1871 687
rect 1905 653 1911 687
rect 1865 615 1911 653
rect 1865 581 1871 615
rect 1905 581 1911 615
rect 1865 543 1911 581
rect 1865 509 1871 543
rect 1905 509 1911 543
rect 1865 471 1911 509
rect 1865 437 1871 471
rect 1905 437 1911 471
rect 1865 399 1911 437
rect 1865 365 1871 399
rect 1905 365 1911 399
rect 1865 327 1911 365
rect 1865 293 1871 327
rect 1905 293 1911 327
rect 1865 255 1911 293
rect 1865 221 1871 255
rect 1905 221 1911 255
rect 1865 183 1911 221
rect 1865 149 1871 183
rect 1905 149 1911 183
rect 1865 118 1911 149
rect 1983 687 2029 718
rect 1983 653 1989 687
rect 2023 653 2029 687
rect 1983 615 2029 653
rect 1983 581 1989 615
rect 2023 581 2029 615
rect 1983 543 2029 581
rect 1983 509 1989 543
rect 2023 509 2029 543
rect 1983 471 2029 509
rect 1983 437 1989 471
rect 2023 437 2029 471
rect 1983 399 2029 437
rect 1983 365 1989 399
rect 2023 365 2029 399
rect 1983 327 2029 365
rect 1983 293 1989 327
rect 2023 293 2029 327
rect 1983 255 2029 293
rect 1983 221 1989 255
rect 2023 221 2029 255
rect 1983 183 2029 221
rect 1983 149 1989 183
rect 2023 149 2029 183
rect 1983 118 2029 149
rect 2101 687 2147 718
rect 2101 653 2107 687
rect 2141 653 2147 687
rect 2101 615 2147 653
rect 2101 581 2107 615
rect 2141 581 2147 615
rect 2101 543 2147 581
rect 2101 509 2107 543
rect 2141 509 2147 543
rect 2101 471 2147 509
rect 2101 437 2107 471
rect 2141 437 2147 471
rect 2101 399 2147 437
rect 2101 365 2107 399
rect 2141 365 2147 399
rect 2101 327 2147 365
rect 2101 293 2107 327
rect 2141 293 2147 327
rect 2101 255 2147 293
rect 2101 221 2107 255
rect 2141 221 2147 255
rect 2101 183 2147 221
rect 2101 149 2107 183
rect 2141 149 2147 183
rect 2101 118 2147 149
rect 2219 687 2265 718
rect 2219 653 2225 687
rect 2259 653 2265 687
rect 2219 615 2265 653
rect 2219 581 2225 615
rect 2259 581 2265 615
rect 2219 543 2265 581
rect 2219 509 2225 543
rect 2259 509 2265 543
rect 2219 471 2265 509
rect 2219 437 2225 471
rect 2259 437 2265 471
rect 2219 399 2265 437
rect 2219 365 2225 399
rect 2259 365 2265 399
rect 2219 327 2265 365
rect 2219 293 2225 327
rect 2259 293 2265 327
rect 2219 255 2265 293
rect 2219 221 2225 255
rect 2259 221 2265 255
rect 2219 183 2265 221
rect 2219 149 2225 183
rect 2259 149 2265 183
rect 2219 118 2265 149
rect 2337 687 2383 718
rect 2337 653 2343 687
rect 2377 653 2383 687
rect 2337 615 2383 653
rect 2337 581 2343 615
rect 2377 581 2383 615
rect 2337 543 2383 581
rect 2337 509 2343 543
rect 2377 509 2383 543
rect 2337 471 2383 509
rect 2337 437 2343 471
rect 2377 437 2383 471
rect 2337 399 2383 437
rect 2337 365 2343 399
rect 2377 365 2383 399
rect 2337 327 2383 365
rect 2337 293 2343 327
rect 2377 293 2383 327
rect 2337 255 2383 293
rect 2337 221 2343 255
rect 2377 221 2383 255
rect 2337 183 2383 221
rect 2337 149 2343 183
rect 2377 149 2383 183
rect 2337 118 2383 149
rect 2455 687 2501 718
rect 2455 653 2461 687
rect 2495 653 2501 687
rect 2455 615 2501 653
rect 2455 581 2461 615
rect 2495 581 2501 615
rect 2455 543 2501 581
rect 2455 509 2461 543
rect 2495 509 2501 543
rect 2455 471 2501 509
rect 2455 437 2461 471
rect 2495 437 2501 471
rect 2455 399 2501 437
rect 2455 365 2461 399
rect 2495 365 2501 399
rect 2455 327 2501 365
rect 2455 293 2461 327
rect 2495 293 2501 327
rect 2455 255 2501 293
rect 2455 221 2461 255
rect 2495 221 2501 255
rect 2455 183 2501 221
rect 2455 149 2461 183
rect 2495 149 2501 183
rect 2455 118 2501 149
rect 2573 687 2619 718
rect 2573 653 2579 687
rect 2613 653 2619 687
rect 2573 615 2619 653
rect 2573 581 2579 615
rect 2613 581 2619 615
rect 2573 543 2619 581
rect 2573 509 2579 543
rect 2613 509 2619 543
rect 2573 471 2619 509
rect 2573 437 2579 471
rect 2613 437 2619 471
rect 2573 399 2619 437
rect 2573 365 2579 399
rect 2613 365 2619 399
rect 2573 327 2619 365
rect 2573 293 2579 327
rect 2613 293 2619 327
rect 2573 255 2619 293
rect 2573 221 2579 255
rect 2613 221 2619 255
rect 2573 183 2619 221
rect 2573 149 2579 183
rect 2613 149 2619 183
rect 2573 118 2619 149
rect 2691 687 2737 718
rect 2691 653 2697 687
rect 2731 653 2737 687
rect 2691 615 2737 653
rect 2691 581 2697 615
rect 2731 581 2737 615
rect 2691 543 2737 581
rect 2691 509 2697 543
rect 2731 509 2737 543
rect 2691 471 2737 509
rect 2691 437 2697 471
rect 2731 437 2737 471
rect 2691 399 2737 437
rect 2691 365 2697 399
rect 2731 365 2737 399
rect 2691 327 2737 365
rect 2691 293 2697 327
rect 2731 293 2737 327
rect 2691 255 2737 293
rect 2691 221 2697 255
rect 2731 221 2737 255
rect 2691 183 2737 221
rect 2691 149 2697 183
rect 2731 149 2737 183
rect 2691 118 2737 149
rect 2809 687 2855 718
rect 2809 653 2815 687
rect 2849 653 2855 687
rect 2809 615 2855 653
rect 2809 581 2815 615
rect 2849 581 2855 615
rect 2809 543 2855 581
rect 2809 509 2815 543
rect 2849 509 2855 543
rect 2809 471 2855 509
rect 2809 437 2815 471
rect 2849 437 2855 471
rect 2809 399 2855 437
rect 2809 365 2815 399
rect 2849 365 2855 399
rect 2809 327 2855 365
rect 2809 293 2815 327
rect 2849 293 2855 327
rect 2809 255 2855 293
rect 2809 221 2815 255
rect 2849 221 2855 255
rect 2809 183 2855 221
rect 2809 149 2815 183
rect 2849 149 2855 183
rect 2809 118 2855 149
rect 2927 687 2973 718
rect 2927 653 2933 687
rect 2967 653 2973 687
rect 2927 615 2973 653
rect 2927 581 2933 615
rect 2967 581 2973 615
rect 2927 543 2973 581
rect 2927 509 2933 543
rect 2967 509 2973 543
rect 2927 471 2973 509
rect 2927 437 2933 471
rect 2967 437 2973 471
rect 2927 399 2973 437
rect 2927 365 2933 399
rect 2967 365 2973 399
rect 2927 327 2973 365
rect 2927 293 2933 327
rect 2967 293 2973 327
rect 2927 255 2973 293
rect 2927 221 2933 255
rect 2967 221 2973 255
rect 2927 183 2973 221
rect 2927 149 2933 183
rect 2967 149 2973 183
rect 2927 118 2973 149
rect -2920 71 -2862 77
rect -2920 37 -2908 71
rect -2874 37 -2862 71
rect -2920 31 -2862 37
rect -2802 71 -2744 77
rect -2802 37 -2790 71
rect -2756 37 -2744 71
rect -2802 31 -2744 37
rect -2684 71 -2626 77
rect -2684 37 -2672 71
rect -2638 37 -2626 71
rect -2684 31 -2626 37
rect -2566 71 -2508 77
rect -2566 37 -2554 71
rect -2520 37 -2508 71
rect -2566 31 -2508 37
rect -2448 71 -2390 77
rect -2448 37 -2436 71
rect -2402 37 -2390 71
rect -2448 31 -2390 37
rect -2330 71 -2272 77
rect -2330 37 -2318 71
rect -2284 37 -2272 71
rect -2330 31 -2272 37
rect -2212 71 -2154 77
rect -2212 37 -2200 71
rect -2166 37 -2154 71
rect -2212 31 -2154 37
rect -2094 71 -2036 77
rect -2094 37 -2082 71
rect -2048 37 -2036 71
rect -2094 31 -2036 37
rect -1976 71 -1918 77
rect -1976 37 -1964 71
rect -1930 37 -1918 71
rect -1976 31 -1918 37
rect -1858 71 -1800 77
rect -1858 37 -1846 71
rect -1812 37 -1800 71
rect -1858 31 -1800 37
rect -1740 71 -1682 77
rect -1740 37 -1728 71
rect -1694 37 -1682 71
rect -1740 31 -1682 37
rect -1622 71 -1564 77
rect -1622 37 -1610 71
rect -1576 37 -1564 71
rect -1622 31 -1564 37
rect -1504 71 -1446 77
rect -1504 37 -1492 71
rect -1458 37 -1446 71
rect -1504 31 -1446 37
rect -1386 71 -1328 77
rect -1386 37 -1374 71
rect -1340 37 -1328 71
rect -1386 31 -1328 37
rect -1268 71 -1210 77
rect -1268 37 -1256 71
rect -1222 37 -1210 71
rect -1268 31 -1210 37
rect -1150 71 -1092 77
rect -1150 37 -1138 71
rect -1104 37 -1092 71
rect -1150 31 -1092 37
rect -1032 71 -974 77
rect -1032 37 -1020 71
rect -986 37 -974 71
rect -1032 31 -974 37
rect -914 71 -856 77
rect -914 37 -902 71
rect -868 37 -856 71
rect -914 31 -856 37
rect -796 71 -738 77
rect -796 37 -784 71
rect -750 37 -738 71
rect -796 31 -738 37
rect -678 71 -620 77
rect -678 37 -666 71
rect -632 37 -620 71
rect -678 31 -620 37
rect -560 71 -502 77
rect -560 37 -548 71
rect -514 37 -502 71
rect -560 31 -502 37
rect -442 71 -384 77
rect -442 37 -430 71
rect -396 37 -384 71
rect -442 31 -384 37
rect -324 71 -266 77
rect -324 37 -312 71
rect -278 37 -266 71
rect -324 31 -266 37
rect -206 71 -148 77
rect -206 37 -194 71
rect -160 37 -148 71
rect -206 31 -148 37
rect -88 71 -30 77
rect -88 37 -76 71
rect -42 37 -30 71
rect -88 31 -30 37
rect 30 71 88 77
rect 30 37 42 71
rect 76 37 88 71
rect 30 31 88 37
rect 148 71 206 77
rect 148 37 160 71
rect 194 37 206 71
rect 148 31 206 37
rect 266 71 324 77
rect 266 37 278 71
rect 312 37 324 71
rect 266 31 324 37
rect 384 71 442 77
rect 384 37 396 71
rect 430 37 442 71
rect 384 31 442 37
rect 502 71 560 77
rect 502 37 514 71
rect 548 37 560 71
rect 502 31 560 37
rect 620 71 678 77
rect 620 37 632 71
rect 666 37 678 71
rect 620 31 678 37
rect 738 71 796 77
rect 738 37 750 71
rect 784 37 796 71
rect 738 31 796 37
rect 856 71 914 77
rect 856 37 868 71
rect 902 37 914 71
rect 856 31 914 37
rect 974 71 1032 77
rect 974 37 986 71
rect 1020 37 1032 71
rect 974 31 1032 37
rect 1092 71 1150 77
rect 1092 37 1104 71
rect 1138 37 1150 71
rect 1092 31 1150 37
rect 1210 71 1268 77
rect 1210 37 1222 71
rect 1256 37 1268 71
rect 1210 31 1268 37
rect 1328 71 1386 77
rect 1328 37 1340 71
rect 1374 37 1386 71
rect 1328 31 1386 37
rect 1446 71 1504 77
rect 1446 37 1458 71
rect 1492 37 1504 71
rect 1446 31 1504 37
rect 1564 71 1622 77
rect 1564 37 1576 71
rect 1610 37 1622 71
rect 1564 31 1622 37
rect 1682 71 1740 77
rect 1682 37 1694 71
rect 1728 37 1740 71
rect 1682 31 1740 37
rect 1800 71 1858 77
rect 1800 37 1812 71
rect 1846 37 1858 71
rect 1800 31 1858 37
rect 1918 71 1976 77
rect 1918 37 1930 71
rect 1964 37 1976 71
rect 1918 31 1976 37
rect 2036 71 2094 77
rect 2036 37 2048 71
rect 2082 37 2094 71
rect 2036 31 2094 37
rect 2154 71 2212 77
rect 2154 37 2166 71
rect 2200 37 2212 71
rect 2154 31 2212 37
rect 2272 71 2330 77
rect 2272 37 2284 71
rect 2318 37 2330 71
rect 2272 31 2330 37
rect 2390 71 2448 77
rect 2390 37 2402 71
rect 2436 37 2448 71
rect 2390 31 2448 37
rect 2508 71 2566 77
rect 2508 37 2520 71
rect 2554 37 2566 71
rect 2508 31 2566 37
rect 2626 71 2684 77
rect 2626 37 2638 71
rect 2672 37 2684 71
rect 2626 31 2684 37
rect 2744 71 2802 77
rect 2744 37 2756 71
rect 2790 37 2802 71
rect 2744 31 2802 37
rect 2862 71 2920 77
rect 2862 37 2874 71
rect 2908 37 2920 71
rect 2862 31 2920 37
rect -2920 -37 -2862 -31
rect -2920 -71 -2908 -37
rect -2874 -71 -2862 -37
rect -2920 -77 -2862 -71
rect -2802 -37 -2744 -31
rect -2802 -71 -2790 -37
rect -2756 -71 -2744 -37
rect -2802 -77 -2744 -71
rect -2684 -37 -2626 -31
rect -2684 -71 -2672 -37
rect -2638 -71 -2626 -37
rect -2684 -77 -2626 -71
rect -2566 -37 -2508 -31
rect -2566 -71 -2554 -37
rect -2520 -71 -2508 -37
rect -2566 -77 -2508 -71
rect -2448 -37 -2390 -31
rect -2448 -71 -2436 -37
rect -2402 -71 -2390 -37
rect -2448 -77 -2390 -71
rect -2330 -37 -2272 -31
rect -2330 -71 -2318 -37
rect -2284 -71 -2272 -37
rect -2330 -77 -2272 -71
rect -2212 -37 -2154 -31
rect -2212 -71 -2200 -37
rect -2166 -71 -2154 -37
rect -2212 -77 -2154 -71
rect -2094 -37 -2036 -31
rect -2094 -71 -2082 -37
rect -2048 -71 -2036 -37
rect -2094 -77 -2036 -71
rect -1976 -37 -1918 -31
rect -1976 -71 -1964 -37
rect -1930 -71 -1918 -37
rect -1976 -77 -1918 -71
rect -1858 -37 -1800 -31
rect -1858 -71 -1846 -37
rect -1812 -71 -1800 -37
rect -1858 -77 -1800 -71
rect -1740 -37 -1682 -31
rect -1740 -71 -1728 -37
rect -1694 -71 -1682 -37
rect -1740 -77 -1682 -71
rect -1622 -37 -1564 -31
rect -1622 -71 -1610 -37
rect -1576 -71 -1564 -37
rect -1622 -77 -1564 -71
rect -1504 -37 -1446 -31
rect -1504 -71 -1492 -37
rect -1458 -71 -1446 -37
rect -1504 -77 -1446 -71
rect -1386 -37 -1328 -31
rect -1386 -71 -1374 -37
rect -1340 -71 -1328 -37
rect -1386 -77 -1328 -71
rect -1268 -37 -1210 -31
rect -1268 -71 -1256 -37
rect -1222 -71 -1210 -37
rect -1268 -77 -1210 -71
rect -1150 -37 -1092 -31
rect -1150 -71 -1138 -37
rect -1104 -71 -1092 -37
rect -1150 -77 -1092 -71
rect -1032 -37 -974 -31
rect -1032 -71 -1020 -37
rect -986 -71 -974 -37
rect -1032 -77 -974 -71
rect -914 -37 -856 -31
rect -914 -71 -902 -37
rect -868 -71 -856 -37
rect -914 -77 -856 -71
rect -796 -37 -738 -31
rect -796 -71 -784 -37
rect -750 -71 -738 -37
rect -796 -77 -738 -71
rect -678 -37 -620 -31
rect -678 -71 -666 -37
rect -632 -71 -620 -37
rect -678 -77 -620 -71
rect -560 -37 -502 -31
rect -560 -71 -548 -37
rect -514 -71 -502 -37
rect -560 -77 -502 -71
rect -442 -37 -384 -31
rect -442 -71 -430 -37
rect -396 -71 -384 -37
rect -442 -77 -384 -71
rect -324 -37 -266 -31
rect -324 -71 -312 -37
rect -278 -71 -266 -37
rect -324 -77 -266 -71
rect -206 -37 -148 -31
rect -206 -71 -194 -37
rect -160 -71 -148 -37
rect -206 -77 -148 -71
rect -88 -37 -30 -31
rect -88 -71 -76 -37
rect -42 -71 -30 -37
rect -88 -77 -30 -71
rect 30 -37 88 -31
rect 30 -71 42 -37
rect 76 -71 88 -37
rect 30 -77 88 -71
rect 148 -37 206 -31
rect 148 -71 160 -37
rect 194 -71 206 -37
rect 148 -77 206 -71
rect 266 -37 324 -31
rect 266 -71 278 -37
rect 312 -71 324 -37
rect 266 -77 324 -71
rect 384 -37 442 -31
rect 384 -71 396 -37
rect 430 -71 442 -37
rect 384 -77 442 -71
rect 502 -37 560 -31
rect 502 -71 514 -37
rect 548 -71 560 -37
rect 502 -77 560 -71
rect 620 -37 678 -31
rect 620 -71 632 -37
rect 666 -71 678 -37
rect 620 -77 678 -71
rect 738 -37 796 -31
rect 738 -71 750 -37
rect 784 -71 796 -37
rect 738 -77 796 -71
rect 856 -37 914 -31
rect 856 -71 868 -37
rect 902 -71 914 -37
rect 856 -77 914 -71
rect 974 -37 1032 -31
rect 974 -71 986 -37
rect 1020 -71 1032 -37
rect 974 -77 1032 -71
rect 1092 -37 1150 -31
rect 1092 -71 1104 -37
rect 1138 -71 1150 -37
rect 1092 -77 1150 -71
rect 1210 -37 1268 -31
rect 1210 -71 1222 -37
rect 1256 -71 1268 -37
rect 1210 -77 1268 -71
rect 1328 -37 1386 -31
rect 1328 -71 1340 -37
rect 1374 -71 1386 -37
rect 1328 -77 1386 -71
rect 1446 -37 1504 -31
rect 1446 -71 1458 -37
rect 1492 -71 1504 -37
rect 1446 -77 1504 -71
rect 1564 -37 1622 -31
rect 1564 -71 1576 -37
rect 1610 -71 1622 -37
rect 1564 -77 1622 -71
rect 1682 -37 1740 -31
rect 1682 -71 1694 -37
rect 1728 -71 1740 -37
rect 1682 -77 1740 -71
rect 1800 -37 1858 -31
rect 1800 -71 1812 -37
rect 1846 -71 1858 -37
rect 1800 -77 1858 -71
rect 1918 -37 1976 -31
rect 1918 -71 1930 -37
rect 1964 -71 1976 -37
rect 1918 -77 1976 -71
rect 2036 -37 2094 -31
rect 2036 -71 2048 -37
rect 2082 -71 2094 -37
rect 2036 -77 2094 -71
rect 2154 -37 2212 -31
rect 2154 -71 2166 -37
rect 2200 -71 2212 -37
rect 2154 -77 2212 -71
rect 2272 -37 2330 -31
rect 2272 -71 2284 -37
rect 2318 -71 2330 -37
rect 2272 -77 2330 -71
rect 2390 -37 2448 -31
rect 2390 -71 2402 -37
rect 2436 -71 2448 -37
rect 2390 -77 2448 -71
rect 2508 -37 2566 -31
rect 2508 -71 2520 -37
rect 2554 -71 2566 -37
rect 2508 -77 2566 -71
rect 2626 -37 2684 -31
rect 2626 -71 2638 -37
rect 2672 -71 2684 -37
rect 2626 -77 2684 -71
rect 2744 -37 2802 -31
rect 2744 -71 2756 -37
rect 2790 -71 2802 -37
rect 2744 -77 2802 -71
rect 2862 -37 2920 -31
rect 2862 -71 2874 -37
rect 2908 -71 2920 -37
rect 2862 -77 2920 -71
rect -2973 -149 -2927 -118
rect -2973 -183 -2967 -149
rect -2933 -183 -2927 -149
rect -2973 -221 -2927 -183
rect -2973 -255 -2967 -221
rect -2933 -255 -2927 -221
rect -2973 -293 -2927 -255
rect -2973 -327 -2967 -293
rect -2933 -327 -2927 -293
rect -2973 -365 -2927 -327
rect -2973 -399 -2967 -365
rect -2933 -399 -2927 -365
rect -2973 -437 -2927 -399
rect -2973 -471 -2967 -437
rect -2933 -471 -2927 -437
rect -2973 -509 -2927 -471
rect -2973 -543 -2967 -509
rect -2933 -543 -2927 -509
rect -2973 -581 -2927 -543
rect -2973 -615 -2967 -581
rect -2933 -615 -2927 -581
rect -2973 -653 -2927 -615
rect -2973 -687 -2967 -653
rect -2933 -687 -2927 -653
rect -2973 -718 -2927 -687
rect -2855 -149 -2809 -118
rect -2855 -183 -2849 -149
rect -2815 -183 -2809 -149
rect -2855 -221 -2809 -183
rect -2855 -255 -2849 -221
rect -2815 -255 -2809 -221
rect -2855 -293 -2809 -255
rect -2855 -327 -2849 -293
rect -2815 -327 -2809 -293
rect -2855 -365 -2809 -327
rect -2855 -399 -2849 -365
rect -2815 -399 -2809 -365
rect -2855 -437 -2809 -399
rect -2855 -471 -2849 -437
rect -2815 -471 -2809 -437
rect -2855 -509 -2809 -471
rect -2855 -543 -2849 -509
rect -2815 -543 -2809 -509
rect -2855 -581 -2809 -543
rect -2855 -615 -2849 -581
rect -2815 -615 -2809 -581
rect -2855 -653 -2809 -615
rect -2855 -687 -2849 -653
rect -2815 -687 -2809 -653
rect -2855 -718 -2809 -687
rect -2737 -149 -2691 -118
rect -2737 -183 -2731 -149
rect -2697 -183 -2691 -149
rect -2737 -221 -2691 -183
rect -2737 -255 -2731 -221
rect -2697 -255 -2691 -221
rect -2737 -293 -2691 -255
rect -2737 -327 -2731 -293
rect -2697 -327 -2691 -293
rect -2737 -365 -2691 -327
rect -2737 -399 -2731 -365
rect -2697 -399 -2691 -365
rect -2737 -437 -2691 -399
rect -2737 -471 -2731 -437
rect -2697 -471 -2691 -437
rect -2737 -509 -2691 -471
rect -2737 -543 -2731 -509
rect -2697 -543 -2691 -509
rect -2737 -581 -2691 -543
rect -2737 -615 -2731 -581
rect -2697 -615 -2691 -581
rect -2737 -653 -2691 -615
rect -2737 -687 -2731 -653
rect -2697 -687 -2691 -653
rect -2737 -718 -2691 -687
rect -2619 -149 -2573 -118
rect -2619 -183 -2613 -149
rect -2579 -183 -2573 -149
rect -2619 -221 -2573 -183
rect -2619 -255 -2613 -221
rect -2579 -255 -2573 -221
rect -2619 -293 -2573 -255
rect -2619 -327 -2613 -293
rect -2579 -327 -2573 -293
rect -2619 -365 -2573 -327
rect -2619 -399 -2613 -365
rect -2579 -399 -2573 -365
rect -2619 -437 -2573 -399
rect -2619 -471 -2613 -437
rect -2579 -471 -2573 -437
rect -2619 -509 -2573 -471
rect -2619 -543 -2613 -509
rect -2579 -543 -2573 -509
rect -2619 -581 -2573 -543
rect -2619 -615 -2613 -581
rect -2579 -615 -2573 -581
rect -2619 -653 -2573 -615
rect -2619 -687 -2613 -653
rect -2579 -687 -2573 -653
rect -2619 -718 -2573 -687
rect -2501 -149 -2455 -118
rect -2501 -183 -2495 -149
rect -2461 -183 -2455 -149
rect -2501 -221 -2455 -183
rect -2501 -255 -2495 -221
rect -2461 -255 -2455 -221
rect -2501 -293 -2455 -255
rect -2501 -327 -2495 -293
rect -2461 -327 -2455 -293
rect -2501 -365 -2455 -327
rect -2501 -399 -2495 -365
rect -2461 -399 -2455 -365
rect -2501 -437 -2455 -399
rect -2501 -471 -2495 -437
rect -2461 -471 -2455 -437
rect -2501 -509 -2455 -471
rect -2501 -543 -2495 -509
rect -2461 -543 -2455 -509
rect -2501 -581 -2455 -543
rect -2501 -615 -2495 -581
rect -2461 -615 -2455 -581
rect -2501 -653 -2455 -615
rect -2501 -687 -2495 -653
rect -2461 -687 -2455 -653
rect -2501 -718 -2455 -687
rect -2383 -149 -2337 -118
rect -2383 -183 -2377 -149
rect -2343 -183 -2337 -149
rect -2383 -221 -2337 -183
rect -2383 -255 -2377 -221
rect -2343 -255 -2337 -221
rect -2383 -293 -2337 -255
rect -2383 -327 -2377 -293
rect -2343 -327 -2337 -293
rect -2383 -365 -2337 -327
rect -2383 -399 -2377 -365
rect -2343 -399 -2337 -365
rect -2383 -437 -2337 -399
rect -2383 -471 -2377 -437
rect -2343 -471 -2337 -437
rect -2383 -509 -2337 -471
rect -2383 -543 -2377 -509
rect -2343 -543 -2337 -509
rect -2383 -581 -2337 -543
rect -2383 -615 -2377 -581
rect -2343 -615 -2337 -581
rect -2383 -653 -2337 -615
rect -2383 -687 -2377 -653
rect -2343 -687 -2337 -653
rect -2383 -718 -2337 -687
rect -2265 -149 -2219 -118
rect -2265 -183 -2259 -149
rect -2225 -183 -2219 -149
rect -2265 -221 -2219 -183
rect -2265 -255 -2259 -221
rect -2225 -255 -2219 -221
rect -2265 -293 -2219 -255
rect -2265 -327 -2259 -293
rect -2225 -327 -2219 -293
rect -2265 -365 -2219 -327
rect -2265 -399 -2259 -365
rect -2225 -399 -2219 -365
rect -2265 -437 -2219 -399
rect -2265 -471 -2259 -437
rect -2225 -471 -2219 -437
rect -2265 -509 -2219 -471
rect -2265 -543 -2259 -509
rect -2225 -543 -2219 -509
rect -2265 -581 -2219 -543
rect -2265 -615 -2259 -581
rect -2225 -615 -2219 -581
rect -2265 -653 -2219 -615
rect -2265 -687 -2259 -653
rect -2225 -687 -2219 -653
rect -2265 -718 -2219 -687
rect -2147 -149 -2101 -118
rect -2147 -183 -2141 -149
rect -2107 -183 -2101 -149
rect -2147 -221 -2101 -183
rect -2147 -255 -2141 -221
rect -2107 -255 -2101 -221
rect -2147 -293 -2101 -255
rect -2147 -327 -2141 -293
rect -2107 -327 -2101 -293
rect -2147 -365 -2101 -327
rect -2147 -399 -2141 -365
rect -2107 -399 -2101 -365
rect -2147 -437 -2101 -399
rect -2147 -471 -2141 -437
rect -2107 -471 -2101 -437
rect -2147 -509 -2101 -471
rect -2147 -543 -2141 -509
rect -2107 -543 -2101 -509
rect -2147 -581 -2101 -543
rect -2147 -615 -2141 -581
rect -2107 -615 -2101 -581
rect -2147 -653 -2101 -615
rect -2147 -687 -2141 -653
rect -2107 -687 -2101 -653
rect -2147 -718 -2101 -687
rect -2029 -149 -1983 -118
rect -2029 -183 -2023 -149
rect -1989 -183 -1983 -149
rect -2029 -221 -1983 -183
rect -2029 -255 -2023 -221
rect -1989 -255 -1983 -221
rect -2029 -293 -1983 -255
rect -2029 -327 -2023 -293
rect -1989 -327 -1983 -293
rect -2029 -365 -1983 -327
rect -2029 -399 -2023 -365
rect -1989 -399 -1983 -365
rect -2029 -437 -1983 -399
rect -2029 -471 -2023 -437
rect -1989 -471 -1983 -437
rect -2029 -509 -1983 -471
rect -2029 -543 -2023 -509
rect -1989 -543 -1983 -509
rect -2029 -581 -1983 -543
rect -2029 -615 -2023 -581
rect -1989 -615 -1983 -581
rect -2029 -653 -1983 -615
rect -2029 -687 -2023 -653
rect -1989 -687 -1983 -653
rect -2029 -718 -1983 -687
rect -1911 -149 -1865 -118
rect -1911 -183 -1905 -149
rect -1871 -183 -1865 -149
rect -1911 -221 -1865 -183
rect -1911 -255 -1905 -221
rect -1871 -255 -1865 -221
rect -1911 -293 -1865 -255
rect -1911 -327 -1905 -293
rect -1871 -327 -1865 -293
rect -1911 -365 -1865 -327
rect -1911 -399 -1905 -365
rect -1871 -399 -1865 -365
rect -1911 -437 -1865 -399
rect -1911 -471 -1905 -437
rect -1871 -471 -1865 -437
rect -1911 -509 -1865 -471
rect -1911 -543 -1905 -509
rect -1871 -543 -1865 -509
rect -1911 -581 -1865 -543
rect -1911 -615 -1905 -581
rect -1871 -615 -1865 -581
rect -1911 -653 -1865 -615
rect -1911 -687 -1905 -653
rect -1871 -687 -1865 -653
rect -1911 -718 -1865 -687
rect -1793 -149 -1747 -118
rect -1793 -183 -1787 -149
rect -1753 -183 -1747 -149
rect -1793 -221 -1747 -183
rect -1793 -255 -1787 -221
rect -1753 -255 -1747 -221
rect -1793 -293 -1747 -255
rect -1793 -327 -1787 -293
rect -1753 -327 -1747 -293
rect -1793 -365 -1747 -327
rect -1793 -399 -1787 -365
rect -1753 -399 -1747 -365
rect -1793 -437 -1747 -399
rect -1793 -471 -1787 -437
rect -1753 -471 -1747 -437
rect -1793 -509 -1747 -471
rect -1793 -543 -1787 -509
rect -1753 -543 -1747 -509
rect -1793 -581 -1747 -543
rect -1793 -615 -1787 -581
rect -1753 -615 -1747 -581
rect -1793 -653 -1747 -615
rect -1793 -687 -1787 -653
rect -1753 -687 -1747 -653
rect -1793 -718 -1747 -687
rect -1675 -149 -1629 -118
rect -1675 -183 -1669 -149
rect -1635 -183 -1629 -149
rect -1675 -221 -1629 -183
rect -1675 -255 -1669 -221
rect -1635 -255 -1629 -221
rect -1675 -293 -1629 -255
rect -1675 -327 -1669 -293
rect -1635 -327 -1629 -293
rect -1675 -365 -1629 -327
rect -1675 -399 -1669 -365
rect -1635 -399 -1629 -365
rect -1675 -437 -1629 -399
rect -1675 -471 -1669 -437
rect -1635 -471 -1629 -437
rect -1675 -509 -1629 -471
rect -1675 -543 -1669 -509
rect -1635 -543 -1629 -509
rect -1675 -581 -1629 -543
rect -1675 -615 -1669 -581
rect -1635 -615 -1629 -581
rect -1675 -653 -1629 -615
rect -1675 -687 -1669 -653
rect -1635 -687 -1629 -653
rect -1675 -718 -1629 -687
rect -1557 -149 -1511 -118
rect -1557 -183 -1551 -149
rect -1517 -183 -1511 -149
rect -1557 -221 -1511 -183
rect -1557 -255 -1551 -221
rect -1517 -255 -1511 -221
rect -1557 -293 -1511 -255
rect -1557 -327 -1551 -293
rect -1517 -327 -1511 -293
rect -1557 -365 -1511 -327
rect -1557 -399 -1551 -365
rect -1517 -399 -1511 -365
rect -1557 -437 -1511 -399
rect -1557 -471 -1551 -437
rect -1517 -471 -1511 -437
rect -1557 -509 -1511 -471
rect -1557 -543 -1551 -509
rect -1517 -543 -1511 -509
rect -1557 -581 -1511 -543
rect -1557 -615 -1551 -581
rect -1517 -615 -1511 -581
rect -1557 -653 -1511 -615
rect -1557 -687 -1551 -653
rect -1517 -687 -1511 -653
rect -1557 -718 -1511 -687
rect -1439 -149 -1393 -118
rect -1439 -183 -1433 -149
rect -1399 -183 -1393 -149
rect -1439 -221 -1393 -183
rect -1439 -255 -1433 -221
rect -1399 -255 -1393 -221
rect -1439 -293 -1393 -255
rect -1439 -327 -1433 -293
rect -1399 -327 -1393 -293
rect -1439 -365 -1393 -327
rect -1439 -399 -1433 -365
rect -1399 -399 -1393 -365
rect -1439 -437 -1393 -399
rect -1439 -471 -1433 -437
rect -1399 -471 -1393 -437
rect -1439 -509 -1393 -471
rect -1439 -543 -1433 -509
rect -1399 -543 -1393 -509
rect -1439 -581 -1393 -543
rect -1439 -615 -1433 -581
rect -1399 -615 -1393 -581
rect -1439 -653 -1393 -615
rect -1439 -687 -1433 -653
rect -1399 -687 -1393 -653
rect -1439 -718 -1393 -687
rect -1321 -149 -1275 -118
rect -1321 -183 -1315 -149
rect -1281 -183 -1275 -149
rect -1321 -221 -1275 -183
rect -1321 -255 -1315 -221
rect -1281 -255 -1275 -221
rect -1321 -293 -1275 -255
rect -1321 -327 -1315 -293
rect -1281 -327 -1275 -293
rect -1321 -365 -1275 -327
rect -1321 -399 -1315 -365
rect -1281 -399 -1275 -365
rect -1321 -437 -1275 -399
rect -1321 -471 -1315 -437
rect -1281 -471 -1275 -437
rect -1321 -509 -1275 -471
rect -1321 -543 -1315 -509
rect -1281 -543 -1275 -509
rect -1321 -581 -1275 -543
rect -1321 -615 -1315 -581
rect -1281 -615 -1275 -581
rect -1321 -653 -1275 -615
rect -1321 -687 -1315 -653
rect -1281 -687 -1275 -653
rect -1321 -718 -1275 -687
rect -1203 -149 -1157 -118
rect -1203 -183 -1197 -149
rect -1163 -183 -1157 -149
rect -1203 -221 -1157 -183
rect -1203 -255 -1197 -221
rect -1163 -255 -1157 -221
rect -1203 -293 -1157 -255
rect -1203 -327 -1197 -293
rect -1163 -327 -1157 -293
rect -1203 -365 -1157 -327
rect -1203 -399 -1197 -365
rect -1163 -399 -1157 -365
rect -1203 -437 -1157 -399
rect -1203 -471 -1197 -437
rect -1163 -471 -1157 -437
rect -1203 -509 -1157 -471
rect -1203 -543 -1197 -509
rect -1163 -543 -1157 -509
rect -1203 -581 -1157 -543
rect -1203 -615 -1197 -581
rect -1163 -615 -1157 -581
rect -1203 -653 -1157 -615
rect -1203 -687 -1197 -653
rect -1163 -687 -1157 -653
rect -1203 -718 -1157 -687
rect -1085 -149 -1039 -118
rect -1085 -183 -1079 -149
rect -1045 -183 -1039 -149
rect -1085 -221 -1039 -183
rect -1085 -255 -1079 -221
rect -1045 -255 -1039 -221
rect -1085 -293 -1039 -255
rect -1085 -327 -1079 -293
rect -1045 -327 -1039 -293
rect -1085 -365 -1039 -327
rect -1085 -399 -1079 -365
rect -1045 -399 -1039 -365
rect -1085 -437 -1039 -399
rect -1085 -471 -1079 -437
rect -1045 -471 -1039 -437
rect -1085 -509 -1039 -471
rect -1085 -543 -1079 -509
rect -1045 -543 -1039 -509
rect -1085 -581 -1039 -543
rect -1085 -615 -1079 -581
rect -1045 -615 -1039 -581
rect -1085 -653 -1039 -615
rect -1085 -687 -1079 -653
rect -1045 -687 -1039 -653
rect -1085 -718 -1039 -687
rect -967 -149 -921 -118
rect -967 -183 -961 -149
rect -927 -183 -921 -149
rect -967 -221 -921 -183
rect -967 -255 -961 -221
rect -927 -255 -921 -221
rect -967 -293 -921 -255
rect -967 -327 -961 -293
rect -927 -327 -921 -293
rect -967 -365 -921 -327
rect -967 -399 -961 -365
rect -927 -399 -921 -365
rect -967 -437 -921 -399
rect -967 -471 -961 -437
rect -927 -471 -921 -437
rect -967 -509 -921 -471
rect -967 -543 -961 -509
rect -927 -543 -921 -509
rect -967 -581 -921 -543
rect -967 -615 -961 -581
rect -927 -615 -921 -581
rect -967 -653 -921 -615
rect -967 -687 -961 -653
rect -927 -687 -921 -653
rect -967 -718 -921 -687
rect -849 -149 -803 -118
rect -849 -183 -843 -149
rect -809 -183 -803 -149
rect -849 -221 -803 -183
rect -849 -255 -843 -221
rect -809 -255 -803 -221
rect -849 -293 -803 -255
rect -849 -327 -843 -293
rect -809 -327 -803 -293
rect -849 -365 -803 -327
rect -849 -399 -843 -365
rect -809 -399 -803 -365
rect -849 -437 -803 -399
rect -849 -471 -843 -437
rect -809 -471 -803 -437
rect -849 -509 -803 -471
rect -849 -543 -843 -509
rect -809 -543 -803 -509
rect -849 -581 -803 -543
rect -849 -615 -843 -581
rect -809 -615 -803 -581
rect -849 -653 -803 -615
rect -849 -687 -843 -653
rect -809 -687 -803 -653
rect -849 -718 -803 -687
rect -731 -149 -685 -118
rect -731 -183 -725 -149
rect -691 -183 -685 -149
rect -731 -221 -685 -183
rect -731 -255 -725 -221
rect -691 -255 -685 -221
rect -731 -293 -685 -255
rect -731 -327 -725 -293
rect -691 -327 -685 -293
rect -731 -365 -685 -327
rect -731 -399 -725 -365
rect -691 -399 -685 -365
rect -731 -437 -685 -399
rect -731 -471 -725 -437
rect -691 -471 -685 -437
rect -731 -509 -685 -471
rect -731 -543 -725 -509
rect -691 -543 -685 -509
rect -731 -581 -685 -543
rect -731 -615 -725 -581
rect -691 -615 -685 -581
rect -731 -653 -685 -615
rect -731 -687 -725 -653
rect -691 -687 -685 -653
rect -731 -718 -685 -687
rect -613 -149 -567 -118
rect -613 -183 -607 -149
rect -573 -183 -567 -149
rect -613 -221 -567 -183
rect -613 -255 -607 -221
rect -573 -255 -567 -221
rect -613 -293 -567 -255
rect -613 -327 -607 -293
rect -573 -327 -567 -293
rect -613 -365 -567 -327
rect -613 -399 -607 -365
rect -573 -399 -567 -365
rect -613 -437 -567 -399
rect -613 -471 -607 -437
rect -573 -471 -567 -437
rect -613 -509 -567 -471
rect -613 -543 -607 -509
rect -573 -543 -567 -509
rect -613 -581 -567 -543
rect -613 -615 -607 -581
rect -573 -615 -567 -581
rect -613 -653 -567 -615
rect -613 -687 -607 -653
rect -573 -687 -567 -653
rect -613 -718 -567 -687
rect -495 -149 -449 -118
rect -495 -183 -489 -149
rect -455 -183 -449 -149
rect -495 -221 -449 -183
rect -495 -255 -489 -221
rect -455 -255 -449 -221
rect -495 -293 -449 -255
rect -495 -327 -489 -293
rect -455 -327 -449 -293
rect -495 -365 -449 -327
rect -495 -399 -489 -365
rect -455 -399 -449 -365
rect -495 -437 -449 -399
rect -495 -471 -489 -437
rect -455 -471 -449 -437
rect -495 -509 -449 -471
rect -495 -543 -489 -509
rect -455 -543 -449 -509
rect -495 -581 -449 -543
rect -495 -615 -489 -581
rect -455 -615 -449 -581
rect -495 -653 -449 -615
rect -495 -687 -489 -653
rect -455 -687 -449 -653
rect -495 -718 -449 -687
rect -377 -149 -331 -118
rect -377 -183 -371 -149
rect -337 -183 -331 -149
rect -377 -221 -331 -183
rect -377 -255 -371 -221
rect -337 -255 -331 -221
rect -377 -293 -331 -255
rect -377 -327 -371 -293
rect -337 -327 -331 -293
rect -377 -365 -331 -327
rect -377 -399 -371 -365
rect -337 -399 -331 -365
rect -377 -437 -331 -399
rect -377 -471 -371 -437
rect -337 -471 -331 -437
rect -377 -509 -331 -471
rect -377 -543 -371 -509
rect -337 -543 -331 -509
rect -377 -581 -331 -543
rect -377 -615 -371 -581
rect -337 -615 -331 -581
rect -377 -653 -331 -615
rect -377 -687 -371 -653
rect -337 -687 -331 -653
rect -377 -718 -331 -687
rect -259 -149 -213 -118
rect -259 -183 -253 -149
rect -219 -183 -213 -149
rect -259 -221 -213 -183
rect -259 -255 -253 -221
rect -219 -255 -213 -221
rect -259 -293 -213 -255
rect -259 -327 -253 -293
rect -219 -327 -213 -293
rect -259 -365 -213 -327
rect -259 -399 -253 -365
rect -219 -399 -213 -365
rect -259 -437 -213 -399
rect -259 -471 -253 -437
rect -219 -471 -213 -437
rect -259 -509 -213 -471
rect -259 -543 -253 -509
rect -219 -543 -213 -509
rect -259 -581 -213 -543
rect -259 -615 -253 -581
rect -219 -615 -213 -581
rect -259 -653 -213 -615
rect -259 -687 -253 -653
rect -219 -687 -213 -653
rect -259 -718 -213 -687
rect -141 -149 -95 -118
rect -141 -183 -135 -149
rect -101 -183 -95 -149
rect -141 -221 -95 -183
rect -141 -255 -135 -221
rect -101 -255 -95 -221
rect -141 -293 -95 -255
rect -141 -327 -135 -293
rect -101 -327 -95 -293
rect -141 -365 -95 -327
rect -141 -399 -135 -365
rect -101 -399 -95 -365
rect -141 -437 -95 -399
rect -141 -471 -135 -437
rect -101 -471 -95 -437
rect -141 -509 -95 -471
rect -141 -543 -135 -509
rect -101 -543 -95 -509
rect -141 -581 -95 -543
rect -141 -615 -135 -581
rect -101 -615 -95 -581
rect -141 -653 -95 -615
rect -141 -687 -135 -653
rect -101 -687 -95 -653
rect -141 -718 -95 -687
rect -23 -149 23 -118
rect -23 -183 -17 -149
rect 17 -183 23 -149
rect -23 -221 23 -183
rect -23 -255 -17 -221
rect 17 -255 23 -221
rect -23 -293 23 -255
rect -23 -327 -17 -293
rect 17 -327 23 -293
rect -23 -365 23 -327
rect -23 -399 -17 -365
rect 17 -399 23 -365
rect -23 -437 23 -399
rect -23 -471 -17 -437
rect 17 -471 23 -437
rect -23 -509 23 -471
rect -23 -543 -17 -509
rect 17 -543 23 -509
rect -23 -581 23 -543
rect -23 -615 -17 -581
rect 17 -615 23 -581
rect -23 -653 23 -615
rect -23 -687 -17 -653
rect 17 -687 23 -653
rect -23 -718 23 -687
rect 95 -149 141 -118
rect 95 -183 101 -149
rect 135 -183 141 -149
rect 95 -221 141 -183
rect 95 -255 101 -221
rect 135 -255 141 -221
rect 95 -293 141 -255
rect 95 -327 101 -293
rect 135 -327 141 -293
rect 95 -365 141 -327
rect 95 -399 101 -365
rect 135 -399 141 -365
rect 95 -437 141 -399
rect 95 -471 101 -437
rect 135 -471 141 -437
rect 95 -509 141 -471
rect 95 -543 101 -509
rect 135 -543 141 -509
rect 95 -581 141 -543
rect 95 -615 101 -581
rect 135 -615 141 -581
rect 95 -653 141 -615
rect 95 -687 101 -653
rect 135 -687 141 -653
rect 95 -718 141 -687
rect 213 -149 259 -118
rect 213 -183 219 -149
rect 253 -183 259 -149
rect 213 -221 259 -183
rect 213 -255 219 -221
rect 253 -255 259 -221
rect 213 -293 259 -255
rect 213 -327 219 -293
rect 253 -327 259 -293
rect 213 -365 259 -327
rect 213 -399 219 -365
rect 253 -399 259 -365
rect 213 -437 259 -399
rect 213 -471 219 -437
rect 253 -471 259 -437
rect 213 -509 259 -471
rect 213 -543 219 -509
rect 253 -543 259 -509
rect 213 -581 259 -543
rect 213 -615 219 -581
rect 253 -615 259 -581
rect 213 -653 259 -615
rect 213 -687 219 -653
rect 253 -687 259 -653
rect 213 -718 259 -687
rect 331 -149 377 -118
rect 331 -183 337 -149
rect 371 -183 377 -149
rect 331 -221 377 -183
rect 331 -255 337 -221
rect 371 -255 377 -221
rect 331 -293 377 -255
rect 331 -327 337 -293
rect 371 -327 377 -293
rect 331 -365 377 -327
rect 331 -399 337 -365
rect 371 -399 377 -365
rect 331 -437 377 -399
rect 331 -471 337 -437
rect 371 -471 377 -437
rect 331 -509 377 -471
rect 331 -543 337 -509
rect 371 -543 377 -509
rect 331 -581 377 -543
rect 331 -615 337 -581
rect 371 -615 377 -581
rect 331 -653 377 -615
rect 331 -687 337 -653
rect 371 -687 377 -653
rect 331 -718 377 -687
rect 449 -149 495 -118
rect 449 -183 455 -149
rect 489 -183 495 -149
rect 449 -221 495 -183
rect 449 -255 455 -221
rect 489 -255 495 -221
rect 449 -293 495 -255
rect 449 -327 455 -293
rect 489 -327 495 -293
rect 449 -365 495 -327
rect 449 -399 455 -365
rect 489 -399 495 -365
rect 449 -437 495 -399
rect 449 -471 455 -437
rect 489 -471 495 -437
rect 449 -509 495 -471
rect 449 -543 455 -509
rect 489 -543 495 -509
rect 449 -581 495 -543
rect 449 -615 455 -581
rect 489 -615 495 -581
rect 449 -653 495 -615
rect 449 -687 455 -653
rect 489 -687 495 -653
rect 449 -718 495 -687
rect 567 -149 613 -118
rect 567 -183 573 -149
rect 607 -183 613 -149
rect 567 -221 613 -183
rect 567 -255 573 -221
rect 607 -255 613 -221
rect 567 -293 613 -255
rect 567 -327 573 -293
rect 607 -327 613 -293
rect 567 -365 613 -327
rect 567 -399 573 -365
rect 607 -399 613 -365
rect 567 -437 613 -399
rect 567 -471 573 -437
rect 607 -471 613 -437
rect 567 -509 613 -471
rect 567 -543 573 -509
rect 607 -543 613 -509
rect 567 -581 613 -543
rect 567 -615 573 -581
rect 607 -615 613 -581
rect 567 -653 613 -615
rect 567 -687 573 -653
rect 607 -687 613 -653
rect 567 -718 613 -687
rect 685 -149 731 -118
rect 685 -183 691 -149
rect 725 -183 731 -149
rect 685 -221 731 -183
rect 685 -255 691 -221
rect 725 -255 731 -221
rect 685 -293 731 -255
rect 685 -327 691 -293
rect 725 -327 731 -293
rect 685 -365 731 -327
rect 685 -399 691 -365
rect 725 -399 731 -365
rect 685 -437 731 -399
rect 685 -471 691 -437
rect 725 -471 731 -437
rect 685 -509 731 -471
rect 685 -543 691 -509
rect 725 -543 731 -509
rect 685 -581 731 -543
rect 685 -615 691 -581
rect 725 -615 731 -581
rect 685 -653 731 -615
rect 685 -687 691 -653
rect 725 -687 731 -653
rect 685 -718 731 -687
rect 803 -149 849 -118
rect 803 -183 809 -149
rect 843 -183 849 -149
rect 803 -221 849 -183
rect 803 -255 809 -221
rect 843 -255 849 -221
rect 803 -293 849 -255
rect 803 -327 809 -293
rect 843 -327 849 -293
rect 803 -365 849 -327
rect 803 -399 809 -365
rect 843 -399 849 -365
rect 803 -437 849 -399
rect 803 -471 809 -437
rect 843 -471 849 -437
rect 803 -509 849 -471
rect 803 -543 809 -509
rect 843 -543 849 -509
rect 803 -581 849 -543
rect 803 -615 809 -581
rect 843 -615 849 -581
rect 803 -653 849 -615
rect 803 -687 809 -653
rect 843 -687 849 -653
rect 803 -718 849 -687
rect 921 -149 967 -118
rect 921 -183 927 -149
rect 961 -183 967 -149
rect 921 -221 967 -183
rect 921 -255 927 -221
rect 961 -255 967 -221
rect 921 -293 967 -255
rect 921 -327 927 -293
rect 961 -327 967 -293
rect 921 -365 967 -327
rect 921 -399 927 -365
rect 961 -399 967 -365
rect 921 -437 967 -399
rect 921 -471 927 -437
rect 961 -471 967 -437
rect 921 -509 967 -471
rect 921 -543 927 -509
rect 961 -543 967 -509
rect 921 -581 967 -543
rect 921 -615 927 -581
rect 961 -615 967 -581
rect 921 -653 967 -615
rect 921 -687 927 -653
rect 961 -687 967 -653
rect 921 -718 967 -687
rect 1039 -149 1085 -118
rect 1039 -183 1045 -149
rect 1079 -183 1085 -149
rect 1039 -221 1085 -183
rect 1039 -255 1045 -221
rect 1079 -255 1085 -221
rect 1039 -293 1085 -255
rect 1039 -327 1045 -293
rect 1079 -327 1085 -293
rect 1039 -365 1085 -327
rect 1039 -399 1045 -365
rect 1079 -399 1085 -365
rect 1039 -437 1085 -399
rect 1039 -471 1045 -437
rect 1079 -471 1085 -437
rect 1039 -509 1085 -471
rect 1039 -543 1045 -509
rect 1079 -543 1085 -509
rect 1039 -581 1085 -543
rect 1039 -615 1045 -581
rect 1079 -615 1085 -581
rect 1039 -653 1085 -615
rect 1039 -687 1045 -653
rect 1079 -687 1085 -653
rect 1039 -718 1085 -687
rect 1157 -149 1203 -118
rect 1157 -183 1163 -149
rect 1197 -183 1203 -149
rect 1157 -221 1203 -183
rect 1157 -255 1163 -221
rect 1197 -255 1203 -221
rect 1157 -293 1203 -255
rect 1157 -327 1163 -293
rect 1197 -327 1203 -293
rect 1157 -365 1203 -327
rect 1157 -399 1163 -365
rect 1197 -399 1203 -365
rect 1157 -437 1203 -399
rect 1157 -471 1163 -437
rect 1197 -471 1203 -437
rect 1157 -509 1203 -471
rect 1157 -543 1163 -509
rect 1197 -543 1203 -509
rect 1157 -581 1203 -543
rect 1157 -615 1163 -581
rect 1197 -615 1203 -581
rect 1157 -653 1203 -615
rect 1157 -687 1163 -653
rect 1197 -687 1203 -653
rect 1157 -718 1203 -687
rect 1275 -149 1321 -118
rect 1275 -183 1281 -149
rect 1315 -183 1321 -149
rect 1275 -221 1321 -183
rect 1275 -255 1281 -221
rect 1315 -255 1321 -221
rect 1275 -293 1321 -255
rect 1275 -327 1281 -293
rect 1315 -327 1321 -293
rect 1275 -365 1321 -327
rect 1275 -399 1281 -365
rect 1315 -399 1321 -365
rect 1275 -437 1321 -399
rect 1275 -471 1281 -437
rect 1315 -471 1321 -437
rect 1275 -509 1321 -471
rect 1275 -543 1281 -509
rect 1315 -543 1321 -509
rect 1275 -581 1321 -543
rect 1275 -615 1281 -581
rect 1315 -615 1321 -581
rect 1275 -653 1321 -615
rect 1275 -687 1281 -653
rect 1315 -687 1321 -653
rect 1275 -718 1321 -687
rect 1393 -149 1439 -118
rect 1393 -183 1399 -149
rect 1433 -183 1439 -149
rect 1393 -221 1439 -183
rect 1393 -255 1399 -221
rect 1433 -255 1439 -221
rect 1393 -293 1439 -255
rect 1393 -327 1399 -293
rect 1433 -327 1439 -293
rect 1393 -365 1439 -327
rect 1393 -399 1399 -365
rect 1433 -399 1439 -365
rect 1393 -437 1439 -399
rect 1393 -471 1399 -437
rect 1433 -471 1439 -437
rect 1393 -509 1439 -471
rect 1393 -543 1399 -509
rect 1433 -543 1439 -509
rect 1393 -581 1439 -543
rect 1393 -615 1399 -581
rect 1433 -615 1439 -581
rect 1393 -653 1439 -615
rect 1393 -687 1399 -653
rect 1433 -687 1439 -653
rect 1393 -718 1439 -687
rect 1511 -149 1557 -118
rect 1511 -183 1517 -149
rect 1551 -183 1557 -149
rect 1511 -221 1557 -183
rect 1511 -255 1517 -221
rect 1551 -255 1557 -221
rect 1511 -293 1557 -255
rect 1511 -327 1517 -293
rect 1551 -327 1557 -293
rect 1511 -365 1557 -327
rect 1511 -399 1517 -365
rect 1551 -399 1557 -365
rect 1511 -437 1557 -399
rect 1511 -471 1517 -437
rect 1551 -471 1557 -437
rect 1511 -509 1557 -471
rect 1511 -543 1517 -509
rect 1551 -543 1557 -509
rect 1511 -581 1557 -543
rect 1511 -615 1517 -581
rect 1551 -615 1557 -581
rect 1511 -653 1557 -615
rect 1511 -687 1517 -653
rect 1551 -687 1557 -653
rect 1511 -718 1557 -687
rect 1629 -149 1675 -118
rect 1629 -183 1635 -149
rect 1669 -183 1675 -149
rect 1629 -221 1675 -183
rect 1629 -255 1635 -221
rect 1669 -255 1675 -221
rect 1629 -293 1675 -255
rect 1629 -327 1635 -293
rect 1669 -327 1675 -293
rect 1629 -365 1675 -327
rect 1629 -399 1635 -365
rect 1669 -399 1675 -365
rect 1629 -437 1675 -399
rect 1629 -471 1635 -437
rect 1669 -471 1675 -437
rect 1629 -509 1675 -471
rect 1629 -543 1635 -509
rect 1669 -543 1675 -509
rect 1629 -581 1675 -543
rect 1629 -615 1635 -581
rect 1669 -615 1675 -581
rect 1629 -653 1675 -615
rect 1629 -687 1635 -653
rect 1669 -687 1675 -653
rect 1629 -718 1675 -687
rect 1747 -149 1793 -118
rect 1747 -183 1753 -149
rect 1787 -183 1793 -149
rect 1747 -221 1793 -183
rect 1747 -255 1753 -221
rect 1787 -255 1793 -221
rect 1747 -293 1793 -255
rect 1747 -327 1753 -293
rect 1787 -327 1793 -293
rect 1747 -365 1793 -327
rect 1747 -399 1753 -365
rect 1787 -399 1793 -365
rect 1747 -437 1793 -399
rect 1747 -471 1753 -437
rect 1787 -471 1793 -437
rect 1747 -509 1793 -471
rect 1747 -543 1753 -509
rect 1787 -543 1793 -509
rect 1747 -581 1793 -543
rect 1747 -615 1753 -581
rect 1787 -615 1793 -581
rect 1747 -653 1793 -615
rect 1747 -687 1753 -653
rect 1787 -687 1793 -653
rect 1747 -718 1793 -687
rect 1865 -149 1911 -118
rect 1865 -183 1871 -149
rect 1905 -183 1911 -149
rect 1865 -221 1911 -183
rect 1865 -255 1871 -221
rect 1905 -255 1911 -221
rect 1865 -293 1911 -255
rect 1865 -327 1871 -293
rect 1905 -327 1911 -293
rect 1865 -365 1911 -327
rect 1865 -399 1871 -365
rect 1905 -399 1911 -365
rect 1865 -437 1911 -399
rect 1865 -471 1871 -437
rect 1905 -471 1911 -437
rect 1865 -509 1911 -471
rect 1865 -543 1871 -509
rect 1905 -543 1911 -509
rect 1865 -581 1911 -543
rect 1865 -615 1871 -581
rect 1905 -615 1911 -581
rect 1865 -653 1911 -615
rect 1865 -687 1871 -653
rect 1905 -687 1911 -653
rect 1865 -718 1911 -687
rect 1983 -149 2029 -118
rect 1983 -183 1989 -149
rect 2023 -183 2029 -149
rect 1983 -221 2029 -183
rect 1983 -255 1989 -221
rect 2023 -255 2029 -221
rect 1983 -293 2029 -255
rect 1983 -327 1989 -293
rect 2023 -327 2029 -293
rect 1983 -365 2029 -327
rect 1983 -399 1989 -365
rect 2023 -399 2029 -365
rect 1983 -437 2029 -399
rect 1983 -471 1989 -437
rect 2023 -471 2029 -437
rect 1983 -509 2029 -471
rect 1983 -543 1989 -509
rect 2023 -543 2029 -509
rect 1983 -581 2029 -543
rect 1983 -615 1989 -581
rect 2023 -615 2029 -581
rect 1983 -653 2029 -615
rect 1983 -687 1989 -653
rect 2023 -687 2029 -653
rect 1983 -718 2029 -687
rect 2101 -149 2147 -118
rect 2101 -183 2107 -149
rect 2141 -183 2147 -149
rect 2101 -221 2147 -183
rect 2101 -255 2107 -221
rect 2141 -255 2147 -221
rect 2101 -293 2147 -255
rect 2101 -327 2107 -293
rect 2141 -327 2147 -293
rect 2101 -365 2147 -327
rect 2101 -399 2107 -365
rect 2141 -399 2147 -365
rect 2101 -437 2147 -399
rect 2101 -471 2107 -437
rect 2141 -471 2147 -437
rect 2101 -509 2147 -471
rect 2101 -543 2107 -509
rect 2141 -543 2147 -509
rect 2101 -581 2147 -543
rect 2101 -615 2107 -581
rect 2141 -615 2147 -581
rect 2101 -653 2147 -615
rect 2101 -687 2107 -653
rect 2141 -687 2147 -653
rect 2101 -718 2147 -687
rect 2219 -149 2265 -118
rect 2219 -183 2225 -149
rect 2259 -183 2265 -149
rect 2219 -221 2265 -183
rect 2219 -255 2225 -221
rect 2259 -255 2265 -221
rect 2219 -293 2265 -255
rect 2219 -327 2225 -293
rect 2259 -327 2265 -293
rect 2219 -365 2265 -327
rect 2219 -399 2225 -365
rect 2259 -399 2265 -365
rect 2219 -437 2265 -399
rect 2219 -471 2225 -437
rect 2259 -471 2265 -437
rect 2219 -509 2265 -471
rect 2219 -543 2225 -509
rect 2259 -543 2265 -509
rect 2219 -581 2265 -543
rect 2219 -615 2225 -581
rect 2259 -615 2265 -581
rect 2219 -653 2265 -615
rect 2219 -687 2225 -653
rect 2259 -687 2265 -653
rect 2219 -718 2265 -687
rect 2337 -149 2383 -118
rect 2337 -183 2343 -149
rect 2377 -183 2383 -149
rect 2337 -221 2383 -183
rect 2337 -255 2343 -221
rect 2377 -255 2383 -221
rect 2337 -293 2383 -255
rect 2337 -327 2343 -293
rect 2377 -327 2383 -293
rect 2337 -365 2383 -327
rect 2337 -399 2343 -365
rect 2377 -399 2383 -365
rect 2337 -437 2383 -399
rect 2337 -471 2343 -437
rect 2377 -471 2383 -437
rect 2337 -509 2383 -471
rect 2337 -543 2343 -509
rect 2377 -543 2383 -509
rect 2337 -581 2383 -543
rect 2337 -615 2343 -581
rect 2377 -615 2383 -581
rect 2337 -653 2383 -615
rect 2337 -687 2343 -653
rect 2377 -687 2383 -653
rect 2337 -718 2383 -687
rect 2455 -149 2501 -118
rect 2455 -183 2461 -149
rect 2495 -183 2501 -149
rect 2455 -221 2501 -183
rect 2455 -255 2461 -221
rect 2495 -255 2501 -221
rect 2455 -293 2501 -255
rect 2455 -327 2461 -293
rect 2495 -327 2501 -293
rect 2455 -365 2501 -327
rect 2455 -399 2461 -365
rect 2495 -399 2501 -365
rect 2455 -437 2501 -399
rect 2455 -471 2461 -437
rect 2495 -471 2501 -437
rect 2455 -509 2501 -471
rect 2455 -543 2461 -509
rect 2495 -543 2501 -509
rect 2455 -581 2501 -543
rect 2455 -615 2461 -581
rect 2495 -615 2501 -581
rect 2455 -653 2501 -615
rect 2455 -687 2461 -653
rect 2495 -687 2501 -653
rect 2455 -718 2501 -687
rect 2573 -149 2619 -118
rect 2573 -183 2579 -149
rect 2613 -183 2619 -149
rect 2573 -221 2619 -183
rect 2573 -255 2579 -221
rect 2613 -255 2619 -221
rect 2573 -293 2619 -255
rect 2573 -327 2579 -293
rect 2613 -327 2619 -293
rect 2573 -365 2619 -327
rect 2573 -399 2579 -365
rect 2613 -399 2619 -365
rect 2573 -437 2619 -399
rect 2573 -471 2579 -437
rect 2613 -471 2619 -437
rect 2573 -509 2619 -471
rect 2573 -543 2579 -509
rect 2613 -543 2619 -509
rect 2573 -581 2619 -543
rect 2573 -615 2579 -581
rect 2613 -615 2619 -581
rect 2573 -653 2619 -615
rect 2573 -687 2579 -653
rect 2613 -687 2619 -653
rect 2573 -718 2619 -687
rect 2691 -149 2737 -118
rect 2691 -183 2697 -149
rect 2731 -183 2737 -149
rect 2691 -221 2737 -183
rect 2691 -255 2697 -221
rect 2731 -255 2737 -221
rect 2691 -293 2737 -255
rect 2691 -327 2697 -293
rect 2731 -327 2737 -293
rect 2691 -365 2737 -327
rect 2691 -399 2697 -365
rect 2731 -399 2737 -365
rect 2691 -437 2737 -399
rect 2691 -471 2697 -437
rect 2731 -471 2737 -437
rect 2691 -509 2737 -471
rect 2691 -543 2697 -509
rect 2731 -543 2737 -509
rect 2691 -581 2737 -543
rect 2691 -615 2697 -581
rect 2731 -615 2737 -581
rect 2691 -653 2737 -615
rect 2691 -687 2697 -653
rect 2731 -687 2737 -653
rect 2691 -718 2737 -687
rect 2809 -149 2855 -118
rect 2809 -183 2815 -149
rect 2849 -183 2855 -149
rect 2809 -221 2855 -183
rect 2809 -255 2815 -221
rect 2849 -255 2855 -221
rect 2809 -293 2855 -255
rect 2809 -327 2815 -293
rect 2849 -327 2855 -293
rect 2809 -365 2855 -327
rect 2809 -399 2815 -365
rect 2849 -399 2855 -365
rect 2809 -437 2855 -399
rect 2809 -471 2815 -437
rect 2849 -471 2855 -437
rect 2809 -509 2855 -471
rect 2809 -543 2815 -509
rect 2849 -543 2855 -509
rect 2809 -581 2855 -543
rect 2809 -615 2815 -581
rect 2849 -615 2855 -581
rect 2809 -653 2855 -615
rect 2809 -687 2815 -653
rect 2849 -687 2855 -653
rect 2809 -718 2855 -687
rect 2927 -149 2973 -118
rect 2927 -183 2933 -149
rect 2967 -183 2973 -149
rect 2927 -221 2973 -183
rect 2927 -255 2933 -221
rect 2967 -255 2973 -221
rect 2927 -293 2973 -255
rect 2927 -327 2933 -293
rect 2967 -327 2973 -293
rect 2927 -365 2973 -327
rect 2927 -399 2933 -365
rect 2967 -399 2973 -365
rect 2927 -437 2973 -399
rect 2927 -471 2933 -437
rect 2967 -471 2973 -437
rect 2927 -509 2973 -471
rect 2927 -543 2933 -509
rect 2967 -543 2973 -509
rect 2927 -581 2973 -543
rect 2927 -615 2933 -581
rect 2967 -615 2973 -581
rect 2927 -653 2973 -615
rect 2927 -687 2933 -653
rect 2967 -687 2973 -653
rect 2927 -718 2973 -687
<< properties >>
string FIXED_BBOX -3064 -884 3064 884
<< end >>
