magic
tech sky130A
magscale 1 2
timestamp 1654715968
<< pwell >>
rect -976 9244 676 10696
rect 254 -1586 1906 -94
<< nmoslvt >>
rect -950 9870 650 10270
rect 280 -850 1880 -450
<< ndiff >>
rect -950 10608 650 10670
rect -950 10302 -915 10608
rect 615 10302 650 10608
rect -950 10270 650 10302
rect -950 9815 650 9870
rect -950 9645 -915 9815
rect 615 9645 650 9815
rect -950 9610 650 9645
rect 280 -161 1880 -120
rect 280 -399 315 -161
rect 1845 -399 1880 -161
rect 280 -450 1880 -399
rect 280 -880 1880 -850
rect 280 -1050 315 -880
rect 1845 -1050 1880 -880
rect 280 -1080 1880 -1050
<< ndiffc >>
rect -915 10302 615 10608
rect -915 9645 615 9815
rect 315 -399 1845 -161
rect 315 -1050 1845 -880
<< psubdiff >>
rect -950 9559 650 9610
rect -950 9321 -915 9559
rect 615 9321 650 9559
rect -950 9270 650 9321
rect 280 -1116 1880 -1080
rect 280 -1354 315 -1116
rect 1845 -1354 1880 -1116
rect 280 -1560 1880 -1354
<< psubdiffcont >>
rect -915 9321 615 9559
rect 315 -1354 1845 -1116
<< poly >>
rect -980 10080 -950 10270
rect -1370 10060 -950 10080
rect -1370 9890 -1325 10060
rect -1155 9890 -950 10060
rect -1370 9870 -950 9890
rect 650 9870 680 10270
rect -110 -240 100 -230
rect -110 -410 -66 -240
rect 36 -410 100 -240
rect -110 -450 100 -410
rect -110 -500 280 -450
rect 250 -850 280 -500
rect 1880 -850 1910 -450
<< polycont >>
rect -1325 9890 -1155 10060
rect -66 -410 36 -240
<< locali >>
rect -950 10616 650 10650
rect -950 10294 -923 10616
rect 623 10294 650 10616
rect -950 10270 650 10294
rect -1690 10028 -1325 10060
rect -1155 10028 -1020 10060
rect -1690 9922 -1660 10028
rect -1050 9922 -1020 10028
rect -1690 9890 -1325 9922
rect -1155 9890 -1020 9922
rect -950 9815 650 9850
rect -950 9768 -915 9815
rect 615 9768 650 9815
rect -950 9302 -923 9768
rect 623 9302 650 9768
rect -950 9270 650 9302
rect 280 53 1880 60
rect -400 -272 -66 -240
rect -400 -378 -375 -272
rect -125 -378 -66 -272
rect -400 -410 -66 -378
rect 36 -410 100 -240
rect 280 -413 307 53
rect 1853 -413 1880 53
rect 280 -430 1880 -413
rect 280 -880 1880 -870
rect 280 -1050 315 -880
rect 1845 -1050 1880 -880
rect 280 -1116 1880 -1050
rect 280 -1326 315 -1116
rect 1845 -1326 1880 -1116
rect 280 -1504 307 -1326
rect 1853 -1504 1880 -1326
rect 280 -1550 1880 -1504
<< viali >>
rect -923 10608 623 10616
rect -923 10302 -915 10608
rect -915 10302 615 10608
rect 615 10302 623 10608
rect -923 10294 623 10302
rect -1660 9922 -1325 10028
rect -1325 9922 -1155 10028
rect -1155 9922 -1050 10028
rect -923 9645 -915 9768
rect -915 9645 615 9768
rect 615 9645 623 9768
rect -923 9559 623 9645
rect -923 9321 -915 9559
rect -915 9321 615 9559
rect 615 9321 623 9559
rect -923 9302 623 9321
rect -375 -378 -125 -272
rect 307 -161 1853 53
rect 307 -399 315 -161
rect 315 -399 1845 -161
rect 1845 -399 1853 -161
rect 307 -413 1853 -399
rect 307 -1354 315 -1326
rect 315 -1354 1845 -1326
rect 1845 -1354 1853 -1326
rect 307 -1504 1853 -1354
<< metal1 >>
rect 23020 11280 26995 11570
rect -950 10616 650 10630
rect -950 10294 -923 10616
rect 623 10294 650 10616
rect -950 10270 650 10294
rect -2210 10040 -1020 10060
rect -2210 9910 -2200 10040
rect -1030 9910 -1020 10040
rect -2210 9890 -1020 9910
rect -960 9768 650 9850
rect -960 9302 -923 9768
rect 623 9302 650 9768
rect -960 9220 650 9302
rect 280 53 1880 180
rect -500 -272 100 -240
rect -500 -388 -486 -272
rect -114 -388 100 -272
rect -500 -410 100 -388
rect 280 -413 307 53
rect 1853 -413 1880 53
rect 280 -430 1880 -413
rect -950 -1298 2500 -1280
rect -950 -1542 -914 -1298
rect 2274 -1542 2500 -1298
rect -950 -1560 2500 -1542
rect 24530 -1570 26980 -1270
<< via1 >>
rect -912 10301 612 10609
rect -2200 10028 -1030 10040
rect -2200 9922 -1660 10028
rect -1660 9922 -1050 10028
rect -1050 9922 -1030 10028
rect -2200 9910 -1030 9922
rect -912 9317 612 9753
rect -486 -378 -375 -272
rect -375 -378 -125 -272
rect -125 -378 -114 -272
rect -486 -388 -114 -378
rect 318 -398 1842 38
rect -914 -1326 2274 -1298
rect -914 -1504 307 -1326
rect 307 -1504 1853 -1326
rect 1853 -1504 2274 -1326
rect -914 -1542 2274 -1504
<< metal2 >>
rect -950 10609 650 10630
rect -950 10301 -912 10609
rect 612 10301 650 10609
rect -950 10270 650 10301
rect -950 10269 529 10270
rect -2280 10040 -1020 10060
rect -2280 9910 -2200 10040
rect -1030 9910 -1020 10040
rect -2280 9890 -1020 9910
rect -960 9763 650 9850
rect -960 9753 -898 9763
rect 598 9753 650 9763
rect -960 9317 -912 9753
rect 612 9317 650 9753
rect -960 9307 -898 9317
rect 598 9307 650 9317
rect -960 9220 650 9307
rect 1300 8348 2520 8450
rect 1300 7732 1357 8348
rect 2453 7732 2520 8348
rect 1300 7620 2520 7732
rect 280 3859 1890 3870
rect -1688 3611 2174 3859
rect 280 38 1890 3611
rect -1925 -260 -100 -240
rect -1925 -390 -1910 -260
rect -1200 -272 -100 -260
rect -1200 -388 -486 -272
rect -114 -388 -100 -272
rect -1200 -390 -100 -388
rect -1925 -410 -100 -390
rect 280 -398 318 38
rect 1842 -398 1890 38
rect 280 -430 1890 -398
rect -950 -1298 2490 -1280
rect -950 -1542 -914 -1298
rect 2274 -1542 2490 -1298
rect -950 -1560 2490 -1542
<< via2 >>
rect -898 9753 598 9763
rect -898 9317 598 9753
rect -898 9307 598 9317
rect 1357 7732 2453 8348
rect -1910 -390 -1200 -260
rect -908 -1528 2268 -1312
<< metal3 >>
rect -960 9763 650 9850
rect -960 9307 -898 9763
rect 598 9307 650 9763
rect -960 9220 650 9307
rect -2280 -260 -1180 -240
rect -2280 -390 -1910 -260
rect -1200 -390 -1180 -260
rect -2280 -410 -1180 -390
rect -950 -1280 -265 9220
rect 1300 8352 2520 8450
rect 1300 7728 1353 8352
rect 2457 7728 2520 8352
rect 1300 7620 2520 7728
rect -950 -1312 2490 -1280
rect -950 -1528 -908 -1312
rect 2268 -1528 2490 -1312
rect -950 -1560 2490 -1528
<< via3 >>
rect 1353 8348 2457 8352
rect 1353 7732 1357 8348
rect 1357 7732 2453 8348
rect 2453 7732 2457 8348
rect 1353 7728 2457 7732
<< metal4 >>
rect -2205 12835 26620 13665
rect -2205 8455 -1375 12835
rect -2205 8352 2515 8455
rect -2205 7728 1353 8352
rect 2457 7728 2515 8352
rect -2205 7625 2515 7728
rect 25795 7690 26620 12835
rect 24850 6830 26620 7690
use opamp_v1  opamp_v1_0 ~/CMOS/TopMetalSe-OpenMPW6/mag/fulgor_opamp
timestamp 1654711683
transform 1 0 -1719 0 1 8419
box 2069 -10028 26971 3199
<< labels >>
rlabel metal1 s 26840 11440 26840 11440 4 VDD
port 1 nsew
rlabel metal4 s 26418 7258 26418 7258 4 AOUT
port 2 nsew
rlabel metal2 s -1078 -314 -1078 -314 4 OUT_IB
port 3 nsew
rlabel metal2 s -1576 3762 -1576 3762 4 ARRAY_OUT
port 5 nsew
rlabel metal1 s 26870 -1360 26870 -1360 4 GND
port 6 nsew
<< end >>
