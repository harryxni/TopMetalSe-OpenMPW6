** sch_path: /home/damic/CMOS/TopmetalSe/xschem/untitled-2.sch
**.subckt untitled-2
V1 VDD GND 1.8
V2 PLUS GND DC=0.60
V5 vbias GND DC=0.9
V6 CSA GND DC=0.35
XM1 NB1 NB1 GND GND sky130_fd_pr__nfet_01v8_lvt L=1.2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
I2 VDD NB1 100n
I3 VDD NB2 100n
XM3 NB2 NB2 GND GND sky130_fd_pr__nfet_01v8_lvt L=1.2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 COL0 COL_SEL0 pix_out GND sky130_fd_pr__nfet_01v8_lvt L=0.8 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vrow0 ROW_SEL0 GND 0 pulse(0.0 1.8 1m 0.1m 0.1m 1m 2m)
Vrow1 ROW_SEL1 GND 0.0 pulse(0.0 1.8 2m 0.1m 0.1m 1m 2m)
Vcol0 COL_SEL0 GND 0 pulse(0.0 1.8 1m 0.1m 0.1m 2m 4m)
Vcol1 COL_SEL1 GND 0.0 pulse(0.0 1.8 3m 0.1m 0.1m 2m 4m)
C1 i_empty GND 10f m=1
I4 sf_ib GND 200n
XM5 sf_ib sf_ib VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 COL1 COL_SEL1 pix_out GND sky130_fd_pr__nfet_01v8_lvt L=0.8 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
R4 pix_out GND 1G m=1
R5 pix_out GND 1G m=1
R1 COL0 GND 2G m=1
R2 COL1 GND 2G m=1
I5 GND itest dc=0 PWL(0 0 9.000000e+04u 0.000000e+00 9.008654e+04u 0.000000e+00 9.017308e+04u
+ 1.848889e-19 9.025962e+04u 1.848889e-19 9.034615e+04u 1.848889e-19 9.043269e+04u 1.848889e-19 9.051923e+04u
+ 3.697778e-19 9.060577e+04u 3.697778e-19 9.069231e+04u 3.697778e-19 9.077885e+04u 3.697778e-19 9.086538e+04u
+ 9.244444e-19 9.095192e+04u 1.294222e-18 9.103846e+04u 1.294222e-18 9.112500e+04u 1.294222e-18 9.121154e+04u
+ 1.109333e-18 9.129808e+04u 1.109333e-18 9.138462e+04u 1.109333e-18 9.147115e+04u 1.109333e-18 9.155769e+04u
+ 9.244444e-19 9.164423e+04u 9.244444e-19 9.173077e+04u 9.244444e-19 9.181731e+04u 9.244444e-19 9.190385e+04u
+ 7.395556e-19 9.199038e+04u 7.395556e-19 9.207692e+04u 7.395556e-19 9.216346e+04u 7.395556e-19 9.225000e+04u
+ 5.546667e-19 9.233654e+04u 5.546667e-19 9.242308e+04u 5.546667e-19 9.250962e+04u 5.546667e-19 9.259615e+04u
+ 3.697778e-19 9.268269e+04u 3.697778e-19 9.276923e+04u 3.697778e-19 9.285577e+04u 3.697778e-19 9.294231e+04u
+ 1.848889e-19 9.302885e+04u 1.848889e-19 9.311538e+04u 1.848889e-19 9.320192e+04u 1.664000e-18 9.328846e+04u
+ 1.664000e-18 9.337500e+04u 1.664000e-18 9.346154e+04u 1.848889e-18 9.354808e+04u 1.848889e-18 9.363462e+04u
+ 1.848889e-18 9.372115e+04u 1.848889e-18 9.380769e+04u 1.848889e-18 9.389423e+04u 2.033778e-18 9.398077e+04u
+ 2.033778e-18 9.406731e+04u 2.033778e-18 9.415385e+04u 2.033778e-18 9.424038e+04u 2.033778e-18 9.432692e+04u
+ 2.218667e-18 9.441346e+04u 2.218667e-18 9.450000e+04u 2.218667e-18 9.458654e+04u 2.218667e-18 9.467308e+04u
+ 2.403556e-18 9.475962e+04u 2.403556e-18 9.484615e+04u 2.403556e-18 9.493269e+04u 2.403556e-18 9.501923e+04u
+ 2.403556e-18 9.510577e+04u 2.588444e-18 9.519231e+04u 3.328000e-18 9.527885e+04u 3.328000e-18 9.536538e+04u
+ 3.328000e-18 9.545192e+04u 3.328000e-18 9.553846e+04u 3.328000e-18 9.562500e+04u 3.328000e-18 9.571154e+04u
+ 3.328000e-18 9.579808e+04u 3.328000e-18 9.588462e+04u 3.328000e-18 9.597115e+04u 3.328000e-18 9.605769e+04u
+ 3.328000e-18 9.614423e+04u 3.328000e-18 9.623077e+04u 3.328000e-18 9.631731e+04u 3.328000e-18 9.640385e+04u
+ 3.328000e-18 9.649038e+04u 3.512889e-18 9.657692e+04u 3.512889e-18 9.666346e+04u 3.512889e-18 9.675000e+04u
+ 3.512889e-18 9.683654e+04u 3.697778e-18 9.692308e+04u 3.882667e-18 9.700962e+04u 3.882667e-18 9.709615e+04u
+ 3.882667e-18 9.718269e+04u 3.882667e-18 9.726923e+04u 3.882667e-18 9.735577e+04u 3.882667e-18 9.744231e+04u
+ 3.697778e-18 9.752885e+04u 3.697778e-18 9.761538e+04u 3.697778e-18 9.770192e+04u 3.697778e-18 9.778846e+04u
+ 3.697778e-18 9.787500e+04u 3.697778e-18 9.796154e+04u 3.697778e-18 9.804808e+04u 3.697778e-18 9.813462e+04u
+ 3.697778e-18 9.822115e+04u 3.697778e-18 9.830769e+04u 3.697778e-18 9.839423e+04u 3.697778e-18 9.848077e+04u
+ 3.697778e-18 9.856731e+04u 3.697778e-18 9.865385e+04u 3.697778e-18 9.874038e+04u 3.697778e-18 9.882692e+04u
+ 3.697778e-18 9.891346e+04u 3.697778e-18 9.900000e+04u 3.697778e-18 9.908654e+04u 3.697778e-18 9.917308e+04u
+ 3.697778e-18 9.925962e+04u 3.697778e-18 9.934615e+04u 3.697778e-18 9.943269e+04u 3.697778e-18 9.951923e+04u
+ 3.697778e-18 9.960577e+04u 3.328000e-18 9.969231e+04u 3.328000e-18 9.977885e+04u 3.328000e-18 9.986538e+04u
+ 3.328000e-18 9.995192e+04u 3.328000e-18 1.000385e+05u 3.328000e-18 1.001250e+05u 3.328000e-18 1.002115e+05u
+ 3.328000e-18 1.002981e+05u 3.328000e-18 1.003846e+05u 3.512889e-18 1.004712e+05u 3.512889e-18 1.005577e+05u
+ 3.512889e-18 1.006442e+05u 3.143111e-18 1.007308e+05u 2.588444e-18 1.008173e+05u 2.588444e-18 1.009038e+05u
+ 2.588444e-18 1.009904e+05u 2.588444e-18 1.010769e+05u 2.588444e-18 1.011635e+05u 2.588444e-18 1.012500e+05u
+ 2.588444e-18 1.013365e+05u 2.588444e-18 1.014231e+05u 2.588444e-18 1.015096e+05u 2.588444e-18 1.015962e+05u
+ 3.328000e-18 1.016827e+05u 3.512889e-18 1.017692e+05u 3.512889e-18 1.018558e+05u 3.512889e-18 1.019423e+05u
+ 3.512889e-18 1.020288e+05u 3.512889e-18 1.021154e+05u 3.512889e-18 1.022019e+05u 3.512889e-18 1.022885e+05u
+ 3.512889e-18 1.023750e+05u 3.882667e-18 1.024615e+05u 4.622222e-18 1.025481e+05u 4.622222e-18 1.026346e+05u
+ 4.622222e-18 1.027212e+05u 4.622222e-18 1.028077e+05u 4.622222e-18 1.028942e+05u 4.622222e-18 1.029808e+05u
+ 4.622222e-18 1.030673e+05u 4.992000e-18 1.031538e+05u 5.361778e-18 1.032404e+05u 5.361778e-18 1.033269e+05u
+ 5.361778e-18 1.034135e+05u 5.361778e-18 1.035000e+05u 5.361778e-18 1.035865e+05u 5.361778e-18 1.036731e+05u
+ 5.731556e-18 1.037596e+05u 5.916444e-18 1.038462e+05u 5.916444e-18 1.039327e+05u 5.916444e-18 1.040192e+05u
+ 5.916444e-18 1.041058e+05u 5.916444e-18 1.041923e+05u 6.101333e-18 1.042788e+05u 6.286222e-18 1.043654e+05u
+ 6.286222e-18 1.044519e+05u 6.286222e-18 1.045385e+05u 6.286222e-18 1.046250e+05u 5.731556e-18 1.047115e+05u
+ 5.361778e-18 1.047981e+05u 5.361778e-18 1.048846e+05u 5.361778e-18 1.049712e+05u 4.807111e-18 1.050577e+05u
+ 3.328000e-18 1.051442e+05u 3.328000e-18 1.052308e+05u 3.328000e-18 1.053173e+05u 2.773333e-18 1.054038e+05u
+ 2.218667e-18 1.054904e+05u 2.218667e-18 1.055769e+05u 2.033778e-18 1.056635e+05u 1.294222e-18 1.057500e+05u
+ 1.294222e-18 1.058365e+05u 3.697778e-19 1.059231e+05u -5.546667e-19 1.060096e+05u -5.546667e-19 1.060962e+05u
+ -5.546667e-19 1.061827e+05u -5.546667e-19 1.062692e+05u 0.000000e+00 1.063558e+05u -1.109333e-17 1.064423e+05u
+ -3.494400e-17 1.065288e+05u -1.872924e-16 1.066154e+05u -7.922489e-16 1.067019e+05u -1.936711e-15 1.067885e+05u
+ -7.567872e-15 1.068750e+05u -2.214507e-14 1.069615e+05u -8.125349e-14 1.070481e+05u -2.706174e-13 1.071346e+05u
+ -9.037204e-13 1.072212e+05u -1.981988e-12 1.072212e+05u 0.000000e+00 1.073077e+05u 0.000000e+00 1.073942e+05u 0)
+

x1 i_empty i_empty i_empty ROW_SEL0 sf_ib GND CSA VDD NB2 NB1 PLUS vbias ROW_SEL1 COL0 COL1 net1
+ array_2x2
C2 itest net1 10f m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /opt/OpenICEDA/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt


**** end user architecture code
**.ends

* expanding   symbol:  /home/damic/CMOS/TopmetalSe/Pixel/Testbench/array_2x2.sym # of pins=16
** sym_path: /home/damic/CMOS/TopmetalSe/Pixel/Testbench/array_2x2.sym
** sch_path: /home/damic/CMOS/TopmetalSe/Pixel/Testbench/array_2x2.sch
.subckt array_2x2  PIX1_IN PIX2_IN PIX3_IN ROW_SEL0 SF_IB GND CSA_VREF VDD NB2 NB1 VREF VBIAS
+ ROW_SEL1 PIX_OUT0 PIX_OUT1 PIX0_IN
Xpixel_5 ROW_SEL0 NB1 CSA_VREF SF_IB NB2 VREF VBIAS PIX3_in PIX_OUT1 VDD GND pixel
Xpixel_6 ROW_SEL0 NB1 CSA_VREF SF_IB NB2 VREF VBIAS PIX2_in PIX_OUT0 VDD GND pixel
Xpixel_7 ROW_SEL1 NB1 CSA_VREF SF_IB NB2 VREF VBIAS PIX1_in PIX_OUT1 VDD GND pixel
Xpixel_8 ROW_SEL1 NB1 CSA_VREF SF_IB NB2 VREF VBIAS PIX0_IN PIX_OUT0 VDD GND pixel
C0 PIX_OUT1 GND 3.53fF
C1 PIX_OUT0 GND 3.53fF
C2 CSA_VREF GND 4.91fF
C3 SF_IB GND 3.80fF
C4 NB2 GND 3.98fF
C5 VREF GND 4.59fF
C6 VBIAS GND 5.46fF
C7 VDD GND 45.33fF
C8 ROW_SEL1 GND 2.43fF
C9 PIX0_IN GND 4.83fF
C10 PIX1_in GND 4.81fF
C11 NB1 GND 6.18fF
C12 ROW_SEL0 GND 2.44fF
C13 PIX2_in GND 4.81fF
C14 PIX3_in GND 4.81fF

.ends

.subckt pixel ROW_SEL NB1 CSA_VREF SF_IB NB2 VREF VBIAS AMP_IN PIX_OUT VDD GND
X0 a_255_n320# a_n315_n320# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=7e+11p pd=5.4e+06u as=1.42e+12p ps=9.2e+06u w=1e+06u l=1.95e+06u
X1 net1 NB2 GND GND sky130_fd_pr__nfet_01v8_lvt ad=5e+11p pd=3e+06u as=7e+11p ps=5.4e+06u w=1e+06u l=1.2e+06u
X2 a_5_n425# VBIAS a_5_n520# GND sky130_fd_pr__nfet_01v8_lvt ad=3.5e+11p pd=2.7e+06u as=1.945e+12p ps=1.71e+07u w=1e+06u l=800000u
X3 a_255_n320# a_n280_n335# a_5_n425# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=3.5e+11p ps=2.7e+06u w=1e+06u l=1.95e+06u
X4 a_495_n465# net1 a_495_n575# GND sky130_fd_pr__nfet_01v8_lvt ad=3.5e+11p pd=2.7e+06u as=3e+11p ps=2.6e+06u w=1e+06u l=800000u
X5 a_n280_n335# a_n280_n335# a_n315_n320# VDD sky130_fd_pr__pfet_01v8_lvt ad=3.5e+11p pd=2.7e+06u as=7e+11p ps=5.4e+06u w=1e+06u l=2e+06u
X6 VDD a_n315_n320# a_n315_n320# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X7 AMP_IN CSA_VREF net1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.25e+11p pd=1.9e+06u as=1.8e+11p ps=1.7e+06u w=450000u l=8e+06u
X8 a_n280_n335# VBIAS a_n125_n520# GND sky130_fd_pr__nfet_01v8_lvt ad=3.5e+11p pd=2.7e+06u as=1.945e+12p ps=1.71e+07u w=1e+06u l=800000u
X9 VDD a_5_n425# net1 GND sky130_fd_pr__nfet_01v8_lvt ad=8.45e+11p pd=5.7e+06u as=0p ps=0u w=1e+06u l=1e+06u
X10 a_n60_n1325# NB1 GND GND sky130_fd_pr__nfet_01v8_lvt ad=3.15e+12p pd=1.75e+07u as=0p ps=0u w=1e+06u l=1.2e+06u
X11 a_n60_n1325# VREF a_n125_n520# GND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=7e+06u l=150000u
X12 a_5_n520# AMP_IN a_n60_n1325# GND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=7e+06u l=150000u
X13 a_495_n575# ROW_SEL PIX_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=800000u
X14 VDD SF_IB a_495_n465# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=5.2e+11p ps=3.4e+06u w=1.3e+06u l=1e+06u
X15 AMP_IN net1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
C0 AMP_IN GND 4.81fF
C1 VDD GND 9.48fF
.ends





.GLOBAL GND
.GLOBAL VDD
**** begin user architecture code


.options savecurrents
.options gmin=0.0000000000000000000001
.control
save all
save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gm]
op
tran 1m 200m
plot v(pix_out)
write pixel_tb.raw
.endc


**** end user architecture code
.end
