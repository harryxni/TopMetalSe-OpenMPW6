magic
tech sky130A
magscale 1 2
timestamp 1654643410
<< error_s >>
rect 200980 681090 201180 681290
rect 201490 681090 201690 681290
rect 200990 680925 201170 681090
rect 201500 680920 201680 681090
rect 198532 675322 198540 675468
rect 198560 675350 198568 675440
rect 198640 675423 198920 675430
rect 198587 675421 198963 675423
rect 198587 675369 198969 675421
rect 198587 675367 198963 675369
rect 198640 675360 198920 675367
rect 198422 674057 198558 674113
rect 198440 674030 198530 674057
rect 198710 673407 198800 673410
rect 198678 673343 198822 673407
rect 198710 673340 198800 673343
rect 198640 672423 198920 672430
rect 198627 672421 198923 672423
rect 198621 672369 198929 672421
rect 198627 672367 198923 672369
rect 198640 672360 198920 672367
rect 198416 671100 198428 671103
rect 198452 671100 198508 671103
rect 198440 671030 198530 671100
rect 198532 671047 198554 671103
rect 198710 670407 198800 670410
rect 198663 670343 198807 670407
rect 198710 670340 198800 670343
rect 198416 668100 198418 668103
rect 198442 668100 198578 668103
rect 198440 668047 198578 668100
rect 198440 668030 198530 668047
<< pwell >>
rect 208934 677354 210586 678576
rect 208554 664744 210206 666016
<< nmoslvt >>
rect 208960 677850 210560 678250
rect 208580 665190 210180 665590
<< ndiff >>
rect 208960 678465 210560 678550
rect 208960 678295 208995 678465
rect 210525 678295 210560 678465
rect 208960 678250 210560 678295
rect 208960 677766 210560 677850
rect 208960 677664 209005 677766
rect 210535 677664 210560 677766
rect 208960 677610 210560 677664
rect 208580 665953 210180 665990
rect 208580 665647 208615 665953
rect 210145 665647 210180 665953
rect 208580 665590 210180 665647
rect 208580 665131 210180 665190
rect 208580 665029 208620 665131
rect 210150 665029 210180 665131
rect 208580 664990 210180 665029
<< ndiffc >>
rect 208995 678295 210525 678465
rect 209005 677664 210535 677766
rect 208615 665647 210145 665953
rect 208620 665029 210150 665131
<< psubdiff >>
rect 208960 677556 210560 677610
rect 208960 677454 208995 677556
rect 210525 677454 210560 677556
rect 208960 677380 210560 677454
rect 208580 664911 210180 664990
rect 208580 664809 208615 664911
rect 210145 664809 210180 664911
rect 208580 664770 210180 664809
<< psubdiffcont >>
rect 208995 677454 210525 677556
rect 208615 664809 210145 664911
<< poly >>
rect 208920 678040 208960 678250
rect 208620 677996 208960 678040
rect 208620 677894 208665 677996
rect 208835 677894 208960 677996
rect 208620 677850 208960 677894
rect 210560 677850 210600 678250
rect 208540 665190 208580 665590
rect 210180 665370 210220 665590
rect 210180 665331 210440 665370
rect 210180 665229 210299 665331
rect 210401 665229 210440 665331
rect 210180 665190 210440 665229
<< polycont >>
rect 208665 677894 208835 677996
rect 210299 665229 210401 665331
<< locali >>
rect 208960 678469 210560 678580
rect 208960 678291 208987 678469
rect 210533 678291 210560 678469
rect 208960 678290 210560 678291
rect 207960 677998 208910 678020
rect 207960 677892 207980 677998
rect 208590 677996 208910 677998
rect 208590 677894 208665 677996
rect 208835 677894 208910 677996
rect 208590 677892 208910 677894
rect 207960 677870 208910 677892
rect 208960 677783 210560 677850
rect 208960 677766 209033 677783
rect 210507 677766 210560 677783
rect 208960 677664 209005 677766
rect 210535 677664 210560 677766
rect 208960 677556 210560 677664
rect 208960 677454 208995 677556
rect 210525 677454 210560 677556
rect 208960 677410 210560 677454
rect 208580 665961 210180 665990
rect 208580 665639 208607 665961
rect 210153 665639 210180 665961
rect 208580 665590 210180 665639
rect 210230 665333 210950 665350
rect 210230 665331 210457 665333
rect 210230 665229 210299 665331
rect 210401 665229 210457 665331
rect 210230 665227 210457 665229
rect 210923 665227 210950 665333
rect 210230 665210 210950 665227
rect 208580 665131 210180 665170
rect 208580 665080 208620 665131
rect 210150 665080 210180 665131
rect 208580 664830 208607 665080
rect 210153 664830 210180 665080
rect 208580 664809 208615 664830
rect 210145 664809 210180 664830
rect 208580 664780 210180 664809
<< viali >>
rect 208987 678465 210533 678469
rect 208987 678295 208995 678465
rect 208995 678295 210525 678465
rect 210525 678295 210533 678465
rect 208987 678291 210533 678295
rect 207980 677892 208590 677998
rect 209033 677766 210507 677783
rect 209033 677677 210507 677766
rect 208607 665953 210153 665961
rect 208607 665647 208615 665953
rect 208615 665647 210145 665953
rect 210145 665647 210153 665953
rect 208607 665639 210153 665647
rect 210457 665227 210923 665333
rect 208607 665029 208620 665080
rect 208620 665029 210150 665080
rect 210150 665029 210153 665080
rect 208607 664911 210153 665029
rect 208607 664830 208615 664911
rect 208615 664830 210145 664911
rect 210145 664830 210153 664911
<< metal1 >>
rect 187620 696780 251410 697300
rect 187620 695320 209762 696780
rect 210518 695320 251410 696780
rect 187620 695300 251410 695320
rect 187620 680451 189620 695300
rect 187620 680399 187877 680451
rect 187929 680399 187941 680451
rect 187993 680399 188005 680451
rect 188057 680399 188069 680451
rect 188121 680399 188133 680451
rect 188185 680399 188197 680451
rect 188249 680399 188261 680451
rect 188313 680399 188325 680451
rect 188377 680399 188389 680451
rect 188441 680399 188453 680451
rect 188505 680399 188517 680451
rect 188569 680399 188581 680451
rect 188633 680399 188645 680451
rect 188697 680399 188709 680451
rect 188761 680399 188773 680451
rect 188825 680399 188837 680451
rect 188889 680399 188901 680451
rect 188953 680399 188965 680451
rect 189017 680399 189029 680451
rect 189081 680399 189093 680451
rect 189145 680399 189157 680451
rect 189209 680399 189221 680451
rect 189273 680399 189285 680451
rect 189337 680399 189349 680451
rect 189401 680399 189413 680451
rect 189465 680399 189477 680451
rect 189529 680399 189541 680451
rect 189593 680399 189620 680451
rect 187620 658480 189620 680399
rect 191760 691140 247870 693140
rect 191760 681370 193760 691140
rect 191760 681220 199630 681370
rect 191760 676840 193760 681220
rect 200990 681105 201170 681120
rect 200990 680910 201170 680925
rect 201500 681100 201680 681110
rect 201500 680910 201680 680920
rect 200160 680493 200400 680500
rect 200160 680377 200190 680493
rect 200370 680377 200400 680493
rect 200160 680370 200400 680377
rect 205720 680360 205800 680460
rect 203600 679850 207450 680010
rect 199670 677990 199760 678000
rect 199160 677985 199910 677990
rect 202670 677985 202760 677990
rect 205670 677985 205760 678000
rect 199160 677971 205775 677985
rect 199160 677919 199689 677971
rect 199741 677966 205689 677971
rect 199741 677919 202689 677966
rect 199160 677914 202689 677919
rect 202741 677919 205689 677966
rect 205741 677919 205775 677971
rect 202741 677914 205775 677919
rect 199160 677900 205775 677914
rect 199670 677890 199760 677900
rect 202670 677890 202760 677900
rect 205670 677890 205760 677900
rect 207290 677460 207450 679850
rect 213860 679590 214570 691140
rect 208960 678470 210560 678730
rect 208960 678469 208998 678470
rect 210522 678469 210560 678470
rect 208960 678291 208987 678469
rect 210533 678291 210560 678469
rect 208960 678290 208998 678291
rect 210522 678290 210560 678291
rect 208960 678270 210560 678290
rect 207960 678003 208620 678040
rect 207960 677887 207971 678003
rect 208599 677887 208620 678003
rect 207960 677850 208620 677887
rect 208960 677800 210560 677830
rect 208960 677783 210570 677800
rect 208960 677667 209008 677783
rect 210532 677667 210570 677783
rect 208960 677660 210570 677667
rect 208960 677620 210560 677660
rect 207290 677300 208990 677460
rect 191760 676680 199270 676840
rect 191760 673840 193760 676680
rect 197782 676670 197939 676680
rect 196600 675421 199070 675440
rect 196600 675369 196621 675421
rect 196673 675369 196685 675421
rect 196737 675369 196749 675421
rect 196801 675369 196813 675421
rect 196865 675369 196877 675421
rect 196929 675369 196941 675421
rect 196993 675369 197005 675421
rect 197057 675369 197069 675421
rect 197121 675369 197133 675421
rect 197185 675369 197197 675421
rect 197249 675369 198597 675421
rect 198649 675369 198661 675421
rect 198713 675369 198725 675421
rect 198777 675369 198789 675421
rect 198841 675369 198853 675421
rect 198905 675369 198917 675421
rect 198969 675369 198981 675421
rect 199033 675369 199070 675421
rect 196600 675350 199070 675369
rect 208830 674640 208990 677300
rect 208830 674480 211090 674640
rect 208180 674009 209210 674050
rect 208180 673900 208861 674009
rect 191760 673680 199240 673840
rect 191760 670825 193760 673680
rect 197130 672421 199020 672440
rect 197130 672369 197169 672421
rect 197221 672369 197233 672421
rect 197285 672369 197297 672421
rect 197349 672369 197361 672421
rect 197413 672369 197425 672421
rect 197477 672369 197489 672421
rect 197541 672369 198557 672421
rect 198609 672369 198621 672421
rect 198673 672369 198685 672421
rect 198737 672369 198749 672421
rect 198801 672369 198813 672421
rect 198865 672369 198877 672421
rect 198929 672369 198941 672421
rect 198993 672369 199020 672421
rect 197130 672350 199020 672369
rect 208810 671050 208861 673900
rect 208180 670900 208861 671050
rect 197255 670825 199185 670840
rect 191760 670670 199185 670825
rect 191760 670668 197640 670670
rect 191760 663130 193760 670668
rect 208810 668050 208861 670900
rect 208170 667941 208861 668050
rect 209169 667941 209210 674009
rect 208170 667900 209210 667941
rect 208810 667880 209210 667900
rect 208580 665961 210180 665990
rect 208580 665639 208607 665961
rect 210153 665639 210180 665961
rect 208580 665590 210180 665639
rect 210930 665370 211090 674480
rect 210440 665333 211090 665370
rect 210440 665227 210457 665333
rect 210923 665227 211090 665333
rect 210440 665190 211090 665227
rect 210940 665180 211090 665190
rect 208580 665080 210180 665170
rect 208580 664830 208607 665080
rect 210153 664830 210180 665080
rect 208580 664770 210180 664830
rect 236140 664885 237090 667020
rect 236140 664065 236173 664885
rect 237057 664065 237090 664885
rect 236140 664040 237090 664065
rect 245870 663130 247870 691140
rect 191730 661020 247870 663130
rect 191760 661010 193760 661020
rect 245870 660130 247870 661020
rect 249410 658480 251410 695300
rect 187620 658443 251410 658480
rect 187620 658387 236178 658443
rect 187620 656863 208822 658387
rect 209578 657047 236178 658387
rect 237062 657047 251410 658443
rect 209578 656863 251410 657047
rect 187620 656480 251410 656863
<< via1 >>
rect 209762 695320 210518 696780
rect 187877 680399 187929 680451
rect 187941 680399 187993 680451
rect 188005 680399 188057 680451
rect 188069 680399 188121 680451
rect 188133 680399 188185 680451
rect 188197 680399 188249 680451
rect 188261 680399 188313 680451
rect 188325 680399 188377 680451
rect 188389 680399 188441 680451
rect 188453 680399 188505 680451
rect 188517 680399 188569 680451
rect 188581 680399 188633 680451
rect 188645 680399 188697 680451
rect 188709 680399 188761 680451
rect 188773 680399 188825 680451
rect 188837 680399 188889 680451
rect 188901 680399 188953 680451
rect 188965 680399 189017 680451
rect 189029 680399 189081 680451
rect 189093 680399 189145 680451
rect 189157 680399 189209 680451
rect 189221 680399 189273 680451
rect 189285 680399 189337 680451
rect 189349 680399 189401 680451
rect 189413 680399 189465 680451
rect 189477 680399 189529 680451
rect 189541 680399 189593 680451
rect 200990 680925 201170 681105
rect 201500 680920 201680 681100
rect 200190 680377 200370 680493
rect 199689 677919 199741 677971
rect 202689 677914 202741 677966
rect 205689 677919 205741 677971
rect 208998 678469 210522 678470
rect 208998 678291 210522 678469
rect 208998 678290 210522 678291
rect 207971 677998 208599 678003
rect 207971 677892 207980 677998
rect 207980 677892 208590 677998
rect 208590 677892 208599 677998
rect 207971 677887 208599 677892
rect 209008 677677 209033 677783
rect 209033 677677 210507 677783
rect 210507 677677 210532 677783
rect 209008 677667 210532 677677
rect 196621 675369 196673 675421
rect 196685 675369 196737 675421
rect 196749 675369 196801 675421
rect 196813 675369 196865 675421
rect 196877 675369 196929 675421
rect 196941 675369 196993 675421
rect 197005 675369 197057 675421
rect 197069 675369 197121 675421
rect 197133 675369 197185 675421
rect 197197 675369 197249 675421
rect 198597 675369 198649 675421
rect 198661 675369 198713 675421
rect 198725 675369 198777 675421
rect 198789 675369 198841 675421
rect 198853 675369 198905 675421
rect 198917 675369 198969 675421
rect 198981 675369 199033 675421
rect 197169 672369 197221 672421
rect 197233 672369 197285 672421
rect 197297 672369 197349 672421
rect 197361 672369 197413 672421
rect 197425 672369 197477 672421
rect 197489 672369 197541 672421
rect 198557 672369 198609 672421
rect 198621 672369 198673 672421
rect 198685 672369 198737 672421
rect 198749 672369 198801 672421
rect 198813 672369 198865 672421
rect 198877 672369 198929 672421
rect 198941 672369 198993 672421
rect 208861 667941 209169 674009
rect 208618 665646 210142 665954
rect 208618 664833 210142 665077
rect 236173 664065 237057 664885
rect 208822 656863 209578 658387
rect 236178 657047 237062 658443
<< metal2 >>
rect 209710 696780 210580 696800
rect 209710 695320 209762 696780
rect 210518 695320 210580 696780
rect 209710 695290 210580 695320
rect 200980 681223 201180 681280
rect 200980 681105 201012 681223
rect 201148 681105 201180 681223
rect 199090 680913 199440 680930
rect 199090 680857 199117 680913
rect 199173 680857 199197 680913
rect 199253 680857 199277 680913
rect 199333 680857 199357 680913
rect 199413 680857 199440 680913
rect 200980 680925 200990 681105
rect 201170 680925 201180 681105
rect 200980 680900 201180 680925
rect 201490 681238 201690 681320
rect 201490 681100 201522 681238
rect 201658 681100 201690 681238
rect 201490 680920 201500 681100
rect 201680 680920 201690 681100
rect 201490 680900 201690 680920
rect 199090 680840 199440 680857
rect 187855 680493 200410 680510
rect 187855 680451 200190 680493
rect 187855 680399 187877 680451
rect 187929 680399 187941 680451
rect 187993 680399 188005 680451
rect 188057 680399 188069 680451
rect 188121 680399 188133 680451
rect 188185 680399 188197 680451
rect 188249 680399 188261 680451
rect 188313 680399 188325 680451
rect 188377 680399 188389 680451
rect 188441 680399 188453 680451
rect 188505 680399 188517 680451
rect 188569 680399 188581 680451
rect 188633 680399 188645 680451
rect 188697 680399 188709 680451
rect 188761 680399 188773 680451
rect 188825 680399 188837 680451
rect 188889 680399 188901 680451
rect 188953 680399 188965 680451
rect 189017 680399 189029 680451
rect 189081 680399 189093 680451
rect 189145 680399 189157 680451
rect 189209 680399 189221 680451
rect 189273 680399 189285 680451
rect 189337 680399 189349 680451
rect 189401 680399 189413 680451
rect 189465 680399 189477 680451
rect 189529 680399 189541 680451
rect 189593 680399 200190 680451
rect 187855 680377 200190 680399
rect 200370 680377 200410 680493
rect 187855 680360 200410 680377
rect 200710 679770 200800 680430
rect 198180 679650 200800 679770
rect 196600 675423 197270 675440
rect 196600 675421 196627 675423
rect 196683 675421 196707 675423
rect 196763 675421 196787 675423
rect 196843 675421 196867 675423
rect 196923 675421 196947 675423
rect 197003 675421 197027 675423
rect 197083 675421 197107 675423
rect 197163 675421 197187 675423
rect 197243 675421 197270 675423
rect 196600 675369 196621 675421
rect 196683 675369 196685 675421
rect 196865 675369 196867 675421
rect 196929 675369 196941 675421
rect 197003 675369 197005 675421
rect 197185 675369 197187 675421
rect 197249 675369 197270 675421
rect 196600 675367 196627 675369
rect 196683 675367 196707 675369
rect 196763 675367 196787 675369
rect 196843 675367 196867 675369
rect 196923 675367 196947 675369
rect 197003 675367 197027 675369
rect 197083 675367 197107 675369
rect 197163 675367 197187 675369
rect 197243 675367 197270 675369
rect 196600 675350 197270 675367
rect 198180 674130 198300 679650
rect 201220 678520 201310 680430
rect 203660 679855 203770 680450
rect 205660 680285 205770 680625
rect 205660 680175 207655 680285
rect 200200 678435 206295 678520
rect 199680 678000 199750 678385
rect 199670 677990 199760 678000
rect 199160 677973 199910 677990
rect 199160 677917 199187 677973
rect 199243 677917 199267 677973
rect 199323 677917 199347 677973
rect 199403 677917 199427 677973
rect 199483 677917 199507 677973
rect 199563 677917 199587 677973
rect 199643 677917 199667 677973
rect 199723 677971 199747 677973
rect 199741 677919 199747 677971
rect 199723 677917 199747 677919
rect 199803 677917 199827 677973
rect 199883 677917 199910 677973
rect 199160 677900 199910 677917
rect 199670 677890 199760 677900
rect 199230 677728 199320 677780
rect 199230 677672 199247 677728
rect 199303 677672 199320 677728
rect 199230 677630 199320 677672
rect 199240 677385 199310 677630
rect 199680 677355 199750 677890
rect 200200 677355 200270 678435
rect 202670 677966 202760 677990
rect 202670 677914 202689 677966
rect 202741 677914 202760 677966
rect 202670 677890 202760 677914
rect 202230 677758 202320 677790
rect 202230 677702 202252 677758
rect 202308 677702 202320 677758
rect 202230 677680 202320 677702
rect 202240 677470 202310 677680
rect 202680 677400 202750 677890
rect 203200 677355 203270 678435
rect 205670 677971 205760 678000
rect 205670 677919 205689 677971
rect 205741 677919 205760 677971
rect 205670 677890 205760 677919
rect 205230 677758 205320 677790
rect 205230 677702 205247 677758
rect 205303 677702 205320 677758
rect 205230 677680 205320 677702
rect 205240 677470 205310 677680
rect 205680 677400 205750 677890
rect 206200 677365 206270 678435
rect 207545 678040 207655 680175
rect 208960 678550 214890 678730
rect 208960 678470 210560 678550
rect 208960 678290 208998 678470
rect 210522 678290 210560 678470
rect 208960 678270 210560 678290
rect 207545 678003 208620 678040
rect 207545 677887 207971 678003
rect 208599 677887 208620 678003
rect 207545 677850 208620 677887
rect 208960 677788 210560 677830
rect 208960 677783 209022 677788
rect 210518 677783 210560 677788
rect 208960 677667 209008 677783
rect 210532 677667 210560 677783
rect 208960 677652 209022 677667
rect 210518 677652 210560 677667
rect 208960 677620 210560 677652
rect 198390 676420 198490 677290
rect 211010 676988 215125 677110
rect 198390 676408 198570 676420
rect 198390 676352 198452 676408
rect 198508 676352 198570 676408
rect 198390 676340 198570 676352
rect 198390 674953 198490 676340
rect 211010 675572 211107 676988
rect 212523 675572 215125 676988
rect 211010 675480 215125 675572
rect 211010 675470 212640 675480
rect 198560 675423 199070 675440
rect 198560 675367 198587 675423
rect 198643 675421 198667 675423
rect 198723 675421 198747 675423
rect 198803 675421 198827 675423
rect 198883 675421 198907 675423
rect 198963 675421 198987 675423
rect 198649 675369 198661 675421
rect 198723 675369 198725 675421
rect 198905 675369 198907 675421
rect 198969 675369 198981 675421
rect 198643 675367 198667 675369
rect 198723 675367 198747 675369
rect 198803 675367 198827 675369
rect 198883 675367 198907 675369
rect 198963 675367 198987 675369
rect 199043 675367 199070 675423
rect 198560 675350 199070 675367
rect 198390 674897 198412 674953
rect 198468 674897 198490 674953
rect 198390 674873 198490 674897
rect 198390 674817 198412 674873
rect 198468 674817 198490 674873
rect 198390 674793 198490 674817
rect 198390 674737 198412 674793
rect 198468 674737 198490 674793
rect 198390 674713 198490 674737
rect 198390 674657 198412 674713
rect 198468 674657 198490 674713
rect 198390 674633 198490 674657
rect 198390 674577 198412 674633
rect 198468 674577 198490 674633
rect 198390 674553 198490 674577
rect 198390 674497 198412 674553
rect 198468 674497 198490 674553
rect 198390 674473 198490 674497
rect 198390 674417 198412 674473
rect 198468 674417 198490 674473
rect 198390 674370 198490 674417
rect 198180 674113 198590 674130
rect 198180 674057 198342 674113
rect 198398 674057 198422 674113
rect 198478 674057 198502 674113
rect 198558 674057 198590 674113
rect 198180 674040 198590 674057
rect 197130 672423 197580 672440
rect 197130 672367 197167 672423
rect 197223 672421 197247 672423
rect 197303 672421 197327 672423
rect 197383 672421 197407 672423
rect 197463 672421 197487 672423
rect 197223 672369 197233 672421
rect 197477 672369 197487 672421
rect 197223 672367 197247 672369
rect 197303 672367 197327 672369
rect 197383 672367 197407 672369
rect 197463 672367 197487 672369
rect 197543 672367 197580 672423
rect 197130 672350 197580 672367
rect 198180 671120 198300 674040
rect 208810 674009 209210 674050
rect 198520 672423 199020 672440
rect 198520 672367 198547 672423
rect 198603 672421 198627 672423
rect 198683 672421 198707 672423
rect 198763 672421 198787 672423
rect 198843 672421 198867 672423
rect 198923 672421 198947 672423
rect 198609 672369 198621 672421
rect 198683 672369 198685 672421
rect 198865 672369 198867 672421
rect 198929 672369 198941 672421
rect 198603 672367 198627 672369
rect 198683 672367 198707 672369
rect 198763 672367 198787 672369
rect 198843 672367 198867 672369
rect 198923 672367 198947 672369
rect 199003 672367 199020 672423
rect 198520 672350 199020 672367
rect 198180 671103 198780 671120
rect 198180 671047 198212 671103
rect 198268 671047 198292 671103
rect 198348 671047 198372 671103
rect 198428 671047 198452 671103
rect 198508 671047 198532 671103
rect 198588 671047 198612 671103
rect 198668 671047 198692 671103
rect 198748 671047 198780 671103
rect 198180 671030 198780 671047
rect 198180 668120 198300 671030
rect 198180 668103 198770 668120
rect 198180 668047 198202 668103
rect 198258 668047 198282 668103
rect 198338 668047 198362 668103
rect 198418 668047 198442 668103
rect 198498 668047 198522 668103
rect 198578 668047 198602 668103
rect 198658 668047 198682 668103
rect 198738 668047 198770 668103
rect 198180 668030 198770 668047
rect 198180 667970 198300 668030
rect 208810 667941 208861 674009
rect 209169 667941 209210 674009
rect 212660 672130 214030 672150
rect 208810 667912 208867 667941
rect 209163 667912 209210 667941
rect 208810 667880 209210 667912
rect 211900 671150 215120 672130
rect 211900 666970 212880 671150
rect 199730 665995 212880 666970
rect 199730 665990 210180 665995
rect 210367 665990 212880 665995
rect 208580 665954 210180 665990
rect 208580 665646 208618 665954
rect 210142 665646 210180 665954
rect 208580 665600 210180 665646
rect 208580 665077 210180 665170
rect 208580 664833 208618 665077
rect 210142 664833 210180 665077
rect 208580 664780 210180 664833
rect 236140 664885 237090 664910
rect 236140 664065 236173 664885
rect 237057 664065 237090 664885
rect 236140 658443 237090 664065
rect 208620 658387 209660 658440
rect 208620 656863 208822 658387
rect 209578 656863 209660 658387
rect 236140 657047 236178 658443
rect 237062 658340 237090 658443
rect 237062 657047 237100 658340
rect 236140 657010 237100 657047
rect 208620 656760 209660 656863
<< via2 >>
rect 209792 695342 210488 696758
rect 201012 681105 201148 681223
rect 199117 680857 199173 680913
rect 199197 680857 199253 680913
rect 199277 680857 199333 680913
rect 199357 680857 199413 680913
rect 201012 680927 201148 681105
rect 201522 681100 201658 681238
rect 201522 680942 201658 681100
rect 196627 675421 196683 675423
rect 196707 675421 196763 675423
rect 196787 675421 196843 675423
rect 196867 675421 196923 675423
rect 196947 675421 197003 675423
rect 197027 675421 197083 675423
rect 197107 675421 197163 675423
rect 197187 675421 197243 675423
rect 196627 675369 196673 675421
rect 196673 675369 196683 675421
rect 196707 675369 196737 675421
rect 196737 675369 196749 675421
rect 196749 675369 196763 675421
rect 196787 675369 196801 675421
rect 196801 675369 196813 675421
rect 196813 675369 196843 675421
rect 196867 675369 196877 675421
rect 196877 675369 196923 675421
rect 196947 675369 196993 675421
rect 196993 675369 197003 675421
rect 197027 675369 197057 675421
rect 197057 675369 197069 675421
rect 197069 675369 197083 675421
rect 197107 675369 197121 675421
rect 197121 675369 197133 675421
rect 197133 675369 197163 675421
rect 197187 675369 197197 675421
rect 197197 675369 197243 675421
rect 196627 675367 196683 675369
rect 196707 675367 196763 675369
rect 196787 675367 196843 675369
rect 196867 675367 196923 675369
rect 196947 675367 197003 675369
rect 197027 675367 197083 675369
rect 197107 675367 197163 675369
rect 197187 675367 197243 675369
rect 199187 677917 199243 677973
rect 199267 677917 199323 677973
rect 199347 677917 199403 677973
rect 199427 677917 199483 677973
rect 199507 677917 199563 677973
rect 199587 677917 199643 677973
rect 199667 677971 199723 677973
rect 199667 677919 199689 677971
rect 199689 677919 199723 677971
rect 199667 677917 199723 677919
rect 199747 677917 199803 677973
rect 199827 677917 199883 677973
rect 199247 677672 199303 677728
rect 202252 677702 202308 677758
rect 205247 677702 205303 677758
rect 209022 677783 210518 677788
rect 209022 677667 210518 677783
rect 209022 677652 210518 677667
rect 198452 676352 198508 676408
rect 211107 675572 212523 676988
rect 198587 675421 198643 675423
rect 198667 675421 198723 675423
rect 198747 675421 198803 675423
rect 198827 675421 198883 675423
rect 198907 675421 198963 675423
rect 198987 675421 199043 675423
rect 198587 675369 198597 675421
rect 198597 675369 198643 675421
rect 198667 675369 198713 675421
rect 198713 675369 198723 675421
rect 198747 675369 198777 675421
rect 198777 675369 198789 675421
rect 198789 675369 198803 675421
rect 198827 675369 198841 675421
rect 198841 675369 198853 675421
rect 198853 675369 198883 675421
rect 198907 675369 198917 675421
rect 198917 675369 198963 675421
rect 198987 675369 199033 675421
rect 199033 675369 199043 675421
rect 198587 675367 198643 675369
rect 198667 675367 198723 675369
rect 198747 675367 198803 675369
rect 198827 675367 198883 675369
rect 198907 675367 198963 675369
rect 198987 675367 199043 675369
rect 198412 674897 198468 674953
rect 198412 674817 198468 674873
rect 198412 674737 198468 674793
rect 198412 674657 198468 674713
rect 198412 674577 198468 674633
rect 198412 674497 198468 674553
rect 198412 674417 198468 674473
rect 198342 674057 198398 674113
rect 198422 674057 198478 674113
rect 198502 674057 198558 674113
rect 197167 672421 197223 672423
rect 197247 672421 197303 672423
rect 197327 672421 197383 672423
rect 197407 672421 197463 672423
rect 197487 672421 197543 672423
rect 197167 672369 197169 672421
rect 197169 672369 197221 672421
rect 197221 672369 197223 672421
rect 197247 672369 197285 672421
rect 197285 672369 197297 672421
rect 197297 672369 197303 672421
rect 197327 672369 197349 672421
rect 197349 672369 197361 672421
rect 197361 672369 197383 672421
rect 197407 672369 197413 672421
rect 197413 672369 197425 672421
rect 197425 672369 197463 672421
rect 197487 672369 197489 672421
rect 197489 672369 197541 672421
rect 197541 672369 197543 672421
rect 197167 672367 197223 672369
rect 197247 672367 197303 672369
rect 197327 672367 197383 672369
rect 197407 672367 197463 672369
rect 197487 672367 197543 672369
rect 198547 672421 198603 672423
rect 198627 672421 198683 672423
rect 198707 672421 198763 672423
rect 198787 672421 198843 672423
rect 198867 672421 198923 672423
rect 198947 672421 199003 672423
rect 198547 672369 198557 672421
rect 198557 672369 198603 672421
rect 198627 672369 198673 672421
rect 198673 672369 198683 672421
rect 198707 672369 198737 672421
rect 198737 672369 198749 672421
rect 198749 672369 198763 672421
rect 198787 672369 198801 672421
rect 198801 672369 198813 672421
rect 198813 672369 198843 672421
rect 198867 672369 198877 672421
rect 198877 672369 198923 672421
rect 198947 672369 198993 672421
rect 198993 672369 199003 672421
rect 198547 672367 198603 672369
rect 198627 672367 198683 672369
rect 198707 672367 198763 672369
rect 198787 672367 198843 672369
rect 198867 672367 198923 672369
rect 198947 672367 199003 672369
rect 198212 671047 198268 671103
rect 198292 671047 198348 671103
rect 198372 671047 198428 671103
rect 198452 671047 198508 671103
rect 198532 671047 198588 671103
rect 198612 671047 198668 671103
rect 198692 671047 198748 671103
rect 198202 668047 198258 668103
rect 198282 668047 198338 668103
rect 198362 668047 198418 668103
rect 198442 668047 198498 668103
rect 198522 668047 198578 668103
rect 198602 668047 198658 668103
rect 198682 668047 198738 668103
rect 208867 667941 209163 668448
rect 208867 667912 209163 667941
rect 208632 664847 210128 665063
rect 208852 656877 209548 658373
<< metal3 >>
rect 200980 681223 201180 701080
rect 201540 700480 201640 700490
rect 187185 680913 199440 680930
rect 187185 680857 199117 680913
rect 199173 680857 199197 680913
rect 199253 680857 199277 680913
rect 199333 680857 199357 680913
rect 199413 680857 199440 680913
rect 200980 680927 201012 681223
rect 201148 680927 201180 681223
rect 200980 680900 201180 680927
rect 201490 681238 201690 700480
rect 201490 680942 201522 681238
rect 201658 680942 201690 681238
rect 201850 681280 203450 700240
rect 201850 681170 203440 681280
rect 203850 681190 205450 700260
rect 209710 696758 210580 696800
rect 209710 695342 209792 696758
rect 210488 695342 210580 696758
rect 209710 695290 210580 695342
rect 201490 680900 201690 680942
rect 187185 680840 199440 680857
rect 200460 679925 200550 680430
rect 197985 679835 200550 679925
rect 198007 676720 198093 679835
rect 199160 677977 199910 677990
rect 199160 677913 199183 677977
rect 199247 677913 199263 677977
rect 199327 677913 199343 677977
rect 199407 677913 199423 677977
rect 199487 677913 199503 677977
rect 199567 677913 199583 677977
rect 199647 677913 199663 677977
rect 199727 677913 199743 677977
rect 199807 677913 199823 677977
rect 199887 677913 199910 677977
rect 199160 677900 199910 677913
rect 209730 677820 210560 695290
rect 199120 677775 199410 677780
rect 202230 677775 202320 677790
rect 205230 677775 205320 677790
rect 208960 677788 210560 677820
rect 199120 677762 205345 677775
rect 199120 677698 199153 677762
rect 199217 677698 199233 677762
rect 199297 677728 199313 677762
rect 199303 677698 199313 677728
rect 199377 677758 205345 677762
rect 199377 677702 202252 677758
rect 202308 677702 205247 677758
rect 205303 677702 205345 677758
rect 199377 677698 205345 677702
rect 199120 677680 199247 677698
rect 199230 677672 199247 677680
rect 199303 677690 205345 677698
rect 199303 677680 199410 677690
rect 202230 677680 202320 677690
rect 205230 677680 205320 677690
rect 199303 677672 199320 677680
rect 199230 677630 199320 677672
rect 208960 677652 209022 677788
rect 210518 677652 210560 677788
rect 208960 677630 210560 677652
rect 209730 677590 210560 677630
rect 211010 676992 212640 677110
rect 198007 676620 198880 676720
rect 198007 676617 198263 676620
rect 198007 676470 198093 676617
rect 198007 676300 198090 676470
rect 198400 676408 198850 676420
rect 198400 676352 198452 676408
rect 198508 676352 198850 676408
rect 198400 676340 198850 676352
rect 186815 675423 197270 675440
rect 186815 675367 196627 675423
rect 196683 675367 196707 675423
rect 196763 675367 196787 675423
rect 196843 675367 196867 675423
rect 196923 675367 196947 675423
rect 197003 675367 197027 675423
rect 197083 675367 197107 675423
rect 197163 675367 197187 675423
rect 197243 675367 197270 675423
rect 186815 675350 197270 675367
rect 198007 673710 198093 676300
rect 211010 675568 211103 676992
rect 212527 675568 212640 676992
rect 211010 675470 212640 675568
rect 198560 675423 199070 675440
rect 198560 675367 198587 675423
rect 198643 675367 198667 675423
rect 198723 675367 198747 675423
rect 198803 675367 198827 675423
rect 198883 675367 198907 675423
rect 198963 675367 198987 675423
rect 199043 675367 199070 675423
rect 198560 675350 199070 675367
rect 198390 674962 198490 675030
rect 198390 674898 198408 674962
rect 198472 674898 198490 674962
rect 198390 674897 198412 674898
rect 198468 674897 198490 674898
rect 198390 674882 198490 674897
rect 198390 674818 198408 674882
rect 198472 674818 198490 674882
rect 198390 674817 198412 674818
rect 198468 674817 198490 674818
rect 198390 674802 198490 674817
rect 198390 674738 198408 674802
rect 198472 674738 198490 674802
rect 198390 674737 198412 674738
rect 198468 674737 198490 674738
rect 198390 674722 198490 674737
rect 198390 674658 198408 674722
rect 198472 674658 198490 674722
rect 198390 674657 198412 674658
rect 198468 674657 198490 674658
rect 198390 674642 198490 674657
rect 198390 674578 198408 674642
rect 198472 674578 198490 674642
rect 198390 674577 198412 674578
rect 198468 674577 198490 674578
rect 198390 674562 198490 674577
rect 198390 674498 198408 674562
rect 198472 674498 198490 674562
rect 198390 674497 198412 674498
rect 198468 674497 198490 674498
rect 198390 674482 198490 674497
rect 198390 674418 198408 674482
rect 198472 674418 198490 674482
rect 198390 674417 198412 674418
rect 198468 674417 198490 674418
rect 198390 674370 198490 674417
rect 198300 674113 198880 674130
rect 198300 674057 198342 674113
rect 198398 674057 198422 674113
rect 198478 674057 198502 674113
rect 198558 674057 198880 674113
rect 198300 674040 198880 674057
rect 198007 673620 198745 673710
rect 186985 672423 197580 672440
rect 186985 672367 197167 672423
rect 197223 672367 197247 672423
rect 197303 672367 197327 672423
rect 197383 672367 197407 672423
rect 197463 672367 197487 672423
rect 197543 672367 197580 672423
rect 186985 672350 197580 672367
rect 198007 671587 198093 673620
rect 198390 673407 198990 673420
rect 198390 673343 198438 673407
rect 198502 673343 198518 673407
rect 198582 673343 198598 673407
rect 198662 673343 198678 673407
rect 198742 673343 198758 673407
rect 198822 673343 198838 673407
rect 198902 673343 198990 673407
rect 198390 673330 198990 673343
rect 198480 672430 198660 672440
rect 198480 672423 199010 672430
rect 198480 672367 198547 672423
rect 198603 672367 198627 672423
rect 198683 672367 198707 672423
rect 198763 672367 198787 672423
rect 198843 672367 198867 672423
rect 198923 672367 198947 672423
rect 199003 672367 199010 672423
rect 198480 672360 199010 672367
rect 198480 672350 198660 672360
rect 198012 670710 198088 671587
rect 198180 671103 198780 671120
rect 198180 671047 198212 671103
rect 198268 671047 198292 671103
rect 198348 671047 198372 671103
rect 198428 671047 198452 671103
rect 198508 671047 198532 671103
rect 198588 671047 198612 671103
rect 198668 671047 198692 671103
rect 198748 671047 198780 671103
rect 198180 671030 198780 671047
rect 198012 670620 198715 670710
rect 198012 670162 198088 670620
rect 198390 670407 199000 670420
rect 198390 670343 198423 670407
rect 198487 670343 198503 670407
rect 198567 670343 198583 670407
rect 198647 670343 198663 670407
rect 198727 670343 198743 670407
rect 198807 670343 198823 670407
rect 198887 670343 198903 670407
rect 198967 670343 199000 670407
rect 198390 670330 199000 670343
rect 186435 669350 199070 669440
rect 208820 668448 209210 668480
rect 198180 668103 198770 668120
rect 198180 668047 198202 668103
rect 198258 668047 198282 668103
rect 198338 668047 198362 668103
rect 198418 668047 198442 668103
rect 198498 668047 198522 668103
rect 198578 668047 198602 668103
rect 198658 668047 198682 668103
rect 198738 668047 198770 668103
rect 198180 668030 198770 668047
rect 208820 667912 208867 668448
rect 209163 667912 209210 668448
rect 208820 667872 209210 667912
rect 208820 667728 208863 667872
rect 209167 667728 209210 667872
rect 208820 667690 209210 667728
rect 208580 665140 209695 665157
rect 208570 665063 210180 665140
rect 208570 664847 208632 665063
rect 210128 664847 210180 665063
rect 208570 664770 210180 664847
rect 208580 658377 209695 664770
rect 208580 657955 208848 658377
rect 208600 656873 208848 657955
rect 209552 658075 209695 658377
rect 209552 656873 209680 658075
rect 208600 656690 209680 656873
<< via3 >>
rect 199183 677973 199247 677977
rect 199183 677917 199187 677973
rect 199187 677917 199243 677973
rect 199243 677917 199247 677973
rect 199183 677913 199247 677917
rect 199263 677973 199327 677977
rect 199263 677917 199267 677973
rect 199267 677917 199323 677973
rect 199323 677917 199327 677973
rect 199263 677913 199327 677917
rect 199343 677973 199407 677977
rect 199343 677917 199347 677973
rect 199347 677917 199403 677973
rect 199403 677917 199407 677973
rect 199343 677913 199407 677917
rect 199423 677973 199487 677977
rect 199423 677917 199427 677973
rect 199427 677917 199483 677973
rect 199483 677917 199487 677973
rect 199423 677913 199487 677917
rect 199503 677973 199567 677977
rect 199503 677917 199507 677973
rect 199507 677917 199563 677973
rect 199563 677917 199567 677973
rect 199503 677913 199567 677917
rect 199583 677973 199647 677977
rect 199583 677917 199587 677973
rect 199587 677917 199643 677973
rect 199643 677917 199647 677973
rect 199583 677913 199647 677917
rect 199663 677973 199727 677977
rect 199663 677917 199667 677973
rect 199667 677917 199723 677973
rect 199723 677917 199727 677973
rect 199663 677913 199727 677917
rect 199743 677973 199807 677977
rect 199743 677917 199747 677973
rect 199747 677917 199803 677973
rect 199803 677917 199807 677973
rect 199743 677913 199807 677917
rect 199823 677973 199887 677977
rect 199823 677917 199827 677973
rect 199827 677917 199883 677973
rect 199883 677917 199887 677973
rect 199823 677913 199887 677917
rect 199153 677698 199217 677762
rect 199233 677728 199297 677762
rect 199233 677698 199247 677728
rect 199247 677698 199297 677728
rect 199313 677698 199377 677762
rect 211103 676988 212527 676992
rect 211103 675572 211107 676988
rect 211107 675572 212523 676988
rect 212523 675572 212527 676988
rect 211103 675568 212527 675572
rect 198408 674953 198472 674962
rect 198408 674898 198412 674953
rect 198412 674898 198468 674953
rect 198468 674898 198472 674953
rect 198408 674873 198472 674882
rect 198408 674818 198412 674873
rect 198412 674818 198468 674873
rect 198468 674818 198472 674873
rect 198408 674793 198472 674802
rect 198408 674738 198412 674793
rect 198412 674738 198468 674793
rect 198468 674738 198472 674793
rect 198408 674713 198472 674722
rect 198408 674658 198412 674713
rect 198412 674658 198468 674713
rect 198468 674658 198472 674713
rect 198408 674633 198472 674642
rect 198408 674578 198412 674633
rect 198412 674578 198468 674633
rect 198468 674578 198472 674633
rect 198408 674553 198472 674562
rect 198408 674498 198412 674553
rect 198412 674498 198468 674553
rect 198468 674498 198472 674553
rect 198408 674473 198472 674482
rect 198408 674418 198412 674473
rect 198412 674418 198468 674473
rect 198468 674418 198472 674473
rect 198438 673343 198502 673407
rect 198518 673343 198582 673407
rect 198598 673343 198662 673407
rect 198678 673343 198742 673407
rect 198758 673343 198822 673407
rect 198838 673343 198902 673407
rect 198423 670343 198487 670407
rect 198503 670343 198567 670407
rect 198583 670343 198647 670407
rect 198663 670343 198727 670407
rect 198743 670343 198807 670407
rect 198823 670343 198887 670407
rect 198903 670343 198967 670407
rect 208863 667728 209167 667872
rect 208848 658373 209552 658377
rect 208848 656877 208852 658373
rect 208852 656877 209548 658373
rect 209548 656877 209552 658373
rect 208848 656873 209552 656877
<< metal4 >>
rect 211005 681705 239800 683335
rect 186835 677977 199910 677990
rect 186835 677913 199183 677977
rect 199247 677913 199263 677977
rect 199327 677913 199343 677977
rect 199407 677913 199423 677977
rect 199487 677913 199503 677977
rect 199567 677913 199583 677977
rect 199647 677913 199663 677977
rect 199727 677913 199743 677977
rect 199807 677913 199823 677977
rect 199887 677913 199910 677977
rect 186835 677900 199910 677913
rect 187270 677762 199410 677780
rect 187270 677698 199153 677762
rect 199217 677698 199233 677762
rect 199297 677698 199313 677762
rect 199377 677698 199410 677762
rect 187270 677680 199410 677698
rect 211005 677110 212635 681705
rect 211005 676992 212640 677110
rect 211005 675975 211103 676992
rect 211010 675568 211103 675975
rect 212527 675568 212640 676992
rect 238170 675970 239800 681705
rect 211010 675470 212640 675568
rect 237430 675074 239800 675970
rect 198390 674962 198490 675030
rect 198390 674898 198408 674962
rect 198472 674898 198490 674962
rect 198390 674882 198490 674898
rect 198390 674818 198408 674882
rect 198472 674818 198490 674882
rect 198390 674802 198490 674818
rect 198390 674738 198408 674802
rect 198472 674738 198490 674802
rect 198390 674722 198490 674738
rect 198390 674658 198408 674722
rect 198472 674658 198490 674722
rect 198390 674642 198490 674658
rect 198390 674578 198408 674642
rect 198472 674578 198490 674642
rect 198390 674562 198490 674578
rect 198390 674498 198408 674562
rect 198472 674498 198490 674562
rect 198390 674482 198490 674498
rect 198390 674418 198408 674482
rect 198472 674418 198490 674482
rect 198390 673420 198490 674418
rect 198390 673407 198990 673420
rect 198390 673343 198438 673407
rect 198502 673343 198518 673407
rect 198582 673343 198598 673407
rect 198662 673343 198678 673407
rect 198742 673343 198758 673407
rect 198822 673343 198838 673407
rect 198902 673343 198990 673407
rect 198390 673330 198990 673343
rect 198390 670420 198490 673330
rect 237412 671740 256224 675074
rect 238170 671690 239800 671740
rect 198390 670407 199000 670420
rect 198390 670343 198423 670407
rect 198487 670343 198503 670407
rect 198567 670343 198583 670407
rect 198647 670343 198663 670407
rect 198727 670343 198743 670407
rect 198807 670343 198823 670407
rect 198887 670343 198903 670407
rect 198967 670343 199000 670407
rect 198390 670330 199000 670343
rect 198390 653670 198490 670330
rect 208820 667872 209210 667910
rect 208820 667728 208863 667872
rect 209167 667728 209210 667872
rect 199400 653670 199620 667050
rect 202400 653670 202620 667160
rect 205400 653670 205620 667110
rect 208820 665171 209210 667728
rect 208820 658460 209210 664359
rect 208630 658377 209660 658460
rect 208630 656873 208848 658377
rect 209552 656873 209660 658377
rect 208630 656800 209660 656873
use bias  bias_0 ~/CMOS/TopmetalSe/magic
timestamp 1654639008
transform 1 0 198620 0 1 681970
box 790 -2236 7180 -220
use pixel_array  pixel_array_0 ~/CMOS/TopmetalSe/magic
timestamp 1654638764
transform 1 0 199180 0 1 673870
box -3000 -7600 9740 5750
use opamp_diego  opamp_diego_0 ~/CMOS/TopmetalSe/magic
timestamp 1654624193
transform 1 0 210841 0 1 676678
box 2069 -10028 26971 3199
<< labels >>
rlabel metal2 s 208860 673370 208860 673370 4 GND
port 1 nsew
rlabel metal1 s 197780 676780 197780 676780 4 VDD
port 2 nsew
rlabel metal1 s 192830 685030 192830 685030 4 VDD
port 2 nsew
rlabel poly s 208560 665370 208560 665370 4 OUT_IB
port 3 nsew
rlabel metal3 s 202930 699380 202930 699380 4 OUT_IB
port 3 nsew
rlabel poly s 208940 678020 208940 678020 4 AMP_IB
port 4 nsew
rlabel metal3 s 204820 699110 204820 699110 4 AMP_IB
port 4 nsew
rlabel metal4 s 239080 677340 239080 677340 4 AOUT
port 5 nsew
rlabel metal4 s 255740 673820 255740 673820 4 AOUT
port 5 nsew
rlabel metal1 s 213860 679590 214570 683520 4 VDD
port 2 nsew
rlabel metal1 s 236140 664040 237090 667020 4 GND
port 1 nsew
rlabel metal1 s 215500 657320 215500 657320 4 GND
port 1 nsew
rlabel metal3 s 198220 676640 198220 676640 4 SF_IB
port 6 nsew
rlabel metal3 s 187260 680880 187260 680880 4 SF_IB
port 6 nsew
rlabel metal2 s 200250 678210 200250 678210 4 NB2
port 7 nsew
rlabel metal3 s 201570 699900 201570 699900 4 NB2
port 7 nsew
rlabel metal3 s 187040 669390 187040 669390 4 ROW_SEL2
port 8 nsew
rlabel metal2 s 199720 678180 199720 678180 4 VBIAS
port 9 nsew
rlabel metal4 s 187050 677950 187050 677950 4 VBIAS
port 9 nsew
rlabel metal3 s 198400 674090 198400 674090 4 NB1
port 10 nsew
rlabel metal3 s 201070 699840 201070 699840 4 NB1
port 10 nsew
rlabel metal4 s 205530 655080 205530 655080 4 COL_SEL2
port 11 nsew
rlabel metal4 s 202530 654980 202530 654980 4 COL_SEL1
port 12 nsew
rlabel metal4 s 199500 654880 199500 654880 4 COL_SEL0
port 13 nsew
rlabel metal4 s 198420 654460 198420 654460 4 CSA_VREF
port 14 nsew
rlabel metal4 s 187400 677730 187400 677730 4 VREF
port 15 nsew
rlabel metal3 s 187290 672420 187290 672420 4 ROW_SEL1
port 16 nsew
rlabel metal3 s 187300 675410 187300 675410 4 ROW_SEL0
port 17 nsew
<< properties >>
string FIXED_BBOX 166434 633669 276225 704000
<< end >>
