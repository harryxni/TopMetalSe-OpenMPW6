magic
tech sky130A
magscale 1 2
timestamp 1654643737
<< pwell >>
rect -5707 -1209 5707 1209
<< nmos >>
rect -5521 109 -5431 1009
rect -5373 109 -5283 1009
rect -5225 109 -5135 1009
rect -5077 109 -4987 1009
rect -4929 109 -4839 1009
rect -4781 109 -4691 1009
rect -4633 109 -4543 1009
rect -4485 109 -4395 1009
rect -4337 109 -4247 1009
rect -4189 109 -4099 1009
rect -4041 109 -3951 1009
rect -3893 109 -3803 1009
rect -3745 109 -3655 1009
rect -3597 109 -3507 1009
rect -3449 109 -3359 1009
rect -3301 109 -3211 1009
rect -3153 109 -3063 1009
rect -3005 109 -2915 1009
rect -2857 109 -2767 1009
rect -2709 109 -2619 1009
rect -2561 109 -2471 1009
rect -2413 109 -2323 1009
rect -2265 109 -2175 1009
rect -2117 109 -2027 1009
rect -1969 109 -1879 1009
rect -1821 109 -1731 1009
rect -1673 109 -1583 1009
rect -1525 109 -1435 1009
rect -1377 109 -1287 1009
rect -1229 109 -1139 1009
rect -1081 109 -991 1009
rect -933 109 -843 1009
rect -785 109 -695 1009
rect -637 109 -547 1009
rect -489 109 -399 1009
rect -341 109 -251 1009
rect -193 109 -103 1009
rect -45 109 45 1009
rect 103 109 193 1009
rect 251 109 341 1009
rect 399 109 489 1009
rect 547 109 637 1009
rect 695 109 785 1009
rect 843 109 933 1009
rect 991 109 1081 1009
rect 1139 109 1229 1009
rect 1287 109 1377 1009
rect 1435 109 1525 1009
rect 1583 109 1673 1009
rect 1731 109 1821 1009
rect 1879 109 1969 1009
rect 2027 109 2117 1009
rect 2175 109 2265 1009
rect 2323 109 2413 1009
rect 2471 109 2561 1009
rect 2619 109 2709 1009
rect 2767 109 2857 1009
rect 2915 109 3005 1009
rect 3063 109 3153 1009
rect 3211 109 3301 1009
rect 3359 109 3449 1009
rect 3507 109 3597 1009
rect 3655 109 3745 1009
rect 3803 109 3893 1009
rect 3951 109 4041 1009
rect 4099 109 4189 1009
rect 4247 109 4337 1009
rect 4395 109 4485 1009
rect 4543 109 4633 1009
rect 4691 109 4781 1009
rect 4839 109 4929 1009
rect 4987 109 5077 1009
rect 5135 109 5225 1009
rect 5283 109 5373 1009
rect 5431 109 5521 1009
rect -5521 -1009 -5431 -109
rect -5373 -1009 -5283 -109
rect -5225 -1009 -5135 -109
rect -5077 -1009 -4987 -109
rect -4929 -1009 -4839 -109
rect -4781 -1009 -4691 -109
rect -4633 -1009 -4543 -109
rect -4485 -1009 -4395 -109
rect -4337 -1009 -4247 -109
rect -4189 -1009 -4099 -109
rect -4041 -1009 -3951 -109
rect -3893 -1009 -3803 -109
rect -3745 -1009 -3655 -109
rect -3597 -1009 -3507 -109
rect -3449 -1009 -3359 -109
rect -3301 -1009 -3211 -109
rect -3153 -1009 -3063 -109
rect -3005 -1009 -2915 -109
rect -2857 -1009 -2767 -109
rect -2709 -1009 -2619 -109
rect -2561 -1009 -2471 -109
rect -2413 -1009 -2323 -109
rect -2265 -1009 -2175 -109
rect -2117 -1009 -2027 -109
rect -1969 -1009 -1879 -109
rect -1821 -1009 -1731 -109
rect -1673 -1009 -1583 -109
rect -1525 -1009 -1435 -109
rect -1377 -1009 -1287 -109
rect -1229 -1009 -1139 -109
rect -1081 -1009 -991 -109
rect -933 -1009 -843 -109
rect -785 -1009 -695 -109
rect -637 -1009 -547 -109
rect -489 -1009 -399 -109
rect -341 -1009 -251 -109
rect -193 -1009 -103 -109
rect -45 -1009 45 -109
rect 103 -1009 193 -109
rect 251 -1009 341 -109
rect 399 -1009 489 -109
rect 547 -1009 637 -109
rect 695 -1009 785 -109
rect 843 -1009 933 -109
rect 991 -1009 1081 -109
rect 1139 -1009 1229 -109
rect 1287 -1009 1377 -109
rect 1435 -1009 1525 -109
rect 1583 -1009 1673 -109
rect 1731 -1009 1821 -109
rect 1879 -1009 1969 -109
rect 2027 -1009 2117 -109
rect 2175 -1009 2265 -109
rect 2323 -1009 2413 -109
rect 2471 -1009 2561 -109
rect 2619 -1009 2709 -109
rect 2767 -1009 2857 -109
rect 2915 -1009 3005 -109
rect 3063 -1009 3153 -109
rect 3211 -1009 3301 -109
rect 3359 -1009 3449 -109
rect 3507 -1009 3597 -109
rect 3655 -1009 3745 -109
rect 3803 -1009 3893 -109
rect 3951 -1009 4041 -109
rect 4099 -1009 4189 -109
rect 4247 -1009 4337 -109
rect 4395 -1009 4485 -109
rect 4543 -1009 4633 -109
rect 4691 -1009 4781 -109
rect 4839 -1009 4929 -109
rect 4987 -1009 5077 -109
rect 5135 -1009 5225 -109
rect 5283 -1009 5373 -109
rect 5431 -1009 5521 -109
<< ndiff >>
rect -5579 984 -5521 1009
rect -5579 950 -5567 984
rect -5533 950 -5521 984
rect -5579 916 -5521 950
rect -5579 882 -5567 916
rect -5533 882 -5521 916
rect -5579 848 -5521 882
rect -5579 814 -5567 848
rect -5533 814 -5521 848
rect -5579 780 -5521 814
rect -5579 746 -5567 780
rect -5533 746 -5521 780
rect -5579 712 -5521 746
rect -5579 678 -5567 712
rect -5533 678 -5521 712
rect -5579 644 -5521 678
rect -5579 610 -5567 644
rect -5533 610 -5521 644
rect -5579 576 -5521 610
rect -5579 542 -5567 576
rect -5533 542 -5521 576
rect -5579 508 -5521 542
rect -5579 474 -5567 508
rect -5533 474 -5521 508
rect -5579 440 -5521 474
rect -5579 406 -5567 440
rect -5533 406 -5521 440
rect -5579 372 -5521 406
rect -5579 338 -5567 372
rect -5533 338 -5521 372
rect -5579 304 -5521 338
rect -5579 270 -5567 304
rect -5533 270 -5521 304
rect -5579 236 -5521 270
rect -5579 202 -5567 236
rect -5533 202 -5521 236
rect -5579 168 -5521 202
rect -5579 134 -5567 168
rect -5533 134 -5521 168
rect -5579 109 -5521 134
rect -5431 984 -5373 1009
rect -5431 950 -5419 984
rect -5385 950 -5373 984
rect -5431 916 -5373 950
rect -5431 882 -5419 916
rect -5385 882 -5373 916
rect -5431 848 -5373 882
rect -5431 814 -5419 848
rect -5385 814 -5373 848
rect -5431 780 -5373 814
rect -5431 746 -5419 780
rect -5385 746 -5373 780
rect -5431 712 -5373 746
rect -5431 678 -5419 712
rect -5385 678 -5373 712
rect -5431 644 -5373 678
rect -5431 610 -5419 644
rect -5385 610 -5373 644
rect -5431 576 -5373 610
rect -5431 542 -5419 576
rect -5385 542 -5373 576
rect -5431 508 -5373 542
rect -5431 474 -5419 508
rect -5385 474 -5373 508
rect -5431 440 -5373 474
rect -5431 406 -5419 440
rect -5385 406 -5373 440
rect -5431 372 -5373 406
rect -5431 338 -5419 372
rect -5385 338 -5373 372
rect -5431 304 -5373 338
rect -5431 270 -5419 304
rect -5385 270 -5373 304
rect -5431 236 -5373 270
rect -5431 202 -5419 236
rect -5385 202 -5373 236
rect -5431 168 -5373 202
rect -5431 134 -5419 168
rect -5385 134 -5373 168
rect -5431 109 -5373 134
rect -5283 984 -5225 1009
rect -5283 950 -5271 984
rect -5237 950 -5225 984
rect -5283 916 -5225 950
rect -5283 882 -5271 916
rect -5237 882 -5225 916
rect -5283 848 -5225 882
rect -5283 814 -5271 848
rect -5237 814 -5225 848
rect -5283 780 -5225 814
rect -5283 746 -5271 780
rect -5237 746 -5225 780
rect -5283 712 -5225 746
rect -5283 678 -5271 712
rect -5237 678 -5225 712
rect -5283 644 -5225 678
rect -5283 610 -5271 644
rect -5237 610 -5225 644
rect -5283 576 -5225 610
rect -5283 542 -5271 576
rect -5237 542 -5225 576
rect -5283 508 -5225 542
rect -5283 474 -5271 508
rect -5237 474 -5225 508
rect -5283 440 -5225 474
rect -5283 406 -5271 440
rect -5237 406 -5225 440
rect -5283 372 -5225 406
rect -5283 338 -5271 372
rect -5237 338 -5225 372
rect -5283 304 -5225 338
rect -5283 270 -5271 304
rect -5237 270 -5225 304
rect -5283 236 -5225 270
rect -5283 202 -5271 236
rect -5237 202 -5225 236
rect -5283 168 -5225 202
rect -5283 134 -5271 168
rect -5237 134 -5225 168
rect -5283 109 -5225 134
rect -5135 984 -5077 1009
rect -5135 950 -5123 984
rect -5089 950 -5077 984
rect -5135 916 -5077 950
rect -5135 882 -5123 916
rect -5089 882 -5077 916
rect -5135 848 -5077 882
rect -5135 814 -5123 848
rect -5089 814 -5077 848
rect -5135 780 -5077 814
rect -5135 746 -5123 780
rect -5089 746 -5077 780
rect -5135 712 -5077 746
rect -5135 678 -5123 712
rect -5089 678 -5077 712
rect -5135 644 -5077 678
rect -5135 610 -5123 644
rect -5089 610 -5077 644
rect -5135 576 -5077 610
rect -5135 542 -5123 576
rect -5089 542 -5077 576
rect -5135 508 -5077 542
rect -5135 474 -5123 508
rect -5089 474 -5077 508
rect -5135 440 -5077 474
rect -5135 406 -5123 440
rect -5089 406 -5077 440
rect -5135 372 -5077 406
rect -5135 338 -5123 372
rect -5089 338 -5077 372
rect -5135 304 -5077 338
rect -5135 270 -5123 304
rect -5089 270 -5077 304
rect -5135 236 -5077 270
rect -5135 202 -5123 236
rect -5089 202 -5077 236
rect -5135 168 -5077 202
rect -5135 134 -5123 168
rect -5089 134 -5077 168
rect -5135 109 -5077 134
rect -4987 984 -4929 1009
rect -4987 950 -4975 984
rect -4941 950 -4929 984
rect -4987 916 -4929 950
rect -4987 882 -4975 916
rect -4941 882 -4929 916
rect -4987 848 -4929 882
rect -4987 814 -4975 848
rect -4941 814 -4929 848
rect -4987 780 -4929 814
rect -4987 746 -4975 780
rect -4941 746 -4929 780
rect -4987 712 -4929 746
rect -4987 678 -4975 712
rect -4941 678 -4929 712
rect -4987 644 -4929 678
rect -4987 610 -4975 644
rect -4941 610 -4929 644
rect -4987 576 -4929 610
rect -4987 542 -4975 576
rect -4941 542 -4929 576
rect -4987 508 -4929 542
rect -4987 474 -4975 508
rect -4941 474 -4929 508
rect -4987 440 -4929 474
rect -4987 406 -4975 440
rect -4941 406 -4929 440
rect -4987 372 -4929 406
rect -4987 338 -4975 372
rect -4941 338 -4929 372
rect -4987 304 -4929 338
rect -4987 270 -4975 304
rect -4941 270 -4929 304
rect -4987 236 -4929 270
rect -4987 202 -4975 236
rect -4941 202 -4929 236
rect -4987 168 -4929 202
rect -4987 134 -4975 168
rect -4941 134 -4929 168
rect -4987 109 -4929 134
rect -4839 984 -4781 1009
rect -4839 950 -4827 984
rect -4793 950 -4781 984
rect -4839 916 -4781 950
rect -4839 882 -4827 916
rect -4793 882 -4781 916
rect -4839 848 -4781 882
rect -4839 814 -4827 848
rect -4793 814 -4781 848
rect -4839 780 -4781 814
rect -4839 746 -4827 780
rect -4793 746 -4781 780
rect -4839 712 -4781 746
rect -4839 678 -4827 712
rect -4793 678 -4781 712
rect -4839 644 -4781 678
rect -4839 610 -4827 644
rect -4793 610 -4781 644
rect -4839 576 -4781 610
rect -4839 542 -4827 576
rect -4793 542 -4781 576
rect -4839 508 -4781 542
rect -4839 474 -4827 508
rect -4793 474 -4781 508
rect -4839 440 -4781 474
rect -4839 406 -4827 440
rect -4793 406 -4781 440
rect -4839 372 -4781 406
rect -4839 338 -4827 372
rect -4793 338 -4781 372
rect -4839 304 -4781 338
rect -4839 270 -4827 304
rect -4793 270 -4781 304
rect -4839 236 -4781 270
rect -4839 202 -4827 236
rect -4793 202 -4781 236
rect -4839 168 -4781 202
rect -4839 134 -4827 168
rect -4793 134 -4781 168
rect -4839 109 -4781 134
rect -4691 984 -4633 1009
rect -4691 950 -4679 984
rect -4645 950 -4633 984
rect -4691 916 -4633 950
rect -4691 882 -4679 916
rect -4645 882 -4633 916
rect -4691 848 -4633 882
rect -4691 814 -4679 848
rect -4645 814 -4633 848
rect -4691 780 -4633 814
rect -4691 746 -4679 780
rect -4645 746 -4633 780
rect -4691 712 -4633 746
rect -4691 678 -4679 712
rect -4645 678 -4633 712
rect -4691 644 -4633 678
rect -4691 610 -4679 644
rect -4645 610 -4633 644
rect -4691 576 -4633 610
rect -4691 542 -4679 576
rect -4645 542 -4633 576
rect -4691 508 -4633 542
rect -4691 474 -4679 508
rect -4645 474 -4633 508
rect -4691 440 -4633 474
rect -4691 406 -4679 440
rect -4645 406 -4633 440
rect -4691 372 -4633 406
rect -4691 338 -4679 372
rect -4645 338 -4633 372
rect -4691 304 -4633 338
rect -4691 270 -4679 304
rect -4645 270 -4633 304
rect -4691 236 -4633 270
rect -4691 202 -4679 236
rect -4645 202 -4633 236
rect -4691 168 -4633 202
rect -4691 134 -4679 168
rect -4645 134 -4633 168
rect -4691 109 -4633 134
rect -4543 984 -4485 1009
rect -4543 950 -4531 984
rect -4497 950 -4485 984
rect -4543 916 -4485 950
rect -4543 882 -4531 916
rect -4497 882 -4485 916
rect -4543 848 -4485 882
rect -4543 814 -4531 848
rect -4497 814 -4485 848
rect -4543 780 -4485 814
rect -4543 746 -4531 780
rect -4497 746 -4485 780
rect -4543 712 -4485 746
rect -4543 678 -4531 712
rect -4497 678 -4485 712
rect -4543 644 -4485 678
rect -4543 610 -4531 644
rect -4497 610 -4485 644
rect -4543 576 -4485 610
rect -4543 542 -4531 576
rect -4497 542 -4485 576
rect -4543 508 -4485 542
rect -4543 474 -4531 508
rect -4497 474 -4485 508
rect -4543 440 -4485 474
rect -4543 406 -4531 440
rect -4497 406 -4485 440
rect -4543 372 -4485 406
rect -4543 338 -4531 372
rect -4497 338 -4485 372
rect -4543 304 -4485 338
rect -4543 270 -4531 304
rect -4497 270 -4485 304
rect -4543 236 -4485 270
rect -4543 202 -4531 236
rect -4497 202 -4485 236
rect -4543 168 -4485 202
rect -4543 134 -4531 168
rect -4497 134 -4485 168
rect -4543 109 -4485 134
rect -4395 984 -4337 1009
rect -4395 950 -4383 984
rect -4349 950 -4337 984
rect -4395 916 -4337 950
rect -4395 882 -4383 916
rect -4349 882 -4337 916
rect -4395 848 -4337 882
rect -4395 814 -4383 848
rect -4349 814 -4337 848
rect -4395 780 -4337 814
rect -4395 746 -4383 780
rect -4349 746 -4337 780
rect -4395 712 -4337 746
rect -4395 678 -4383 712
rect -4349 678 -4337 712
rect -4395 644 -4337 678
rect -4395 610 -4383 644
rect -4349 610 -4337 644
rect -4395 576 -4337 610
rect -4395 542 -4383 576
rect -4349 542 -4337 576
rect -4395 508 -4337 542
rect -4395 474 -4383 508
rect -4349 474 -4337 508
rect -4395 440 -4337 474
rect -4395 406 -4383 440
rect -4349 406 -4337 440
rect -4395 372 -4337 406
rect -4395 338 -4383 372
rect -4349 338 -4337 372
rect -4395 304 -4337 338
rect -4395 270 -4383 304
rect -4349 270 -4337 304
rect -4395 236 -4337 270
rect -4395 202 -4383 236
rect -4349 202 -4337 236
rect -4395 168 -4337 202
rect -4395 134 -4383 168
rect -4349 134 -4337 168
rect -4395 109 -4337 134
rect -4247 984 -4189 1009
rect -4247 950 -4235 984
rect -4201 950 -4189 984
rect -4247 916 -4189 950
rect -4247 882 -4235 916
rect -4201 882 -4189 916
rect -4247 848 -4189 882
rect -4247 814 -4235 848
rect -4201 814 -4189 848
rect -4247 780 -4189 814
rect -4247 746 -4235 780
rect -4201 746 -4189 780
rect -4247 712 -4189 746
rect -4247 678 -4235 712
rect -4201 678 -4189 712
rect -4247 644 -4189 678
rect -4247 610 -4235 644
rect -4201 610 -4189 644
rect -4247 576 -4189 610
rect -4247 542 -4235 576
rect -4201 542 -4189 576
rect -4247 508 -4189 542
rect -4247 474 -4235 508
rect -4201 474 -4189 508
rect -4247 440 -4189 474
rect -4247 406 -4235 440
rect -4201 406 -4189 440
rect -4247 372 -4189 406
rect -4247 338 -4235 372
rect -4201 338 -4189 372
rect -4247 304 -4189 338
rect -4247 270 -4235 304
rect -4201 270 -4189 304
rect -4247 236 -4189 270
rect -4247 202 -4235 236
rect -4201 202 -4189 236
rect -4247 168 -4189 202
rect -4247 134 -4235 168
rect -4201 134 -4189 168
rect -4247 109 -4189 134
rect -4099 984 -4041 1009
rect -4099 950 -4087 984
rect -4053 950 -4041 984
rect -4099 916 -4041 950
rect -4099 882 -4087 916
rect -4053 882 -4041 916
rect -4099 848 -4041 882
rect -4099 814 -4087 848
rect -4053 814 -4041 848
rect -4099 780 -4041 814
rect -4099 746 -4087 780
rect -4053 746 -4041 780
rect -4099 712 -4041 746
rect -4099 678 -4087 712
rect -4053 678 -4041 712
rect -4099 644 -4041 678
rect -4099 610 -4087 644
rect -4053 610 -4041 644
rect -4099 576 -4041 610
rect -4099 542 -4087 576
rect -4053 542 -4041 576
rect -4099 508 -4041 542
rect -4099 474 -4087 508
rect -4053 474 -4041 508
rect -4099 440 -4041 474
rect -4099 406 -4087 440
rect -4053 406 -4041 440
rect -4099 372 -4041 406
rect -4099 338 -4087 372
rect -4053 338 -4041 372
rect -4099 304 -4041 338
rect -4099 270 -4087 304
rect -4053 270 -4041 304
rect -4099 236 -4041 270
rect -4099 202 -4087 236
rect -4053 202 -4041 236
rect -4099 168 -4041 202
rect -4099 134 -4087 168
rect -4053 134 -4041 168
rect -4099 109 -4041 134
rect -3951 984 -3893 1009
rect -3951 950 -3939 984
rect -3905 950 -3893 984
rect -3951 916 -3893 950
rect -3951 882 -3939 916
rect -3905 882 -3893 916
rect -3951 848 -3893 882
rect -3951 814 -3939 848
rect -3905 814 -3893 848
rect -3951 780 -3893 814
rect -3951 746 -3939 780
rect -3905 746 -3893 780
rect -3951 712 -3893 746
rect -3951 678 -3939 712
rect -3905 678 -3893 712
rect -3951 644 -3893 678
rect -3951 610 -3939 644
rect -3905 610 -3893 644
rect -3951 576 -3893 610
rect -3951 542 -3939 576
rect -3905 542 -3893 576
rect -3951 508 -3893 542
rect -3951 474 -3939 508
rect -3905 474 -3893 508
rect -3951 440 -3893 474
rect -3951 406 -3939 440
rect -3905 406 -3893 440
rect -3951 372 -3893 406
rect -3951 338 -3939 372
rect -3905 338 -3893 372
rect -3951 304 -3893 338
rect -3951 270 -3939 304
rect -3905 270 -3893 304
rect -3951 236 -3893 270
rect -3951 202 -3939 236
rect -3905 202 -3893 236
rect -3951 168 -3893 202
rect -3951 134 -3939 168
rect -3905 134 -3893 168
rect -3951 109 -3893 134
rect -3803 984 -3745 1009
rect -3803 950 -3791 984
rect -3757 950 -3745 984
rect -3803 916 -3745 950
rect -3803 882 -3791 916
rect -3757 882 -3745 916
rect -3803 848 -3745 882
rect -3803 814 -3791 848
rect -3757 814 -3745 848
rect -3803 780 -3745 814
rect -3803 746 -3791 780
rect -3757 746 -3745 780
rect -3803 712 -3745 746
rect -3803 678 -3791 712
rect -3757 678 -3745 712
rect -3803 644 -3745 678
rect -3803 610 -3791 644
rect -3757 610 -3745 644
rect -3803 576 -3745 610
rect -3803 542 -3791 576
rect -3757 542 -3745 576
rect -3803 508 -3745 542
rect -3803 474 -3791 508
rect -3757 474 -3745 508
rect -3803 440 -3745 474
rect -3803 406 -3791 440
rect -3757 406 -3745 440
rect -3803 372 -3745 406
rect -3803 338 -3791 372
rect -3757 338 -3745 372
rect -3803 304 -3745 338
rect -3803 270 -3791 304
rect -3757 270 -3745 304
rect -3803 236 -3745 270
rect -3803 202 -3791 236
rect -3757 202 -3745 236
rect -3803 168 -3745 202
rect -3803 134 -3791 168
rect -3757 134 -3745 168
rect -3803 109 -3745 134
rect -3655 984 -3597 1009
rect -3655 950 -3643 984
rect -3609 950 -3597 984
rect -3655 916 -3597 950
rect -3655 882 -3643 916
rect -3609 882 -3597 916
rect -3655 848 -3597 882
rect -3655 814 -3643 848
rect -3609 814 -3597 848
rect -3655 780 -3597 814
rect -3655 746 -3643 780
rect -3609 746 -3597 780
rect -3655 712 -3597 746
rect -3655 678 -3643 712
rect -3609 678 -3597 712
rect -3655 644 -3597 678
rect -3655 610 -3643 644
rect -3609 610 -3597 644
rect -3655 576 -3597 610
rect -3655 542 -3643 576
rect -3609 542 -3597 576
rect -3655 508 -3597 542
rect -3655 474 -3643 508
rect -3609 474 -3597 508
rect -3655 440 -3597 474
rect -3655 406 -3643 440
rect -3609 406 -3597 440
rect -3655 372 -3597 406
rect -3655 338 -3643 372
rect -3609 338 -3597 372
rect -3655 304 -3597 338
rect -3655 270 -3643 304
rect -3609 270 -3597 304
rect -3655 236 -3597 270
rect -3655 202 -3643 236
rect -3609 202 -3597 236
rect -3655 168 -3597 202
rect -3655 134 -3643 168
rect -3609 134 -3597 168
rect -3655 109 -3597 134
rect -3507 984 -3449 1009
rect -3507 950 -3495 984
rect -3461 950 -3449 984
rect -3507 916 -3449 950
rect -3507 882 -3495 916
rect -3461 882 -3449 916
rect -3507 848 -3449 882
rect -3507 814 -3495 848
rect -3461 814 -3449 848
rect -3507 780 -3449 814
rect -3507 746 -3495 780
rect -3461 746 -3449 780
rect -3507 712 -3449 746
rect -3507 678 -3495 712
rect -3461 678 -3449 712
rect -3507 644 -3449 678
rect -3507 610 -3495 644
rect -3461 610 -3449 644
rect -3507 576 -3449 610
rect -3507 542 -3495 576
rect -3461 542 -3449 576
rect -3507 508 -3449 542
rect -3507 474 -3495 508
rect -3461 474 -3449 508
rect -3507 440 -3449 474
rect -3507 406 -3495 440
rect -3461 406 -3449 440
rect -3507 372 -3449 406
rect -3507 338 -3495 372
rect -3461 338 -3449 372
rect -3507 304 -3449 338
rect -3507 270 -3495 304
rect -3461 270 -3449 304
rect -3507 236 -3449 270
rect -3507 202 -3495 236
rect -3461 202 -3449 236
rect -3507 168 -3449 202
rect -3507 134 -3495 168
rect -3461 134 -3449 168
rect -3507 109 -3449 134
rect -3359 984 -3301 1009
rect -3359 950 -3347 984
rect -3313 950 -3301 984
rect -3359 916 -3301 950
rect -3359 882 -3347 916
rect -3313 882 -3301 916
rect -3359 848 -3301 882
rect -3359 814 -3347 848
rect -3313 814 -3301 848
rect -3359 780 -3301 814
rect -3359 746 -3347 780
rect -3313 746 -3301 780
rect -3359 712 -3301 746
rect -3359 678 -3347 712
rect -3313 678 -3301 712
rect -3359 644 -3301 678
rect -3359 610 -3347 644
rect -3313 610 -3301 644
rect -3359 576 -3301 610
rect -3359 542 -3347 576
rect -3313 542 -3301 576
rect -3359 508 -3301 542
rect -3359 474 -3347 508
rect -3313 474 -3301 508
rect -3359 440 -3301 474
rect -3359 406 -3347 440
rect -3313 406 -3301 440
rect -3359 372 -3301 406
rect -3359 338 -3347 372
rect -3313 338 -3301 372
rect -3359 304 -3301 338
rect -3359 270 -3347 304
rect -3313 270 -3301 304
rect -3359 236 -3301 270
rect -3359 202 -3347 236
rect -3313 202 -3301 236
rect -3359 168 -3301 202
rect -3359 134 -3347 168
rect -3313 134 -3301 168
rect -3359 109 -3301 134
rect -3211 984 -3153 1009
rect -3211 950 -3199 984
rect -3165 950 -3153 984
rect -3211 916 -3153 950
rect -3211 882 -3199 916
rect -3165 882 -3153 916
rect -3211 848 -3153 882
rect -3211 814 -3199 848
rect -3165 814 -3153 848
rect -3211 780 -3153 814
rect -3211 746 -3199 780
rect -3165 746 -3153 780
rect -3211 712 -3153 746
rect -3211 678 -3199 712
rect -3165 678 -3153 712
rect -3211 644 -3153 678
rect -3211 610 -3199 644
rect -3165 610 -3153 644
rect -3211 576 -3153 610
rect -3211 542 -3199 576
rect -3165 542 -3153 576
rect -3211 508 -3153 542
rect -3211 474 -3199 508
rect -3165 474 -3153 508
rect -3211 440 -3153 474
rect -3211 406 -3199 440
rect -3165 406 -3153 440
rect -3211 372 -3153 406
rect -3211 338 -3199 372
rect -3165 338 -3153 372
rect -3211 304 -3153 338
rect -3211 270 -3199 304
rect -3165 270 -3153 304
rect -3211 236 -3153 270
rect -3211 202 -3199 236
rect -3165 202 -3153 236
rect -3211 168 -3153 202
rect -3211 134 -3199 168
rect -3165 134 -3153 168
rect -3211 109 -3153 134
rect -3063 984 -3005 1009
rect -3063 950 -3051 984
rect -3017 950 -3005 984
rect -3063 916 -3005 950
rect -3063 882 -3051 916
rect -3017 882 -3005 916
rect -3063 848 -3005 882
rect -3063 814 -3051 848
rect -3017 814 -3005 848
rect -3063 780 -3005 814
rect -3063 746 -3051 780
rect -3017 746 -3005 780
rect -3063 712 -3005 746
rect -3063 678 -3051 712
rect -3017 678 -3005 712
rect -3063 644 -3005 678
rect -3063 610 -3051 644
rect -3017 610 -3005 644
rect -3063 576 -3005 610
rect -3063 542 -3051 576
rect -3017 542 -3005 576
rect -3063 508 -3005 542
rect -3063 474 -3051 508
rect -3017 474 -3005 508
rect -3063 440 -3005 474
rect -3063 406 -3051 440
rect -3017 406 -3005 440
rect -3063 372 -3005 406
rect -3063 338 -3051 372
rect -3017 338 -3005 372
rect -3063 304 -3005 338
rect -3063 270 -3051 304
rect -3017 270 -3005 304
rect -3063 236 -3005 270
rect -3063 202 -3051 236
rect -3017 202 -3005 236
rect -3063 168 -3005 202
rect -3063 134 -3051 168
rect -3017 134 -3005 168
rect -3063 109 -3005 134
rect -2915 984 -2857 1009
rect -2915 950 -2903 984
rect -2869 950 -2857 984
rect -2915 916 -2857 950
rect -2915 882 -2903 916
rect -2869 882 -2857 916
rect -2915 848 -2857 882
rect -2915 814 -2903 848
rect -2869 814 -2857 848
rect -2915 780 -2857 814
rect -2915 746 -2903 780
rect -2869 746 -2857 780
rect -2915 712 -2857 746
rect -2915 678 -2903 712
rect -2869 678 -2857 712
rect -2915 644 -2857 678
rect -2915 610 -2903 644
rect -2869 610 -2857 644
rect -2915 576 -2857 610
rect -2915 542 -2903 576
rect -2869 542 -2857 576
rect -2915 508 -2857 542
rect -2915 474 -2903 508
rect -2869 474 -2857 508
rect -2915 440 -2857 474
rect -2915 406 -2903 440
rect -2869 406 -2857 440
rect -2915 372 -2857 406
rect -2915 338 -2903 372
rect -2869 338 -2857 372
rect -2915 304 -2857 338
rect -2915 270 -2903 304
rect -2869 270 -2857 304
rect -2915 236 -2857 270
rect -2915 202 -2903 236
rect -2869 202 -2857 236
rect -2915 168 -2857 202
rect -2915 134 -2903 168
rect -2869 134 -2857 168
rect -2915 109 -2857 134
rect -2767 984 -2709 1009
rect -2767 950 -2755 984
rect -2721 950 -2709 984
rect -2767 916 -2709 950
rect -2767 882 -2755 916
rect -2721 882 -2709 916
rect -2767 848 -2709 882
rect -2767 814 -2755 848
rect -2721 814 -2709 848
rect -2767 780 -2709 814
rect -2767 746 -2755 780
rect -2721 746 -2709 780
rect -2767 712 -2709 746
rect -2767 678 -2755 712
rect -2721 678 -2709 712
rect -2767 644 -2709 678
rect -2767 610 -2755 644
rect -2721 610 -2709 644
rect -2767 576 -2709 610
rect -2767 542 -2755 576
rect -2721 542 -2709 576
rect -2767 508 -2709 542
rect -2767 474 -2755 508
rect -2721 474 -2709 508
rect -2767 440 -2709 474
rect -2767 406 -2755 440
rect -2721 406 -2709 440
rect -2767 372 -2709 406
rect -2767 338 -2755 372
rect -2721 338 -2709 372
rect -2767 304 -2709 338
rect -2767 270 -2755 304
rect -2721 270 -2709 304
rect -2767 236 -2709 270
rect -2767 202 -2755 236
rect -2721 202 -2709 236
rect -2767 168 -2709 202
rect -2767 134 -2755 168
rect -2721 134 -2709 168
rect -2767 109 -2709 134
rect -2619 984 -2561 1009
rect -2619 950 -2607 984
rect -2573 950 -2561 984
rect -2619 916 -2561 950
rect -2619 882 -2607 916
rect -2573 882 -2561 916
rect -2619 848 -2561 882
rect -2619 814 -2607 848
rect -2573 814 -2561 848
rect -2619 780 -2561 814
rect -2619 746 -2607 780
rect -2573 746 -2561 780
rect -2619 712 -2561 746
rect -2619 678 -2607 712
rect -2573 678 -2561 712
rect -2619 644 -2561 678
rect -2619 610 -2607 644
rect -2573 610 -2561 644
rect -2619 576 -2561 610
rect -2619 542 -2607 576
rect -2573 542 -2561 576
rect -2619 508 -2561 542
rect -2619 474 -2607 508
rect -2573 474 -2561 508
rect -2619 440 -2561 474
rect -2619 406 -2607 440
rect -2573 406 -2561 440
rect -2619 372 -2561 406
rect -2619 338 -2607 372
rect -2573 338 -2561 372
rect -2619 304 -2561 338
rect -2619 270 -2607 304
rect -2573 270 -2561 304
rect -2619 236 -2561 270
rect -2619 202 -2607 236
rect -2573 202 -2561 236
rect -2619 168 -2561 202
rect -2619 134 -2607 168
rect -2573 134 -2561 168
rect -2619 109 -2561 134
rect -2471 984 -2413 1009
rect -2471 950 -2459 984
rect -2425 950 -2413 984
rect -2471 916 -2413 950
rect -2471 882 -2459 916
rect -2425 882 -2413 916
rect -2471 848 -2413 882
rect -2471 814 -2459 848
rect -2425 814 -2413 848
rect -2471 780 -2413 814
rect -2471 746 -2459 780
rect -2425 746 -2413 780
rect -2471 712 -2413 746
rect -2471 678 -2459 712
rect -2425 678 -2413 712
rect -2471 644 -2413 678
rect -2471 610 -2459 644
rect -2425 610 -2413 644
rect -2471 576 -2413 610
rect -2471 542 -2459 576
rect -2425 542 -2413 576
rect -2471 508 -2413 542
rect -2471 474 -2459 508
rect -2425 474 -2413 508
rect -2471 440 -2413 474
rect -2471 406 -2459 440
rect -2425 406 -2413 440
rect -2471 372 -2413 406
rect -2471 338 -2459 372
rect -2425 338 -2413 372
rect -2471 304 -2413 338
rect -2471 270 -2459 304
rect -2425 270 -2413 304
rect -2471 236 -2413 270
rect -2471 202 -2459 236
rect -2425 202 -2413 236
rect -2471 168 -2413 202
rect -2471 134 -2459 168
rect -2425 134 -2413 168
rect -2471 109 -2413 134
rect -2323 984 -2265 1009
rect -2323 950 -2311 984
rect -2277 950 -2265 984
rect -2323 916 -2265 950
rect -2323 882 -2311 916
rect -2277 882 -2265 916
rect -2323 848 -2265 882
rect -2323 814 -2311 848
rect -2277 814 -2265 848
rect -2323 780 -2265 814
rect -2323 746 -2311 780
rect -2277 746 -2265 780
rect -2323 712 -2265 746
rect -2323 678 -2311 712
rect -2277 678 -2265 712
rect -2323 644 -2265 678
rect -2323 610 -2311 644
rect -2277 610 -2265 644
rect -2323 576 -2265 610
rect -2323 542 -2311 576
rect -2277 542 -2265 576
rect -2323 508 -2265 542
rect -2323 474 -2311 508
rect -2277 474 -2265 508
rect -2323 440 -2265 474
rect -2323 406 -2311 440
rect -2277 406 -2265 440
rect -2323 372 -2265 406
rect -2323 338 -2311 372
rect -2277 338 -2265 372
rect -2323 304 -2265 338
rect -2323 270 -2311 304
rect -2277 270 -2265 304
rect -2323 236 -2265 270
rect -2323 202 -2311 236
rect -2277 202 -2265 236
rect -2323 168 -2265 202
rect -2323 134 -2311 168
rect -2277 134 -2265 168
rect -2323 109 -2265 134
rect -2175 984 -2117 1009
rect -2175 950 -2163 984
rect -2129 950 -2117 984
rect -2175 916 -2117 950
rect -2175 882 -2163 916
rect -2129 882 -2117 916
rect -2175 848 -2117 882
rect -2175 814 -2163 848
rect -2129 814 -2117 848
rect -2175 780 -2117 814
rect -2175 746 -2163 780
rect -2129 746 -2117 780
rect -2175 712 -2117 746
rect -2175 678 -2163 712
rect -2129 678 -2117 712
rect -2175 644 -2117 678
rect -2175 610 -2163 644
rect -2129 610 -2117 644
rect -2175 576 -2117 610
rect -2175 542 -2163 576
rect -2129 542 -2117 576
rect -2175 508 -2117 542
rect -2175 474 -2163 508
rect -2129 474 -2117 508
rect -2175 440 -2117 474
rect -2175 406 -2163 440
rect -2129 406 -2117 440
rect -2175 372 -2117 406
rect -2175 338 -2163 372
rect -2129 338 -2117 372
rect -2175 304 -2117 338
rect -2175 270 -2163 304
rect -2129 270 -2117 304
rect -2175 236 -2117 270
rect -2175 202 -2163 236
rect -2129 202 -2117 236
rect -2175 168 -2117 202
rect -2175 134 -2163 168
rect -2129 134 -2117 168
rect -2175 109 -2117 134
rect -2027 984 -1969 1009
rect -2027 950 -2015 984
rect -1981 950 -1969 984
rect -2027 916 -1969 950
rect -2027 882 -2015 916
rect -1981 882 -1969 916
rect -2027 848 -1969 882
rect -2027 814 -2015 848
rect -1981 814 -1969 848
rect -2027 780 -1969 814
rect -2027 746 -2015 780
rect -1981 746 -1969 780
rect -2027 712 -1969 746
rect -2027 678 -2015 712
rect -1981 678 -1969 712
rect -2027 644 -1969 678
rect -2027 610 -2015 644
rect -1981 610 -1969 644
rect -2027 576 -1969 610
rect -2027 542 -2015 576
rect -1981 542 -1969 576
rect -2027 508 -1969 542
rect -2027 474 -2015 508
rect -1981 474 -1969 508
rect -2027 440 -1969 474
rect -2027 406 -2015 440
rect -1981 406 -1969 440
rect -2027 372 -1969 406
rect -2027 338 -2015 372
rect -1981 338 -1969 372
rect -2027 304 -1969 338
rect -2027 270 -2015 304
rect -1981 270 -1969 304
rect -2027 236 -1969 270
rect -2027 202 -2015 236
rect -1981 202 -1969 236
rect -2027 168 -1969 202
rect -2027 134 -2015 168
rect -1981 134 -1969 168
rect -2027 109 -1969 134
rect -1879 984 -1821 1009
rect -1879 950 -1867 984
rect -1833 950 -1821 984
rect -1879 916 -1821 950
rect -1879 882 -1867 916
rect -1833 882 -1821 916
rect -1879 848 -1821 882
rect -1879 814 -1867 848
rect -1833 814 -1821 848
rect -1879 780 -1821 814
rect -1879 746 -1867 780
rect -1833 746 -1821 780
rect -1879 712 -1821 746
rect -1879 678 -1867 712
rect -1833 678 -1821 712
rect -1879 644 -1821 678
rect -1879 610 -1867 644
rect -1833 610 -1821 644
rect -1879 576 -1821 610
rect -1879 542 -1867 576
rect -1833 542 -1821 576
rect -1879 508 -1821 542
rect -1879 474 -1867 508
rect -1833 474 -1821 508
rect -1879 440 -1821 474
rect -1879 406 -1867 440
rect -1833 406 -1821 440
rect -1879 372 -1821 406
rect -1879 338 -1867 372
rect -1833 338 -1821 372
rect -1879 304 -1821 338
rect -1879 270 -1867 304
rect -1833 270 -1821 304
rect -1879 236 -1821 270
rect -1879 202 -1867 236
rect -1833 202 -1821 236
rect -1879 168 -1821 202
rect -1879 134 -1867 168
rect -1833 134 -1821 168
rect -1879 109 -1821 134
rect -1731 984 -1673 1009
rect -1731 950 -1719 984
rect -1685 950 -1673 984
rect -1731 916 -1673 950
rect -1731 882 -1719 916
rect -1685 882 -1673 916
rect -1731 848 -1673 882
rect -1731 814 -1719 848
rect -1685 814 -1673 848
rect -1731 780 -1673 814
rect -1731 746 -1719 780
rect -1685 746 -1673 780
rect -1731 712 -1673 746
rect -1731 678 -1719 712
rect -1685 678 -1673 712
rect -1731 644 -1673 678
rect -1731 610 -1719 644
rect -1685 610 -1673 644
rect -1731 576 -1673 610
rect -1731 542 -1719 576
rect -1685 542 -1673 576
rect -1731 508 -1673 542
rect -1731 474 -1719 508
rect -1685 474 -1673 508
rect -1731 440 -1673 474
rect -1731 406 -1719 440
rect -1685 406 -1673 440
rect -1731 372 -1673 406
rect -1731 338 -1719 372
rect -1685 338 -1673 372
rect -1731 304 -1673 338
rect -1731 270 -1719 304
rect -1685 270 -1673 304
rect -1731 236 -1673 270
rect -1731 202 -1719 236
rect -1685 202 -1673 236
rect -1731 168 -1673 202
rect -1731 134 -1719 168
rect -1685 134 -1673 168
rect -1731 109 -1673 134
rect -1583 984 -1525 1009
rect -1583 950 -1571 984
rect -1537 950 -1525 984
rect -1583 916 -1525 950
rect -1583 882 -1571 916
rect -1537 882 -1525 916
rect -1583 848 -1525 882
rect -1583 814 -1571 848
rect -1537 814 -1525 848
rect -1583 780 -1525 814
rect -1583 746 -1571 780
rect -1537 746 -1525 780
rect -1583 712 -1525 746
rect -1583 678 -1571 712
rect -1537 678 -1525 712
rect -1583 644 -1525 678
rect -1583 610 -1571 644
rect -1537 610 -1525 644
rect -1583 576 -1525 610
rect -1583 542 -1571 576
rect -1537 542 -1525 576
rect -1583 508 -1525 542
rect -1583 474 -1571 508
rect -1537 474 -1525 508
rect -1583 440 -1525 474
rect -1583 406 -1571 440
rect -1537 406 -1525 440
rect -1583 372 -1525 406
rect -1583 338 -1571 372
rect -1537 338 -1525 372
rect -1583 304 -1525 338
rect -1583 270 -1571 304
rect -1537 270 -1525 304
rect -1583 236 -1525 270
rect -1583 202 -1571 236
rect -1537 202 -1525 236
rect -1583 168 -1525 202
rect -1583 134 -1571 168
rect -1537 134 -1525 168
rect -1583 109 -1525 134
rect -1435 984 -1377 1009
rect -1435 950 -1423 984
rect -1389 950 -1377 984
rect -1435 916 -1377 950
rect -1435 882 -1423 916
rect -1389 882 -1377 916
rect -1435 848 -1377 882
rect -1435 814 -1423 848
rect -1389 814 -1377 848
rect -1435 780 -1377 814
rect -1435 746 -1423 780
rect -1389 746 -1377 780
rect -1435 712 -1377 746
rect -1435 678 -1423 712
rect -1389 678 -1377 712
rect -1435 644 -1377 678
rect -1435 610 -1423 644
rect -1389 610 -1377 644
rect -1435 576 -1377 610
rect -1435 542 -1423 576
rect -1389 542 -1377 576
rect -1435 508 -1377 542
rect -1435 474 -1423 508
rect -1389 474 -1377 508
rect -1435 440 -1377 474
rect -1435 406 -1423 440
rect -1389 406 -1377 440
rect -1435 372 -1377 406
rect -1435 338 -1423 372
rect -1389 338 -1377 372
rect -1435 304 -1377 338
rect -1435 270 -1423 304
rect -1389 270 -1377 304
rect -1435 236 -1377 270
rect -1435 202 -1423 236
rect -1389 202 -1377 236
rect -1435 168 -1377 202
rect -1435 134 -1423 168
rect -1389 134 -1377 168
rect -1435 109 -1377 134
rect -1287 984 -1229 1009
rect -1287 950 -1275 984
rect -1241 950 -1229 984
rect -1287 916 -1229 950
rect -1287 882 -1275 916
rect -1241 882 -1229 916
rect -1287 848 -1229 882
rect -1287 814 -1275 848
rect -1241 814 -1229 848
rect -1287 780 -1229 814
rect -1287 746 -1275 780
rect -1241 746 -1229 780
rect -1287 712 -1229 746
rect -1287 678 -1275 712
rect -1241 678 -1229 712
rect -1287 644 -1229 678
rect -1287 610 -1275 644
rect -1241 610 -1229 644
rect -1287 576 -1229 610
rect -1287 542 -1275 576
rect -1241 542 -1229 576
rect -1287 508 -1229 542
rect -1287 474 -1275 508
rect -1241 474 -1229 508
rect -1287 440 -1229 474
rect -1287 406 -1275 440
rect -1241 406 -1229 440
rect -1287 372 -1229 406
rect -1287 338 -1275 372
rect -1241 338 -1229 372
rect -1287 304 -1229 338
rect -1287 270 -1275 304
rect -1241 270 -1229 304
rect -1287 236 -1229 270
rect -1287 202 -1275 236
rect -1241 202 -1229 236
rect -1287 168 -1229 202
rect -1287 134 -1275 168
rect -1241 134 -1229 168
rect -1287 109 -1229 134
rect -1139 984 -1081 1009
rect -1139 950 -1127 984
rect -1093 950 -1081 984
rect -1139 916 -1081 950
rect -1139 882 -1127 916
rect -1093 882 -1081 916
rect -1139 848 -1081 882
rect -1139 814 -1127 848
rect -1093 814 -1081 848
rect -1139 780 -1081 814
rect -1139 746 -1127 780
rect -1093 746 -1081 780
rect -1139 712 -1081 746
rect -1139 678 -1127 712
rect -1093 678 -1081 712
rect -1139 644 -1081 678
rect -1139 610 -1127 644
rect -1093 610 -1081 644
rect -1139 576 -1081 610
rect -1139 542 -1127 576
rect -1093 542 -1081 576
rect -1139 508 -1081 542
rect -1139 474 -1127 508
rect -1093 474 -1081 508
rect -1139 440 -1081 474
rect -1139 406 -1127 440
rect -1093 406 -1081 440
rect -1139 372 -1081 406
rect -1139 338 -1127 372
rect -1093 338 -1081 372
rect -1139 304 -1081 338
rect -1139 270 -1127 304
rect -1093 270 -1081 304
rect -1139 236 -1081 270
rect -1139 202 -1127 236
rect -1093 202 -1081 236
rect -1139 168 -1081 202
rect -1139 134 -1127 168
rect -1093 134 -1081 168
rect -1139 109 -1081 134
rect -991 984 -933 1009
rect -991 950 -979 984
rect -945 950 -933 984
rect -991 916 -933 950
rect -991 882 -979 916
rect -945 882 -933 916
rect -991 848 -933 882
rect -991 814 -979 848
rect -945 814 -933 848
rect -991 780 -933 814
rect -991 746 -979 780
rect -945 746 -933 780
rect -991 712 -933 746
rect -991 678 -979 712
rect -945 678 -933 712
rect -991 644 -933 678
rect -991 610 -979 644
rect -945 610 -933 644
rect -991 576 -933 610
rect -991 542 -979 576
rect -945 542 -933 576
rect -991 508 -933 542
rect -991 474 -979 508
rect -945 474 -933 508
rect -991 440 -933 474
rect -991 406 -979 440
rect -945 406 -933 440
rect -991 372 -933 406
rect -991 338 -979 372
rect -945 338 -933 372
rect -991 304 -933 338
rect -991 270 -979 304
rect -945 270 -933 304
rect -991 236 -933 270
rect -991 202 -979 236
rect -945 202 -933 236
rect -991 168 -933 202
rect -991 134 -979 168
rect -945 134 -933 168
rect -991 109 -933 134
rect -843 984 -785 1009
rect -843 950 -831 984
rect -797 950 -785 984
rect -843 916 -785 950
rect -843 882 -831 916
rect -797 882 -785 916
rect -843 848 -785 882
rect -843 814 -831 848
rect -797 814 -785 848
rect -843 780 -785 814
rect -843 746 -831 780
rect -797 746 -785 780
rect -843 712 -785 746
rect -843 678 -831 712
rect -797 678 -785 712
rect -843 644 -785 678
rect -843 610 -831 644
rect -797 610 -785 644
rect -843 576 -785 610
rect -843 542 -831 576
rect -797 542 -785 576
rect -843 508 -785 542
rect -843 474 -831 508
rect -797 474 -785 508
rect -843 440 -785 474
rect -843 406 -831 440
rect -797 406 -785 440
rect -843 372 -785 406
rect -843 338 -831 372
rect -797 338 -785 372
rect -843 304 -785 338
rect -843 270 -831 304
rect -797 270 -785 304
rect -843 236 -785 270
rect -843 202 -831 236
rect -797 202 -785 236
rect -843 168 -785 202
rect -843 134 -831 168
rect -797 134 -785 168
rect -843 109 -785 134
rect -695 984 -637 1009
rect -695 950 -683 984
rect -649 950 -637 984
rect -695 916 -637 950
rect -695 882 -683 916
rect -649 882 -637 916
rect -695 848 -637 882
rect -695 814 -683 848
rect -649 814 -637 848
rect -695 780 -637 814
rect -695 746 -683 780
rect -649 746 -637 780
rect -695 712 -637 746
rect -695 678 -683 712
rect -649 678 -637 712
rect -695 644 -637 678
rect -695 610 -683 644
rect -649 610 -637 644
rect -695 576 -637 610
rect -695 542 -683 576
rect -649 542 -637 576
rect -695 508 -637 542
rect -695 474 -683 508
rect -649 474 -637 508
rect -695 440 -637 474
rect -695 406 -683 440
rect -649 406 -637 440
rect -695 372 -637 406
rect -695 338 -683 372
rect -649 338 -637 372
rect -695 304 -637 338
rect -695 270 -683 304
rect -649 270 -637 304
rect -695 236 -637 270
rect -695 202 -683 236
rect -649 202 -637 236
rect -695 168 -637 202
rect -695 134 -683 168
rect -649 134 -637 168
rect -695 109 -637 134
rect -547 984 -489 1009
rect -547 950 -535 984
rect -501 950 -489 984
rect -547 916 -489 950
rect -547 882 -535 916
rect -501 882 -489 916
rect -547 848 -489 882
rect -547 814 -535 848
rect -501 814 -489 848
rect -547 780 -489 814
rect -547 746 -535 780
rect -501 746 -489 780
rect -547 712 -489 746
rect -547 678 -535 712
rect -501 678 -489 712
rect -547 644 -489 678
rect -547 610 -535 644
rect -501 610 -489 644
rect -547 576 -489 610
rect -547 542 -535 576
rect -501 542 -489 576
rect -547 508 -489 542
rect -547 474 -535 508
rect -501 474 -489 508
rect -547 440 -489 474
rect -547 406 -535 440
rect -501 406 -489 440
rect -547 372 -489 406
rect -547 338 -535 372
rect -501 338 -489 372
rect -547 304 -489 338
rect -547 270 -535 304
rect -501 270 -489 304
rect -547 236 -489 270
rect -547 202 -535 236
rect -501 202 -489 236
rect -547 168 -489 202
rect -547 134 -535 168
rect -501 134 -489 168
rect -547 109 -489 134
rect -399 984 -341 1009
rect -399 950 -387 984
rect -353 950 -341 984
rect -399 916 -341 950
rect -399 882 -387 916
rect -353 882 -341 916
rect -399 848 -341 882
rect -399 814 -387 848
rect -353 814 -341 848
rect -399 780 -341 814
rect -399 746 -387 780
rect -353 746 -341 780
rect -399 712 -341 746
rect -399 678 -387 712
rect -353 678 -341 712
rect -399 644 -341 678
rect -399 610 -387 644
rect -353 610 -341 644
rect -399 576 -341 610
rect -399 542 -387 576
rect -353 542 -341 576
rect -399 508 -341 542
rect -399 474 -387 508
rect -353 474 -341 508
rect -399 440 -341 474
rect -399 406 -387 440
rect -353 406 -341 440
rect -399 372 -341 406
rect -399 338 -387 372
rect -353 338 -341 372
rect -399 304 -341 338
rect -399 270 -387 304
rect -353 270 -341 304
rect -399 236 -341 270
rect -399 202 -387 236
rect -353 202 -341 236
rect -399 168 -341 202
rect -399 134 -387 168
rect -353 134 -341 168
rect -399 109 -341 134
rect -251 984 -193 1009
rect -251 950 -239 984
rect -205 950 -193 984
rect -251 916 -193 950
rect -251 882 -239 916
rect -205 882 -193 916
rect -251 848 -193 882
rect -251 814 -239 848
rect -205 814 -193 848
rect -251 780 -193 814
rect -251 746 -239 780
rect -205 746 -193 780
rect -251 712 -193 746
rect -251 678 -239 712
rect -205 678 -193 712
rect -251 644 -193 678
rect -251 610 -239 644
rect -205 610 -193 644
rect -251 576 -193 610
rect -251 542 -239 576
rect -205 542 -193 576
rect -251 508 -193 542
rect -251 474 -239 508
rect -205 474 -193 508
rect -251 440 -193 474
rect -251 406 -239 440
rect -205 406 -193 440
rect -251 372 -193 406
rect -251 338 -239 372
rect -205 338 -193 372
rect -251 304 -193 338
rect -251 270 -239 304
rect -205 270 -193 304
rect -251 236 -193 270
rect -251 202 -239 236
rect -205 202 -193 236
rect -251 168 -193 202
rect -251 134 -239 168
rect -205 134 -193 168
rect -251 109 -193 134
rect -103 984 -45 1009
rect -103 950 -91 984
rect -57 950 -45 984
rect -103 916 -45 950
rect -103 882 -91 916
rect -57 882 -45 916
rect -103 848 -45 882
rect -103 814 -91 848
rect -57 814 -45 848
rect -103 780 -45 814
rect -103 746 -91 780
rect -57 746 -45 780
rect -103 712 -45 746
rect -103 678 -91 712
rect -57 678 -45 712
rect -103 644 -45 678
rect -103 610 -91 644
rect -57 610 -45 644
rect -103 576 -45 610
rect -103 542 -91 576
rect -57 542 -45 576
rect -103 508 -45 542
rect -103 474 -91 508
rect -57 474 -45 508
rect -103 440 -45 474
rect -103 406 -91 440
rect -57 406 -45 440
rect -103 372 -45 406
rect -103 338 -91 372
rect -57 338 -45 372
rect -103 304 -45 338
rect -103 270 -91 304
rect -57 270 -45 304
rect -103 236 -45 270
rect -103 202 -91 236
rect -57 202 -45 236
rect -103 168 -45 202
rect -103 134 -91 168
rect -57 134 -45 168
rect -103 109 -45 134
rect 45 984 103 1009
rect 45 950 57 984
rect 91 950 103 984
rect 45 916 103 950
rect 45 882 57 916
rect 91 882 103 916
rect 45 848 103 882
rect 45 814 57 848
rect 91 814 103 848
rect 45 780 103 814
rect 45 746 57 780
rect 91 746 103 780
rect 45 712 103 746
rect 45 678 57 712
rect 91 678 103 712
rect 45 644 103 678
rect 45 610 57 644
rect 91 610 103 644
rect 45 576 103 610
rect 45 542 57 576
rect 91 542 103 576
rect 45 508 103 542
rect 45 474 57 508
rect 91 474 103 508
rect 45 440 103 474
rect 45 406 57 440
rect 91 406 103 440
rect 45 372 103 406
rect 45 338 57 372
rect 91 338 103 372
rect 45 304 103 338
rect 45 270 57 304
rect 91 270 103 304
rect 45 236 103 270
rect 45 202 57 236
rect 91 202 103 236
rect 45 168 103 202
rect 45 134 57 168
rect 91 134 103 168
rect 45 109 103 134
rect 193 984 251 1009
rect 193 950 205 984
rect 239 950 251 984
rect 193 916 251 950
rect 193 882 205 916
rect 239 882 251 916
rect 193 848 251 882
rect 193 814 205 848
rect 239 814 251 848
rect 193 780 251 814
rect 193 746 205 780
rect 239 746 251 780
rect 193 712 251 746
rect 193 678 205 712
rect 239 678 251 712
rect 193 644 251 678
rect 193 610 205 644
rect 239 610 251 644
rect 193 576 251 610
rect 193 542 205 576
rect 239 542 251 576
rect 193 508 251 542
rect 193 474 205 508
rect 239 474 251 508
rect 193 440 251 474
rect 193 406 205 440
rect 239 406 251 440
rect 193 372 251 406
rect 193 338 205 372
rect 239 338 251 372
rect 193 304 251 338
rect 193 270 205 304
rect 239 270 251 304
rect 193 236 251 270
rect 193 202 205 236
rect 239 202 251 236
rect 193 168 251 202
rect 193 134 205 168
rect 239 134 251 168
rect 193 109 251 134
rect 341 984 399 1009
rect 341 950 353 984
rect 387 950 399 984
rect 341 916 399 950
rect 341 882 353 916
rect 387 882 399 916
rect 341 848 399 882
rect 341 814 353 848
rect 387 814 399 848
rect 341 780 399 814
rect 341 746 353 780
rect 387 746 399 780
rect 341 712 399 746
rect 341 678 353 712
rect 387 678 399 712
rect 341 644 399 678
rect 341 610 353 644
rect 387 610 399 644
rect 341 576 399 610
rect 341 542 353 576
rect 387 542 399 576
rect 341 508 399 542
rect 341 474 353 508
rect 387 474 399 508
rect 341 440 399 474
rect 341 406 353 440
rect 387 406 399 440
rect 341 372 399 406
rect 341 338 353 372
rect 387 338 399 372
rect 341 304 399 338
rect 341 270 353 304
rect 387 270 399 304
rect 341 236 399 270
rect 341 202 353 236
rect 387 202 399 236
rect 341 168 399 202
rect 341 134 353 168
rect 387 134 399 168
rect 341 109 399 134
rect 489 984 547 1009
rect 489 950 501 984
rect 535 950 547 984
rect 489 916 547 950
rect 489 882 501 916
rect 535 882 547 916
rect 489 848 547 882
rect 489 814 501 848
rect 535 814 547 848
rect 489 780 547 814
rect 489 746 501 780
rect 535 746 547 780
rect 489 712 547 746
rect 489 678 501 712
rect 535 678 547 712
rect 489 644 547 678
rect 489 610 501 644
rect 535 610 547 644
rect 489 576 547 610
rect 489 542 501 576
rect 535 542 547 576
rect 489 508 547 542
rect 489 474 501 508
rect 535 474 547 508
rect 489 440 547 474
rect 489 406 501 440
rect 535 406 547 440
rect 489 372 547 406
rect 489 338 501 372
rect 535 338 547 372
rect 489 304 547 338
rect 489 270 501 304
rect 535 270 547 304
rect 489 236 547 270
rect 489 202 501 236
rect 535 202 547 236
rect 489 168 547 202
rect 489 134 501 168
rect 535 134 547 168
rect 489 109 547 134
rect 637 984 695 1009
rect 637 950 649 984
rect 683 950 695 984
rect 637 916 695 950
rect 637 882 649 916
rect 683 882 695 916
rect 637 848 695 882
rect 637 814 649 848
rect 683 814 695 848
rect 637 780 695 814
rect 637 746 649 780
rect 683 746 695 780
rect 637 712 695 746
rect 637 678 649 712
rect 683 678 695 712
rect 637 644 695 678
rect 637 610 649 644
rect 683 610 695 644
rect 637 576 695 610
rect 637 542 649 576
rect 683 542 695 576
rect 637 508 695 542
rect 637 474 649 508
rect 683 474 695 508
rect 637 440 695 474
rect 637 406 649 440
rect 683 406 695 440
rect 637 372 695 406
rect 637 338 649 372
rect 683 338 695 372
rect 637 304 695 338
rect 637 270 649 304
rect 683 270 695 304
rect 637 236 695 270
rect 637 202 649 236
rect 683 202 695 236
rect 637 168 695 202
rect 637 134 649 168
rect 683 134 695 168
rect 637 109 695 134
rect 785 984 843 1009
rect 785 950 797 984
rect 831 950 843 984
rect 785 916 843 950
rect 785 882 797 916
rect 831 882 843 916
rect 785 848 843 882
rect 785 814 797 848
rect 831 814 843 848
rect 785 780 843 814
rect 785 746 797 780
rect 831 746 843 780
rect 785 712 843 746
rect 785 678 797 712
rect 831 678 843 712
rect 785 644 843 678
rect 785 610 797 644
rect 831 610 843 644
rect 785 576 843 610
rect 785 542 797 576
rect 831 542 843 576
rect 785 508 843 542
rect 785 474 797 508
rect 831 474 843 508
rect 785 440 843 474
rect 785 406 797 440
rect 831 406 843 440
rect 785 372 843 406
rect 785 338 797 372
rect 831 338 843 372
rect 785 304 843 338
rect 785 270 797 304
rect 831 270 843 304
rect 785 236 843 270
rect 785 202 797 236
rect 831 202 843 236
rect 785 168 843 202
rect 785 134 797 168
rect 831 134 843 168
rect 785 109 843 134
rect 933 984 991 1009
rect 933 950 945 984
rect 979 950 991 984
rect 933 916 991 950
rect 933 882 945 916
rect 979 882 991 916
rect 933 848 991 882
rect 933 814 945 848
rect 979 814 991 848
rect 933 780 991 814
rect 933 746 945 780
rect 979 746 991 780
rect 933 712 991 746
rect 933 678 945 712
rect 979 678 991 712
rect 933 644 991 678
rect 933 610 945 644
rect 979 610 991 644
rect 933 576 991 610
rect 933 542 945 576
rect 979 542 991 576
rect 933 508 991 542
rect 933 474 945 508
rect 979 474 991 508
rect 933 440 991 474
rect 933 406 945 440
rect 979 406 991 440
rect 933 372 991 406
rect 933 338 945 372
rect 979 338 991 372
rect 933 304 991 338
rect 933 270 945 304
rect 979 270 991 304
rect 933 236 991 270
rect 933 202 945 236
rect 979 202 991 236
rect 933 168 991 202
rect 933 134 945 168
rect 979 134 991 168
rect 933 109 991 134
rect 1081 984 1139 1009
rect 1081 950 1093 984
rect 1127 950 1139 984
rect 1081 916 1139 950
rect 1081 882 1093 916
rect 1127 882 1139 916
rect 1081 848 1139 882
rect 1081 814 1093 848
rect 1127 814 1139 848
rect 1081 780 1139 814
rect 1081 746 1093 780
rect 1127 746 1139 780
rect 1081 712 1139 746
rect 1081 678 1093 712
rect 1127 678 1139 712
rect 1081 644 1139 678
rect 1081 610 1093 644
rect 1127 610 1139 644
rect 1081 576 1139 610
rect 1081 542 1093 576
rect 1127 542 1139 576
rect 1081 508 1139 542
rect 1081 474 1093 508
rect 1127 474 1139 508
rect 1081 440 1139 474
rect 1081 406 1093 440
rect 1127 406 1139 440
rect 1081 372 1139 406
rect 1081 338 1093 372
rect 1127 338 1139 372
rect 1081 304 1139 338
rect 1081 270 1093 304
rect 1127 270 1139 304
rect 1081 236 1139 270
rect 1081 202 1093 236
rect 1127 202 1139 236
rect 1081 168 1139 202
rect 1081 134 1093 168
rect 1127 134 1139 168
rect 1081 109 1139 134
rect 1229 984 1287 1009
rect 1229 950 1241 984
rect 1275 950 1287 984
rect 1229 916 1287 950
rect 1229 882 1241 916
rect 1275 882 1287 916
rect 1229 848 1287 882
rect 1229 814 1241 848
rect 1275 814 1287 848
rect 1229 780 1287 814
rect 1229 746 1241 780
rect 1275 746 1287 780
rect 1229 712 1287 746
rect 1229 678 1241 712
rect 1275 678 1287 712
rect 1229 644 1287 678
rect 1229 610 1241 644
rect 1275 610 1287 644
rect 1229 576 1287 610
rect 1229 542 1241 576
rect 1275 542 1287 576
rect 1229 508 1287 542
rect 1229 474 1241 508
rect 1275 474 1287 508
rect 1229 440 1287 474
rect 1229 406 1241 440
rect 1275 406 1287 440
rect 1229 372 1287 406
rect 1229 338 1241 372
rect 1275 338 1287 372
rect 1229 304 1287 338
rect 1229 270 1241 304
rect 1275 270 1287 304
rect 1229 236 1287 270
rect 1229 202 1241 236
rect 1275 202 1287 236
rect 1229 168 1287 202
rect 1229 134 1241 168
rect 1275 134 1287 168
rect 1229 109 1287 134
rect 1377 984 1435 1009
rect 1377 950 1389 984
rect 1423 950 1435 984
rect 1377 916 1435 950
rect 1377 882 1389 916
rect 1423 882 1435 916
rect 1377 848 1435 882
rect 1377 814 1389 848
rect 1423 814 1435 848
rect 1377 780 1435 814
rect 1377 746 1389 780
rect 1423 746 1435 780
rect 1377 712 1435 746
rect 1377 678 1389 712
rect 1423 678 1435 712
rect 1377 644 1435 678
rect 1377 610 1389 644
rect 1423 610 1435 644
rect 1377 576 1435 610
rect 1377 542 1389 576
rect 1423 542 1435 576
rect 1377 508 1435 542
rect 1377 474 1389 508
rect 1423 474 1435 508
rect 1377 440 1435 474
rect 1377 406 1389 440
rect 1423 406 1435 440
rect 1377 372 1435 406
rect 1377 338 1389 372
rect 1423 338 1435 372
rect 1377 304 1435 338
rect 1377 270 1389 304
rect 1423 270 1435 304
rect 1377 236 1435 270
rect 1377 202 1389 236
rect 1423 202 1435 236
rect 1377 168 1435 202
rect 1377 134 1389 168
rect 1423 134 1435 168
rect 1377 109 1435 134
rect 1525 984 1583 1009
rect 1525 950 1537 984
rect 1571 950 1583 984
rect 1525 916 1583 950
rect 1525 882 1537 916
rect 1571 882 1583 916
rect 1525 848 1583 882
rect 1525 814 1537 848
rect 1571 814 1583 848
rect 1525 780 1583 814
rect 1525 746 1537 780
rect 1571 746 1583 780
rect 1525 712 1583 746
rect 1525 678 1537 712
rect 1571 678 1583 712
rect 1525 644 1583 678
rect 1525 610 1537 644
rect 1571 610 1583 644
rect 1525 576 1583 610
rect 1525 542 1537 576
rect 1571 542 1583 576
rect 1525 508 1583 542
rect 1525 474 1537 508
rect 1571 474 1583 508
rect 1525 440 1583 474
rect 1525 406 1537 440
rect 1571 406 1583 440
rect 1525 372 1583 406
rect 1525 338 1537 372
rect 1571 338 1583 372
rect 1525 304 1583 338
rect 1525 270 1537 304
rect 1571 270 1583 304
rect 1525 236 1583 270
rect 1525 202 1537 236
rect 1571 202 1583 236
rect 1525 168 1583 202
rect 1525 134 1537 168
rect 1571 134 1583 168
rect 1525 109 1583 134
rect 1673 984 1731 1009
rect 1673 950 1685 984
rect 1719 950 1731 984
rect 1673 916 1731 950
rect 1673 882 1685 916
rect 1719 882 1731 916
rect 1673 848 1731 882
rect 1673 814 1685 848
rect 1719 814 1731 848
rect 1673 780 1731 814
rect 1673 746 1685 780
rect 1719 746 1731 780
rect 1673 712 1731 746
rect 1673 678 1685 712
rect 1719 678 1731 712
rect 1673 644 1731 678
rect 1673 610 1685 644
rect 1719 610 1731 644
rect 1673 576 1731 610
rect 1673 542 1685 576
rect 1719 542 1731 576
rect 1673 508 1731 542
rect 1673 474 1685 508
rect 1719 474 1731 508
rect 1673 440 1731 474
rect 1673 406 1685 440
rect 1719 406 1731 440
rect 1673 372 1731 406
rect 1673 338 1685 372
rect 1719 338 1731 372
rect 1673 304 1731 338
rect 1673 270 1685 304
rect 1719 270 1731 304
rect 1673 236 1731 270
rect 1673 202 1685 236
rect 1719 202 1731 236
rect 1673 168 1731 202
rect 1673 134 1685 168
rect 1719 134 1731 168
rect 1673 109 1731 134
rect 1821 984 1879 1009
rect 1821 950 1833 984
rect 1867 950 1879 984
rect 1821 916 1879 950
rect 1821 882 1833 916
rect 1867 882 1879 916
rect 1821 848 1879 882
rect 1821 814 1833 848
rect 1867 814 1879 848
rect 1821 780 1879 814
rect 1821 746 1833 780
rect 1867 746 1879 780
rect 1821 712 1879 746
rect 1821 678 1833 712
rect 1867 678 1879 712
rect 1821 644 1879 678
rect 1821 610 1833 644
rect 1867 610 1879 644
rect 1821 576 1879 610
rect 1821 542 1833 576
rect 1867 542 1879 576
rect 1821 508 1879 542
rect 1821 474 1833 508
rect 1867 474 1879 508
rect 1821 440 1879 474
rect 1821 406 1833 440
rect 1867 406 1879 440
rect 1821 372 1879 406
rect 1821 338 1833 372
rect 1867 338 1879 372
rect 1821 304 1879 338
rect 1821 270 1833 304
rect 1867 270 1879 304
rect 1821 236 1879 270
rect 1821 202 1833 236
rect 1867 202 1879 236
rect 1821 168 1879 202
rect 1821 134 1833 168
rect 1867 134 1879 168
rect 1821 109 1879 134
rect 1969 984 2027 1009
rect 1969 950 1981 984
rect 2015 950 2027 984
rect 1969 916 2027 950
rect 1969 882 1981 916
rect 2015 882 2027 916
rect 1969 848 2027 882
rect 1969 814 1981 848
rect 2015 814 2027 848
rect 1969 780 2027 814
rect 1969 746 1981 780
rect 2015 746 2027 780
rect 1969 712 2027 746
rect 1969 678 1981 712
rect 2015 678 2027 712
rect 1969 644 2027 678
rect 1969 610 1981 644
rect 2015 610 2027 644
rect 1969 576 2027 610
rect 1969 542 1981 576
rect 2015 542 2027 576
rect 1969 508 2027 542
rect 1969 474 1981 508
rect 2015 474 2027 508
rect 1969 440 2027 474
rect 1969 406 1981 440
rect 2015 406 2027 440
rect 1969 372 2027 406
rect 1969 338 1981 372
rect 2015 338 2027 372
rect 1969 304 2027 338
rect 1969 270 1981 304
rect 2015 270 2027 304
rect 1969 236 2027 270
rect 1969 202 1981 236
rect 2015 202 2027 236
rect 1969 168 2027 202
rect 1969 134 1981 168
rect 2015 134 2027 168
rect 1969 109 2027 134
rect 2117 984 2175 1009
rect 2117 950 2129 984
rect 2163 950 2175 984
rect 2117 916 2175 950
rect 2117 882 2129 916
rect 2163 882 2175 916
rect 2117 848 2175 882
rect 2117 814 2129 848
rect 2163 814 2175 848
rect 2117 780 2175 814
rect 2117 746 2129 780
rect 2163 746 2175 780
rect 2117 712 2175 746
rect 2117 678 2129 712
rect 2163 678 2175 712
rect 2117 644 2175 678
rect 2117 610 2129 644
rect 2163 610 2175 644
rect 2117 576 2175 610
rect 2117 542 2129 576
rect 2163 542 2175 576
rect 2117 508 2175 542
rect 2117 474 2129 508
rect 2163 474 2175 508
rect 2117 440 2175 474
rect 2117 406 2129 440
rect 2163 406 2175 440
rect 2117 372 2175 406
rect 2117 338 2129 372
rect 2163 338 2175 372
rect 2117 304 2175 338
rect 2117 270 2129 304
rect 2163 270 2175 304
rect 2117 236 2175 270
rect 2117 202 2129 236
rect 2163 202 2175 236
rect 2117 168 2175 202
rect 2117 134 2129 168
rect 2163 134 2175 168
rect 2117 109 2175 134
rect 2265 984 2323 1009
rect 2265 950 2277 984
rect 2311 950 2323 984
rect 2265 916 2323 950
rect 2265 882 2277 916
rect 2311 882 2323 916
rect 2265 848 2323 882
rect 2265 814 2277 848
rect 2311 814 2323 848
rect 2265 780 2323 814
rect 2265 746 2277 780
rect 2311 746 2323 780
rect 2265 712 2323 746
rect 2265 678 2277 712
rect 2311 678 2323 712
rect 2265 644 2323 678
rect 2265 610 2277 644
rect 2311 610 2323 644
rect 2265 576 2323 610
rect 2265 542 2277 576
rect 2311 542 2323 576
rect 2265 508 2323 542
rect 2265 474 2277 508
rect 2311 474 2323 508
rect 2265 440 2323 474
rect 2265 406 2277 440
rect 2311 406 2323 440
rect 2265 372 2323 406
rect 2265 338 2277 372
rect 2311 338 2323 372
rect 2265 304 2323 338
rect 2265 270 2277 304
rect 2311 270 2323 304
rect 2265 236 2323 270
rect 2265 202 2277 236
rect 2311 202 2323 236
rect 2265 168 2323 202
rect 2265 134 2277 168
rect 2311 134 2323 168
rect 2265 109 2323 134
rect 2413 984 2471 1009
rect 2413 950 2425 984
rect 2459 950 2471 984
rect 2413 916 2471 950
rect 2413 882 2425 916
rect 2459 882 2471 916
rect 2413 848 2471 882
rect 2413 814 2425 848
rect 2459 814 2471 848
rect 2413 780 2471 814
rect 2413 746 2425 780
rect 2459 746 2471 780
rect 2413 712 2471 746
rect 2413 678 2425 712
rect 2459 678 2471 712
rect 2413 644 2471 678
rect 2413 610 2425 644
rect 2459 610 2471 644
rect 2413 576 2471 610
rect 2413 542 2425 576
rect 2459 542 2471 576
rect 2413 508 2471 542
rect 2413 474 2425 508
rect 2459 474 2471 508
rect 2413 440 2471 474
rect 2413 406 2425 440
rect 2459 406 2471 440
rect 2413 372 2471 406
rect 2413 338 2425 372
rect 2459 338 2471 372
rect 2413 304 2471 338
rect 2413 270 2425 304
rect 2459 270 2471 304
rect 2413 236 2471 270
rect 2413 202 2425 236
rect 2459 202 2471 236
rect 2413 168 2471 202
rect 2413 134 2425 168
rect 2459 134 2471 168
rect 2413 109 2471 134
rect 2561 984 2619 1009
rect 2561 950 2573 984
rect 2607 950 2619 984
rect 2561 916 2619 950
rect 2561 882 2573 916
rect 2607 882 2619 916
rect 2561 848 2619 882
rect 2561 814 2573 848
rect 2607 814 2619 848
rect 2561 780 2619 814
rect 2561 746 2573 780
rect 2607 746 2619 780
rect 2561 712 2619 746
rect 2561 678 2573 712
rect 2607 678 2619 712
rect 2561 644 2619 678
rect 2561 610 2573 644
rect 2607 610 2619 644
rect 2561 576 2619 610
rect 2561 542 2573 576
rect 2607 542 2619 576
rect 2561 508 2619 542
rect 2561 474 2573 508
rect 2607 474 2619 508
rect 2561 440 2619 474
rect 2561 406 2573 440
rect 2607 406 2619 440
rect 2561 372 2619 406
rect 2561 338 2573 372
rect 2607 338 2619 372
rect 2561 304 2619 338
rect 2561 270 2573 304
rect 2607 270 2619 304
rect 2561 236 2619 270
rect 2561 202 2573 236
rect 2607 202 2619 236
rect 2561 168 2619 202
rect 2561 134 2573 168
rect 2607 134 2619 168
rect 2561 109 2619 134
rect 2709 984 2767 1009
rect 2709 950 2721 984
rect 2755 950 2767 984
rect 2709 916 2767 950
rect 2709 882 2721 916
rect 2755 882 2767 916
rect 2709 848 2767 882
rect 2709 814 2721 848
rect 2755 814 2767 848
rect 2709 780 2767 814
rect 2709 746 2721 780
rect 2755 746 2767 780
rect 2709 712 2767 746
rect 2709 678 2721 712
rect 2755 678 2767 712
rect 2709 644 2767 678
rect 2709 610 2721 644
rect 2755 610 2767 644
rect 2709 576 2767 610
rect 2709 542 2721 576
rect 2755 542 2767 576
rect 2709 508 2767 542
rect 2709 474 2721 508
rect 2755 474 2767 508
rect 2709 440 2767 474
rect 2709 406 2721 440
rect 2755 406 2767 440
rect 2709 372 2767 406
rect 2709 338 2721 372
rect 2755 338 2767 372
rect 2709 304 2767 338
rect 2709 270 2721 304
rect 2755 270 2767 304
rect 2709 236 2767 270
rect 2709 202 2721 236
rect 2755 202 2767 236
rect 2709 168 2767 202
rect 2709 134 2721 168
rect 2755 134 2767 168
rect 2709 109 2767 134
rect 2857 984 2915 1009
rect 2857 950 2869 984
rect 2903 950 2915 984
rect 2857 916 2915 950
rect 2857 882 2869 916
rect 2903 882 2915 916
rect 2857 848 2915 882
rect 2857 814 2869 848
rect 2903 814 2915 848
rect 2857 780 2915 814
rect 2857 746 2869 780
rect 2903 746 2915 780
rect 2857 712 2915 746
rect 2857 678 2869 712
rect 2903 678 2915 712
rect 2857 644 2915 678
rect 2857 610 2869 644
rect 2903 610 2915 644
rect 2857 576 2915 610
rect 2857 542 2869 576
rect 2903 542 2915 576
rect 2857 508 2915 542
rect 2857 474 2869 508
rect 2903 474 2915 508
rect 2857 440 2915 474
rect 2857 406 2869 440
rect 2903 406 2915 440
rect 2857 372 2915 406
rect 2857 338 2869 372
rect 2903 338 2915 372
rect 2857 304 2915 338
rect 2857 270 2869 304
rect 2903 270 2915 304
rect 2857 236 2915 270
rect 2857 202 2869 236
rect 2903 202 2915 236
rect 2857 168 2915 202
rect 2857 134 2869 168
rect 2903 134 2915 168
rect 2857 109 2915 134
rect 3005 984 3063 1009
rect 3005 950 3017 984
rect 3051 950 3063 984
rect 3005 916 3063 950
rect 3005 882 3017 916
rect 3051 882 3063 916
rect 3005 848 3063 882
rect 3005 814 3017 848
rect 3051 814 3063 848
rect 3005 780 3063 814
rect 3005 746 3017 780
rect 3051 746 3063 780
rect 3005 712 3063 746
rect 3005 678 3017 712
rect 3051 678 3063 712
rect 3005 644 3063 678
rect 3005 610 3017 644
rect 3051 610 3063 644
rect 3005 576 3063 610
rect 3005 542 3017 576
rect 3051 542 3063 576
rect 3005 508 3063 542
rect 3005 474 3017 508
rect 3051 474 3063 508
rect 3005 440 3063 474
rect 3005 406 3017 440
rect 3051 406 3063 440
rect 3005 372 3063 406
rect 3005 338 3017 372
rect 3051 338 3063 372
rect 3005 304 3063 338
rect 3005 270 3017 304
rect 3051 270 3063 304
rect 3005 236 3063 270
rect 3005 202 3017 236
rect 3051 202 3063 236
rect 3005 168 3063 202
rect 3005 134 3017 168
rect 3051 134 3063 168
rect 3005 109 3063 134
rect 3153 984 3211 1009
rect 3153 950 3165 984
rect 3199 950 3211 984
rect 3153 916 3211 950
rect 3153 882 3165 916
rect 3199 882 3211 916
rect 3153 848 3211 882
rect 3153 814 3165 848
rect 3199 814 3211 848
rect 3153 780 3211 814
rect 3153 746 3165 780
rect 3199 746 3211 780
rect 3153 712 3211 746
rect 3153 678 3165 712
rect 3199 678 3211 712
rect 3153 644 3211 678
rect 3153 610 3165 644
rect 3199 610 3211 644
rect 3153 576 3211 610
rect 3153 542 3165 576
rect 3199 542 3211 576
rect 3153 508 3211 542
rect 3153 474 3165 508
rect 3199 474 3211 508
rect 3153 440 3211 474
rect 3153 406 3165 440
rect 3199 406 3211 440
rect 3153 372 3211 406
rect 3153 338 3165 372
rect 3199 338 3211 372
rect 3153 304 3211 338
rect 3153 270 3165 304
rect 3199 270 3211 304
rect 3153 236 3211 270
rect 3153 202 3165 236
rect 3199 202 3211 236
rect 3153 168 3211 202
rect 3153 134 3165 168
rect 3199 134 3211 168
rect 3153 109 3211 134
rect 3301 984 3359 1009
rect 3301 950 3313 984
rect 3347 950 3359 984
rect 3301 916 3359 950
rect 3301 882 3313 916
rect 3347 882 3359 916
rect 3301 848 3359 882
rect 3301 814 3313 848
rect 3347 814 3359 848
rect 3301 780 3359 814
rect 3301 746 3313 780
rect 3347 746 3359 780
rect 3301 712 3359 746
rect 3301 678 3313 712
rect 3347 678 3359 712
rect 3301 644 3359 678
rect 3301 610 3313 644
rect 3347 610 3359 644
rect 3301 576 3359 610
rect 3301 542 3313 576
rect 3347 542 3359 576
rect 3301 508 3359 542
rect 3301 474 3313 508
rect 3347 474 3359 508
rect 3301 440 3359 474
rect 3301 406 3313 440
rect 3347 406 3359 440
rect 3301 372 3359 406
rect 3301 338 3313 372
rect 3347 338 3359 372
rect 3301 304 3359 338
rect 3301 270 3313 304
rect 3347 270 3359 304
rect 3301 236 3359 270
rect 3301 202 3313 236
rect 3347 202 3359 236
rect 3301 168 3359 202
rect 3301 134 3313 168
rect 3347 134 3359 168
rect 3301 109 3359 134
rect 3449 984 3507 1009
rect 3449 950 3461 984
rect 3495 950 3507 984
rect 3449 916 3507 950
rect 3449 882 3461 916
rect 3495 882 3507 916
rect 3449 848 3507 882
rect 3449 814 3461 848
rect 3495 814 3507 848
rect 3449 780 3507 814
rect 3449 746 3461 780
rect 3495 746 3507 780
rect 3449 712 3507 746
rect 3449 678 3461 712
rect 3495 678 3507 712
rect 3449 644 3507 678
rect 3449 610 3461 644
rect 3495 610 3507 644
rect 3449 576 3507 610
rect 3449 542 3461 576
rect 3495 542 3507 576
rect 3449 508 3507 542
rect 3449 474 3461 508
rect 3495 474 3507 508
rect 3449 440 3507 474
rect 3449 406 3461 440
rect 3495 406 3507 440
rect 3449 372 3507 406
rect 3449 338 3461 372
rect 3495 338 3507 372
rect 3449 304 3507 338
rect 3449 270 3461 304
rect 3495 270 3507 304
rect 3449 236 3507 270
rect 3449 202 3461 236
rect 3495 202 3507 236
rect 3449 168 3507 202
rect 3449 134 3461 168
rect 3495 134 3507 168
rect 3449 109 3507 134
rect 3597 984 3655 1009
rect 3597 950 3609 984
rect 3643 950 3655 984
rect 3597 916 3655 950
rect 3597 882 3609 916
rect 3643 882 3655 916
rect 3597 848 3655 882
rect 3597 814 3609 848
rect 3643 814 3655 848
rect 3597 780 3655 814
rect 3597 746 3609 780
rect 3643 746 3655 780
rect 3597 712 3655 746
rect 3597 678 3609 712
rect 3643 678 3655 712
rect 3597 644 3655 678
rect 3597 610 3609 644
rect 3643 610 3655 644
rect 3597 576 3655 610
rect 3597 542 3609 576
rect 3643 542 3655 576
rect 3597 508 3655 542
rect 3597 474 3609 508
rect 3643 474 3655 508
rect 3597 440 3655 474
rect 3597 406 3609 440
rect 3643 406 3655 440
rect 3597 372 3655 406
rect 3597 338 3609 372
rect 3643 338 3655 372
rect 3597 304 3655 338
rect 3597 270 3609 304
rect 3643 270 3655 304
rect 3597 236 3655 270
rect 3597 202 3609 236
rect 3643 202 3655 236
rect 3597 168 3655 202
rect 3597 134 3609 168
rect 3643 134 3655 168
rect 3597 109 3655 134
rect 3745 984 3803 1009
rect 3745 950 3757 984
rect 3791 950 3803 984
rect 3745 916 3803 950
rect 3745 882 3757 916
rect 3791 882 3803 916
rect 3745 848 3803 882
rect 3745 814 3757 848
rect 3791 814 3803 848
rect 3745 780 3803 814
rect 3745 746 3757 780
rect 3791 746 3803 780
rect 3745 712 3803 746
rect 3745 678 3757 712
rect 3791 678 3803 712
rect 3745 644 3803 678
rect 3745 610 3757 644
rect 3791 610 3803 644
rect 3745 576 3803 610
rect 3745 542 3757 576
rect 3791 542 3803 576
rect 3745 508 3803 542
rect 3745 474 3757 508
rect 3791 474 3803 508
rect 3745 440 3803 474
rect 3745 406 3757 440
rect 3791 406 3803 440
rect 3745 372 3803 406
rect 3745 338 3757 372
rect 3791 338 3803 372
rect 3745 304 3803 338
rect 3745 270 3757 304
rect 3791 270 3803 304
rect 3745 236 3803 270
rect 3745 202 3757 236
rect 3791 202 3803 236
rect 3745 168 3803 202
rect 3745 134 3757 168
rect 3791 134 3803 168
rect 3745 109 3803 134
rect 3893 984 3951 1009
rect 3893 950 3905 984
rect 3939 950 3951 984
rect 3893 916 3951 950
rect 3893 882 3905 916
rect 3939 882 3951 916
rect 3893 848 3951 882
rect 3893 814 3905 848
rect 3939 814 3951 848
rect 3893 780 3951 814
rect 3893 746 3905 780
rect 3939 746 3951 780
rect 3893 712 3951 746
rect 3893 678 3905 712
rect 3939 678 3951 712
rect 3893 644 3951 678
rect 3893 610 3905 644
rect 3939 610 3951 644
rect 3893 576 3951 610
rect 3893 542 3905 576
rect 3939 542 3951 576
rect 3893 508 3951 542
rect 3893 474 3905 508
rect 3939 474 3951 508
rect 3893 440 3951 474
rect 3893 406 3905 440
rect 3939 406 3951 440
rect 3893 372 3951 406
rect 3893 338 3905 372
rect 3939 338 3951 372
rect 3893 304 3951 338
rect 3893 270 3905 304
rect 3939 270 3951 304
rect 3893 236 3951 270
rect 3893 202 3905 236
rect 3939 202 3951 236
rect 3893 168 3951 202
rect 3893 134 3905 168
rect 3939 134 3951 168
rect 3893 109 3951 134
rect 4041 984 4099 1009
rect 4041 950 4053 984
rect 4087 950 4099 984
rect 4041 916 4099 950
rect 4041 882 4053 916
rect 4087 882 4099 916
rect 4041 848 4099 882
rect 4041 814 4053 848
rect 4087 814 4099 848
rect 4041 780 4099 814
rect 4041 746 4053 780
rect 4087 746 4099 780
rect 4041 712 4099 746
rect 4041 678 4053 712
rect 4087 678 4099 712
rect 4041 644 4099 678
rect 4041 610 4053 644
rect 4087 610 4099 644
rect 4041 576 4099 610
rect 4041 542 4053 576
rect 4087 542 4099 576
rect 4041 508 4099 542
rect 4041 474 4053 508
rect 4087 474 4099 508
rect 4041 440 4099 474
rect 4041 406 4053 440
rect 4087 406 4099 440
rect 4041 372 4099 406
rect 4041 338 4053 372
rect 4087 338 4099 372
rect 4041 304 4099 338
rect 4041 270 4053 304
rect 4087 270 4099 304
rect 4041 236 4099 270
rect 4041 202 4053 236
rect 4087 202 4099 236
rect 4041 168 4099 202
rect 4041 134 4053 168
rect 4087 134 4099 168
rect 4041 109 4099 134
rect 4189 984 4247 1009
rect 4189 950 4201 984
rect 4235 950 4247 984
rect 4189 916 4247 950
rect 4189 882 4201 916
rect 4235 882 4247 916
rect 4189 848 4247 882
rect 4189 814 4201 848
rect 4235 814 4247 848
rect 4189 780 4247 814
rect 4189 746 4201 780
rect 4235 746 4247 780
rect 4189 712 4247 746
rect 4189 678 4201 712
rect 4235 678 4247 712
rect 4189 644 4247 678
rect 4189 610 4201 644
rect 4235 610 4247 644
rect 4189 576 4247 610
rect 4189 542 4201 576
rect 4235 542 4247 576
rect 4189 508 4247 542
rect 4189 474 4201 508
rect 4235 474 4247 508
rect 4189 440 4247 474
rect 4189 406 4201 440
rect 4235 406 4247 440
rect 4189 372 4247 406
rect 4189 338 4201 372
rect 4235 338 4247 372
rect 4189 304 4247 338
rect 4189 270 4201 304
rect 4235 270 4247 304
rect 4189 236 4247 270
rect 4189 202 4201 236
rect 4235 202 4247 236
rect 4189 168 4247 202
rect 4189 134 4201 168
rect 4235 134 4247 168
rect 4189 109 4247 134
rect 4337 984 4395 1009
rect 4337 950 4349 984
rect 4383 950 4395 984
rect 4337 916 4395 950
rect 4337 882 4349 916
rect 4383 882 4395 916
rect 4337 848 4395 882
rect 4337 814 4349 848
rect 4383 814 4395 848
rect 4337 780 4395 814
rect 4337 746 4349 780
rect 4383 746 4395 780
rect 4337 712 4395 746
rect 4337 678 4349 712
rect 4383 678 4395 712
rect 4337 644 4395 678
rect 4337 610 4349 644
rect 4383 610 4395 644
rect 4337 576 4395 610
rect 4337 542 4349 576
rect 4383 542 4395 576
rect 4337 508 4395 542
rect 4337 474 4349 508
rect 4383 474 4395 508
rect 4337 440 4395 474
rect 4337 406 4349 440
rect 4383 406 4395 440
rect 4337 372 4395 406
rect 4337 338 4349 372
rect 4383 338 4395 372
rect 4337 304 4395 338
rect 4337 270 4349 304
rect 4383 270 4395 304
rect 4337 236 4395 270
rect 4337 202 4349 236
rect 4383 202 4395 236
rect 4337 168 4395 202
rect 4337 134 4349 168
rect 4383 134 4395 168
rect 4337 109 4395 134
rect 4485 984 4543 1009
rect 4485 950 4497 984
rect 4531 950 4543 984
rect 4485 916 4543 950
rect 4485 882 4497 916
rect 4531 882 4543 916
rect 4485 848 4543 882
rect 4485 814 4497 848
rect 4531 814 4543 848
rect 4485 780 4543 814
rect 4485 746 4497 780
rect 4531 746 4543 780
rect 4485 712 4543 746
rect 4485 678 4497 712
rect 4531 678 4543 712
rect 4485 644 4543 678
rect 4485 610 4497 644
rect 4531 610 4543 644
rect 4485 576 4543 610
rect 4485 542 4497 576
rect 4531 542 4543 576
rect 4485 508 4543 542
rect 4485 474 4497 508
rect 4531 474 4543 508
rect 4485 440 4543 474
rect 4485 406 4497 440
rect 4531 406 4543 440
rect 4485 372 4543 406
rect 4485 338 4497 372
rect 4531 338 4543 372
rect 4485 304 4543 338
rect 4485 270 4497 304
rect 4531 270 4543 304
rect 4485 236 4543 270
rect 4485 202 4497 236
rect 4531 202 4543 236
rect 4485 168 4543 202
rect 4485 134 4497 168
rect 4531 134 4543 168
rect 4485 109 4543 134
rect 4633 984 4691 1009
rect 4633 950 4645 984
rect 4679 950 4691 984
rect 4633 916 4691 950
rect 4633 882 4645 916
rect 4679 882 4691 916
rect 4633 848 4691 882
rect 4633 814 4645 848
rect 4679 814 4691 848
rect 4633 780 4691 814
rect 4633 746 4645 780
rect 4679 746 4691 780
rect 4633 712 4691 746
rect 4633 678 4645 712
rect 4679 678 4691 712
rect 4633 644 4691 678
rect 4633 610 4645 644
rect 4679 610 4691 644
rect 4633 576 4691 610
rect 4633 542 4645 576
rect 4679 542 4691 576
rect 4633 508 4691 542
rect 4633 474 4645 508
rect 4679 474 4691 508
rect 4633 440 4691 474
rect 4633 406 4645 440
rect 4679 406 4691 440
rect 4633 372 4691 406
rect 4633 338 4645 372
rect 4679 338 4691 372
rect 4633 304 4691 338
rect 4633 270 4645 304
rect 4679 270 4691 304
rect 4633 236 4691 270
rect 4633 202 4645 236
rect 4679 202 4691 236
rect 4633 168 4691 202
rect 4633 134 4645 168
rect 4679 134 4691 168
rect 4633 109 4691 134
rect 4781 984 4839 1009
rect 4781 950 4793 984
rect 4827 950 4839 984
rect 4781 916 4839 950
rect 4781 882 4793 916
rect 4827 882 4839 916
rect 4781 848 4839 882
rect 4781 814 4793 848
rect 4827 814 4839 848
rect 4781 780 4839 814
rect 4781 746 4793 780
rect 4827 746 4839 780
rect 4781 712 4839 746
rect 4781 678 4793 712
rect 4827 678 4839 712
rect 4781 644 4839 678
rect 4781 610 4793 644
rect 4827 610 4839 644
rect 4781 576 4839 610
rect 4781 542 4793 576
rect 4827 542 4839 576
rect 4781 508 4839 542
rect 4781 474 4793 508
rect 4827 474 4839 508
rect 4781 440 4839 474
rect 4781 406 4793 440
rect 4827 406 4839 440
rect 4781 372 4839 406
rect 4781 338 4793 372
rect 4827 338 4839 372
rect 4781 304 4839 338
rect 4781 270 4793 304
rect 4827 270 4839 304
rect 4781 236 4839 270
rect 4781 202 4793 236
rect 4827 202 4839 236
rect 4781 168 4839 202
rect 4781 134 4793 168
rect 4827 134 4839 168
rect 4781 109 4839 134
rect 4929 984 4987 1009
rect 4929 950 4941 984
rect 4975 950 4987 984
rect 4929 916 4987 950
rect 4929 882 4941 916
rect 4975 882 4987 916
rect 4929 848 4987 882
rect 4929 814 4941 848
rect 4975 814 4987 848
rect 4929 780 4987 814
rect 4929 746 4941 780
rect 4975 746 4987 780
rect 4929 712 4987 746
rect 4929 678 4941 712
rect 4975 678 4987 712
rect 4929 644 4987 678
rect 4929 610 4941 644
rect 4975 610 4987 644
rect 4929 576 4987 610
rect 4929 542 4941 576
rect 4975 542 4987 576
rect 4929 508 4987 542
rect 4929 474 4941 508
rect 4975 474 4987 508
rect 4929 440 4987 474
rect 4929 406 4941 440
rect 4975 406 4987 440
rect 4929 372 4987 406
rect 4929 338 4941 372
rect 4975 338 4987 372
rect 4929 304 4987 338
rect 4929 270 4941 304
rect 4975 270 4987 304
rect 4929 236 4987 270
rect 4929 202 4941 236
rect 4975 202 4987 236
rect 4929 168 4987 202
rect 4929 134 4941 168
rect 4975 134 4987 168
rect 4929 109 4987 134
rect 5077 984 5135 1009
rect 5077 950 5089 984
rect 5123 950 5135 984
rect 5077 916 5135 950
rect 5077 882 5089 916
rect 5123 882 5135 916
rect 5077 848 5135 882
rect 5077 814 5089 848
rect 5123 814 5135 848
rect 5077 780 5135 814
rect 5077 746 5089 780
rect 5123 746 5135 780
rect 5077 712 5135 746
rect 5077 678 5089 712
rect 5123 678 5135 712
rect 5077 644 5135 678
rect 5077 610 5089 644
rect 5123 610 5135 644
rect 5077 576 5135 610
rect 5077 542 5089 576
rect 5123 542 5135 576
rect 5077 508 5135 542
rect 5077 474 5089 508
rect 5123 474 5135 508
rect 5077 440 5135 474
rect 5077 406 5089 440
rect 5123 406 5135 440
rect 5077 372 5135 406
rect 5077 338 5089 372
rect 5123 338 5135 372
rect 5077 304 5135 338
rect 5077 270 5089 304
rect 5123 270 5135 304
rect 5077 236 5135 270
rect 5077 202 5089 236
rect 5123 202 5135 236
rect 5077 168 5135 202
rect 5077 134 5089 168
rect 5123 134 5135 168
rect 5077 109 5135 134
rect 5225 984 5283 1009
rect 5225 950 5237 984
rect 5271 950 5283 984
rect 5225 916 5283 950
rect 5225 882 5237 916
rect 5271 882 5283 916
rect 5225 848 5283 882
rect 5225 814 5237 848
rect 5271 814 5283 848
rect 5225 780 5283 814
rect 5225 746 5237 780
rect 5271 746 5283 780
rect 5225 712 5283 746
rect 5225 678 5237 712
rect 5271 678 5283 712
rect 5225 644 5283 678
rect 5225 610 5237 644
rect 5271 610 5283 644
rect 5225 576 5283 610
rect 5225 542 5237 576
rect 5271 542 5283 576
rect 5225 508 5283 542
rect 5225 474 5237 508
rect 5271 474 5283 508
rect 5225 440 5283 474
rect 5225 406 5237 440
rect 5271 406 5283 440
rect 5225 372 5283 406
rect 5225 338 5237 372
rect 5271 338 5283 372
rect 5225 304 5283 338
rect 5225 270 5237 304
rect 5271 270 5283 304
rect 5225 236 5283 270
rect 5225 202 5237 236
rect 5271 202 5283 236
rect 5225 168 5283 202
rect 5225 134 5237 168
rect 5271 134 5283 168
rect 5225 109 5283 134
rect 5373 984 5431 1009
rect 5373 950 5385 984
rect 5419 950 5431 984
rect 5373 916 5431 950
rect 5373 882 5385 916
rect 5419 882 5431 916
rect 5373 848 5431 882
rect 5373 814 5385 848
rect 5419 814 5431 848
rect 5373 780 5431 814
rect 5373 746 5385 780
rect 5419 746 5431 780
rect 5373 712 5431 746
rect 5373 678 5385 712
rect 5419 678 5431 712
rect 5373 644 5431 678
rect 5373 610 5385 644
rect 5419 610 5431 644
rect 5373 576 5431 610
rect 5373 542 5385 576
rect 5419 542 5431 576
rect 5373 508 5431 542
rect 5373 474 5385 508
rect 5419 474 5431 508
rect 5373 440 5431 474
rect 5373 406 5385 440
rect 5419 406 5431 440
rect 5373 372 5431 406
rect 5373 338 5385 372
rect 5419 338 5431 372
rect 5373 304 5431 338
rect 5373 270 5385 304
rect 5419 270 5431 304
rect 5373 236 5431 270
rect 5373 202 5385 236
rect 5419 202 5431 236
rect 5373 168 5431 202
rect 5373 134 5385 168
rect 5419 134 5431 168
rect 5373 109 5431 134
rect 5521 984 5579 1009
rect 5521 950 5533 984
rect 5567 950 5579 984
rect 5521 916 5579 950
rect 5521 882 5533 916
rect 5567 882 5579 916
rect 5521 848 5579 882
rect 5521 814 5533 848
rect 5567 814 5579 848
rect 5521 780 5579 814
rect 5521 746 5533 780
rect 5567 746 5579 780
rect 5521 712 5579 746
rect 5521 678 5533 712
rect 5567 678 5579 712
rect 5521 644 5579 678
rect 5521 610 5533 644
rect 5567 610 5579 644
rect 5521 576 5579 610
rect 5521 542 5533 576
rect 5567 542 5579 576
rect 5521 508 5579 542
rect 5521 474 5533 508
rect 5567 474 5579 508
rect 5521 440 5579 474
rect 5521 406 5533 440
rect 5567 406 5579 440
rect 5521 372 5579 406
rect 5521 338 5533 372
rect 5567 338 5579 372
rect 5521 304 5579 338
rect 5521 270 5533 304
rect 5567 270 5579 304
rect 5521 236 5579 270
rect 5521 202 5533 236
rect 5567 202 5579 236
rect 5521 168 5579 202
rect 5521 134 5533 168
rect 5567 134 5579 168
rect 5521 109 5579 134
rect -5579 -134 -5521 -109
rect -5579 -168 -5567 -134
rect -5533 -168 -5521 -134
rect -5579 -202 -5521 -168
rect -5579 -236 -5567 -202
rect -5533 -236 -5521 -202
rect -5579 -270 -5521 -236
rect -5579 -304 -5567 -270
rect -5533 -304 -5521 -270
rect -5579 -338 -5521 -304
rect -5579 -372 -5567 -338
rect -5533 -372 -5521 -338
rect -5579 -406 -5521 -372
rect -5579 -440 -5567 -406
rect -5533 -440 -5521 -406
rect -5579 -474 -5521 -440
rect -5579 -508 -5567 -474
rect -5533 -508 -5521 -474
rect -5579 -542 -5521 -508
rect -5579 -576 -5567 -542
rect -5533 -576 -5521 -542
rect -5579 -610 -5521 -576
rect -5579 -644 -5567 -610
rect -5533 -644 -5521 -610
rect -5579 -678 -5521 -644
rect -5579 -712 -5567 -678
rect -5533 -712 -5521 -678
rect -5579 -746 -5521 -712
rect -5579 -780 -5567 -746
rect -5533 -780 -5521 -746
rect -5579 -814 -5521 -780
rect -5579 -848 -5567 -814
rect -5533 -848 -5521 -814
rect -5579 -882 -5521 -848
rect -5579 -916 -5567 -882
rect -5533 -916 -5521 -882
rect -5579 -950 -5521 -916
rect -5579 -984 -5567 -950
rect -5533 -984 -5521 -950
rect -5579 -1009 -5521 -984
rect -5431 -134 -5373 -109
rect -5431 -168 -5419 -134
rect -5385 -168 -5373 -134
rect -5431 -202 -5373 -168
rect -5431 -236 -5419 -202
rect -5385 -236 -5373 -202
rect -5431 -270 -5373 -236
rect -5431 -304 -5419 -270
rect -5385 -304 -5373 -270
rect -5431 -338 -5373 -304
rect -5431 -372 -5419 -338
rect -5385 -372 -5373 -338
rect -5431 -406 -5373 -372
rect -5431 -440 -5419 -406
rect -5385 -440 -5373 -406
rect -5431 -474 -5373 -440
rect -5431 -508 -5419 -474
rect -5385 -508 -5373 -474
rect -5431 -542 -5373 -508
rect -5431 -576 -5419 -542
rect -5385 -576 -5373 -542
rect -5431 -610 -5373 -576
rect -5431 -644 -5419 -610
rect -5385 -644 -5373 -610
rect -5431 -678 -5373 -644
rect -5431 -712 -5419 -678
rect -5385 -712 -5373 -678
rect -5431 -746 -5373 -712
rect -5431 -780 -5419 -746
rect -5385 -780 -5373 -746
rect -5431 -814 -5373 -780
rect -5431 -848 -5419 -814
rect -5385 -848 -5373 -814
rect -5431 -882 -5373 -848
rect -5431 -916 -5419 -882
rect -5385 -916 -5373 -882
rect -5431 -950 -5373 -916
rect -5431 -984 -5419 -950
rect -5385 -984 -5373 -950
rect -5431 -1009 -5373 -984
rect -5283 -134 -5225 -109
rect -5283 -168 -5271 -134
rect -5237 -168 -5225 -134
rect -5283 -202 -5225 -168
rect -5283 -236 -5271 -202
rect -5237 -236 -5225 -202
rect -5283 -270 -5225 -236
rect -5283 -304 -5271 -270
rect -5237 -304 -5225 -270
rect -5283 -338 -5225 -304
rect -5283 -372 -5271 -338
rect -5237 -372 -5225 -338
rect -5283 -406 -5225 -372
rect -5283 -440 -5271 -406
rect -5237 -440 -5225 -406
rect -5283 -474 -5225 -440
rect -5283 -508 -5271 -474
rect -5237 -508 -5225 -474
rect -5283 -542 -5225 -508
rect -5283 -576 -5271 -542
rect -5237 -576 -5225 -542
rect -5283 -610 -5225 -576
rect -5283 -644 -5271 -610
rect -5237 -644 -5225 -610
rect -5283 -678 -5225 -644
rect -5283 -712 -5271 -678
rect -5237 -712 -5225 -678
rect -5283 -746 -5225 -712
rect -5283 -780 -5271 -746
rect -5237 -780 -5225 -746
rect -5283 -814 -5225 -780
rect -5283 -848 -5271 -814
rect -5237 -848 -5225 -814
rect -5283 -882 -5225 -848
rect -5283 -916 -5271 -882
rect -5237 -916 -5225 -882
rect -5283 -950 -5225 -916
rect -5283 -984 -5271 -950
rect -5237 -984 -5225 -950
rect -5283 -1009 -5225 -984
rect -5135 -134 -5077 -109
rect -5135 -168 -5123 -134
rect -5089 -168 -5077 -134
rect -5135 -202 -5077 -168
rect -5135 -236 -5123 -202
rect -5089 -236 -5077 -202
rect -5135 -270 -5077 -236
rect -5135 -304 -5123 -270
rect -5089 -304 -5077 -270
rect -5135 -338 -5077 -304
rect -5135 -372 -5123 -338
rect -5089 -372 -5077 -338
rect -5135 -406 -5077 -372
rect -5135 -440 -5123 -406
rect -5089 -440 -5077 -406
rect -5135 -474 -5077 -440
rect -5135 -508 -5123 -474
rect -5089 -508 -5077 -474
rect -5135 -542 -5077 -508
rect -5135 -576 -5123 -542
rect -5089 -576 -5077 -542
rect -5135 -610 -5077 -576
rect -5135 -644 -5123 -610
rect -5089 -644 -5077 -610
rect -5135 -678 -5077 -644
rect -5135 -712 -5123 -678
rect -5089 -712 -5077 -678
rect -5135 -746 -5077 -712
rect -5135 -780 -5123 -746
rect -5089 -780 -5077 -746
rect -5135 -814 -5077 -780
rect -5135 -848 -5123 -814
rect -5089 -848 -5077 -814
rect -5135 -882 -5077 -848
rect -5135 -916 -5123 -882
rect -5089 -916 -5077 -882
rect -5135 -950 -5077 -916
rect -5135 -984 -5123 -950
rect -5089 -984 -5077 -950
rect -5135 -1009 -5077 -984
rect -4987 -134 -4929 -109
rect -4987 -168 -4975 -134
rect -4941 -168 -4929 -134
rect -4987 -202 -4929 -168
rect -4987 -236 -4975 -202
rect -4941 -236 -4929 -202
rect -4987 -270 -4929 -236
rect -4987 -304 -4975 -270
rect -4941 -304 -4929 -270
rect -4987 -338 -4929 -304
rect -4987 -372 -4975 -338
rect -4941 -372 -4929 -338
rect -4987 -406 -4929 -372
rect -4987 -440 -4975 -406
rect -4941 -440 -4929 -406
rect -4987 -474 -4929 -440
rect -4987 -508 -4975 -474
rect -4941 -508 -4929 -474
rect -4987 -542 -4929 -508
rect -4987 -576 -4975 -542
rect -4941 -576 -4929 -542
rect -4987 -610 -4929 -576
rect -4987 -644 -4975 -610
rect -4941 -644 -4929 -610
rect -4987 -678 -4929 -644
rect -4987 -712 -4975 -678
rect -4941 -712 -4929 -678
rect -4987 -746 -4929 -712
rect -4987 -780 -4975 -746
rect -4941 -780 -4929 -746
rect -4987 -814 -4929 -780
rect -4987 -848 -4975 -814
rect -4941 -848 -4929 -814
rect -4987 -882 -4929 -848
rect -4987 -916 -4975 -882
rect -4941 -916 -4929 -882
rect -4987 -950 -4929 -916
rect -4987 -984 -4975 -950
rect -4941 -984 -4929 -950
rect -4987 -1009 -4929 -984
rect -4839 -134 -4781 -109
rect -4839 -168 -4827 -134
rect -4793 -168 -4781 -134
rect -4839 -202 -4781 -168
rect -4839 -236 -4827 -202
rect -4793 -236 -4781 -202
rect -4839 -270 -4781 -236
rect -4839 -304 -4827 -270
rect -4793 -304 -4781 -270
rect -4839 -338 -4781 -304
rect -4839 -372 -4827 -338
rect -4793 -372 -4781 -338
rect -4839 -406 -4781 -372
rect -4839 -440 -4827 -406
rect -4793 -440 -4781 -406
rect -4839 -474 -4781 -440
rect -4839 -508 -4827 -474
rect -4793 -508 -4781 -474
rect -4839 -542 -4781 -508
rect -4839 -576 -4827 -542
rect -4793 -576 -4781 -542
rect -4839 -610 -4781 -576
rect -4839 -644 -4827 -610
rect -4793 -644 -4781 -610
rect -4839 -678 -4781 -644
rect -4839 -712 -4827 -678
rect -4793 -712 -4781 -678
rect -4839 -746 -4781 -712
rect -4839 -780 -4827 -746
rect -4793 -780 -4781 -746
rect -4839 -814 -4781 -780
rect -4839 -848 -4827 -814
rect -4793 -848 -4781 -814
rect -4839 -882 -4781 -848
rect -4839 -916 -4827 -882
rect -4793 -916 -4781 -882
rect -4839 -950 -4781 -916
rect -4839 -984 -4827 -950
rect -4793 -984 -4781 -950
rect -4839 -1009 -4781 -984
rect -4691 -134 -4633 -109
rect -4691 -168 -4679 -134
rect -4645 -168 -4633 -134
rect -4691 -202 -4633 -168
rect -4691 -236 -4679 -202
rect -4645 -236 -4633 -202
rect -4691 -270 -4633 -236
rect -4691 -304 -4679 -270
rect -4645 -304 -4633 -270
rect -4691 -338 -4633 -304
rect -4691 -372 -4679 -338
rect -4645 -372 -4633 -338
rect -4691 -406 -4633 -372
rect -4691 -440 -4679 -406
rect -4645 -440 -4633 -406
rect -4691 -474 -4633 -440
rect -4691 -508 -4679 -474
rect -4645 -508 -4633 -474
rect -4691 -542 -4633 -508
rect -4691 -576 -4679 -542
rect -4645 -576 -4633 -542
rect -4691 -610 -4633 -576
rect -4691 -644 -4679 -610
rect -4645 -644 -4633 -610
rect -4691 -678 -4633 -644
rect -4691 -712 -4679 -678
rect -4645 -712 -4633 -678
rect -4691 -746 -4633 -712
rect -4691 -780 -4679 -746
rect -4645 -780 -4633 -746
rect -4691 -814 -4633 -780
rect -4691 -848 -4679 -814
rect -4645 -848 -4633 -814
rect -4691 -882 -4633 -848
rect -4691 -916 -4679 -882
rect -4645 -916 -4633 -882
rect -4691 -950 -4633 -916
rect -4691 -984 -4679 -950
rect -4645 -984 -4633 -950
rect -4691 -1009 -4633 -984
rect -4543 -134 -4485 -109
rect -4543 -168 -4531 -134
rect -4497 -168 -4485 -134
rect -4543 -202 -4485 -168
rect -4543 -236 -4531 -202
rect -4497 -236 -4485 -202
rect -4543 -270 -4485 -236
rect -4543 -304 -4531 -270
rect -4497 -304 -4485 -270
rect -4543 -338 -4485 -304
rect -4543 -372 -4531 -338
rect -4497 -372 -4485 -338
rect -4543 -406 -4485 -372
rect -4543 -440 -4531 -406
rect -4497 -440 -4485 -406
rect -4543 -474 -4485 -440
rect -4543 -508 -4531 -474
rect -4497 -508 -4485 -474
rect -4543 -542 -4485 -508
rect -4543 -576 -4531 -542
rect -4497 -576 -4485 -542
rect -4543 -610 -4485 -576
rect -4543 -644 -4531 -610
rect -4497 -644 -4485 -610
rect -4543 -678 -4485 -644
rect -4543 -712 -4531 -678
rect -4497 -712 -4485 -678
rect -4543 -746 -4485 -712
rect -4543 -780 -4531 -746
rect -4497 -780 -4485 -746
rect -4543 -814 -4485 -780
rect -4543 -848 -4531 -814
rect -4497 -848 -4485 -814
rect -4543 -882 -4485 -848
rect -4543 -916 -4531 -882
rect -4497 -916 -4485 -882
rect -4543 -950 -4485 -916
rect -4543 -984 -4531 -950
rect -4497 -984 -4485 -950
rect -4543 -1009 -4485 -984
rect -4395 -134 -4337 -109
rect -4395 -168 -4383 -134
rect -4349 -168 -4337 -134
rect -4395 -202 -4337 -168
rect -4395 -236 -4383 -202
rect -4349 -236 -4337 -202
rect -4395 -270 -4337 -236
rect -4395 -304 -4383 -270
rect -4349 -304 -4337 -270
rect -4395 -338 -4337 -304
rect -4395 -372 -4383 -338
rect -4349 -372 -4337 -338
rect -4395 -406 -4337 -372
rect -4395 -440 -4383 -406
rect -4349 -440 -4337 -406
rect -4395 -474 -4337 -440
rect -4395 -508 -4383 -474
rect -4349 -508 -4337 -474
rect -4395 -542 -4337 -508
rect -4395 -576 -4383 -542
rect -4349 -576 -4337 -542
rect -4395 -610 -4337 -576
rect -4395 -644 -4383 -610
rect -4349 -644 -4337 -610
rect -4395 -678 -4337 -644
rect -4395 -712 -4383 -678
rect -4349 -712 -4337 -678
rect -4395 -746 -4337 -712
rect -4395 -780 -4383 -746
rect -4349 -780 -4337 -746
rect -4395 -814 -4337 -780
rect -4395 -848 -4383 -814
rect -4349 -848 -4337 -814
rect -4395 -882 -4337 -848
rect -4395 -916 -4383 -882
rect -4349 -916 -4337 -882
rect -4395 -950 -4337 -916
rect -4395 -984 -4383 -950
rect -4349 -984 -4337 -950
rect -4395 -1009 -4337 -984
rect -4247 -134 -4189 -109
rect -4247 -168 -4235 -134
rect -4201 -168 -4189 -134
rect -4247 -202 -4189 -168
rect -4247 -236 -4235 -202
rect -4201 -236 -4189 -202
rect -4247 -270 -4189 -236
rect -4247 -304 -4235 -270
rect -4201 -304 -4189 -270
rect -4247 -338 -4189 -304
rect -4247 -372 -4235 -338
rect -4201 -372 -4189 -338
rect -4247 -406 -4189 -372
rect -4247 -440 -4235 -406
rect -4201 -440 -4189 -406
rect -4247 -474 -4189 -440
rect -4247 -508 -4235 -474
rect -4201 -508 -4189 -474
rect -4247 -542 -4189 -508
rect -4247 -576 -4235 -542
rect -4201 -576 -4189 -542
rect -4247 -610 -4189 -576
rect -4247 -644 -4235 -610
rect -4201 -644 -4189 -610
rect -4247 -678 -4189 -644
rect -4247 -712 -4235 -678
rect -4201 -712 -4189 -678
rect -4247 -746 -4189 -712
rect -4247 -780 -4235 -746
rect -4201 -780 -4189 -746
rect -4247 -814 -4189 -780
rect -4247 -848 -4235 -814
rect -4201 -848 -4189 -814
rect -4247 -882 -4189 -848
rect -4247 -916 -4235 -882
rect -4201 -916 -4189 -882
rect -4247 -950 -4189 -916
rect -4247 -984 -4235 -950
rect -4201 -984 -4189 -950
rect -4247 -1009 -4189 -984
rect -4099 -134 -4041 -109
rect -4099 -168 -4087 -134
rect -4053 -168 -4041 -134
rect -4099 -202 -4041 -168
rect -4099 -236 -4087 -202
rect -4053 -236 -4041 -202
rect -4099 -270 -4041 -236
rect -4099 -304 -4087 -270
rect -4053 -304 -4041 -270
rect -4099 -338 -4041 -304
rect -4099 -372 -4087 -338
rect -4053 -372 -4041 -338
rect -4099 -406 -4041 -372
rect -4099 -440 -4087 -406
rect -4053 -440 -4041 -406
rect -4099 -474 -4041 -440
rect -4099 -508 -4087 -474
rect -4053 -508 -4041 -474
rect -4099 -542 -4041 -508
rect -4099 -576 -4087 -542
rect -4053 -576 -4041 -542
rect -4099 -610 -4041 -576
rect -4099 -644 -4087 -610
rect -4053 -644 -4041 -610
rect -4099 -678 -4041 -644
rect -4099 -712 -4087 -678
rect -4053 -712 -4041 -678
rect -4099 -746 -4041 -712
rect -4099 -780 -4087 -746
rect -4053 -780 -4041 -746
rect -4099 -814 -4041 -780
rect -4099 -848 -4087 -814
rect -4053 -848 -4041 -814
rect -4099 -882 -4041 -848
rect -4099 -916 -4087 -882
rect -4053 -916 -4041 -882
rect -4099 -950 -4041 -916
rect -4099 -984 -4087 -950
rect -4053 -984 -4041 -950
rect -4099 -1009 -4041 -984
rect -3951 -134 -3893 -109
rect -3951 -168 -3939 -134
rect -3905 -168 -3893 -134
rect -3951 -202 -3893 -168
rect -3951 -236 -3939 -202
rect -3905 -236 -3893 -202
rect -3951 -270 -3893 -236
rect -3951 -304 -3939 -270
rect -3905 -304 -3893 -270
rect -3951 -338 -3893 -304
rect -3951 -372 -3939 -338
rect -3905 -372 -3893 -338
rect -3951 -406 -3893 -372
rect -3951 -440 -3939 -406
rect -3905 -440 -3893 -406
rect -3951 -474 -3893 -440
rect -3951 -508 -3939 -474
rect -3905 -508 -3893 -474
rect -3951 -542 -3893 -508
rect -3951 -576 -3939 -542
rect -3905 -576 -3893 -542
rect -3951 -610 -3893 -576
rect -3951 -644 -3939 -610
rect -3905 -644 -3893 -610
rect -3951 -678 -3893 -644
rect -3951 -712 -3939 -678
rect -3905 -712 -3893 -678
rect -3951 -746 -3893 -712
rect -3951 -780 -3939 -746
rect -3905 -780 -3893 -746
rect -3951 -814 -3893 -780
rect -3951 -848 -3939 -814
rect -3905 -848 -3893 -814
rect -3951 -882 -3893 -848
rect -3951 -916 -3939 -882
rect -3905 -916 -3893 -882
rect -3951 -950 -3893 -916
rect -3951 -984 -3939 -950
rect -3905 -984 -3893 -950
rect -3951 -1009 -3893 -984
rect -3803 -134 -3745 -109
rect -3803 -168 -3791 -134
rect -3757 -168 -3745 -134
rect -3803 -202 -3745 -168
rect -3803 -236 -3791 -202
rect -3757 -236 -3745 -202
rect -3803 -270 -3745 -236
rect -3803 -304 -3791 -270
rect -3757 -304 -3745 -270
rect -3803 -338 -3745 -304
rect -3803 -372 -3791 -338
rect -3757 -372 -3745 -338
rect -3803 -406 -3745 -372
rect -3803 -440 -3791 -406
rect -3757 -440 -3745 -406
rect -3803 -474 -3745 -440
rect -3803 -508 -3791 -474
rect -3757 -508 -3745 -474
rect -3803 -542 -3745 -508
rect -3803 -576 -3791 -542
rect -3757 -576 -3745 -542
rect -3803 -610 -3745 -576
rect -3803 -644 -3791 -610
rect -3757 -644 -3745 -610
rect -3803 -678 -3745 -644
rect -3803 -712 -3791 -678
rect -3757 -712 -3745 -678
rect -3803 -746 -3745 -712
rect -3803 -780 -3791 -746
rect -3757 -780 -3745 -746
rect -3803 -814 -3745 -780
rect -3803 -848 -3791 -814
rect -3757 -848 -3745 -814
rect -3803 -882 -3745 -848
rect -3803 -916 -3791 -882
rect -3757 -916 -3745 -882
rect -3803 -950 -3745 -916
rect -3803 -984 -3791 -950
rect -3757 -984 -3745 -950
rect -3803 -1009 -3745 -984
rect -3655 -134 -3597 -109
rect -3655 -168 -3643 -134
rect -3609 -168 -3597 -134
rect -3655 -202 -3597 -168
rect -3655 -236 -3643 -202
rect -3609 -236 -3597 -202
rect -3655 -270 -3597 -236
rect -3655 -304 -3643 -270
rect -3609 -304 -3597 -270
rect -3655 -338 -3597 -304
rect -3655 -372 -3643 -338
rect -3609 -372 -3597 -338
rect -3655 -406 -3597 -372
rect -3655 -440 -3643 -406
rect -3609 -440 -3597 -406
rect -3655 -474 -3597 -440
rect -3655 -508 -3643 -474
rect -3609 -508 -3597 -474
rect -3655 -542 -3597 -508
rect -3655 -576 -3643 -542
rect -3609 -576 -3597 -542
rect -3655 -610 -3597 -576
rect -3655 -644 -3643 -610
rect -3609 -644 -3597 -610
rect -3655 -678 -3597 -644
rect -3655 -712 -3643 -678
rect -3609 -712 -3597 -678
rect -3655 -746 -3597 -712
rect -3655 -780 -3643 -746
rect -3609 -780 -3597 -746
rect -3655 -814 -3597 -780
rect -3655 -848 -3643 -814
rect -3609 -848 -3597 -814
rect -3655 -882 -3597 -848
rect -3655 -916 -3643 -882
rect -3609 -916 -3597 -882
rect -3655 -950 -3597 -916
rect -3655 -984 -3643 -950
rect -3609 -984 -3597 -950
rect -3655 -1009 -3597 -984
rect -3507 -134 -3449 -109
rect -3507 -168 -3495 -134
rect -3461 -168 -3449 -134
rect -3507 -202 -3449 -168
rect -3507 -236 -3495 -202
rect -3461 -236 -3449 -202
rect -3507 -270 -3449 -236
rect -3507 -304 -3495 -270
rect -3461 -304 -3449 -270
rect -3507 -338 -3449 -304
rect -3507 -372 -3495 -338
rect -3461 -372 -3449 -338
rect -3507 -406 -3449 -372
rect -3507 -440 -3495 -406
rect -3461 -440 -3449 -406
rect -3507 -474 -3449 -440
rect -3507 -508 -3495 -474
rect -3461 -508 -3449 -474
rect -3507 -542 -3449 -508
rect -3507 -576 -3495 -542
rect -3461 -576 -3449 -542
rect -3507 -610 -3449 -576
rect -3507 -644 -3495 -610
rect -3461 -644 -3449 -610
rect -3507 -678 -3449 -644
rect -3507 -712 -3495 -678
rect -3461 -712 -3449 -678
rect -3507 -746 -3449 -712
rect -3507 -780 -3495 -746
rect -3461 -780 -3449 -746
rect -3507 -814 -3449 -780
rect -3507 -848 -3495 -814
rect -3461 -848 -3449 -814
rect -3507 -882 -3449 -848
rect -3507 -916 -3495 -882
rect -3461 -916 -3449 -882
rect -3507 -950 -3449 -916
rect -3507 -984 -3495 -950
rect -3461 -984 -3449 -950
rect -3507 -1009 -3449 -984
rect -3359 -134 -3301 -109
rect -3359 -168 -3347 -134
rect -3313 -168 -3301 -134
rect -3359 -202 -3301 -168
rect -3359 -236 -3347 -202
rect -3313 -236 -3301 -202
rect -3359 -270 -3301 -236
rect -3359 -304 -3347 -270
rect -3313 -304 -3301 -270
rect -3359 -338 -3301 -304
rect -3359 -372 -3347 -338
rect -3313 -372 -3301 -338
rect -3359 -406 -3301 -372
rect -3359 -440 -3347 -406
rect -3313 -440 -3301 -406
rect -3359 -474 -3301 -440
rect -3359 -508 -3347 -474
rect -3313 -508 -3301 -474
rect -3359 -542 -3301 -508
rect -3359 -576 -3347 -542
rect -3313 -576 -3301 -542
rect -3359 -610 -3301 -576
rect -3359 -644 -3347 -610
rect -3313 -644 -3301 -610
rect -3359 -678 -3301 -644
rect -3359 -712 -3347 -678
rect -3313 -712 -3301 -678
rect -3359 -746 -3301 -712
rect -3359 -780 -3347 -746
rect -3313 -780 -3301 -746
rect -3359 -814 -3301 -780
rect -3359 -848 -3347 -814
rect -3313 -848 -3301 -814
rect -3359 -882 -3301 -848
rect -3359 -916 -3347 -882
rect -3313 -916 -3301 -882
rect -3359 -950 -3301 -916
rect -3359 -984 -3347 -950
rect -3313 -984 -3301 -950
rect -3359 -1009 -3301 -984
rect -3211 -134 -3153 -109
rect -3211 -168 -3199 -134
rect -3165 -168 -3153 -134
rect -3211 -202 -3153 -168
rect -3211 -236 -3199 -202
rect -3165 -236 -3153 -202
rect -3211 -270 -3153 -236
rect -3211 -304 -3199 -270
rect -3165 -304 -3153 -270
rect -3211 -338 -3153 -304
rect -3211 -372 -3199 -338
rect -3165 -372 -3153 -338
rect -3211 -406 -3153 -372
rect -3211 -440 -3199 -406
rect -3165 -440 -3153 -406
rect -3211 -474 -3153 -440
rect -3211 -508 -3199 -474
rect -3165 -508 -3153 -474
rect -3211 -542 -3153 -508
rect -3211 -576 -3199 -542
rect -3165 -576 -3153 -542
rect -3211 -610 -3153 -576
rect -3211 -644 -3199 -610
rect -3165 -644 -3153 -610
rect -3211 -678 -3153 -644
rect -3211 -712 -3199 -678
rect -3165 -712 -3153 -678
rect -3211 -746 -3153 -712
rect -3211 -780 -3199 -746
rect -3165 -780 -3153 -746
rect -3211 -814 -3153 -780
rect -3211 -848 -3199 -814
rect -3165 -848 -3153 -814
rect -3211 -882 -3153 -848
rect -3211 -916 -3199 -882
rect -3165 -916 -3153 -882
rect -3211 -950 -3153 -916
rect -3211 -984 -3199 -950
rect -3165 -984 -3153 -950
rect -3211 -1009 -3153 -984
rect -3063 -134 -3005 -109
rect -3063 -168 -3051 -134
rect -3017 -168 -3005 -134
rect -3063 -202 -3005 -168
rect -3063 -236 -3051 -202
rect -3017 -236 -3005 -202
rect -3063 -270 -3005 -236
rect -3063 -304 -3051 -270
rect -3017 -304 -3005 -270
rect -3063 -338 -3005 -304
rect -3063 -372 -3051 -338
rect -3017 -372 -3005 -338
rect -3063 -406 -3005 -372
rect -3063 -440 -3051 -406
rect -3017 -440 -3005 -406
rect -3063 -474 -3005 -440
rect -3063 -508 -3051 -474
rect -3017 -508 -3005 -474
rect -3063 -542 -3005 -508
rect -3063 -576 -3051 -542
rect -3017 -576 -3005 -542
rect -3063 -610 -3005 -576
rect -3063 -644 -3051 -610
rect -3017 -644 -3005 -610
rect -3063 -678 -3005 -644
rect -3063 -712 -3051 -678
rect -3017 -712 -3005 -678
rect -3063 -746 -3005 -712
rect -3063 -780 -3051 -746
rect -3017 -780 -3005 -746
rect -3063 -814 -3005 -780
rect -3063 -848 -3051 -814
rect -3017 -848 -3005 -814
rect -3063 -882 -3005 -848
rect -3063 -916 -3051 -882
rect -3017 -916 -3005 -882
rect -3063 -950 -3005 -916
rect -3063 -984 -3051 -950
rect -3017 -984 -3005 -950
rect -3063 -1009 -3005 -984
rect -2915 -134 -2857 -109
rect -2915 -168 -2903 -134
rect -2869 -168 -2857 -134
rect -2915 -202 -2857 -168
rect -2915 -236 -2903 -202
rect -2869 -236 -2857 -202
rect -2915 -270 -2857 -236
rect -2915 -304 -2903 -270
rect -2869 -304 -2857 -270
rect -2915 -338 -2857 -304
rect -2915 -372 -2903 -338
rect -2869 -372 -2857 -338
rect -2915 -406 -2857 -372
rect -2915 -440 -2903 -406
rect -2869 -440 -2857 -406
rect -2915 -474 -2857 -440
rect -2915 -508 -2903 -474
rect -2869 -508 -2857 -474
rect -2915 -542 -2857 -508
rect -2915 -576 -2903 -542
rect -2869 -576 -2857 -542
rect -2915 -610 -2857 -576
rect -2915 -644 -2903 -610
rect -2869 -644 -2857 -610
rect -2915 -678 -2857 -644
rect -2915 -712 -2903 -678
rect -2869 -712 -2857 -678
rect -2915 -746 -2857 -712
rect -2915 -780 -2903 -746
rect -2869 -780 -2857 -746
rect -2915 -814 -2857 -780
rect -2915 -848 -2903 -814
rect -2869 -848 -2857 -814
rect -2915 -882 -2857 -848
rect -2915 -916 -2903 -882
rect -2869 -916 -2857 -882
rect -2915 -950 -2857 -916
rect -2915 -984 -2903 -950
rect -2869 -984 -2857 -950
rect -2915 -1009 -2857 -984
rect -2767 -134 -2709 -109
rect -2767 -168 -2755 -134
rect -2721 -168 -2709 -134
rect -2767 -202 -2709 -168
rect -2767 -236 -2755 -202
rect -2721 -236 -2709 -202
rect -2767 -270 -2709 -236
rect -2767 -304 -2755 -270
rect -2721 -304 -2709 -270
rect -2767 -338 -2709 -304
rect -2767 -372 -2755 -338
rect -2721 -372 -2709 -338
rect -2767 -406 -2709 -372
rect -2767 -440 -2755 -406
rect -2721 -440 -2709 -406
rect -2767 -474 -2709 -440
rect -2767 -508 -2755 -474
rect -2721 -508 -2709 -474
rect -2767 -542 -2709 -508
rect -2767 -576 -2755 -542
rect -2721 -576 -2709 -542
rect -2767 -610 -2709 -576
rect -2767 -644 -2755 -610
rect -2721 -644 -2709 -610
rect -2767 -678 -2709 -644
rect -2767 -712 -2755 -678
rect -2721 -712 -2709 -678
rect -2767 -746 -2709 -712
rect -2767 -780 -2755 -746
rect -2721 -780 -2709 -746
rect -2767 -814 -2709 -780
rect -2767 -848 -2755 -814
rect -2721 -848 -2709 -814
rect -2767 -882 -2709 -848
rect -2767 -916 -2755 -882
rect -2721 -916 -2709 -882
rect -2767 -950 -2709 -916
rect -2767 -984 -2755 -950
rect -2721 -984 -2709 -950
rect -2767 -1009 -2709 -984
rect -2619 -134 -2561 -109
rect -2619 -168 -2607 -134
rect -2573 -168 -2561 -134
rect -2619 -202 -2561 -168
rect -2619 -236 -2607 -202
rect -2573 -236 -2561 -202
rect -2619 -270 -2561 -236
rect -2619 -304 -2607 -270
rect -2573 -304 -2561 -270
rect -2619 -338 -2561 -304
rect -2619 -372 -2607 -338
rect -2573 -372 -2561 -338
rect -2619 -406 -2561 -372
rect -2619 -440 -2607 -406
rect -2573 -440 -2561 -406
rect -2619 -474 -2561 -440
rect -2619 -508 -2607 -474
rect -2573 -508 -2561 -474
rect -2619 -542 -2561 -508
rect -2619 -576 -2607 -542
rect -2573 -576 -2561 -542
rect -2619 -610 -2561 -576
rect -2619 -644 -2607 -610
rect -2573 -644 -2561 -610
rect -2619 -678 -2561 -644
rect -2619 -712 -2607 -678
rect -2573 -712 -2561 -678
rect -2619 -746 -2561 -712
rect -2619 -780 -2607 -746
rect -2573 -780 -2561 -746
rect -2619 -814 -2561 -780
rect -2619 -848 -2607 -814
rect -2573 -848 -2561 -814
rect -2619 -882 -2561 -848
rect -2619 -916 -2607 -882
rect -2573 -916 -2561 -882
rect -2619 -950 -2561 -916
rect -2619 -984 -2607 -950
rect -2573 -984 -2561 -950
rect -2619 -1009 -2561 -984
rect -2471 -134 -2413 -109
rect -2471 -168 -2459 -134
rect -2425 -168 -2413 -134
rect -2471 -202 -2413 -168
rect -2471 -236 -2459 -202
rect -2425 -236 -2413 -202
rect -2471 -270 -2413 -236
rect -2471 -304 -2459 -270
rect -2425 -304 -2413 -270
rect -2471 -338 -2413 -304
rect -2471 -372 -2459 -338
rect -2425 -372 -2413 -338
rect -2471 -406 -2413 -372
rect -2471 -440 -2459 -406
rect -2425 -440 -2413 -406
rect -2471 -474 -2413 -440
rect -2471 -508 -2459 -474
rect -2425 -508 -2413 -474
rect -2471 -542 -2413 -508
rect -2471 -576 -2459 -542
rect -2425 -576 -2413 -542
rect -2471 -610 -2413 -576
rect -2471 -644 -2459 -610
rect -2425 -644 -2413 -610
rect -2471 -678 -2413 -644
rect -2471 -712 -2459 -678
rect -2425 -712 -2413 -678
rect -2471 -746 -2413 -712
rect -2471 -780 -2459 -746
rect -2425 -780 -2413 -746
rect -2471 -814 -2413 -780
rect -2471 -848 -2459 -814
rect -2425 -848 -2413 -814
rect -2471 -882 -2413 -848
rect -2471 -916 -2459 -882
rect -2425 -916 -2413 -882
rect -2471 -950 -2413 -916
rect -2471 -984 -2459 -950
rect -2425 -984 -2413 -950
rect -2471 -1009 -2413 -984
rect -2323 -134 -2265 -109
rect -2323 -168 -2311 -134
rect -2277 -168 -2265 -134
rect -2323 -202 -2265 -168
rect -2323 -236 -2311 -202
rect -2277 -236 -2265 -202
rect -2323 -270 -2265 -236
rect -2323 -304 -2311 -270
rect -2277 -304 -2265 -270
rect -2323 -338 -2265 -304
rect -2323 -372 -2311 -338
rect -2277 -372 -2265 -338
rect -2323 -406 -2265 -372
rect -2323 -440 -2311 -406
rect -2277 -440 -2265 -406
rect -2323 -474 -2265 -440
rect -2323 -508 -2311 -474
rect -2277 -508 -2265 -474
rect -2323 -542 -2265 -508
rect -2323 -576 -2311 -542
rect -2277 -576 -2265 -542
rect -2323 -610 -2265 -576
rect -2323 -644 -2311 -610
rect -2277 -644 -2265 -610
rect -2323 -678 -2265 -644
rect -2323 -712 -2311 -678
rect -2277 -712 -2265 -678
rect -2323 -746 -2265 -712
rect -2323 -780 -2311 -746
rect -2277 -780 -2265 -746
rect -2323 -814 -2265 -780
rect -2323 -848 -2311 -814
rect -2277 -848 -2265 -814
rect -2323 -882 -2265 -848
rect -2323 -916 -2311 -882
rect -2277 -916 -2265 -882
rect -2323 -950 -2265 -916
rect -2323 -984 -2311 -950
rect -2277 -984 -2265 -950
rect -2323 -1009 -2265 -984
rect -2175 -134 -2117 -109
rect -2175 -168 -2163 -134
rect -2129 -168 -2117 -134
rect -2175 -202 -2117 -168
rect -2175 -236 -2163 -202
rect -2129 -236 -2117 -202
rect -2175 -270 -2117 -236
rect -2175 -304 -2163 -270
rect -2129 -304 -2117 -270
rect -2175 -338 -2117 -304
rect -2175 -372 -2163 -338
rect -2129 -372 -2117 -338
rect -2175 -406 -2117 -372
rect -2175 -440 -2163 -406
rect -2129 -440 -2117 -406
rect -2175 -474 -2117 -440
rect -2175 -508 -2163 -474
rect -2129 -508 -2117 -474
rect -2175 -542 -2117 -508
rect -2175 -576 -2163 -542
rect -2129 -576 -2117 -542
rect -2175 -610 -2117 -576
rect -2175 -644 -2163 -610
rect -2129 -644 -2117 -610
rect -2175 -678 -2117 -644
rect -2175 -712 -2163 -678
rect -2129 -712 -2117 -678
rect -2175 -746 -2117 -712
rect -2175 -780 -2163 -746
rect -2129 -780 -2117 -746
rect -2175 -814 -2117 -780
rect -2175 -848 -2163 -814
rect -2129 -848 -2117 -814
rect -2175 -882 -2117 -848
rect -2175 -916 -2163 -882
rect -2129 -916 -2117 -882
rect -2175 -950 -2117 -916
rect -2175 -984 -2163 -950
rect -2129 -984 -2117 -950
rect -2175 -1009 -2117 -984
rect -2027 -134 -1969 -109
rect -2027 -168 -2015 -134
rect -1981 -168 -1969 -134
rect -2027 -202 -1969 -168
rect -2027 -236 -2015 -202
rect -1981 -236 -1969 -202
rect -2027 -270 -1969 -236
rect -2027 -304 -2015 -270
rect -1981 -304 -1969 -270
rect -2027 -338 -1969 -304
rect -2027 -372 -2015 -338
rect -1981 -372 -1969 -338
rect -2027 -406 -1969 -372
rect -2027 -440 -2015 -406
rect -1981 -440 -1969 -406
rect -2027 -474 -1969 -440
rect -2027 -508 -2015 -474
rect -1981 -508 -1969 -474
rect -2027 -542 -1969 -508
rect -2027 -576 -2015 -542
rect -1981 -576 -1969 -542
rect -2027 -610 -1969 -576
rect -2027 -644 -2015 -610
rect -1981 -644 -1969 -610
rect -2027 -678 -1969 -644
rect -2027 -712 -2015 -678
rect -1981 -712 -1969 -678
rect -2027 -746 -1969 -712
rect -2027 -780 -2015 -746
rect -1981 -780 -1969 -746
rect -2027 -814 -1969 -780
rect -2027 -848 -2015 -814
rect -1981 -848 -1969 -814
rect -2027 -882 -1969 -848
rect -2027 -916 -2015 -882
rect -1981 -916 -1969 -882
rect -2027 -950 -1969 -916
rect -2027 -984 -2015 -950
rect -1981 -984 -1969 -950
rect -2027 -1009 -1969 -984
rect -1879 -134 -1821 -109
rect -1879 -168 -1867 -134
rect -1833 -168 -1821 -134
rect -1879 -202 -1821 -168
rect -1879 -236 -1867 -202
rect -1833 -236 -1821 -202
rect -1879 -270 -1821 -236
rect -1879 -304 -1867 -270
rect -1833 -304 -1821 -270
rect -1879 -338 -1821 -304
rect -1879 -372 -1867 -338
rect -1833 -372 -1821 -338
rect -1879 -406 -1821 -372
rect -1879 -440 -1867 -406
rect -1833 -440 -1821 -406
rect -1879 -474 -1821 -440
rect -1879 -508 -1867 -474
rect -1833 -508 -1821 -474
rect -1879 -542 -1821 -508
rect -1879 -576 -1867 -542
rect -1833 -576 -1821 -542
rect -1879 -610 -1821 -576
rect -1879 -644 -1867 -610
rect -1833 -644 -1821 -610
rect -1879 -678 -1821 -644
rect -1879 -712 -1867 -678
rect -1833 -712 -1821 -678
rect -1879 -746 -1821 -712
rect -1879 -780 -1867 -746
rect -1833 -780 -1821 -746
rect -1879 -814 -1821 -780
rect -1879 -848 -1867 -814
rect -1833 -848 -1821 -814
rect -1879 -882 -1821 -848
rect -1879 -916 -1867 -882
rect -1833 -916 -1821 -882
rect -1879 -950 -1821 -916
rect -1879 -984 -1867 -950
rect -1833 -984 -1821 -950
rect -1879 -1009 -1821 -984
rect -1731 -134 -1673 -109
rect -1731 -168 -1719 -134
rect -1685 -168 -1673 -134
rect -1731 -202 -1673 -168
rect -1731 -236 -1719 -202
rect -1685 -236 -1673 -202
rect -1731 -270 -1673 -236
rect -1731 -304 -1719 -270
rect -1685 -304 -1673 -270
rect -1731 -338 -1673 -304
rect -1731 -372 -1719 -338
rect -1685 -372 -1673 -338
rect -1731 -406 -1673 -372
rect -1731 -440 -1719 -406
rect -1685 -440 -1673 -406
rect -1731 -474 -1673 -440
rect -1731 -508 -1719 -474
rect -1685 -508 -1673 -474
rect -1731 -542 -1673 -508
rect -1731 -576 -1719 -542
rect -1685 -576 -1673 -542
rect -1731 -610 -1673 -576
rect -1731 -644 -1719 -610
rect -1685 -644 -1673 -610
rect -1731 -678 -1673 -644
rect -1731 -712 -1719 -678
rect -1685 -712 -1673 -678
rect -1731 -746 -1673 -712
rect -1731 -780 -1719 -746
rect -1685 -780 -1673 -746
rect -1731 -814 -1673 -780
rect -1731 -848 -1719 -814
rect -1685 -848 -1673 -814
rect -1731 -882 -1673 -848
rect -1731 -916 -1719 -882
rect -1685 -916 -1673 -882
rect -1731 -950 -1673 -916
rect -1731 -984 -1719 -950
rect -1685 -984 -1673 -950
rect -1731 -1009 -1673 -984
rect -1583 -134 -1525 -109
rect -1583 -168 -1571 -134
rect -1537 -168 -1525 -134
rect -1583 -202 -1525 -168
rect -1583 -236 -1571 -202
rect -1537 -236 -1525 -202
rect -1583 -270 -1525 -236
rect -1583 -304 -1571 -270
rect -1537 -304 -1525 -270
rect -1583 -338 -1525 -304
rect -1583 -372 -1571 -338
rect -1537 -372 -1525 -338
rect -1583 -406 -1525 -372
rect -1583 -440 -1571 -406
rect -1537 -440 -1525 -406
rect -1583 -474 -1525 -440
rect -1583 -508 -1571 -474
rect -1537 -508 -1525 -474
rect -1583 -542 -1525 -508
rect -1583 -576 -1571 -542
rect -1537 -576 -1525 -542
rect -1583 -610 -1525 -576
rect -1583 -644 -1571 -610
rect -1537 -644 -1525 -610
rect -1583 -678 -1525 -644
rect -1583 -712 -1571 -678
rect -1537 -712 -1525 -678
rect -1583 -746 -1525 -712
rect -1583 -780 -1571 -746
rect -1537 -780 -1525 -746
rect -1583 -814 -1525 -780
rect -1583 -848 -1571 -814
rect -1537 -848 -1525 -814
rect -1583 -882 -1525 -848
rect -1583 -916 -1571 -882
rect -1537 -916 -1525 -882
rect -1583 -950 -1525 -916
rect -1583 -984 -1571 -950
rect -1537 -984 -1525 -950
rect -1583 -1009 -1525 -984
rect -1435 -134 -1377 -109
rect -1435 -168 -1423 -134
rect -1389 -168 -1377 -134
rect -1435 -202 -1377 -168
rect -1435 -236 -1423 -202
rect -1389 -236 -1377 -202
rect -1435 -270 -1377 -236
rect -1435 -304 -1423 -270
rect -1389 -304 -1377 -270
rect -1435 -338 -1377 -304
rect -1435 -372 -1423 -338
rect -1389 -372 -1377 -338
rect -1435 -406 -1377 -372
rect -1435 -440 -1423 -406
rect -1389 -440 -1377 -406
rect -1435 -474 -1377 -440
rect -1435 -508 -1423 -474
rect -1389 -508 -1377 -474
rect -1435 -542 -1377 -508
rect -1435 -576 -1423 -542
rect -1389 -576 -1377 -542
rect -1435 -610 -1377 -576
rect -1435 -644 -1423 -610
rect -1389 -644 -1377 -610
rect -1435 -678 -1377 -644
rect -1435 -712 -1423 -678
rect -1389 -712 -1377 -678
rect -1435 -746 -1377 -712
rect -1435 -780 -1423 -746
rect -1389 -780 -1377 -746
rect -1435 -814 -1377 -780
rect -1435 -848 -1423 -814
rect -1389 -848 -1377 -814
rect -1435 -882 -1377 -848
rect -1435 -916 -1423 -882
rect -1389 -916 -1377 -882
rect -1435 -950 -1377 -916
rect -1435 -984 -1423 -950
rect -1389 -984 -1377 -950
rect -1435 -1009 -1377 -984
rect -1287 -134 -1229 -109
rect -1287 -168 -1275 -134
rect -1241 -168 -1229 -134
rect -1287 -202 -1229 -168
rect -1287 -236 -1275 -202
rect -1241 -236 -1229 -202
rect -1287 -270 -1229 -236
rect -1287 -304 -1275 -270
rect -1241 -304 -1229 -270
rect -1287 -338 -1229 -304
rect -1287 -372 -1275 -338
rect -1241 -372 -1229 -338
rect -1287 -406 -1229 -372
rect -1287 -440 -1275 -406
rect -1241 -440 -1229 -406
rect -1287 -474 -1229 -440
rect -1287 -508 -1275 -474
rect -1241 -508 -1229 -474
rect -1287 -542 -1229 -508
rect -1287 -576 -1275 -542
rect -1241 -576 -1229 -542
rect -1287 -610 -1229 -576
rect -1287 -644 -1275 -610
rect -1241 -644 -1229 -610
rect -1287 -678 -1229 -644
rect -1287 -712 -1275 -678
rect -1241 -712 -1229 -678
rect -1287 -746 -1229 -712
rect -1287 -780 -1275 -746
rect -1241 -780 -1229 -746
rect -1287 -814 -1229 -780
rect -1287 -848 -1275 -814
rect -1241 -848 -1229 -814
rect -1287 -882 -1229 -848
rect -1287 -916 -1275 -882
rect -1241 -916 -1229 -882
rect -1287 -950 -1229 -916
rect -1287 -984 -1275 -950
rect -1241 -984 -1229 -950
rect -1287 -1009 -1229 -984
rect -1139 -134 -1081 -109
rect -1139 -168 -1127 -134
rect -1093 -168 -1081 -134
rect -1139 -202 -1081 -168
rect -1139 -236 -1127 -202
rect -1093 -236 -1081 -202
rect -1139 -270 -1081 -236
rect -1139 -304 -1127 -270
rect -1093 -304 -1081 -270
rect -1139 -338 -1081 -304
rect -1139 -372 -1127 -338
rect -1093 -372 -1081 -338
rect -1139 -406 -1081 -372
rect -1139 -440 -1127 -406
rect -1093 -440 -1081 -406
rect -1139 -474 -1081 -440
rect -1139 -508 -1127 -474
rect -1093 -508 -1081 -474
rect -1139 -542 -1081 -508
rect -1139 -576 -1127 -542
rect -1093 -576 -1081 -542
rect -1139 -610 -1081 -576
rect -1139 -644 -1127 -610
rect -1093 -644 -1081 -610
rect -1139 -678 -1081 -644
rect -1139 -712 -1127 -678
rect -1093 -712 -1081 -678
rect -1139 -746 -1081 -712
rect -1139 -780 -1127 -746
rect -1093 -780 -1081 -746
rect -1139 -814 -1081 -780
rect -1139 -848 -1127 -814
rect -1093 -848 -1081 -814
rect -1139 -882 -1081 -848
rect -1139 -916 -1127 -882
rect -1093 -916 -1081 -882
rect -1139 -950 -1081 -916
rect -1139 -984 -1127 -950
rect -1093 -984 -1081 -950
rect -1139 -1009 -1081 -984
rect -991 -134 -933 -109
rect -991 -168 -979 -134
rect -945 -168 -933 -134
rect -991 -202 -933 -168
rect -991 -236 -979 -202
rect -945 -236 -933 -202
rect -991 -270 -933 -236
rect -991 -304 -979 -270
rect -945 -304 -933 -270
rect -991 -338 -933 -304
rect -991 -372 -979 -338
rect -945 -372 -933 -338
rect -991 -406 -933 -372
rect -991 -440 -979 -406
rect -945 -440 -933 -406
rect -991 -474 -933 -440
rect -991 -508 -979 -474
rect -945 -508 -933 -474
rect -991 -542 -933 -508
rect -991 -576 -979 -542
rect -945 -576 -933 -542
rect -991 -610 -933 -576
rect -991 -644 -979 -610
rect -945 -644 -933 -610
rect -991 -678 -933 -644
rect -991 -712 -979 -678
rect -945 -712 -933 -678
rect -991 -746 -933 -712
rect -991 -780 -979 -746
rect -945 -780 -933 -746
rect -991 -814 -933 -780
rect -991 -848 -979 -814
rect -945 -848 -933 -814
rect -991 -882 -933 -848
rect -991 -916 -979 -882
rect -945 -916 -933 -882
rect -991 -950 -933 -916
rect -991 -984 -979 -950
rect -945 -984 -933 -950
rect -991 -1009 -933 -984
rect -843 -134 -785 -109
rect -843 -168 -831 -134
rect -797 -168 -785 -134
rect -843 -202 -785 -168
rect -843 -236 -831 -202
rect -797 -236 -785 -202
rect -843 -270 -785 -236
rect -843 -304 -831 -270
rect -797 -304 -785 -270
rect -843 -338 -785 -304
rect -843 -372 -831 -338
rect -797 -372 -785 -338
rect -843 -406 -785 -372
rect -843 -440 -831 -406
rect -797 -440 -785 -406
rect -843 -474 -785 -440
rect -843 -508 -831 -474
rect -797 -508 -785 -474
rect -843 -542 -785 -508
rect -843 -576 -831 -542
rect -797 -576 -785 -542
rect -843 -610 -785 -576
rect -843 -644 -831 -610
rect -797 -644 -785 -610
rect -843 -678 -785 -644
rect -843 -712 -831 -678
rect -797 -712 -785 -678
rect -843 -746 -785 -712
rect -843 -780 -831 -746
rect -797 -780 -785 -746
rect -843 -814 -785 -780
rect -843 -848 -831 -814
rect -797 -848 -785 -814
rect -843 -882 -785 -848
rect -843 -916 -831 -882
rect -797 -916 -785 -882
rect -843 -950 -785 -916
rect -843 -984 -831 -950
rect -797 -984 -785 -950
rect -843 -1009 -785 -984
rect -695 -134 -637 -109
rect -695 -168 -683 -134
rect -649 -168 -637 -134
rect -695 -202 -637 -168
rect -695 -236 -683 -202
rect -649 -236 -637 -202
rect -695 -270 -637 -236
rect -695 -304 -683 -270
rect -649 -304 -637 -270
rect -695 -338 -637 -304
rect -695 -372 -683 -338
rect -649 -372 -637 -338
rect -695 -406 -637 -372
rect -695 -440 -683 -406
rect -649 -440 -637 -406
rect -695 -474 -637 -440
rect -695 -508 -683 -474
rect -649 -508 -637 -474
rect -695 -542 -637 -508
rect -695 -576 -683 -542
rect -649 -576 -637 -542
rect -695 -610 -637 -576
rect -695 -644 -683 -610
rect -649 -644 -637 -610
rect -695 -678 -637 -644
rect -695 -712 -683 -678
rect -649 -712 -637 -678
rect -695 -746 -637 -712
rect -695 -780 -683 -746
rect -649 -780 -637 -746
rect -695 -814 -637 -780
rect -695 -848 -683 -814
rect -649 -848 -637 -814
rect -695 -882 -637 -848
rect -695 -916 -683 -882
rect -649 -916 -637 -882
rect -695 -950 -637 -916
rect -695 -984 -683 -950
rect -649 -984 -637 -950
rect -695 -1009 -637 -984
rect -547 -134 -489 -109
rect -547 -168 -535 -134
rect -501 -168 -489 -134
rect -547 -202 -489 -168
rect -547 -236 -535 -202
rect -501 -236 -489 -202
rect -547 -270 -489 -236
rect -547 -304 -535 -270
rect -501 -304 -489 -270
rect -547 -338 -489 -304
rect -547 -372 -535 -338
rect -501 -372 -489 -338
rect -547 -406 -489 -372
rect -547 -440 -535 -406
rect -501 -440 -489 -406
rect -547 -474 -489 -440
rect -547 -508 -535 -474
rect -501 -508 -489 -474
rect -547 -542 -489 -508
rect -547 -576 -535 -542
rect -501 -576 -489 -542
rect -547 -610 -489 -576
rect -547 -644 -535 -610
rect -501 -644 -489 -610
rect -547 -678 -489 -644
rect -547 -712 -535 -678
rect -501 -712 -489 -678
rect -547 -746 -489 -712
rect -547 -780 -535 -746
rect -501 -780 -489 -746
rect -547 -814 -489 -780
rect -547 -848 -535 -814
rect -501 -848 -489 -814
rect -547 -882 -489 -848
rect -547 -916 -535 -882
rect -501 -916 -489 -882
rect -547 -950 -489 -916
rect -547 -984 -535 -950
rect -501 -984 -489 -950
rect -547 -1009 -489 -984
rect -399 -134 -341 -109
rect -399 -168 -387 -134
rect -353 -168 -341 -134
rect -399 -202 -341 -168
rect -399 -236 -387 -202
rect -353 -236 -341 -202
rect -399 -270 -341 -236
rect -399 -304 -387 -270
rect -353 -304 -341 -270
rect -399 -338 -341 -304
rect -399 -372 -387 -338
rect -353 -372 -341 -338
rect -399 -406 -341 -372
rect -399 -440 -387 -406
rect -353 -440 -341 -406
rect -399 -474 -341 -440
rect -399 -508 -387 -474
rect -353 -508 -341 -474
rect -399 -542 -341 -508
rect -399 -576 -387 -542
rect -353 -576 -341 -542
rect -399 -610 -341 -576
rect -399 -644 -387 -610
rect -353 -644 -341 -610
rect -399 -678 -341 -644
rect -399 -712 -387 -678
rect -353 -712 -341 -678
rect -399 -746 -341 -712
rect -399 -780 -387 -746
rect -353 -780 -341 -746
rect -399 -814 -341 -780
rect -399 -848 -387 -814
rect -353 -848 -341 -814
rect -399 -882 -341 -848
rect -399 -916 -387 -882
rect -353 -916 -341 -882
rect -399 -950 -341 -916
rect -399 -984 -387 -950
rect -353 -984 -341 -950
rect -399 -1009 -341 -984
rect -251 -134 -193 -109
rect -251 -168 -239 -134
rect -205 -168 -193 -134
rect -251 -202 -193 -168
rect -251 -236 -239 -202
rect -205 -236 -193 -202
rect -251 -270 -193 -236
rect -251 -304 -239 -270
rect -205 -304 -193 -270
rect -251 -338 -193 -304
rect -251 -372 -239 -338
rect -205 -372 -193 -338
rect -251 -406 -193 -372
rect -251 -440 -239 -406
rect -205 -440 -193 -406
rect -251 -474 -193 -440
rect -251 -508 -239 -474
rect -205 -508 -193 -474
rect -251 -542 -193 -508
rect -251 -576 -239 -542
rect -205 -576 -193 -542
rect -251 -610 -193 -576
rect -251 -644 -239 -610
rect -205 -644 -193 -610
rect -251 -678 -193 -644
rect -251 -712 -239 -678
rect -205 -712 -193 -678
rect -251 -746 -193 -712
rect -251 -780 -239 -746
rect -205 -780 -193 -746
rect -251 -814 -193 -780
rect -251 -848 -239 -814
rect -205 -848 -193 -814
rect -251 -882 -193 -848
rect -251 -916 -239 -882
rect -205 -916 -193 -882
rect -251 -950 -193 -916
rect -251 -984 -239 -950
rect -205 -984 -193 -950
rect -251 -1009 -193 -984
rect -103 -134 -45 -109
rect -103 -168 -91 -134
rect -57 -168 -45 -134
rect -103 -202 -45 -168
rect -103 -236 -91 -202
rect -57 -236 -45 -202
rect -103 -270 -45 -236
rect -103 -304 -91 -270
rect -57 -304 -45 -270
rect -103 -338 -45 -304
rect -103 -372 -91 -338
rect -57 -372 -45 -338
rect -103 -406 -45 -372
rect -103 -440 -91 -406
rect -57 -440 -45 -406
rect -103 -474 -45 -440
rect -103 -508 -91 -474
rect -57 -508 -45 -474
rect -103 -542 -45 -508
rect -103 -576 -91 -542
rect -57 -576 -45 -542
rect -103 -610 -45 -576
rect -103 -644 -91 -610
rect -57 -644 -45 -610
rect -103 -678 -45 -644
rect -103 -712 -91 -678
rect -57 -712 -45 -678
rect -103 -746 -45 -712
rect -103 -780 -91 -746
rect -57 -780 -45 -746
rect -103 -814 -45 -780
rect -103 -848 -91 -814
rect -57 -848 -45 -814
rect -103 -882 -45 -848
rect -103 -916 -91 -882
rect -57 -916 -45 -882
rect -103 -950 -45 -916
rect -103 -984 -91 -950
rect -57 -984 -45 -950
rect -103 -1009 -45 -984
rect 45 -134 103 -109
rect 45 -168 57 -134
rect 91 -168 103 -134
rect 45 -202 103 -168
rect 45 -236 57 -202
rect 91 -236 103 -202
rect 45 -270 103 -236
rect 45 -304 57 -270
rect 91 -304 103 -270
rect 45 -338 103 -304
rect 45 -372 57 -338
rect 91 -372 103 -338
rect 45 -406 103 -372
rect 45 -440 57 -406
rect 91 -440 103 -406
rect 45 -474 103 -440
rect 45 -508 57 -474
rect 91 -508 103 -474
rect 45 -542 103 -508
rect 45 -576 57 -542
rect 91 -576 103 -542
rect 45 -610 103 -576
rect 45 -644 57 -610
rect 91 -644 103 -610
rect 45 -678 103 -644
rect 45 -712 57 -678
rect 91 -712 103 -678
rect 45 -746 103 -712
rect 45 -780 57 -746
rect 91 -780 103 -746
rect 45 -814 103 -780
rect 45 -848 57 -814
rect 91 -848 103 -814
rect 45 -882 103 -848
rect 45 -916 57 -882
rect 91 -916 103 -882
rect 45 -950 103 -916
rect 45 -984 57 -950
rect 91 -984 103 -950
rect 45 -1009 103 -984
rect 193 -134 251 -109
rect 193 -168 205 -134
rect 239 -168 251 -134
rect 193 -202 251 -168
rect 193 -236 205 -202
rect 239 -236 251 -202
rect 193 -270 251 -236
rect 193 -304 205 -270
rect 239 -304 251 -270
rect 193 -338 251 -304
rect 193 -372 205 -338
rect 239 -372 251 -338
rect 193 -406 251 -372
rect 193 -440 205 -406
rect 239 -440 251 -406
rect 193 -474 251 -440
rect 193 -508 205 -474
rect 239 -508 251 -474
rect 193 -542 251 -508
rect 193 -576 205 -542
rect 239 -576 251 -542
rect 193 -610 251 -576
rect 193 -644 205 -610
rect 239 -644 251 -610
rect 193 -678 251 -644
rect 193 -712 205 -678
rect 239 -712 251 -678
rect 193 -746 251 -712
rect 193 -780 205 -746
rect 239 -780 251 -746
rect 193 -814 251 -780
rect 193 -848 205 -814
rect 239 -848 251 -814
rect 193 -882 251 -848
rect 193 -916 205 -882
rect 239 -916 251 -882
rect 193 -950 251 -916
rect 193 -984 205 -950
rect 239 -984 251 -950
rect 193 -1009 251 -984
rect 341 -134 399 -109
rect 341 -168 353 -134
rect 387 -168 399 -134
rect 341 -202 399 -168
rect 341 -236 353 -202
rect 387 -236 399 -202
rect 341 -270 399 -236
rect 341 -304 353 -270
rect 387 -304 399 -270
rect 341 -338 399 -304
rect 341 -372 353 -338
rect 387 -372 399 -338
rect 341 -406 399 -372
rect 341 -440 353 -406
rect 387 -440 399 -406
rect 341 -474 399 -440
rect 341 -508 353 -474
rect 387 -508 399 -474
rect 341 -542 399 -508
rect 341 -576 353 -542
rect 387 -576 399 -542
rect 341 -610 399 -576
rect 341 -644 353 -610
rect 387 -644 399 -610
rect 341 -678 399 -644
rect 341 -712 353 -678
rect 387 -712 399 -678
rect 341 -746 399 -712
rect 341 -780 353 -746
rect 387 -780 399 -746
rect 341 -814 399 -780
rect 341 -848 353 -814
rect 387 -848 399 -814
rect 341 -882 399 -848
rect 341 -916 353 -882
rect 387 -916 399 -882
rect 341 -950 399 -916
rect 341 -984 353 -950
rect 387 -984 399 -950
rect 341 -1009 399 -984
rect 489 -134 547 -109
rect 489 -168 501 -134
rect 535 -168 547 -134
rect 489 -202 547 -168
rect 489 -236 501 -202
rect 535 -236 547 -202
rect 489 -270 547 -236
rect 489 -304 501 -270
rect 535 -304 547 -270
rect 489 -338 547 -304
rect 489 -372 501 -338
rect 535 -372 547 -338
rect 489 -406 547 -372
rect 489 -440 501 -406
rect 535 -440 547 -406
rect 489 -474 547 -440
rect 489 -508 501 -474
rect 535 -508 547 -474
rect 489 -542 547 -508
rect 489 -576 501 -542
rect 535 -576 547 -542
rect 489 -610 547 -576
rect 489 -644 501 -610
rect 535 -644 547 -610
rect 489 -678 547 -644
rect 489 -712 501 -678
rect 535 -712 547 -678
rect 489 -746 547 -712
rect 489 -780 501 -746
rect 535 -780 547 -746
rect 489 -814 547 -780
rect 489 -848 501 -814
rect 535 -848 547 -814
rect 489 -882 547 -848
rect 489 -916 501 -882
rect 535 -916 547 -882
rect 489 -950 547 -916
rect 489 -984 501 -950
rect 535 -984 547 -950
rect 489 -1009 547 -984
rect 637 -134 695 -109
rect 637 -168 649 -134
rect 683 -168 695 -134
rect 637 -202 695 -168
rect 637 -236 649 -202
rect 683 -236 695 -202
rect 637 -270 695 -236
rect 637 -304 649 -270
rect 683 -304 695 -270
rect 637 -338 695 -304
rect 637 -372 649 -338
rect 683 -372 695 -338
rect 637 -406 695 -372
rect 637 -440 649 -406
rect 683 -440 695 -406
rect 637 -474 695 -440
rect 637 -508 649 -474
rect 683 -508 695 -474
rect 637 -542 695 -508
rect 637 -576 649 -542
rect 683 -576 695 -542
rect 637 -610 695 -576
rect 637 -644 649 -610
rect 683 -644 695 -610
rect 637 -678 695 -644
rect 637 -712 649 -678
rect 683 -712 695 -678
rect 637 -746 695 -712
rect 637 -780 649 -746
rect 683 -780 695 -746
rect 637 -814 695 -780
rect 637 -848 649 -814
rect 683 -848 695 -814
rect 637 -882 695 -848
rect 637 -916 649 -882
rect 683 -916 695 -882
rect 637 -950 695 -916
rect 637 -984 649 -950
rect 683 -984 695 -950
rect 637 -1009 695 -984
rect 785 -134 843 -109
rect 785 -168 797 -134
rect 831 -168 843 -134
rect 785 -202 843 -168
rect 785 -236 797 -202
rect 831 -236 843 -202
rect 785 -270 843 -236
rect 785 -304 797 -270
rect 831 -304 843 -270
rect 785 -338 843 -304
rect 785 -372 797 -338
rect 831 -372 843 -338
rect 785 -406 843 -372
rect 785 -440 797 -406
rect 831 -440 843 -406
rect 785 -474 843 -440
rect 785 -508 797 -474
rect 831 -508 843 -474
rect 785 -542 843 -508
rect 785 -576 797 -542
rect 831 -576 843 -542
rect 785 -610 843 -576
rect 785 -644 797 -610
rect 831 -644 843 -610
rect 785 -678 843 -644
rect 785 -712 797 -678
rect 831 -712 843 -678
rect 785 -746 843 -712
rect 785 -780 797 -746
rect 831 -780 843 -746
rect 785 -814 843 -780
rect 785 -848 797 -814
rect 831 -848 843 -814
rect 785 -882 843 -848
rect 785 -916 797 -882
rect 831 -916 843 -882
rect 785 -950 843 -916
rect 785 -984 797 -950
rect 831 -984 843 -950
rect 785 -1009 843 -984
rect 933 -134 991 -109
rect 933 -168 945 -134
rect 979 -168 991 -134
rect 933 -202 991 -168
rect 933 -236 945 -202
rect 979 -236 991 -202
rect 933 -270 991 -236
rect 933 -304 945 -270
rect 979 -304 991 -270
rect 933 -338 991 -304
rect 933 -372 945 -338
rect 979 -372 991 -338
rect 933 -406 991 -372
rect 933 -440 945 -406
rect 979 -440 991 -406
rect 933 -474 991 -440
rect 933 -508 945 -474
rect 979 -508 991 -474
rect 933 -542 991 -508
rect 933 -576 945 -542
rect 979 -576 991 -542
rect 933 -610 991 -576
rect 933 -644 945 -610
rect 979 -644 991 -610
rect 933 -678 991 -644
rect 933 -712 945 -678
rect 979 -712 991 -678
rect 933 -746 991 -712
rect 933 -780 945 -746
rect 979 -780 991 -746
rect 933 -814 991 -780
rect 933 -848 945 -814
rect 979 -848 991 -814
rect 933 -882 991 -848
rect 933 -916 945 -882
rect 979 -916 991 -882
rect 933 -950 991 -916
rect 933 -984 945 -950
rect 979 -984 991 -950
rect 933 -1009 991 -984
rect 1081 -134 1139 -109
rect 1081 -168 1093 -134
rect 1127 -168 1139 -134
rect 1081 -202 1139 -168
rect 1081 -236 1093 -202
rect 1127 -236 1139 -202
rect 1081 -270 1139 -236
rect 1081 -304 1093 -270
rect 1127 -304 1139 -270
rect 1081 -338 1139 -304
rect 1081 -372 1093 -338
rect 1127 -372 1139 -338
rect 1081 -406 1139 -372
rect 1081 -440 1093 -406
rect 1127 -440 1139 -406
rect 1081 -474 1139 -440
rect 1081 -508 1093 -474
rect 1127 -508 1139 -474
rect 1081 -542 1139 -508
rect 1081 -576 1093 -542
rect 1127 -576 1139 -542
rect 1081 -610 1139 -576
rect 1081 -644 1093 -610
rect 1127 -644 1139 -610
rect 1081 -678 1139 -644
rect 1081 -712 1093 -678
rect 1127 -712 1139 -678
rect 1081 -746 1139 -712
rect 1081 -780 1093 -746
rect 1127 -780 1139 -746
rect 1081 -814 1139 -780
rect 1081 -848 1093 -814
rect 1127 -848 1139 -814
rect 1081 -882 1139 -848
rect 1081 -916 1093 -882
rect 1127 -916 1139 -882
rect 1081 -950 1139 -916
rect 1081 -984 1093 -950
rect 1127 -984 1139 -950
rect 1081 -1009 1139 -984
rect 1229 -134 1287 -109
rect 1229 -168 1241 -134
rect 1275 -168 1287 -134
rect 1229 -202 1287 -168
rect 1229 -236 1241 -202
rect 1275 -236 1287 -202
rect 1229 -270 1287 -236
rect 1229 -304 1241 -270
rect 1275 -304 1287 -270
rect 1229 -338 1287 -304
rect 1229 -372 1241 -338
rect 1275 -372 1287 -338
rect 1229 -406 1287 -372
rect 1229 -440 1241 -406
rect 1275 -440 1287 -406
rect 1229 -474 1287 -440
rect 1229 -508 1241 -474
rect 1275 -508 1287 -474
rect 1229 -542 1287 -508
rect 1229 -576 1241 -542
rect 1275 -576 1287 -542
rect 1229 -610 1287 -576
rect 1229 -644 1241 -610
rect 1275 -644 1287 -610
rect 1229 -678 1287 -644
rect 1229 -712 1241 -678
rect 1275 -712 1287 -678
rect 1229 -746 1287 -712
rect 1229 -780 1241 -746
rect 1275 -780 1287 -746
rect 1229 -814 1287 -780
rect 1229 -848 1241 -814
rect 1275 -848 1287 -814
rect 1229 -882 1287 -848
rect 1229 -916 1241 -882
rect 1275 -916 1287 -882
rect 1229 -950 1287 -916
rect 1229 -984 1241 -950
rect 1275 -984 1287 -950
rect 1229 -1009 1287 -984
rect 1377 -134 1435 -109
rect 1377 -168 1389 -134
rect 1423 -168 1435 -134
rect 1377 -202 1435 -168
rect 1377 -236 1389 -202
rect 1423 -236 1435 -202
rect 1377 -270 1435 -236
rect 1377 -304 1389 -270
rect 1423 -304 1435 -270
rect 1377 -338 1435 -304
rect 1377 -372 1389 -338
rect 1423 -372 1435 -338
rect 1377 -406 1435 -372
rect 1377 -440 1389 -406
rect 1423 -440 1435 -406
rect 1377 -474 1435 -440
rect 1377 -508 1389 -474
rect 1423 -508 1435 -474
rect 1377 -542 1435 -508
rect 1377 -576 1389 -542
rect 1423 -576 1435 -542
rect 1377 -610 1435 -576
rect 1377 -644 1389 -610
rect 1423 -644 1435 -610
rect 1377 -678 1435 -644
rect 1377 -712 1389 -678
rect 1423 -712 1435 -678
rect 1377 -746 1435 -712
rect 1377 -780 1389 -746
rect 1423 -780 1435 -746
rect 1377 -814 1435 -780
rect 1377 -848 1389 -814
rect 1423 -848 1435 -814
rect 1377 -882 1435 -848
rect 1377 -916 1389 -882
rect 1423 -916 1435 -882
rect 1377 -950 1435 -916
rect 1377 -984 1389 -950
rect 1423 -984 1435 -950
rect 1377 -1009 1435 -984
rect 1525 -134 1583 -109
rect 1525 -168 1537 -134
rect 1571 -168 1583 -134
rect 1525 -202 1583 -168
rect 1525 -236 1537 -202
rect 1571 -236 1583 -202
rect 1525 -270 1583 -236
rect 1525 -304 1537 -270
rect 1571 -304 1583 -270
rect 1525 -338 1583 -304
rect 1525 -372 1537 -338
rect 1571 -372 1583 -338
rect 1525 -406 1583 -372
rect 1525 -440 1537 -406
rect 1571 -440 1583 -406
rect 1525 -474 1583 -440
rect 1525 -508 1537 -474
rect 1571 -508 1583 -474
rect 1525 -542 1583 -508
rect 1525 -576 1537 -542
rect 1571 -576 1583 -542
rect 1525 -610 1583 -576
rect 1525 -644 1537 -610
rect 1571 -644 1583 -610
rect 1525 -678 1583 -644
rect 1525 -712 1537 -678
rect 1571 -712 1583 -678
rect 1525 -746 1583 -712
rect 1525 -780 1537 -746
rect 1571 -780 1583 -746
rect 1525 -814 1583 -780
rect 1525 -848 1537 -814
rect 1571 -848 1583 -814
rect 1525 -882 1583 -848
rect 1525 -916 1537 -882
rect 1571 -916 1583 -882
rect 1525 -950 1583 -916
rect 1525 -984 1537 -950
rect 1571 -984 1583 -950
rect 1525 -1009 1583 -984
rect 1673 -134 1731 -109
rect 1673 -168 1685 -134
rect 1719 -168 1731 -134
rect 1673 -202 1731 -168
rect 1673 -236 1685 -202
rect 1719 -236 1731 -202
rect 1673 -270 1731 -236
rect 1673 -304 1685 -270
rect 1719 -304 1731 -270
rect 1673 -338 1731 -304
rect 1673 -372 1685 -338
rect 1719 -372 1731 -338
rect 1673 -406 1731 -372
rect 1673 -440 1685 -406
rect 1719 -440 1731 -406
rect 1673 -474 1731 -440
rect 1673 -508 1685 -474
rect 1719 -508 1731 -474
rect 1673 -542 1731 -508
rect 1673 -576 1685 -542
rect 1719 -576 1731 -542
rect 1673 -610 1731 -576
rect 1673 -644 1685 -610
rect 1719 -644 1731 -610
rect 1673 -678 1731 -644
rect 1673 -712 1685 -678
rect 1719 -712 1731 -678
rect 1673 -746 1731 -712
rect 1673 -780 1685 -746
rect 1719 -780 1731 -746
rect 1673 -814 1731 -780
rect 1673 -848 1685 -814
rect 1719 -848 1731 -814
rect 1673 -882 1731 -848
rect 1673 -916 1685 -882
rect 1719 -916 1731 -882
rect 1673 -950 1731 -916
rect 1673 -984 1685 -950
rect 1719 -984 1731 -950
rect 1673 -1009 1731 -984
rect 1821 -134 1879 -109
rect 1821 -168 1833 -134
rect 1867 -168 1879 -134
rect 1821 -202 1879 -168
rect 1821 -236 1833 -202
rect 1867 -236 1879 -202
rect 1821 -270 1879 -236
rect 1821 -304 1833 -270
rect 1867 -304 1879 -270
rect 1821 -338 1879 -304
rect 1821 -372 1833 -338
rect 1867 -372 1879 -338
rect 1821 -406 1879 -372
rect 1821 -440 1833 -406
rect 1867 -440 1879 -406
rect 1821 -474 1879 -440
rect 1821 -508 1833 -474
rect 1867 -508 1879 -474
rect 1821 -542 1879 -508
rect 1821 -576 1833 -542
rect 1867 -576 1879 -542
rect 1821 -610 1879 -576
rect 1821 -644 1833 -610
rect 1867 -644 1879 -610
rect 1821 -678 1879 -644
rect 1821 -712 1833 -678
rect 1867 -712 1879 -678
rect 1821 -746 1879 -712
rect 1821 -780 1833 -746
rect 1867 -780 1879 -746
rect 1821 -814 1879 -780
rect 1821 -848 1833 -814
rect 1867 -848 1879 -814
rect 1821 -882 1879 -848
rect 1821 -916 1833 -882
rect 1867 -916 1879 -882
rect 1821 -950 1879 -916
rect 1821 -984 1833 -950
rect 1867 -984 1879 -950
rect 1821 -1009 1879 -984
rect 1969 -134 2027 -109
rect 1969 -168 1981 -134
rect 2015 -168 2027 -134
rect 1969 -202 2027 -168
rect 1969 -236 1981 -202
rect 2015 -236 2027 -202
rect 1969 -270 2027 -236
rect 1969 -304 1981 -270
rect 2015 -304 2027 -270
rect 1969 -338 2027 -304
rect 1969 -372 1981 -338
rect 2015 -372 2027 -338
rect 1969 -406 2027 -372
rect 1969 -440 1981 -406
rect 2015 -440 2027 -406
rect 1969 -474 2027 -440
rect 1969 -508 1981 -474
rect 2015 -508 2027 -474
rect 1969 -542 2027 -508
rect 1969 -576 1981 -542
rect 2015 -576 2027 -542
rect 1969 -610 2027 -576
rect 1969 -644 1981 -610
rect 2015 -644 2027 -610
rect 1969 -678 2027 -644
rect 1969 -712 1981 -678
rect 2015 -712 2027 -678
rect 1969 -746 2027 -712
rect 1969 -780 1981 -746
rect 2015 -780 2027 -746
rect 1969 -814 2027 -780
rect 1969 -848 1981 -814
rect 2015 -848 2027 -814
rect 1969 -882 2027 -848
rect 1969 -916 1981 -882
rect 2015 -916 2027 -882
rect 1969 -950 2027 -916
rect 1969 -984 1981 -950
rect 2015 -984 2027 -950
rect 1969 -1009 2027 -984
rect 2117 -134 2175 -109
rect 2117 -168 2129 -134
rect 2163 -168 2175 -134
rect 2117 -202 2175 -168
rect 2117 -236 2129 -202
rect 2163 -236 2175 -202
rect 2117 -270 2175 -236
rect 2117 -304 2129 -270
rect 2163 -304 2175 -270
rect 2117 -338 2175 -304
rect 2117 -372 2129 -338
rect 2163 -372 2175 -338
rect 2117 -406 2175 -372
rect 2117 -440 2129 -406
rect 2163 -440 2175 -406
rect 2117 -474 2175 -440
rect 2117 -508 2129 -474
rect 2163 -508 2175 -474
rect 2117 -542 2175 -508
rect 2117 -576 2129 -542
rect 2163 -576 2175 -542
rect 2117 -610 2175 -576
rect 2117 -644 2129 -610
rect 2163 -644 2175 -610
rect 2117 -678 2175 -644
rect 2117 -712 2129 -678
rect 2163 -712 2175 -678
rect 2117 -746 2175 -712
rect 2117 -780 2129 -746
rect 2163 -780 2175 -746
rect 2117 -814 2175 -780
rect 2117 -848 2129 -814
rect 2163 -848 2175 -814
rect 2117 -882 2175 -848
rect 2117 -916 2129 -882
rect 2163 -916 2175 -882
rect 2117 -950 2175 -916
rect 2117 -984 2129 -950
rect 2163 -984 2175 -950
rect 2117 -1009 2175 -984
rect 2265 -134 2323 -109
rect 2265 -168 2277 -134
rect 2311 -168 2323 -134
rect 2265 -202 2323 -168
rect 2265 -236 2277 -202
rect 2311 -236 2323 -202
rect 2265 -270 2323 -236
rect 2265 -304 2277 -270
rect 2311 -304 2323 -270
rect 2265 -338 2323 -304
rect 2265 -372 2277 -338
rect 2311 -372 2323 -338
rect 2265 -406 2323 -372
rect 2265 -440 2277 -406
rect 2311 -440 2323 -406
rect 2265 -474 2323 -440
rect 2265 -508 2277 -474
rect 2311 -508 2323 -474
rect 2265 -542 2323 -508
rect 2265 -576 2277 -542
rect 2311 -576 2323 -542
rect 2265 -610 2323 -576
rect 2265 -644 2277 -610
rect 2311 -644 2323 -610
rect 2265 -678 2323 -644
rect 2265 -712 2277 -678
rect 2311 -712 2323 -678
rect 2265 -746 2323 -712
rect 2265 -780 2277 -746
rect 2311 -780 2323 -746
rect 2265 -814 2323 -780
rect 2265 -848 2277 -814
rect 2311 -848 2323 -814
rect 2265 -882 2323 -848
rect 2265 -916 2277 -882
rect 2311 -916 2323 -882
rect 2265 -950 2323 -916
rect 2265 -984 2277 -950
rect 2311 -984 2323 -950
rect 2265 -1009 2323 -984
rect 2413 -134 2471 -109
rect 2413 -168 2425 -134
rect 2459 -168 2471 -134
rect 2413 -202 2471 -168
rect 2413 -236 2425 -202
rect 2459 -236 2471 -202
rect 2413 -270 2471 -236
rect 2413 -304 2425 -270
rect 2459 -304 2471 -270
rect 2413 -338 2471 -304
rect 2413 -372 2425 -338
rect 2459 -372 2471 -338
rect 2413 -406 2471 -372
rect 2413 -440 2425 -406
rect 2459 -440 2471 -406
rect 2413 -474 2471 -440
rect 2413 -508 2425 -474
rect 2459 -508 2471 -474
rect 2413 -542 2471 -508
rect 2413 -576 2425 -542
rect 2459 -576 2471 -542
rect 2413 -610 2471 -576
rect 2413 -644 2425 -610
rect 2459 -644 2471 -610
rect 2413 -678 2471 -644
rect 2413 -712 2425 -678
rect 2459 -712 2471 -678
rect 2413 -746 2471 -712
rect 2413 -780 2425 -746
rect 2459 -780 2471 -746
rect 2413 -814 2471 -780
rect 2413 -848 2425 -814
rect 2459 -848 2471 -814
rect 2413 -882 2471 -848
rect 2413 -916 2425 -882
rect 2459 -916 2471 -882
rect 2413 -950 2471 -916
rect 2413 -984 2425 -950
rect 2459 -984 2471 -950
rect 2413 -1009 2471 -984
rect 2561 -134 2619 -109
rect 2561 -168 2573 -134
rect 2607 -168 2619 -134
rect 2561 -202 2619 -168
rect 2561 -236 2573 -202
rect 2607 -236 2619 -202
rect 2561 -270 2619 -236
rect 2561 -304 2573 -270
rect 2607 -304 2619 -270
rect 2561 -338 2619 -304
rect 2561 -372 2573 -338
rect 2607 -372 2619 -338
rect 2561 -406 2619 -372
rect 2561 -440 2573 -406
rect 2607 -440 2619 -406
rect 2561 -474 2619 -440
rect 2561 -508 2573 -474
rect 2607 -508 2619 -474
rect 2561 -542 2619 -508
rect 2561 -576 2573 -542
rect 2607 -576 2619 -542
rect 2561 -610 2619 -576
rect 2561 -644 2573 -610
rect 2607 -644 2619 -610
rect 2561 -678 2619 -644
rect 2561 -712 2573 -678
rect 2607 -712 2619 -678
rect 2561 -746 2619 -712
rect 2561 -780 2573 -746
rect 2607 -780 2619 -746
rect 2561 -814 2619 -780
rect 2561 -848 2573 -814
rect 2607 -848 2619 -814
rect 2561 -882 2619 -848
rect 2561 -916 2573 -882
rect 2607 -916 2619 -882
rect 2561 -950 2619 -916
rect 2561 -984 2573 -950
rect 2607 -984 2619 -950
rect 2561 -1009 2619 -984
rect 2709 -134 2767 -109
rect 2709 -168 2721 -134
rect 2755 -168 2767 -134
rect 2709 -202 2767 -168
rect 2709 -236 2721 -202
rect 2755 -236 2767 -202
rect 2709 -270 2767 -236
rect 2709 -304 2721 -270
rect 2755 -304 2767 -270
rect 2709 -338 2767 -304
rect 2709 -372 2721 -338
rect 2755 -372 2767 -338
rect 2709 -406 2767 -372
rect 2709 -440 2721 -406
rect 2755 -440 2767 -406
rect 2709 -474 2767 -440
rect 2709 -508 2721 -474
rect 2755 -508 2767 -474
rect 2709 -542 2767 -508
rect 2709 -576 2721 -542
rect 2755 -576 2767 -542
rect 2709 -610 2767 -576
rect 2709 -644 2721 -610
rect 2755 -644 2767 -610
rect 2709 -678 2767 -644
rect 2709 -712 2721 -678
rect 2755 -712 2767 -678
rect 2709 -746 2767 -712
rect 2709 -780 2721 -746
rect 2755 -780 2767 -746
rect 2709 -814 2767 -780
rect 2709 -848 2721 -814
rect 2755 -848 2767 -814
rect 2709 -882 2767 -848
rect 2709 -916 2721 -882
rect 2755 -916 2767 -882
rect 2709 -950 2767 -916
rect 2709 -984 2721 -950
rect 2755 -984 2767 -950
rect 2709 -1009 2767 -984
rect 2857 -134 2915 -109
rect 2857 -168 2869 -134
rect 2903 -168 2915 -134
rect 2857 -202 2915 -168
rect 2857 -236 2869 -202
rect 2903 -236 2915 -202
rect 2857 -270 2915 -236
rect 2857 -304 2869 -270
rect 2903 -304 2915 -270
rect 2857 -338 2915 -304
rect 2857 -372 2869 -338
rect 2903 -372 2915 -338
rect 2857 -406 2915 -372
rect 2857 -440 2869 -406
rect 2903 -440 2915 -406
rect 2857 -474 2915 -440
rect 2857 -508 2869 -474
rect 2903 -508 2915 -474
rect 2857 -542 2915 -508
rect 2857 -576 2869 -542
rect 2903 -576 2915 -542
rect 2857 -610 2915 -576
rect 2857 -644 2869 -610
rect 2903 -644 2915 -610
rect 2857 -678 2915 -644
rect 2857 -712 2869 -678
rect 2903 -712 2915 -678
rect 2857 -746 2915 -712
rect 2857 -780 2869 -746
rect 2903 -780 2915 -746
rect 2857 -814 2915 -780
rect 2857 -848 2869 -814
rect 2903 -848 2915 -814
rect 2857 -882 2915 -848
rect 2857 -916 2869 -882
rect 2903 -916 2915 -882
rect 2857 -950 2915 -916
rect 2857 -984 2869 -950
rect 2903 -984 2915 -950
rect 2857 -1009 2915 -984
rect 3005 -134 3063 -109
rect 3005 -168 3017 -134
rect 3051 -168 3063 -134
rect 3005 -202 3063 -168
rect 3005 -236 3017 -202
rect 3051 -236 3063 -202
rect 3005 -270 3063 -236
rect 3005 -304 3017 -270
rect 3051 -304 3063 -270
rect 3005 -338 3063 -304
rect 3005 -372 3017 -338
rect 3051 -372 3063 -338
rect 3005 -406 3063 -372
rect 3005 -440 3017 -406
rect 3051 -440 3063 -406
rect 3005 -474 3063 -440
rect 3005 -508 3017 -474
rect 3051 -508 3063 -474
rect 3005 -542 3063 -508
rect 3005 -576 3017 -542
rect 3051 -576 3063 -542
rect 3005 -610 3063 -576
rect 3005 -644 3017 -610
rect 3051 -644 3063 -610
rect 3005 -678 3063 -644
rect 3005 -712 3017 -678
rect 3051 -712 3063 -678
rect 3005 -746 3063 -712
rect 3005 -780 3017 -746
rect 3051 -780 3063 -746
rect 3005 -814 3063 -780
rect 3005 -848 3017 -814
rect 3051 -848 3063 -814
rect 3005 -882 3063 -848
rect 3005 -916 3017 -882
rect 3051 -916 3063 -882
rect 3005 -950 3063 -916
rect 3005 -984 3017 -950
rect 3051 -984 3063 -950
rect 3005 -1009 3063 -984
rect 3153 -134 3211 -109
rect 3153 -168 3165 -134
rect 3199 -168 3211 -134
rect 3153 -202 3211 -168
rect 3153 -236 3165 -202
rect 3199 -236 3211 -202
rect 3153 -270 3211 -236
rect 3153 -304 3165 -270
rect 3199 -304 3211 -270
rect 3153 -338 3211 -304
rect 3153 -372 3165 -338
rect 3199 -372 3211 -338
rect 3153 -406 3211 -372
rect 3153 -440 3165 -406
rect 3199 -440 3211 -406
rect 3153 -474 3211 -440
rect 3153 -508 3165 -474
rect 3199 -508 3211 -474
rect 3153 -542 3211 -508
rect 3153 -576 3165 -542
rect 3199 -576 3211 -542
rect 3153 -610 3211 -576
rect 3153 -644 3165 -610
rect 3199 -644 3211 -610
rect 3153 -678 3211 -644
rect 3153 -712 3165 -678
rect 3199 -712 3211 -678
rect 3153 -746 3211 -712
rect 3153 -780 3165 -746
rect 3199 -780 3211 -746
rect 3153 -814 3211 -780
rect 3153 -848 3165 -814
rect 3199 -848 3211 -814
rect 3153 -882 3211 -848
rect 3153 -916 3165 -882
rect 3199 -916 3211 -882
rect 3153 -950 3211 -916
rect 3153 -984 3165 -950
rect 3199 -984 3211 -950
rect 3153 -1009 3211 -984
rect 3301 -134 3359 -109
rect 3301 -168 3313 -134
rect 3347 -168 3359 -134
rect 3301 -202 3359 -168
rect 3301 -236 3313 -202
rect 3347 -236 3359 -202
rect 3301 -270 3359 -236
rect 3301 -304 3313 -270
rect 3347 -304 3359 -270
rect 3301 -338 3359 -304
rect 3301 -372 3313 -338
rect 3347 -372 3359 -338
rect 3301 -406 3359 -372
rect 3301 -440 3313 -406
rect 3347 -440 3359 -406
rect 3301 -474 3359 -440
rect 3301 -508 3313 -474
rect 3347 -508 3359 -474
rect 3301 -542 3359 -508
rect 3301 -576 3313 -542
rect 3347 -576 3359 -542
rect 3301 -610 3359 -576
rect 3301 -644 3313 -610
rect 3347 -644 3359 -610
rect 3301 -678 3359 -644
rect 3301 -712 3313 -678
rect 3347 -712 3359 -678
rect 3301 -746 3359 -712
rect 3301 -780 3313 -746
rect 3347 -780 3359 -746
rect 3301 -814 3359 -780
rect 3301 -848 3313 -814
rect 3347 -848 3359 -814
rect 3301 -882 3359 -848
rect 3301 -916 3313 -882
rect 3347 -916 3359 -882
rect 3301 -950 3359 -916
rect 3301 -984 3313 -950
rect 3347 -984 3359 -950
rect 3301 -1009 3359 -984
rect 3449 -134 3507 -109
rect 3449 -168 3461 -134
rect 3495 -168 3507 -134
rect 3449 -202 3507 -168
rect 3449 -236 3461 -202
rect 3495 -236 3507 -202
rect 3449 -270 3507 -236
rect 3449 -304 3461 -270
rect 3495 -304 3507 -270
rect 3449 -338 3507 -304
rect 3449 -372 3461 -338
rect 3495 -372 3507 -338
rect 3449 -406 3507 -372
rect 3449 -440 3461 -406
rect 3495 -440 3507 -406
rect 3449 -474 3507 -440
rect 3449 -508 3461 -474
rect 3495 -508 3507 -474
rect 3449 -542 3507 -508
rect 3449 -576 3461 -542
rect 3495 -576 3507 -542
rect 3449 -610 3507 -576
rect 3449 -644 3461 -610
rect 3495 -644 3507 -610
rect 3449 -678 3507 -644
rect 3449 -712 3461 -678
rect 3495 -712 3507 -678
rect 3449 -746 3507 -712
rect 3449 -780 3461 -746
rect 3495 -780 3507 -746
rect 3449 -814 3507 -780
rect 3449 -848 3461 -814
rect 3495 -848 3507 -814
rect 3449 -882 3507 -848
rect 3449 -916 3461 -882
rect 3495 -916 3507 -882
rect 3449 -950 3507 -916
rect 3449 -984 3461 -950
rect 3495 -984 3507 -950
rect 3449 -1009 3507 -984
rect 3597 -134 3655 -109
rect 3597 -168 3609 -134
rect 3643 -168 3655 -134
rect 3597 -202 3655 -168
rect 3597 -236 3609 -202
rect 3643 -236 3655 -202
rect 3597 -270 3655 -236
rect 3597 -304 3609 -270
rect 3643 -304 3655 -270
rect 3597 -338 3655 -304
rect 3597 -372 3609 -338
rect 3643 -372 3655 -338
rect 3597 -406 3655 -372
rect 3597 -440 3609 -406
rect 3643 -440 3655 -406
rect 3597 -474 3655 -440
rect 3597 -508 3609 -474
rect 3643 -508 3655 -474
rect 3597 -542 3655 -508
rect 3597 -576 3609 -542
rect 3643 -576 3655 -542
rect 3597 -610 3655 -576
rect 3597 -644 3609 -610
rect 3643 -644 3655 -610
rect 3597 -678 3655 -644
rect 3597 -712 3609 -678
rect 3643 -712 3655 -678
rect 3597 -746 3655 -712
rect 3597 -780 3609 -746
rect 3643 -780 3655 -746
rect 3597 -814 3655 -780
rect 3597 -848 3609 -814
rect 3643 -848 3655 -814
rect 3597 -882 3655 -848
rect 3597 -916 3609 -882
rect 3643 -916 3655 -882
rect 3597 -950 3655 -916
rect 3597 -984 3609 -950
rect 3643 -984 3655 -950
rect 3597 -1009 3655 -984
rect 3745 -134 3803 -109
rect 3745 -168 3757 -134
rect 3791 -168 3803 -134
rect 3745 -202 3803 -168
rect 3745 -236 3757 -202
rect 3791 -236 3803 -202
rect 3745 -270 3803 -236
rect 3745 -304 3757 -270
rect 3791 -304 3803 -270
rect 3745 -338 3803 -304
rect 3745 -372 3757 -338
rect 3791 -372 3803 -338
rect 3745 -406 3803 -372
rect 3745 -440 3757 -406
rect 3791 -440 3803 -406
rect 3745 -474 3803 -440
rect 3745 -508 3757 -474
rect 3791 -508 3803 -474
rect 3745 -542 3803 -508
rect 3745 -576 3757 -542
rect 3791 -576 3803 -542
rect 3745 -610 3803 -576
rect 3745 -644 3757 -610
rect 3791 -644 3803 -610
rect 3745 -678 3803 -644
rect 3745 -712 3757 -678
rect 3791 -712 3803 -678
rect 3745 -746 3803 -712
rect 3745 -780 3757 -746
rect 3791 -780 3803 -746
rect 3745 -814 3803 -780
rect 3745 -848 3757 -814
rect 3791 -848 3803 -814
rect 3745 -882 3803 -848
rect 3745 -916 3757 -882
rect 3791 -916 3803 -882
rect 3745 -950 3803 -916
rect 3745 -984 3757 -950
rect 3791 -984 3803 -950
rect 3745 -1009 3803 -984
rect 3893 -134 3951 -109
rect 3893 -168 3905 -134
rect 3939 -168 3951 -134
rect 3893 -202 3951 -168
rect 3893 -236 3905 -202
rect 3939 -236 3951 -202
rect 3893 -270 3951 -236
rect 3893 -304 3905 -270
rect 3939 -304 3951 -270
rect 3893 -338 3951 -304
rect 3893 -372 3905 -338
rect 3939 -372 3951 -338
rect 3893 -406 3951 -372
rect 3893 -440 3905 -406
rect 3939 -440 3951 -406
rect 3893 -474 3951 -440
rect 3893 -508 3905 -474
rect 3939 -508 3951 -474
rect 3893 -542 3951 -508
rect 3893 -576 3905 -542
rect 3939 -576 3951 -542
rect 3893 -610 3951 -576
rect 3893 -644 3905 -610
rect 3939 -644 3951 -610
rect 3893 -678 3951 -644
rect 3893 -712 3905 -678
rect 3939 -712 3951 -678
rect 3893 -746 3951 -712
rect 3893 -780 3905 -746
rect 3939 -780 3951 -746
rect 3893 -814 3951 -780
rect 3893 -848 3905 -814
rect 3939 -848 3951 -814
rect 3893 -882 3951 -848
rect 3893 -916 3905 -882
rect 3939 -916 3951 -882
rect 3893 -950 3951 -916
rect 3893 -984 3905 -950
rect 3939 -984 3951 -950
rect 3893 -1009 3951 -984
rect 4041 -134 4099 -109
rect 4041 -168 4053 -134
rect 4087 -168 4099 -134
rect 4041 -202 4099 -168
rect 4041 -236 4053 -202
rect 4087 -236 4099 -202
rect 4041 -270 4099 -236
rect 4041 -304 4053 -270
rect 4087 -304 4099 -270
rect 4041 -338 4099 -304
rect 4041 -372 4053 -338
rect 4087 -372 4099 -338
rect 4041 -406 4099 -372
rect 4041 -440 4053 -406
rect 4087 -440 4099 -406
rect 4041 -474 4099 -440
rect 4041 -508 4053 -474
rect 4087 -508 4099 -474
rect 4041 -542 4099 -508
rect 4041 -576 4053 -542
rect 4087 -576 4099 -542
rect 4041 -610 4099 -576
rect 4041 -644 4053 -610
rect 4087 -644 4099 -610
rect 4041 -678 4099 -644
rect 4041 -712 4053 -678
rect 4087 -712 4099 -678
rect 4041 -746 4099 -712
rect 4041 -780 4053 -746
rect 4087 -780 4099 -746
rect 4041 -814 4099 -780
rect 4041 -848 4053 -814
rect 4087 -848 4099 -814
rect 4041 -882 4099 -848
rect 4041 -916 4053 -882
rect 4087 -916 4099 -882
rect 4041 -950 4099 -916
rect 4041 -984 4053 -950
rect 4087 -984 4099 -950
rect 4041 -1009 4099 -984
rect 4189 -134 4247 -109
rect 4189 -168 4201 -134
rect 4235 -168 4247 -134
rect 4189 -202 4247 -168
rect 4189 -236 4201 -202
rect 4235 -236 4247 -202
rect 4189 -270 4247 -236
rect 4189 -304 4201 -270
rect 4235 -304 4247 -270
rect 4189 -338 4247 -304
rect 4189 -372 4201 -338
rect 4235 -372 4247 -338
rect 4189 -406 4247 -372
rect 4189 -440 4201 -406
rect 4235 -440 4247 -406
rect 4189 -474 4247 -440
rect 4189 -508 4201 -474
rect 4235 -508 4247 -474
rect 4189 -542 4247 -508
rect 4189 -576 4201 -542
rect 4235 -576 4247 -542
rect 4189 -610 4247 -576
rect 4189 -644 4201 -610
rect 4235 -644 4247 -610
rect 4189 -678 4247 -644
rect 4189 -712 4201 -678
rect 4235 -712 4247 -678
rect 4189 -746 4247 -712
rect 4189 -780 4201 -746
rect 4235 -780 4247 -746
rect 4189 -814 4247 -780
rect 4189 -848 4201 -814
rect 4235 -848 4247 -814
rect 4189 -882 4247 -848
rect 4189 -916 4201 -882
rect 4235 -916 4247 -882
rect 4189 -950 4247 -916
rect 4189 -984 4201 -950
rect 4235 -984 4247 -950
rect 4189 -1009 4247 -984
rect 4337 -134 4395 -109
rect 4337 -168 4349 -134
rect 4383 -168 4395 -134
rect 4337 -202 4395 -168
rect 4337 -236 4349 -202
rect 4383 -236 4395 -202
rect 4337 -270 4395 -236
rect 4337 -304 4349 -270
rect 4383 -304 4395 -270
rect 4337 -338 4395 -304
rect 4337 -372 4349 -338
rect 4383 -372 4395 -338
rect 4337 -406 4395 -372
rect 4337 -440 4349 -406
rect 4383 -440 4395 -406
rect 4337 -474 4395 -440
rect 4337 -508 4349 -474
rect 4383 -508 4395 -474
rect 4337 -542 4395 -508
rect 4337 -576 4349 -542
rect 4383 -576 4395 -542
rect 4337 -610 4395 -576
rect 4337 -644 4349 -610
rect 4383 -644 4395 -610
rect 4337 -678 4395 -644
rect 4337 -712 4349 -678
rect 4383 -712 4395 -678
rect 4337 -746 4395 -712
rect 4337 -780 4349 -746
rect 4383 -780 4395 -746
rect 4337 -814 4395 -780
rect 4337 -848 4349 -814
rect 4383 -848 4395 -814
rect 4337 -882 4395 -848
rect 4337 -916 4349 -882
rect 4383 -916 4395 -882
rect 4337 -950 4395 -916
rect 4337 -984 4349 -950
rect 4383 -984 4395 -950
rect 4337 -1009 4395 -984
rect 4485 -134 4543 -109
rect 4485 -168 4497 -134
rect 4531 -168 4543 -134
rect 4485 -202 4543 -168
rect 4485 -236 4497 -202
rect 4531 -236 4543 -202
rect 4485 -270 4543 -236
rect 4485 -304 4497 -270
rect 4531 -304 4543 -270
rect 4485 -338 4543 -304
rect 4485 -372 4497 -338
rect 4531 -372 4543 -338
rect 4485 -406 4543 -372
rect 4485 -440 4497 -406
rect 4531 -440 4543 -406
rect 4485 -474 4543 -440
rect 4485 -508 4497 -474
rect 4531 -508 4543 -474
rect 4485 -542 4543 -508
rect 4485 -576 4497 -542
rect 4531 -576 4543 -542
rect 4485 -610 4543 -576
rect 4485 -644 4497 -610
rect 4531 -644 4543 -610
rect 4485 -678 4543 -644
rect 4485 -712 4497 -678
rect 4531 -712 4543 -678
rect 4485 -746 4543 -712
rect 4485 -780 4497 -746
rect 4531 -780 4543 -746
rect 4485 -814 4543 -780
rect 4485 -848 4497 -814
rect 4531 -848 4543 -814
rect 4485 -882 4543 -848
rect 4485 -916 4497 -882
rect 4531 -916 4543 -882
rect 4485 -950 4543 -916
rect 4485 -984 4497 -950
rect 4531 -984 4543 -950
rect 4485 -1009 4543 -984
rect 4633 -134 4691 -109
rect 4633 -168 4645 -134
rect 4679 -168 4691 -134
rect 4633 -202 4691 -168
rect 4633 -236 4645 -202
rect 4679 -236 4691 -202
rect 4633 -270 4691 -236
rect 4633 -304 4645 -270
rect 4679 -304 4691 -270
rect 4633 -338 4691 -304
rect 4633 -372 4645 -338
rect 4679 -372 4691 -338
rect 4633 -406 4691 -372
rect 4633 -440 4645 -406
rect 4679 -440 4691 -406
rect 4633 -474 4691 -440
rect 4633 -508 4645 -474
rect 4679 -508 4691 -474
rect 4633 -542 4691 -508
rect 4633 -576 4645 -542
rect 4679 -576 4691 -542
rect 4633 -610 4691 -576
rect 4633 -644 4645 -610
rect 4679 -644 4691 -610
rect 4633 -678 4691 -644
rect 4633 -712 4645 -678
rect 4679 -712 4691 -678
rect 4633 -746 4691 -712
rect 4633 -780 4645 -746
rect 4679 -780 4691 -746
rect 4633 -814 4691 -780
rect 4633 -848 4645 -814
rect 4679 -848 4691 -814
rect 4633 -882 4691 -848
rect 4633 -916 4645 -882
rect 4679 -916 4691 -882
rect 4633 -950 4691 -916
rect 4633 -984 4645 -950
rect 4679 -984 4691 -950
rect 4633 -1009 4691 -984
rect 4781 -134 4839 -109
rect 4781 -168 4793 -134
rect 4827 -168 4839 -134
rect 4781 -202 4839 -168
rect 4781 -236 4793 -202
rect 4827 -236 4839 -202
rect 4781 -270 4839 -236
rect 4781 -304 4793 -270
rect 4827 -304 4839 -270
rect 4781 -338 4839 -304
rect 4781 -372 4793 -338
rect 4827 -372 4839 -338
rect 4781 -406 4839 -372
rect 4781 -440 4793 -406
rect 4827 -440 4839 -406
rect 4781 -474 4839 -440
rect 4781 -508 4793 -474
rect 4827 -508 4839 -474
rect 4781 -542 4839 -508
rect 4781 -576 4793 -542
rect 4827 -576 4839 -542
rect 4781 -610 4839 -576
rect 4781 -644 4793 -610
rect 4827 -644 4839 -610
rect 4781 -678 4839 -644
rect 4781 -712 4793 -678
rect 4827 -712 4839 -678
rect 4781 -746 4839 -712
rect 4781 -780 4793 -746
rect 4827 -780 4839 -746
rect 4781 -814 4839 -780
rect 4781 -848 4793 -814
rect 4827 -848 4839 -814
rect 4781 -882 4839 -848
rect 4781 -916 4793 -882
rect 4827 -916 4839 -882
rect 4781 -950 4839 -916
rect 4781 -984 4793 -950
rect 4827 -984 4839 -950
rect 4781 -1009 4839 -984
rect 4929 -134 4987 -109
rect 4929 -168 4941 -134
rect 4975 -168 4987 -134
rect 4929 -202 4987 -168
rect 4929 -236 4941 -202
rect 4975 -236 4987 -202
rect 4929 -270 4987 -236
rect 4929 -304 4941 -270
rect 4975 -304 4987 -270
rect 4929 -338 4987 -304
rect 4929 -372 4941 -338
rect 4975 -372 4987 -338
rect 4929 -406 4987 -372
rect 4929 -440 4941 -406
rect 4975 -440 4987 -406
rect 4929 -474 4987 -440
rect 4929 -508 4941 -474
rect 4975 -508 4987 -474
rect 4929 -542 4987 -508
rect 4929 -576 4941 -542
rect 4975 -576 4987 -542
rect 4929 -610 4987 -576
rect 4929 -644 4941 -610
rect 4975 -644 4987 -610
rect 4929 -678 4987 -644
rect 4929 -712 4941 -678
rect 4975 -712 4987 -678
rect 4929 -746 4987 -712
rect 4929 -780 4941 -746
rect 4975 -780 4987 -746
rect 4929 -814 4987 -780
rect 4929 -848 4941 -814
rect 4975 -848 4987 -814
rect 4929 -882 4987 -848
rect 4929 -916 4941 -882
rect 4975 -916 4987 -882
rect 4929 -950 4987 -916
rect 4929 -984 4941 -950
rect 4975 -984 4987 -950
rect 4929 -1009 4987 -984
rect 5077 -134 5135 -109
rect 5077 -168 5089 -134
rect 5123 -168 5135 -134
rect 5077 -202 5135 -168
rect 5077 -236 5089 -202
rect 5123 -236 5135 -202
rect 5077 -270 5135 -236
rect 5077 -304 5089 -270
rect 5123 -304 5135 -270
rect 5077 -338 5135 -304
rect 5077 -372 5089 -338
rect 5123 -372 5135 -338
rect 5077 -406 5135 -372
rect 5077 -440 5089 -406
rect 5123 -440 5135 -406
rect 5077 -474 5135 -440
rect 5077 -508 5089 -474
rect 5123 -508 5135 -474
rect 5077 -542 5135 -508
rect 5077 -576 5089 -542
rect 5123 -576 5135 -542
rect 5077 -610 5135 -576
rect 5077 -644 5089 -610
rect 5123 -644 5135 -610
rect 5077 -678 5135 -644
rect 5077 -712 5089 -678
rect 5123 -712 5135 -678
rect 5077 -746 5135 -712
rect 5077 -780 5089 -746
rect 5123 -780 5135 -746
rect 5077 -814 5135 -780
rect 5077 -848 5089 -814
rect 5123 -848 5135 -814
rect 5077 -882 5135 -848
rect 5077 -916 5089 -882
rect 5123 -916 5135 -882
rect 5077 -950 5135 -916
rect 5077 -984 5089 -950
rect 5123 -984 5135 -950
rect 5077 -1009 5135 -984
rect 5225 -134 5283 -109
rect 5225 -168 5237 -134
rect 5271 -168 5283 -134
rect 5225 -202 5283 -168
rect 5225 -236 5237 -202
rect 5271 -236 5283 -202
rect 5225 -270 5283 -236
rect 5225 -304 5237 -270
rect 5271 -304 5283 -270
rect 5225 -338 5283 -304
rect 5225 -372 5237 -338
rect 5271 -372 5283 -338
rect 5225 -406 5283 -372
rect 5225 -440 5237 -406
rect 5271 -440 5283 -406
rect 5225 -474 5283 -440
rect 5225 -508 5237 -474
rect 5271 -508 5283 -474
rect 5225 -542 5283 -508
rect 5225 -576 5237 -542
rect 5271 -576 5283 -542
rect 5225 -610 5283 -576
rect 5225 -644 5237 -610
rect 5271 -644 5283 -610
rect 5225 -678 5283 -644
rect 5225 -712 5237 -678
rect 5271 -712 5283 -678
rect 5225 -746 5283 -712
rect 5225 -780 5237 -746
rect 5271 -780 5283 -746
rect 5225 -814 5283 -780
rect 5225 -848 5237 -814
rect 5271 -848 5283 -814
rect 5225 -882 5283 -848
rect 5225 -916 5237 -882
rect 5271 -916 5283 -882
rect 5225 -950 5283 -916
rect 5225 -984 5237 -950
rect 5271 -984 5283 -950
rect 5225 -1009 5283 -984
rect 5373 -134 5431 -109
rect 5373 -168 5385 -134
rect 5419 -168 5431 -134
rect 5373 -202 5431 -168
rect 5373 -236 5385 -202
rect 5419 -236 5431 -202
rect 5373 -270 5431 -236
rect 5373 -304 5385 -270
rect 5419 -304 5431 -270
rect 5373 -338 5431 -304
rect 5373 -372 5385 -338
rect 5419 -372 5431 -338
rect 5373 -406 5431 -372
rect 5373 -440 5385 -406
rect 5419 -440 5431 -406
rect 5373 -474 5431 -440
rect 5373 -508 5385 -474
rect 5419 -508 5431 -474
rect 5373 -542 5431 -508
rect 5373 -576 5385 -542
rect 5419 -576 5431 -542
rect 5373 -610 5431 -576
rect 5373 -644 5385 -610
rect 5419 -644 5431 -610
rect 5373 -678 5431 -644
rect 5373 -712 5385 -678
rect 5419 -712 5431 -678
rect 5373 -746 5431 -712
rect 5373 -780 5385 -746
rect 5419 -780 5431 -746
rect 5373 -814 5431 -780
rect 5373 -848 5385 -814
rect 5419 -848 5431 -814
rect 5373 -882 5431 -848
rect 5373 -916 5385 -882
rect 5419 -916 5431 -882
rect 5373 -950 5431 -916
rect 5373 -984 5385 -950
rect 5419 -984 5431 -950
rect 5373 -1009 5431 -984
rect 5521 -134 5579 -109
rect 5521 -168 5533 -134
rect 5567 -168 5579 -134
rect 5521 -202 5579 -168
rect 5521 -236 5533 -202
rect 5567 -236 5579 -202
rect 5521 -270 5579 -236
rect 5521 -304 5533 -270
rect 5567 -304 5579 -270
rect 5521 -338 5579 -304
rect 5521 -372 5533 -338
rect 5567 -372 5579 -338
rect 5521 -406 5579 -372
rect 5521 -440 5533 -406
rect 5567 -440 5579 -406
rect 5521 -474 5579 -440
rect 5521 -508 5533 -474
rect 5567 -508 5579 -474
rect 5521 -542 5579 -508
rect 5521 -576 5533 -542
rect 5567 -576 5579 -542
rect 5521 -610 5579 -576
rect 5521 -644 5533 -610
rect 5567 -644 5579 -610
rect 5521 -678 5579 -644
rect 5521 -712 5533 -678
rect 5567 -712 5579 -678
rect 5521 -746 5579 -712
rect 5521 -780 5533 -746
rect 5567 -780 5579 -746
rect 5521 -814 5579 -780
rect 5521 -848 5533 -814
rect 5567 -848 5579 -814
rect 5521 -882 5579 -848
rect 5521 -916 5533 -882
rect 5567 -916 5579 -882
rect 5521 -950 5579 -916
rect 5521 -984 5533 -950
rect 5567 -984 5579 -950
rect 5521 -1009 5579 -984
<< ndiffc >>
rect -5567 950 -5533 984
rect -5567 882 -5533 916
rect -5567 814 -5533 848
rect -5567 746 -5533 780
rect -5567 678 -5533 712
rect -5567 610 -5533 644
rect -5567 542 -5533 576
rect -5567 474 -5533 508
rect -5567 406 -5533 440
rect -5567 338 -5533 372
rect -5567 270 -5533 304
rect -5567 202 -5533 236
rect -5567 134 -5533 168
rect -5419 950 -5385 984
rect -5419 882 -5385 916
rect -5419 814 -5385 848
rect -5419 746 -5385 780
rect -5419 678 -5385 712
rect -5419 610 -5385 644
rect -5419 542 -5385 576
rect -5419 474 -5385 508
rect -5419 406 -5385 440
rect -5419 338 -5385 372
rect -5419 270 -5385 304
rect -5419 202 -5385 236
rect -5419 134 -5385 168
rect -5271 950 -5237 984
rect -5271 882 -5237 916
rect -5271 814 -5237 848
rect -5271 746 -5237 780
rect -5271 678 -5237 712
rect -5271 610 -5237 644
rect -5271 542 -5237 576
rect -5271 474 -5237 508
rect -5271 406 -5237 440
rect -5271 338 -5237 372
rect -5271 270 -5237 304
rect -5271 202 -5237 236
rect -5271 134 -5237 168
rect -5123 950 -5089 984
rect -5123 882 -5089 916
rect -5123 814 -5089 848
rect -5123 746 -5089 780
rect -5123 678 -5089 712
rect -5123 610 -5089 644
rect -5123 542 -5089 576
rect -5123 474 -5089 508
rect -5123 406 -5089 440
rect -5123 338 -5089 372
rect -5123 270 -5089 304
rect -5123 202 -5089 236
rect -5123 134 -5089 168
rect -4975 950 -4941 984
rect -4975 882 -4941 916
rect -4975 814 -4941 848
rect -4975 746 -4941 780
rect -4975 678 -4941 712
rect -4975 610 -4941 644
rect -4975 542 -4941 576
rect -4975 474 -4941 508
rect -4975 406 -4941 440
rect -4975 338 -4941 372
rect -4975 270 -4941 304
rect -4975 202 -4941 236
rect -4975 134 -4941 168
rect -4827 950 -4793 984
rect -4827 882 -4793 916
rect -4827 814 -4793 848
rect -4827 746 -4793 780
rect -4827 678 -4793 712
rect -4827 610 -4793 644
rect -4827 542 -4793 576
rect -4827 474 -4793 508
rect -4827 406 -4793 440
rect -4827 338 -4793 372
rect -4827 270 -4793 304
rect -4827 202 -4793 236
rect -4827 134 -4793 168
rect -4679 950 -4645 984
rect -4679 882 -4645 916
rect -4679 814 -4645 848
rect -4679 746 -4645 780
rect -4679 678 -4645 712
rect -4679 610 -4645 644
rect -4679 542 -4645 576
rect -4679 474 -4645 508
rect -4679 406 -4645 440
rect -4679 338 -4645 372
rect -4679 270 -4645 304
rect -4679 202 -4645 236
rect -4679 134 -4645 168
rect -4531 950 -4497 984
rect -4531 882 -4497 916
rect -4531 814 -4497 848
rect -4531 746 -4497 780
rect -4531 678 -4497 712
rect -4531 610 -4497 644
rect -4531 542 -4497 576
rect -4531 474 -4497 508
rect -4531 406 -4497 440
rect -4531 338 -4497 372
rect -4531 270 -4497 304
rect -4531 202 -4497 236
rect -4531 134 -4497 168
rect -4383 950 -4349 984
rect -4383 882 -4349 916
rect -4383 814 -4349 848
rect -4383 746 -4349 780
rect -4383 678 -4349 712
rect -4383 610 -4349 644
rect -4383 542 -4349 576
rect -4383 474 -4349 508
rect -4383 406 -4349 440
rect -4383 338 -4349 372
rect -4383 270 -4349 304
rect -4383 202 -4349 236
rect -4383 134 -4349 168
rect -4235 950 -4201 984
rect -4235 882 -4201 916
rect -4235 814 -4201 848
rect -4235 746 -4201 780
rect -4235 678 -4201 712
rect -4235 610 -4201 644
rect -4235 542 -4201 576
rect -4235 474 -4201 508
rect -4235 406 -4201 440
rect -4235 338 -4201 372
rect -4235 270 -4201 304
rect -4235 202 -4201 236
rect -4235 134 -4201 168
rect -4087 950 -4053 984
rect -4087 882 -4053 916
rect -4087 814 -4053 848
rect -4087 746 -4053 780
rect -4087 678 -4053 712
rect -4087 610 -4053 644
rect -4087 542 -4053 576
rect -4087 474 -4053 508
rect -4087 406 -4053 440
rect -4087 338 -4053 372
rect -4087 270 -4053 304
rect -4087 202 -4053 236
rect -4087 134 -4053 168
rect -3939 950 -3905 984
rect -3939 882 -3905 916
rect -3939 814 -3905 848
rect -3939 746 -3905 780
rect -3939 678 -3905 712
rect -3939 610 -3905 644
rect -3939 542 -3905 576
rect -3939 474 -3905 508
rect -3939 406 -3905 440
rect -3939 338 -3905 372
rect -3939 270 -3905 304
rect -3939 202 -3905 236
rect -3939 134 -3905 168
rect -3791 950 -3757 984
rect -3791 882 -3757 916
rect -3791 814 -3757 848
rect -3791 746 -3757 780
rect -3791 678 -3757 712
rect -3791 610 -3757 644
rect -3791 542 -3757 576
rect -3791 474 -3757 508
rect -3791 406 -3757 440
rect -3791 338 -3757 372
rect -3791 270 -3757 304
rect -3791 202 -3757 236
rect -3791 134 -3757 168
rect -3643 950 -3609 984
rect -3643 882 -3609 916
rect -3643 814 -3609 848
rect -3643 746 -3609 780
rect -3643 678 -3609 712
rect -3643 610 -3609 644
rect -3643 542 -3609 576
rect -3643 474 -3609 508
rect -3643 406 -3609 440
rect -3643 338 -3609 372
rect -3643 270 -3609 304
rect -3643 202 -3609 236
rect -3643 134 -3609 168
rect -3495 950 -3461 984
rect -3495 882 -3461 916
rect -3495 814 -3461 848
rect -3495 746 -3461 780
rect -3495 678 -3461 712
rect -3495 610 -3461 644
rect -3495 542 -3461 576
rect -3495 474 -3461 508
rect -3495 406 -3461 440
rect -3495 338 -3461 372
rect -3495 270 -3461 304
rect -3495 202 -3461 236
rect -3495 134 -3461 168
rect -3347 950 -3313 984
rect -3347 882 -3313 916
rect -3347 814 -3313 848
rect -3347 746 -3313 780
rect -3347 678 -3313 712
rect -3347 610 -3313 644
rect -3347 542 -3313 576
rect -3347 474 -3313 508
rect -3347 406 -3313 440
rect -3347 338 -3313 372
rect -3347 270 -3313 304
rect -3347 202 -3313 236
rect -3347 134 -3313 168
rect -3199 950 -3165 984
rect -3199 882 -3165 916
rect -3199 814 -3165 848
rect -3199 746 -3165 780
rect -3199 678 -3165 712
rect -3199 610 -3165 644
rect -3199 542 -3165 576
rect -3199 474 -3165 508
rect -3199 406 -3165 440
rect -3199 338 -3165 372
rect -3199 270 -3165 304
rect -3199 202 -3165 236
rect -3199 134 -3165 168
rect -3051 950 -3017 984
rect -3051 882 -3017 916
rect -3051 814 -3017 848
rect -3051 746 -3017 780
rect -3051 678 -3017 712
rect -3051 610 -3017 644
rect -3051 542 -3017 576
rect -3051 474 -3017 508
rect -3051 406 -3017 440
rect -3051 338 -3017 372
rect -3051 270 -3017 304
rect -3051 202 -3017 236
rect -3051 134 -3017 168
rect -2903 950 -2869 984
rect -2903 882 -2869 916
rect -2903 814 -2869 848
rect -2903 746 -2869 780
rect -2903 678 -2869 712
rect -2903 610 -2869 644
rect -2903 542 -2869 576
rect -2903 474 -2869 508
rect -2903 406 -2869 440
rect -2903 338 -2869 372
rect -2903 270 -2869 304
rect -2903 202 -2869 236
rect -2903 134 -2869 168
rect -2755 950 -2721 984
rect -2755 882 -2721 916
rect -2755 814 -2721 848
rect -2755 746 -2721 780
rect -2755 678 -2721 712
rect -2755 610 -2721 644
rect -2755 542 -2721 576
rect -2755 474 -2721 508
rect -2755 406 -2721 440
rect -2755 338 -2721 372
rect -2755 270 -2721 304
rect -2755 202 -2721 236
rect -2755 134 -2721 168
rect -2607 950 -2573 984
rect -2607 882 -2573 916
rect -2607 814 -2573 848
rect -2607 746 -2573 780
rect -2607 678 -2573 712
rect -2607 610 -2573 644
rect -2607 542 -2573 576
rect -2607 474 -2573 508
rect -2607 406 -2573 440
rect -2607 338 -2573 372
rect -2607 270 -2573 304
rect -2607 202 -2573 236
rect -2607 134 -2573 168
rect -2459 950 -2425 984
rect -2459 882 -2425 916
rect -2459 814 -2425 848
rect -2459 746 -2425 780
rect -2459 678 -2425 712
rect -2459 610 -2425 644
rect -2459 542 -2425 576
rect -2459 474 -2425 508
rect -2459 406 -2425 440
rect -2459 338 -2425 372
rect -2459 270 -2425 304
rect -2459 202 -2425 236
rect -2459 134 -2425 168
rect -2311 950 -2277 984
rect -2311 882 -2277 916
rect -2311 814 -2277 848
rect -2311 746 -2277 780
rect -2311 678 -2277 712
rect -2311 610 -2277 644
rect -2311 542 -2277 576
rect -2311 474 -2277 508
rect -2311 406 -2277 440
rect -2311 338 -2277 372
rect -2311 270 -2277 304
rect -2311 202 -2277 236
rect -2311 134 -2277 168
rect -2163 950 -2129 984
rect -2163 882 -2129 916
rect -2163 814 -2129 848
rect -2163 746 -2129 780
rect -2163 678 -2129 712
rect -2163 610 -2129 644
rect -2163 542 -2129 576
rect -2163 474 -2129 508
rect -2163 406 -2129 440
rect -2163 338 -2129 372
rect -2163 270 -2129 304
rect -2163 202 -2129 236
rect -2163 134 -2129 168
rect -2015 950 -1981 984
rect -2015 882 -1981 916
rect -2015 814 -1981 848
rect -2015 746 -1981 780
rect -2015 678 -1981 712
rect -2015 610 -1981 644
rect -2015 542 -1981 576
rect -2015 474 -1981 508
rect -2015 406 -1981 440
rect -2015 338 -1981 372
rect -2015 270 -1981 304
rect -2015 202 -1981 236
rect -2015 134 -1981 168
rect -1867 950 -1833 984
rect -1867 882 -1833 916
rect -1867 814 -1833 848
rect -1867 746 -1833 780
rect -1867 678 -1833 712
rect -1867 610 -1833 644
rect -1867 542 -1833 576
rect -1867 474 -1833 508
rect -1867 406 -1833 440
rect -1867 338 -1833 372
rect -1867 270 -1833 304
rect -1867 202 -1833 236
rect -1867 134 -1833 168
rect -1719 950 -1685 984
rect -1719 882 -1685 916
rect -1719 814 -1685 848
rect -1719 746 -1685 780
rect -1719 678 -1685 712
rect -1719 610 -1685 644
rect -1719 542 -1685 576
rect -1719 474 -1685 508
rect -1719 406 -1685 440
rect -1719 338 -1685 372
rect -1719 270 -1685 304
rect -1719 202 -1685 236
rect -1719 134 -1685 168
rect -1571 950 -1537 984
rect -1571 882 -1537 916
rect -1571 814 -1537 848
rect -1571 746 -1537 780
rect -1571 678 -1537 712
rect -1571 610 -1537 644
rect -1571 542 -1537 576
rect -1571 474 -1537 508
rect -1571 406 -1537 440
rect -1571 338 -1537 372
rect -1571 270 -1537 304
rect -1571 202 -1537 236
rect -1571 134 -1537 168
rect -1423 950 -1389 984
rect -1423 882 -1389 916
rect -1423 814 -1389 848
rect -1423 746 -1389 780
rect -1423 678 -1389 712
rect -1423 610 -1389 644
rect -1423 542 -1389 576
rect -1423 474 -1389 508
rect -1423 406 -1389 440
rect -1423 338 -1389 372
rect -1423 270 -1389 304
rect -1423 202 -1389 236
rect -1423 134 -1389 168
rect -1275 950 -1241 984
rect -1275 882 -1241 916
rect -1275 814 -1241 848
rect -1275 746 -1241 780
rect -1275 678 -1241 712
rect -1275 610 -1241 644
rect -1275 542 -1241 576
rect -1275 474 -1241 508
rect -1275 406 -1241 440
rect -1275 338 -1241 372
rect -1275 270 -1241 304
rect -1275 202 -1241 236
rect -1275 134 -1241 168
rect -1127 950 -1093 984
rect -1127 882 -1093 916
rect -1127 814 -1093 848
rect -1127 746 -1093 780
rect -1127 678 -1093 712
rect -1127 610 -1093 644
rect -1127 542 -1093 576
rect -1127 474 -1093 508
rect -1127 406 -1093 440
rect -1127 338 -1093 372
rect -1127 270 -1093 304
rect -1127 202 -1093 236
rect -1127 134 -1093 168
rect -979 950 -945 984
rect -979 882 -945 916
rect -979 814 -945 848
rect -979 746 -945 780
rect -979 678 -945 712
rect -979 610 -945 644
rect -979 542 -945 576
rect -979 474 -945 508
rect -979 406 -945 440
rect -979 338 -945 372
rect -979 270 -945 304
rect -979 202 -945 236
rect -979 134 -945 168
rect -831 950 -797 984
rect -831 882 -797 916
rect -831 814 -797 848
rect -831 746 -797 780
rect -831 678 -797 712
rect -831 610 -797 644
rect -831 542 -797 576
rect -831 474 -797 508
rect -831 406 -797 440
rect -831 338 -797 372
rect -831 270 -797 304
rect -831 202 -797 236
rect -831 134 -797 168
rect -683 950 -649 984
rect -683 882 -649 916
rect -683 814 -649 848
rect -683 746 -649 780
rect -683 678 -649 712
rect -683 610 -649 644
rect -683 542 -649 576
rect -683 474 -649 508
rect -683 406 -649 440
rect -683 338 -649 372
rect -683 270 -649 304
rect -683 202 -649 236
rect -683 134 -649 168
rect -535 950 -501 984
rect -535 882 -501 916
rect -535 814 -501 848
rect -535 746 -501 780
rect -535 678 -501 712
rect -535 610 -501 644
rect -535 542 -501 576
rect -535 474 -501 508
rect -535 406 -501 440
rect -535 338 -501 372
rect -535 270 -501 304
rect -535 202 -501 236
rect -535 134 -501 168
rect -387 950 -353 984
rect -387 882 -353 916
rect -387 814 -353 848
rect -387 746 -353 780
rect -387 678 -353 712
rect -387 610 -353 644
rect -387 542 -353 576
rect -387 474 -353 508
rect -387 406 -353 440
rect -387 338 -353 372
rect -387 270 -353 304
rect -387 202 -353 236
rect -387 134 -353 168
rect -239 950 -205 984
rect -239 882 -205 916
rect -239 814 -205 848
rect -239 746 -205 780
rect -239 678 -205 712
rect -239 610 -205 644
rect -239 542 -205 576
rect -239 474 -205 508
rect -239 406 -205 440
rect -239 338 -205 372
rect -239 270 -205 304
rect -239 202 -205 236
rect -239 134 -205 168
rect -91 950 -57 984
rect -91 882 -57 916
rect -91 814 -57 848
rect -91 746 -57 780
rect -91 678 -57 712
rect -91 610 -57 644
rect -91 542 -57 576
rect -91 474 -57 508
rect -91 406 -57 440
rect -91 338 -57 372
rect -91 270 -57 304
rect -91 202 -57 236
rect -91 134 -57 168
rect 57 950 91 984
rect 57 882 91 916
rect 57 814 91 848
rect 57 746 91 780
rect 57 678 91 712
rect 57 610 91 644
rect 57 542 91 576
rect 57 474 91 508
rect 57 406 91 440
rect 57 338 91 372
rect 57 270 91 304
rect 57 202 91 236
rect 57 134 91 168
rect 205 950 239 984
rect 205 882 239 916
rect 205 814 239 848
rect 205 746 239 780
rect 205 678 239 712
rect 205 610 239 644
rect 205 542 239 576
rect 205 474 239 508
rect 205 406 239 440
rect 205 338 239 372
rect 205 270 239 304
rect 205 202 239 236
rect 205 134 239 168
rect 353 950 387 984
rect 353 882 387 916
rect 353 814 387 848
rect 353 746 387 780
rect 353 678 387 712
rect 353 610 387 644
rect 353 542 387 576
rect 353 474 387 508
rect 353 406 387 440
rect 353 338 387 372
rect 353 270 387 304
rect 353 202 387 236
rect 353 134 387 168
rect 501 950 535 984
rect 501 882 535 916
rect 501 814 535 848
rect 501 746 535 780
rect 501 678 535 712
rect 501 610 535 644
rect 501 542 535 576
rect 501 474 535 508
rect 501 406 535 440
rect 501 338 535 372
rect 501 270 535 304
rect 501 202 535 236
rect 501 134 535 168
rect 649 950 683 984
rect 649 882 683 916
rect 649 814 683 848
rect 649 746 683 780
rect 649 678 683 712
rect 649 610 683 644
rect 649 542 683 576
rect 649 474 683 508
rect 649 406 683 440
rect 649 338 683 372
rect 649 270 683 304
rect 649 202 683 236
rect 649 134 683 168
rect 797 950 831 984
rect 797 882 831 916
rect 797 814 831 848
rect 797 746 831 780
rect 797 678 831 712
rect 797 610 831 644
rect 797 542 831 576
rect 797 474 831 508
rect 797 406 831 440
rect 797 338 831 372
rect 797 270 831 304
rect 797 202 831 236
rect 797 134 831 168
rect 945 950 979 984
rect 945 882 979 916
rect 945 814 979 848
rect 945 746 979 780
rect 945 678 979 712
rect 945 610 979 644
rect 945 542 979 576
rect 945 474 979 508
rect 945 406 979 440
rect 945 338 979 372
rect 945 270 979 304
rect 945 202 979 236
rect 945 134 979 168
rect 1093 950 1127 984
rect 1093 882 1127 916
rect 1093 814 1127 848
rect 1093 746 1127 780
rect 1093 678 1127 712
rect 1093 610 1127 644
rect 1093 542 1127 576
rect 1093 474 1127 508
rect 1093 406 1127 440
rect 1093 338 1127 372
rect 1093 270 1127 304
rect 1093 202 1127 236
rect 1093 134 1127 168
rect 1241 950 1275 984
rect 1241 882 1275 916
rect 1241 814 1275 848
rect 1241 746 1275 780
rect 1241 678 1275 712
rect 1241 610 1275 644
rect 1241 542 1275 576
rect 1241 474 1275 508
rect 1241 406 1275 440
rect 1241 338 1275 372
rect 1241 270 1275 304
rect 1241 202 1275 236
rect 1241 134 1275 168
rect 1389 950 1423 984
rect 1389 882 1423 916
rect 1389 814 1423 848
rect 1389 746 1423 780
rect 1389 678 1423 712
rect 1389 610 1423 644
rect 1389 542 1423 576
rect 1389 474 1423 508
rect 1389 406 1423 440
rect 1389 338 1423 372
rect 1389 270 1423 304
rect 1389 202 1423 236
rect 1389 134 1423 168
rect 1537 950 1571 984
rect 1537 882 1571 916
rect 1537 814 1571 848
rect 1537 746 1571 780
rect 1537 678 1571 712
rect 1537 610 1571 644
rect 1537 542 1571 576
rect 1537 474 1571 508
rect 1537 406 1571 440
rect 1537 338 1571 372
rect 1537 270 1571 304
rect 1537 202 1571 236
rect 1537 134 1571 168
rect 1685 950 1719 984
rect 1685 882 1719 916
rect 1685 814 1719 848
rect 1685 746 1719 780
rect 1685 678 1719 712
rect 1685 610 1719 644
rect 1685 542 1719 576
rect 1685 474 1719 508
rect 1685 406 1719 440
rect 1685 338 1719 372
rect 1685 270 1719 304
rect 1685 202 1719 236
rect 1685 134 1719 168
rect 1833 950 1867 984
rect 1833 882 1867 916
rect 1833 814 1867 848
rect 1833 746 1867 780
rect 1833 678 1867 712
rect 1833 610 1867 644
rect 1833 542 1867 576
rect 1833 474 1867 508
rect 1833 406 1867 440
rect 1833 338 1867 372
rect 1833 270 1867 304
rect 1833 202 1867 236
rect 1833 134 1867 168
rect 1981 950 2015 984
rect 1981 882 2015 916
rect 1981 814 2015 848
rect 1981 746 2015 780
rect 1981 678 2015 712
rect 1981 610 2015 644
rect 1981 542 2015 576
rect 1981 474 2015 508
rect 1981 406 2015 440
rect 1981 338 2015 372
rect 1981 270 2015 304
rect 1981 202 2015 236
rect 1981 134 2015 168
rect 2129 950 2163 984
rect 2129 882 2163 916
rect 2129 814 2163 848
rect 2129 746 2163 780
rect 2129 678 2163 712
rect 2129 610 2163 644
rect 2129 542 2163 576
rect 2129 474 2163 508
rect 2129 406 2163 440
rect 2129 338 2163 372
rect 2129 270 2163 304
rect 2129 202 2163 236
rect 2129 134 2163 168
rect 2277 950 2311 984
rect 2277 882 2311 916
rect 2277 814 2311 848
rect 2277 746 2311 780
rect 2277 678 2311 712
rect 2277 610 2311 644
rect 2277 542 2311 576
rect 2277 474 2311 508
rect 2277 406 2311 440
rect 2277 338 2311 372
rect 2277 270 2311 304
rect 2277 202 2311 236
rect 2277 134 2311 168
rect 2425 950 2459 984
rect 2425 882 2459 916
rect 2425 814 2459 848
rect 2425 746 2459 780
rect 2425 678 2459 712
rect 2425 610 2459 644
rect 2425 542 2459 576
rect 2425 474 2459 508
rect 2425 406 2459 440
rect 2425 338 2459 372
rect 2425 270 2459 304
rect 2425 202 2459 236
rect 2425 134 2459 168
rect 2573 950 2607 984
rect 2573 882 2607 916
rect 2573 814 2607 848
rect 2573 746 2607 780
rect 2573 678 2607 712
rect 2573 610 2607 644
rect 2573 542 2607 576
rect 2573 474 2607 508
rect 2573 406 2607 440
rect 2573 338 2607 372
rect 2573 270 2607 304
rect 2573 202 2607 236
rect 2573 134 2607 168
rect 2721 950 2755 984
rect 2721 882 2755 916
rect 2721 814 2755 848
rect 2721 746 2755 780
rect 2721 678 2755 712
rect 2721 610 2755 644
rect 2721 542 2755 576
rect 2721 474 2755 508
rect 2721 406 2755 440
rect 2721 338 2755 372
rect 2721 270 2755 304
rect 2721 202 2755 236
rect 2721 134 2755 168
rect 2869 950 2903 984
rect 2869 882 2903 916
rect 2869 814 2903 848
rect 2869 746 2903 780
rect 2869 678 2903 712
rect 2869 610 2903 644
rect 2869 542 2903 576
rect 2869 474 2903 508
rect 2869 406 2903 440
rect 2869 338 2903 372
rect 2869 270 2903 304
rect 2869 202 2903 236
rect 2869 134 2903 168
rect 3017 950 3051 984
rect 3017 882 3051 916
rect 3017 814 3051 848
rect 3017 746 3051 780
rect 3017 678 3051 712
rect 3017 610 3051 644
rect 3017 542 3051 576
rect 3017 474 3051 508
rect 3017 406 3051 440
rect 3017 338 3051 372
rect 3017 270 3051 304
rect 3017 202 3051 236
rect 3017 134 3051 168
rect 3165 950 3199 984
rect 3165 882 3199 916
rect 3165 814 3199 848
rect 3165 746 3199 780
rect 3165 678 3199 712
rect 3165 610 3199 644
rect 3165 542 3199 576
rect 3165 474 3199 508
rect 3165 406 3199 440
rect 3165 338 3199 372
rect 3165 270 3199 304
rect 3165 202 3199 236
rect 3165 134 3199 168
rect 3313 950 3347 984
rect 3313 882 3347 916
rect 3313 814 3347 848
rect 3313 746 3347 780
rect 3313 678 3347 712
rect 3313 610 3347 644
rect 3313 542 3347 576
rect 3313 474 3347 508
rect 3313 406 3347 440
rect 3313 338 3347 372
rect 3313 270 3347 304
rect 3313 202 3347 236
rect 3313 134 3347 168
rect 3461 950 3495 984
rect 3461 882 3495 916
rect 3461 814 3495 848
rect 3461 746 3495 780
rect 3461 678 3495 712
rect 3461 610 3495 644
rect 3461 542 3495 576
rect 3461 474 3495 508
rect 3461 406 3495 440
rect 3461 338 3495 372
rect 3461 270 3495 304
rect 3461 202 3495 236
rect 3461 134 3495 168
rect 3609 950 3643 984
rect 3609 882 3643 916
rect 3609 814 3643 848
rect 3609 746 3643 780
rect 3609 678 3643 712
rect 3609 610 3643 644
rect 3609 542 3643 576
rect 3609 474 3643 508
rect 3609 406 3643 440
rect 3609 338 3643 372
rect 3609 270 3643 304
rect 3609 202 3643 236
rect 3609 134 3643 168
rect 3757 950 3791 984
rect 3757 882 3791 916
rect 3757 814 3791 848
rect 3757 746 3791 780
rect 3757 678 3791 712
rect 3757 610 3791 644
rect 3757 542 3791 576
rect 3757 474 3791 508
rect 3757 406 3791 440
rect 3757 338 3791 372
rect 3757 270 3791 304
rect 3757 202 3791 236
rect 3757 134 3791 168
rect 3905 950 3939 984
rect 3905 882 3939 916
rect 3905 814 3939 848
rect 3905 746 3939 780
rect 3905 678 3939 712
rect 3905 610 3939 644
rect 3905 542 3939 576
rect 3905 474 3939 508
rect 3905 406 3939 440
rect 3905 338 3939 372
rect 3905 270 3939 304
rect 3905 202 3939 236
rect 3905 134 3939 168
rect 4053 950 4087 984
rect 4053 882 4087 916
rect 4053 814 4087 848
rect 4053 746 4087 780
rect 4053 678 4087 712
rect 4053 610 4087 644
rect 4053 542 4087 576
rect 4053 474 4087 508
rect 4053 406 4087 440
rect 4053 338 4087 372
rect 4053 270 4087 304
rect 4053 202 4087 236
rect 4053 134 4087 168
rect 4201 950 4235 984
rect 4201 882 4235 916
rect 4201 814 4235 848
rect 4201 746 4235 780
rect 4201 678 4235 712
rect 4201 610 4235 644
rect 4201 542 4235 576
rect 4201 474 4235 508
rect 4201 406 4235 440
rect 4201 338 4235 372
rect 4201 270 4235 304
rect 4201 202 4235 236
rect 4201 134 4235 168
rect 4349 950 4383 984
rect 4349 882 4383 916
rect 4349 814 4383 848
rect 4349 746 4383 780
rect 4349 678 4383 712
rect 4349 610 4383 644
rect 4349 542 4383 576
rect 4349 474 4383 508
rect 4349 406 4383 440
rect 4349 338 4383 372
rect 4349 270 4383 304
rect 4349 202 4383 236
rect 4349 134 4383 168
rect 4497 950 4531 984
rect 4497 882 4531 916
rect 4497 814 4531 848
rect 4497 746 4531 780
rect 4497 678 4531 712
rect 4497 610 4531 644
rect 4497 542 4531 576
rect 4497 474 4531 508
rect 4497 406 4531 440
rect 4497 338 4531 372
rect 4497 270 4531 304
rect 4497 202 4531 236
rect 4497 134 4531 168
rect 4645 950 4679 984
rect 4645 882 4679 916
rect 4645 814 4679 848
rect 4645 746 4679 780
rect 4645 678 4679 712
rect 4645 610 4679 644
rect 4645 542 4679 576
rect 4645 474 4679 508
rect 4645 406 4679 440
rect 4645 338 4679 372
rect 4645 270 4679 304
rect 4645 202 4679 236
rect 4645 134 4679 168
rect 4793 950 4827 984
rect 4793 882 4827 916
rect 4793 814 4827 848
rect 4793 746 4827 780
rect 4793 678 4827 712
rect 4793 610 4827 644
rect 4793 542 4827 576
rect 4793 474 4827 508
rect 4793 406 4827 440
rect 4793 338 4827 372
rect 4793 270 4827 304
rect 4793 202 4827 236
rect 4793 134 4827 168
rect 4941 950 4975 984
rect 4941 882 4975 916
rect 4941 814 4975 848
rect 4941 746 4975 780
rect 4941 678 4975 712
rect 4941 610 4975 644
rect 4941 542 4975 576
rect 4941 474 4975 508
rect 4941 406 4975 440
rect 4941 338 4975 372
rect 4941 270 4975 304
rect 4941 202 4975 236
rect 4941 134 4975 168
rect 5089 950 5123 984
rect 5089 882 5123 916
rect 5089 814 5123 848
rect 5089 746 5123 780
rect 5089 678 5123 712
rect 5089 610 5123 644
rect 5089 542 5123 576
rect 5089 474 5123 508
rect 5089 406 5123 440
rect 5089 338 5123 372
rect 5089 270 5123 304
rect 5089 202 5123 236
rect 5089 134 5123 168
rect 5237 950 5271 984
rect 5237 882 5271 916
rect 5237 814 5271 848
rect 5237 746 5271 780
rect 5237 678 5271 712
rect 5237 610 5271 644
rect 5237 542 5271 576
rect 5237 474 5271 508
rect 5237 406 5271 440
rect 5237 338 5271 372
rect 5237 270 5271 304
rect 5237 202 5271 236
rect 5237 134 5271 168
rect 5385 950 5419 984
rect 5385 882 5419 916
rect 5385 814 5419 848
rect 5385 746 5419 780
rect 5385 678 5419 712
rect 5385 610 5419 644
rect 5385 542 5419 576
rect 5385 474 5419 508
rect 5385 406 5419 440
rect 5385 338 5419 372
rect 5385 270 5419 304
rect 5385 202 5419 236
rect 5385 134 5419 168
rect 5533 950 5567 984
rect 5533 882 5567 916
rect 5533 814 5567 848
rect 5533 746 5567 780
rect 5533 678 5567 712
rect 5533 610 5567 644
rect 5533 542 5567 576
rect 5533 474 5567 508
rect 5533 406 5567 440
rect 5533 338 5567 372
rect 5533 270 5567 304
rect 5533 202 5567 236
rect 5533 134 5567 168
rect -5567 -168 -5533 -134
rect -5567 -236 -5533 -202
rect -5567 -304 -5533 -270
rect -5567 -372 -5533 -338
rect -5567 -440 -5533 -406
rect -5567 -508 -5533 -474
rect -5567 -576 -5533 -542
rect -5567 -644 -5533 -610
rect -5567 -712 -5533 -678
rect -5567 -780 -5533 -746
rect -5567 -848 -5533 -814
rect -5567 -916 -5533 -882
rect -5567 -984 -5533 -950
rect -5419 -168 -5385 -134
rect -5419 -236 -5385 -202
rect -5419 -304 -5385 -270
rect -5419 -372 -5385 -338
rect -5419 -440 -5385 -406
rect -5419 -508 -5385 -474
rect -5419 -576 -5385 -542
rect -5419 -644 -5385 -610
rect -5419 -712 -5385 -678
rect -5419 -780 -5385 -746
rect -5419 -848 -5385 -814
rect -5419 -916 -5385 -882
rect -5419 -984 -5385 -950
rect -5271 -168 -5237 -134
rect -5271 -236 -5237 -202
rect -5271 -304 -5237 -270
rect -5271 -372 -5237 -338
rect -5271 -440 -5237 -406
rect -5271 -508 -5237 -474
rect -5271 -576 -5237 -542
rect -5271 -644 -5237 -610
rect -5271 -712 -5237 -678
rect -5271 -780 -5237 -746
rect -5271 -848 -5237 -814
rect -5271 -916 -5237 -882
rect -5271 -984 -5237 -950
rect -5123 -168 -5089 -134
rect -5123 -236 -5089 -202
rect -5123 -304 -5089 -270
rect -5123 -372 -5089 -338
rect -5123 -440 -5089 -406
rect -5123 -508 -5089 -474
rect -5123 -576 -5089 -542
rect -5123 -644 -5089 -610
rect -5123 -712 -5089 -678
rect -5123 -780 -5089 -746
rect -5123 -848 -5089 -814
rect -5123 -916 -5089 -882
rect -5123 -984 -5089 -950
rect -4975 -168 -4941 -134
rect -4975 -236 -4941 -202
rect -4975 -304 -4941 -270
rect -4975 -372 -4941 -338
rect -4975 -440 -4941 -406
rect -4975 -508 -4941 -474
rect -4975 -576 -4941 -542
rect -4975 -644 -4941 -610
rect -4975 -712 -4941 -678
rect -4975 -780 -4941 -746
rect -4975 -848 -4941 -814
rect -4975 -916 -4941 -882
rect -4975 -984 -4941 -950
rect -4827 -168 -4793 -134
rect -4827 -236 -4793 -202
rect -4827 -304 -4793 -270
rect -4827 -372 -4793 -338
rect -4827 -440 -4793 -406
rect -4827 -508 -4793 -474
rect -4827 -576 -4793 -542
rect -4827 -644 -4793 -610
rect -4827 -712 -4793 -678
rect -4827 -780 -4793 -746
rect -4827 -848 -4793 -814
rect -4827 -916 -4793 -882
rect -4827 -984 -4793 -950
rect -4679 -168 -4645 -134
rect -4679 -236 -4645 -202
rect -4679 -304 -4645 -270
rect -4679 -372 -4645 -338
rect -4679 -440 -4645 -406
rect -4679 -508 -4645 -474
rect -4679 -576 -4645 -542
rect -4679 -644 -4645 -610
rect -4679 -712 -4645 -678
rect -4679 -780 -4645 -746
rect -4679 -848 -4645 -814
rect -4679 -916 -4645 -882
rect -4679 -984 -4645 -950
rect -4531 -168 -4497 -134
rect -4531 -236 -4497 -202
rect -4531 -304 -4497 -270
rect -4531 -372 -4497 -338
rect -4531 -440 -4497 -406
rect -4531 -508 -4497 -474
rect -4531 -576 -4497 -542
rect -4531 -644 -4497 -610
rect -4531 -712 -4497 -678
rect -4531 -780 -4497 -746
rect -4531 -848 -4497 -814
rect -4531 -916 -4497 -882
rect -4531 -984 -4497 -950
rect -4383 -168 -4349 -134
rect -4383 -236 -4349 -202
rect -4383 -304 -4349 -270
rect -4383 -372 -4349 -338
rect -4383 -440 -4349 -406
rect -4383 -508 -4349 -474
rect -4383 -576 -4349 -542
rect -4383 -644 -4349 -610
rect -4383 -712 -4349 -678
rect -4383 -780 -4349 -746
rect -4383 -848 -4349 -814
rect -4383 -916 -4349 -882
rect -4383 -984 -4349 -950
rect -4235 -168 -4201 -134
rect -4235 -236 -4201 -202
rect -4235 -304 -4201 -270
rect -4235 -372 -4201 -338
rect -4235 -440 -4201 -406
rect -4235 -508 -4201 -474
rect -4235 -576 -4201 -542
rect -4235 -644 -4201 -610
rect -4235 -712 -4201 -678
rect -4235 -780 -4201 -746
rect -4235 -848 -4201 -814
rect -4235 -916 -4201 -882
rect -4235 -984 -4201 -950
rect -4087 -168 -4053 -134
rect -4087 -236 -4053 -202
rect -4087 -304 -4053 -270
rect -4087 -372 -4053 -338
rect -4087 -440 -4053 -406
rect -4087 -508 -4053 -474
rect -4087 -576 -4053 -542
rect -4087 -644 -4053 -610
rect -4087 -712 -4053 -678
rect -4087 -780 -4053 -746
rect -4087 -848 -4053 -814
rect -4087 -916 -4053 -882
rect -4087 -984 -4053 -950
rect -3939 -168 -3905 -134
rect -3939 -236 -3905 -202
rect -3939 -304 -3905 -270
rect -3939 -372 -3905 -338
rect -3939 -440 -3905 -406
rect -3939 -508 -3905 -474
rect -3939 -576 -3905 -542
rect -3939 -644 -3905 -610
rect -3939 -712 -3905 -678
rect -3939 -780 -3905 -746
rect -3939 -848 -3905 -814
rect -3939 -916 -3905 -882
rect -3939 -984 -3905 -950
rect -3791 -168 -3757 -134
rect -3791 -236 -3757 -202
rect -3791 -304 -3757 -270
rect -3791 -372 -3757 -338
rect -3791 -440 -3757 -406
rect -3791 -508 -3757 -474
rect -3791 -576 -3757 -542
rect -3791 -644 -3757 -610
rect -3791 -712 -3757 -678
rect -3791 -780 -3757 -746
rect -3791 -848 -3757 -814
rect -3791 -916 -3757 -882
rect -3791 -984 -3757 -950
rect -3643 -168 -3609 -134
rect -3643 -236 -3609 -202
rect -3643 -304 -3609 -270
rect -3643 -372 -3609 -338
rect -3643 -440 -3609 -406
rect -3643 -508 -3609 -474
rect -3643 -576 -3609 -542
rect -3643 -644 -3609 -610
rect -3643 -712 -3609 -678
rect -3643 -780 -3609 -746
rect -3643 -848 -3609 -814
rect -3643 -916 -3609 -882
rect -3643 -984 -3609 -950
rect -3495 -168 -3461 -134
rect -3495 -236 -3461 -202
rect -3495 -304 -3461 -270
rect -3495 -372 -3461 -338
rect -3495 -440 -3461 -406
rect -3495 -508 -3461 -474
rect -3495 -576 -3461 -542
rect -3495 -644 -3461 -610
rect -3495 -712 -3461 -678
rect -3495 -780 -3461 -746
rect -3495 -848 -3461 -814
rect -3495 -916 -3461 -882
rect -3495 -984 -3461 -950
rect -3347 -168 -3313 -134
rect -3347 -236 -3313 -202
rect -3347 -304 -3313 -270
rect -3347 -372 -3313 -338
rect -3347 -440 -3313 -406
rect -3347 -508 -3313 -474
rect -3347 -576 -3313 -542
rect -3347 -644 -3313 -610
rect -3347 -712 -3313 -678
rect -3347 -780 -3313 -746
rect -3347 -848 -3313 -814
rect -3347 -916 -3313 -882
rect -3347 -984 -3313 -950
rect -3199 -168 -3165 -134
rect -3199 -236 -3165 -202
rect -3199 -304 -3165 -270
rect -3199 -372 -3165 -338
rect -3199 -440 -3165 -406
rect -3199 -508 -3165 -474
rect -3199 -576 -3165 -542
rect -3199 -644 -3165 -610
rect -3199 -712 -3165 -678
rect -3199 -780 -3165 -746
rect -3199 -848 -3165 -814
rect -3199 -916 -3165 -882
rect -3199 -984 -3165 -950
rect -3051 -168 -3017 -134
rect -3051 -236 -3017 -202
rect -3051 -304 -3017 -270
rect -3051 -372 -3017 -338
rect -3051 -440 -3017 -406
rect -3051 -508 -3017 -474
rect -3051 -576 -3017 -542
rect -3051 -644 -3017 -610
rect -3051 -712 -3017 -678
rect -3051 -780 -3017 -746
rect -3051 -848 -3017 -814
rect -3051 -916 -3017 -882
rect -3051 -984 -3017 -950
rect -2903 -168 -2869 -134
rect -2903 -236 -2869 -202
rect -2903 -304 -2869 -270
rect -2903 -372 -2869 -338
rect -2903 -440 -2869 -406
rect -2903 -508 -2869 -474
rect -2903 -576 -2869 -542
rect -2903 -644 -2869 -610
rect -2903 -712 -2869 -678
rect -2903 -780 -2869 -746
rect -2903 -848 -2869 -814
rect -2903 -916 -2869 -882
rect -2903 -984 -2869 -950
rect -2755 -168 -2721 -134
rect -2755 -236 -2721 -202
rect -2755 -304 -2721 -270
rect -2755 -372 -2721 -338
rect -2755 -440 -2721 -406
rect -2755 -508 -2721 -474
rect -2755 -576 -2721 -542
rect -2755 -644 -2721 -610
rect -2755 -712 -2721 -678
rect -2755 -780 -2721 -746
rect -2755 -848 -2721 -814
rect -2755 -916 -2721 -882
rect -2755 -984 -2721 -950
rect -2607 -168 -2573 -134
rect -2607 -236 -2573 -202
rect -2607 -304 -2573 -270
rect -2607 -372 -2573 -338
rect -2607 -440 -2573 -406
rect -2607 -508 -2573 -474
rect -2607 -576 -2573 -542
rect -2607 -644 -2573 -610
rect -2607 -712 -2573 -678
rect -2607 -780 -2573 -746
rect -2607 -848 -2573 -814
rect -2607 -916 -2573 -882
rect -2607 -984 -2573 -950
rect -2459 -168 -2425 -134
rect -2459 -236 -2425 -202
rect -2459 -304 -2425 -270
rect -2459 -372 -2425 -338
rect -2459 -440 -2425 -406
rect -2459 -508 -2425 -474
rect -2459 -576 -2425 -542
rect -2459 -644 -2425 -610
rect -2459 -712 -2425 -678
rect -2459 -780 -2425 -746
rect -2459 -848 -2425 -814
rect -2459 -916 -2425 -882
rect -2459 -984 -2425 -950
rect -2311 -168 -2277 -134
rect -2311 -236 -2277 -202
rect -2311 -304 -2277 -270
rect -2311 -372 -2277 -338
rect -2311 -440 -2277 -406
rect -2311 -508 -2277 -474
rect -2311 -576 -2277 -542
rect -2311 -644 -2277 -610
rect -2311 -712 -2277 -678
rect -2311 -780 -2277 -746
rect -2311 -848 -2277 -814
rect -2311 -916 -2277 -882
rect -2311 -984 -2277 -950
rect -2163 -168 -2129 -134
rect -2163 -236 -2129 -202
rect -2163 -304 -2129 -270
rect -2163 -372 -2129 -338
rect -2163 -440 -2129 -406
rect -2163 -508 -2129 -474
rect -2163 -576 -2129 -542
rect -2163 -644 -2129 -610
rect -2163 -712 -2129 -678
rect -2163 -780 -2129 -746
rect -2163 -848 -2129 -814
rect -2163 -916 -2129 -882
rect -2163 -984 -2129 -950
rect -2015 -168 -1981 -134
rect -2015 -236 -1981 -202
rect -2015 -304 -1981 -270
rect -2015 -372 -1981 -338
rect -2015 -440 -1981 -406
rect -2015 -508 -1981 -474
rect -2015 -576 -1981 -542
rect -2015 -644 -1981 -610
rect -2015 -712 -1981 -678
rect -2015 -780 -1981 -746
rect -2015 -848 -1981 -814
rect -2015 -916 -1981 -882
rect -2015 -984 -1981 -950
rect -1867 -168 -1833 -134
rect -1867 -236 -1833 -202
rect -1867 -304 -1833 -270
rect -1867 -372 -1833 -338
rect -1867 -440 -1833 -406
rect -1867 -508 -1833 -474
rect -1867 -576 -1833 -542
rect -1867 -644 -1833 -610
rect -1867 -712 -1833 -678
rect -1867 -780 -1833 -746
rect -1867 -848 -1833 -814
rect -1867 -916 -1833 -882
rect -1867 -984 -1833 -950
rect -1719 -168 -1685 -134
rect -1719 -236 -1685 -202
rect -1719 -304 -1685 -270
rect -1719 -372 -1685 -338
rect -1719 -440 -1685 -406
rect -1719 -508 -1685 -474
rect -1719 -576 -1685 -542
rect -1719 -644 -1685 -610
rect -1719 -712 -1685 -678
rect -1719 -780 -1685 -746
rect -1719 -848 -1685 -814
rect -1719 -916 -1685 -882
rect -1719 -984 -1685 -950
rect -1571 -168 -1537 -134
rect -1571 -236 -1537 -202
rect -1571 -304 -1537 -270
rect -1571 -372 -1537 -338
rect -1571 -440 -1537 -406
rect -1571 -508 -1537 -474
rect -1571 -576 -1537 -542
rect -1571 -644 -1537 -610
rect -1571 -712 -1537 -678
rect -1571 -780 -1537 -746
rect -1571 -848 -1537 -814
rect -1571 -916 -1537 -882
rect -1571 -984 -1537 -950
rect -1423 -168 -1389 -134
rect -1423 -236 -1389 -202
rect -1423 -304 -1389 -270
rect -1423 -372 -1389 -338
rect -1423 -440 -1389 -406
rect -1423 -508 -1389 -474
rect -1423 -576 -1389 -542
rect -1423 -644 -1389 -610
rect -1423 -712 -1389 -678
rect -1423 -780 -1389 -746
rect -1423 -848 -1389 -814
rect -1423 -916 -1389 -882
rect -1423 -984 -1389 -950
rect -1275 -168 -1241 -134
rect -1275 -236 -1241 -202
rect -1275 -304 -1241 -270
rect -1275 -372 -1241 -338
rect -1275 -440 -1241 -406
rect -1275 -508 -1241 -474
rect -1275 -576 -1241 -542
rect -1275 -644 -1241 -610
rect -1275 -712 -1241 -678
rect -1275 -780 -1241 -746
rect -1275 -848 -1241 -814
rect -1275 -916 -1241 -882
rect -1275 -984 -1241 -950
rect -1127 -168 -1093 -134
rect -1127 -236 -1093 -202
rect -1127 -304 -1093 -270
rect -1127 -372 -1093 -338
rect -1127 -440 -1093 -406
rect -1127 -508 -1093 -474
rect -1127 -576 -1093 -542
rect -1127 -644 -1093 -610
rect -1127 -712 -1093 -678
rect -1127 -780 -1093 -746
rect -1127 -848 -1093 -814
rect -1127 -916 -1093 -882
rect -1127 -984 -1093 -950
rect -979 -168 -945 -134
rect -979 -236 -945 -202
rect -979 -304 -945 -270
rect -979 -372 -945 -338
rect -979 -440 -945 -406
rect -979 -508 -945 -474
rect -979 -576 -945 -542
rect -979 -644 -945 -610
rect -979 -712 -945 -678
rect -979 -780 -945 -746
rect -979 -848 -945 -814
rect -979 -916 -945 -882
rect -979 -984 -945 -950
rect -831 -168 -797 -134
rect -831 -236 -797 -202
rect -831 -304 -797 -270
rect -831 -372 -797 -338
rect -831 -440 -797 -406
rect -831 -508 -797 -474
rect -831 -576 -797 -542
rect -831 -644 -797 -610
rect -831 -712 -797 -678
rect -831 -780 -797 -746
rect -831 -848 -797 -814
rect -831 -916 -797 -882
rect -831 -984 -797 -950
rect -683 -168 -649 -134
rect -683 -236 -649 -202
rect -683 -304 -649 -270
rect -683 -372 -649 -338
rect -683 -440 -649 -406
rect -683 -508 -649 -474
rect -683 -576 -649 -542
rect -683 -644 -649 -610
rect -683 -712 -649 -678
rect -683 -780 -649 -746
rect -683 -848 -649 -814
rect -683 -916 -649 -882
rect -683 -984 -649 -950
rect -535 -168 -501 -134
rect -535 -236 -501 -202
rect -535 -304 -501 -270
rect -535 -372 -501 -338
rect -535 -440 -501 -406
rect -535 -508 -501 -474
rect -535 -576 -501 -542
rect -535 -644 -501 -610
rect -535 -712 -501 -678
rect -535 -780 -501 -746
rect -535 -848 -501 -814
rect -535 -916 -501 -882
rect -535 -984 -501 -950
rect -387 -168 -353 -134
rect -387 -236 -353 -202
rect -387 -304 -353 -270
rect -387 -372 -353 -338
rect -387 -440 -353 -406
rect -387 -508 -353 -474
rect -387 -576 -353 -542
rect -387 -644 -353 -610
rect -387 -712 -353 -678
rect -387 -780 -353 -746
rect -387 -848 -353 -814
rect -387 -916 -353 -882
rect -387 -984 -353 -950
rect -239 -168 -205 -134
rect -239 -236 -205 -202
rect -239 -304 -205 -270
rect -239 -372 -205 -338
rect -239 -440 -205 -406
rect -239 -508 -205 -474
rect -239 -576 -205 -542
rect -239 -644 -205 -610
rect -239 -712 -205 -678
rect -239 -780 -205 -746
rect -239 -848 -205 -814
rect -239 -916 -205 -882
rect -239 -984 -205 -950
rect -91 -168 -57 -134
rect -91 -236 -57 -202
rect -91 -304 -57 -270
rect -91 -372 -57 -338
rect -91 -440 -57 -406
rect -91 -508 -57 -474
rect -91 -576 -57 -542
rect -91 -644 -57 -610
rect -91 -712 -57 -678
rect -91 -780 -57 -746
rect -91 -848 -57 -814
rect -91 -916 -57 -882
rect -91 -984 -57 -950
rect 57 -168 91 -134
rect 57 -236 91 -202
rect 57 -304 91 -270
rect 57 -372 91 -338
rect 57 -440 91 -406
rect 57 -508 91 -474
rect 57 -576 91 -542
rect 57 -644 91 -610
rect 57 -712 91 -678
rect 57 -780 91 -746
rect 57 -848 91 -814
rect 57 -916 91 -882
rect 57 -984 91 -950
rect 205 -168 239 -134
rect 205 -236 239 -202
rect 205 -304 239 -270
rect 205 -372 239 -338
rect 205 -440 239 -406
rect 205 -508 239 -474
rect 205 -576 239 -542
rect 205 -644 239 -610
rect 205 -712 239 -678
rect 205 -780 239 -746
rect 205 -848 239 -814
rect 205 -916 239 -882
rect 205 -984 239 -950
rect 353 -168 387 -134
rect 353 -236 387 -202
rect 353 -304 387 -270
rect 353 -372 387 -338
rect 353 -440 387 -406
rect 353 -508 387 -474
rect 353 -576 387 -542
rect 353 -644 387 -610
rect 353 -712 387 -678
rect 353 -780 387 -746
rect 353 -848 387 -814
rect 353 -916 387 -882
rect 353 -984 387 -950
rect 501 -168 535 -134
rect 501 -236 535 -202
rect 501 -304 535 -270
rect 501 -372 535 -338
rect 501 -440 535 -406
rect 501 -508 535 -474
rect 501 -576 535 -542
rect 501 -644 535 -610
rect 501 -712 535 -678
rect 501 -780 535 -746
rect 501 -848 535 -814
rect 501 -916 535 -882
rect 501 -984 535 -950
rect 649 -168 683 -134
rect 649 -236 683 -202
rect 649 -304 683 -270
rect 649 -372 683 -338
rect 649 -440 683 -406
rect 649 -508 683 -474
rect 649 -576 683 -542
rect 649 -644 683 -610
rect 649 -712 683 -678
rect 649 -780 683 -746
rect 649 -848 683 -814
rect 649 -916 683 -882
rect 649 -984 683 -950
rect 797 -168 831 -134
rect 797 -236 831 -202
rect 797 -304 831 -270
rect 797 -372 831 -338
rect 797 -440 831 -406
rect 797 -508 831 -474
rect 797 -576 831 -542
rect 797 -644 831 -610
rect 797 -712 831 -678
rect 797 -780 831 -746
rect 797 -848 831 -814
rect 797 -916 831 -882
rect 797 -984 831 -950
rect 945 -168 979 -134
rect 945 -236 979 -202
rect 945 -304 979 -270
rect 945 -372 979 -338
rect 945 -440 979 -406
rect 945 -508 979 -474
rect 945 -576 979 -542
rect 945 -644 979 -610
rect 945 -712 979 -678
rect 945 -780 979 -746
rect 945 -848 979 -814
rect 945 -916 979 -882
rect 945 -984 979 -950
rect 1093 -168 1127 -134
rect 1093 -236 1127 -202
rect 1093 -304 1127 -270
rect 1093 -372 1127 -338
rect 1093 -440 1127 -406
rect 1093 -508 1127 -474
rect 1093 -576 1127 -542
rect 1093 -644 1127 -610
rect 1093 -712 1127 -678
rect 1093 -780 1127 -746
rect 1093 -848 1127 -814
rect 1093 -916 1127 -882
rect 1093 -984 1127 -950
rect 1241 -168 1275 -134
rect 1241 -236 1275 -202
rect 1241 -304 1275 -270
rect 1241 -372 1275 -338
rect 1241 -440 1275 -406
rect 1241 -508 1275 -474
rect 1241 -576 1275 -542
rect 1241 -644 1275 -610
rect 1241 -712 1275 -678
rect 1241 -780 1275 -746
rect 1241 -848 1275 -814
rect 1241 -916 1275 -882
rect 1241 -984 1275 -950
rect 1389 -168 1423 -134
rect 1389 -236 1423 -202
rect 1389 -304 1423 -270
rect 1389 -372 1423 -338
rect 1389 -440 1423 -406
rect 1389 -508 1423 -474
rect 1389 -576 1423 -542
rect 1389 -644 1423 -610
rect 1389 -712 1423 -678
rect 1389 -780 1423 -746
rect 1389 -848 1423 -814
rect 1389 -916 1423 -882
rect 1389 -984 1423 -950
rect 1537 -168 1571 -134
rect 1537 -236 1571 -202
rect 1537 -304 1571 -270
rect 1537 -372 1571 -338
rect 1537 -440 1571 -406
rect 1537 -508 1571 -474
rect 1537 -576 1571 -542
rect 1537 -644 1571 -610
rect 1537 -712 1571 -678
rect 1537 -780 1571 -746
rect 1537 -848 1571 -814
rect 1537 -916 1571 -882
rect 1537 -984 1571 -950
rect 1685 -168 1719 -134
rect 1685 -236 1719 -202
rect 1685 -304 1719 -270
rect 1685 -372 1719 -338
rect 1685 -440 1719 -406
rect 1685 -508 1719 -474
rect 1685 -576 1719 -542
rect 1685 -644 1719 -610
rect 1685 -712 1719 -678
rect 1685 -780 1719 -746
rect 1685 -848 1719 -814
rect 1685 -916 1719 -882
rect 1685 -984 1719 -950
rect 1833 -168 1867 -134
rect 1833 -236 1867 -202
rect 1833 -304 1867 -270
rect 1833 -372 1867 -338
rect 1833 -440 1867 -406
rect 1833 -508 1867 -474
rect 1833 -576 1867 -542
rect 1833 -644 1867 -610
rect 1833 -712 1867 -678
rect 1833 -780 1867 -746
rect 1833 -848 1867 -814
rect 1833 -916 1867 -882
rect 1833 -984 1867 -950
rect 1981 -168 2015 -134
rect 1981 -236 2015 -202
rect 1981 -304 2015 -270
rect 1981 -372 2015 -338
rect 1981 -440 2015 -406
rect 1981 -508 2015 -474
rect 1981 -576 2015 -542
rect 1981 -644 2015 -610
rect 1981 -712 2015 -678
rect 1981 -780 2015 -746
rect 1981 -848 2015 -814
rect 1981 -916 2015 -882
rect 1981 -984 2015 -950
rect 2129 -168 2163 -134
rect 2129 -236 2163 -202
rect 2129 -304 2163 -270
rect 2129 -372 2163 -338
rect 2129 -440 2163 -406
rect 2129 -508 2163 -474
rect 2129 -576 2163 -542
rect 2129 -644 2163 -610
rect 2129 -712 2163 -678
rect 2129 -780 2163 -746
rect 2129 -848 2163 -814
rect 2129 -916 2163 -882
rect 2129 -984 2163 -950
rect 2277 -168 2311 -134
rect 2277 -236 2311 -202
rect 2277 -304 2311 -270
rect 2277 -372 2311 -338
rect 2277 -440 2311 -406
rect 2277 -508 2311 -474
rect 2277 -576 2311 -542
rect 2277 -644 2311 -610
rect 2277 -712 2311 -678
rect 2277 -780 2311 -746
rect 2277 -848 2311 -814
rect 2277 -916 2311 -882
rect 2277 -984 2311 -950
rect 2425 -168 2459 -134
rect 2425 -236 2459 -202
rect 2425 -304 2459 -270
rect 2425 -372 2459 -338
rect 2425 -440 2459 -406
rect 2425 -508 2459 -474
rect 2425 -576 2459 -542
rect 2425 -644 2459 -610
rect 2425 -712 2459 -678
rect 2425 -780 2459 -746
rect 2425 -848 2459 -814
rect 2425 -916 2459 -882
rect 2425 -984 2459 -950
rect 2573 -168 2607 -134
rect 2573 -236 2607 -202
rect 2573 -304 2607 -270
rect 2573 -372 2607 -338
rect 2573 -440 2607 -406
rect 2573 -508 2607 -474
rect 2573 -576 2607 -542
rect 2573 -644 2607 -610
rect 2573 -712 2607 -678
rect 2573 -780 2607 -746
rect 2573 -848 2607 -814
rect 2573 -916 2607 -882
rect 2573 -984 2607 -950
rect 2721 -168 2755 -134
rect 2721 -236 2755 -202
rect 2721 -304 2755 -270
rect 2721 -372 2755 -338
rect 2721 -440 2755 -406
rect 2721 -508 2755 -474
rect 2721 -576 2755 -542
rect 2721 -644 2755 -610
rect 2721 -712 2755 -678
rect 2721 -780 2755 -746
rect 2721 -848 2755 -814
rect 2721 -916 2755 -882
rect 2721 -984 2755 -950
rect 2869 -168 2903 -134
rect 2869 -236 2903 -202
rect 2869 -304 2903 -270
rect 2869 -372 2903 -338
rect 2869 -440 2903 -406
rect 2869 -508 2903 -474
rect 2869 -576 2903 -542
rect 2869 -644 2903 -610
rect 2869 -712 2903 -678
rect 2869 -780 2903 -746
rect 2869 -848 2903 -814
rect 2869 -916 2903 -882
rect 2869 -984 2903 -950
rect 3017 -168 3051 -134
rect 3017 -236 3051 -202
rect 3017 -304 3051 -270
rect 3017 -372 3051 -338
rect 3017 -440 3051 -406
rect 3017 -508 3051 -474
rect 3017 -576 3051 -542
rect 3017 -644 3051 -610
rect 3017 -712 3051 -678
rect 3017 -780 3051 -746
rect 3017 -848 3051 -814
rect 3017 -916 3051 -882
rect 3017 -984 3051 -950
rect 3165 -168 3199 -134
rect 3165 -236 3199 -202
rect 3165 -304 3199 -270
rect 3165 -372 3199 -338
rect 3165 -440 3199 -406
rect 3165 -508 3199 -474
rect 3165 -576 3199 -542
rect 3165 -644 3199 -610
rect 3165 -712 3199 -678
rect 3165 -780 3199 -746
rect 3165 -848 3199 -814
rect 3165 -916 3199 -882
rect 3165 -984 3199 -950
rect 3313 -168 3347 -134
rect 3313 -236 3347 -202
rect 3313 -304 3347 -270
rect 3313 -372 3347 -338
rect 3313 -440 3347 -406
rect 3313 -508 3347 -474
rect 3313 -576 3347 -542
rect 3313 -644 3347 -610
rect 3313 -712 3347 -678
rect 3313 -780 3347 -746
rect 3313 -848 3347 -814
rect 3313 -916 3347 -882
rect 3313 -984 3347 -950
rect 3461 -168 3495 -134
rect 3461 -236 3495 -202
rect 3461 -304 3495 -270
rect 3461 -372 3495 -338
rect 3461 -440 3495 -406
rect 3461 -508 3495 -474
rect 3461 -576 3495 -542
rect 3461 -644 3495 -610
rect 3461 -712 3495 -678
rect 3461 -780 3495 -746
rect 3461 -848 3495 -814
rect 3461 -916 3495 -882
rect 3461 -984 3495 -950
rect 3609 -168 3643 -134
rect 3609 -236 3643 -202
rect 3609 -304 3643 -270
rect 3609 -372 3643 -338
rect 3609 -440 3643 -406
rect 3609 -508 3643 -474
rect 3609 -576 3643 -542
rect 3609 -644 3643 -610
rect 3609 -712 3643 -678
rect 3609 -780 3643 -746
rect 3609 -848 3643 -814
rect 3609 -916 3643 -882
rect 3609 -984 3643 -950
rect 3757 -168 3791 -134
rect 3757 -236 3791 -202
rect 3757 -304 3791 -270
rect 3757 -372 3791 -338
rect 3757 -440 3791 -406
rect 3757 -508 3791 -474
rect 3757 -576 3791 -542
rect 3757 -644 3791 -610
rect 3757 -712 3791 -678
rect 3757 -780 3791 -746
rect 3757 -848 3791 -814
rect 3757 -916 3791 -882
rect 3757 -984 3791 -950
rect 3905 -168 3939 -134
rect 3905 -236 3939 -202
rect 3905 -304 3939 -270
rect 3905 -372 3939 -338
rect 3905 -440 3939 -406
rect 3905 -508 3939 -474
rect 3905 -576 3939 -542
rect 3905 -644 3939 -610
rect 3905 -712 3939 -678
rect 3905 -780 3939 -746
rect 3905 -848 3939 -814
rect 3905 -916 3939 -882
rect 3905 -984 3939 -950
rect 4053 -168 4087 -134
rect 4053 -236 4087 -202
rect 4053 -304 4087 -270
rect 4053 -372 4087 -338
rect 4053 -440 4087 -406
rect 4053 -508 4087 -474
rect 4053 -576 4087 -542
rect 4053 -644 4087 -610
rect 4053 -712 4087 -678
rect 4053 -780 4087 -746
rect 4053 -848 4087 -814
rect 4053 -916 4087 -882
rect 4053 -984 4087 -950
rect 4201 -168 4235 -134
rect 4201 -236 4235 -202
rect 4201 -304 4235 -270
rect 4201 -372 4235 -338
rect 4201 -440 4235 -406
rect 4201 -508 4235 -474
rect 4201 -576 4235 -542
rect 4201 -644 4235 -610
rect 4201 -712 4235 -678
rect 4201 -780 4235 -746
rect 4201 -848 4235 -814
rect 4201 -916 4235 -882
rect 4201 -984 4235 -950
rect 4349 -168 4383 -134
rect 4349 -236 4383 -202
rect 4349 -304 4383 -270
rect 4349 -372 4383 -338
rect 4349 -440 4383 -406
rect 4349 -508 4383 -474
rect 4349 -576 4383 -542
rect 4349 -644 4383 -610
rect 4349 -712 4383 -678
rect 4349 -780 4383 -746
rect 4349 -848 4383 -814
rect 4349 -916 4383 -882
rect 4349 -984 4383 -950
rect 4497 -168 4531 -134
rect 4497 -236 4531 -202
rect 4497 -304 4531 -270
rect 4497 -372 4531 -338
rect 4497 -440 4531 -406
rect 4497 -508 4531 -474
rect 4497 -576 4531 -542
rect 4497 -644 4531 -610
rect 4497 -712 4531 -678
rect 4497 -780 4531 -746
rect 4497 -848 4531 -814
rect 4497 -916 4531 -882
rect 4497 -984 4531 -950
rect 4645 -168 4679 -134
rect 4645 -236 4679 -202
rect 4645 -304 4679 -270
rect 4645 -372 4679 -338
rect 4645 -440 4679 -406
rect 4645 -508 4679 -474
rect 4645 -576 4679 -542
rect 4645 -644 4679 -610
rect 4645 -712 4679 -678
rect 4645 -780 4679 -746
rect 4645 -848 4679 -814
rect 4645 -916 4679 -882
rect 4645 -984 4679 -950
rect 4793 -168 4827 -134
rect 4793 -236 4827 -202
rect 4793 -304 4827 -270
rect 4793 -372 4827 -338
rect 4793 -440 4827 -406
rect 4793 -508 4827 -474
rect 4793 -576 4827 -542
rect 4793 -644 4827 -610
rect 4793 -712 4827 -678
rect 4793 -780 4827 -746
rect 4793 -848 4827 -814
rect 4793 -916 4827 -882
rect 4793 -984 4827 -950
rect 4941 -168 4975 -134
rect 4941 -236 4975 -202
rect 4941 -304 4975 -270
rect 4941 -372 4975 -338
rect 4941 -440 4975 -406
rect 4941 -508 4975 -474
rect 4941 -576 4975 -542
rect 4941 -644 4975 -610
rect 4941 -712 4975 -678
rect 4941 -780 4975 -746
rect 4941 -848 4975 -814
rect 4941 -916 4975 -882
rect 4941 -984 4975 -950
rect 5089 -168 5123 -134
rect 5089 -236 5123 -202
rect 5089 -304 5123 -270
rect 5089 -372 5123 -338
rect 5089 -440 5123 -406
rect 5089 -508 5123 -474
rect 5089 -576 5123 -542
rect 5089 -644 5123 -610
rect 5089 -712 5123 -678
rect 5089 -780 5123 -746
rect 5089 -848 5123 -814
rect 5089 -916 5123 -882
rect 5089 -984 5123 -950
rect 5237 -168 5271 -134
rect 5237 -236 5271 -202
rect 5237 -304 5271 -270
rect 5237 -372 5271 -338
rect 5237 -440 5271 -406
rect 5237 -508 5271 -474
rect 5237 -576 5271 -542
rect 5237 -644 5271 -610
rect 5237 -712 5271 -678
rect 5237 -780 5271 -746
rect 5237 -848 5271 -814
rect 5237 -916 5271 -882
rect 5237 -984 5271 -950
rect 5385 -168 5419 -134
rect 5385 -236 5419 -202
rect 5385 -304 5419 -270
rect 5385 -372 5419 -338
rect 5385 -440 5419 -406
rect 5385 -508 5419 -474
rect 5385 -576 5419 -542
rect 5385 -644 5419 -610
rect 5385 -712 5419 -678
rect 5385 -780 5419 -746
rect 5385 -848 5419 -814
rect 5385 -916 5419 -882
rect 5385 -984 5419 -950
rect 5533 -168 5567 -134
rect 5533 -236 5567 -202
rect 5533 -304 5567 -270
rect 5533 -372 5567 -338
rect 5533 -440 5567 -406
rect 5533 -508 5567 -474
rect 5533 -576 5567 -542
rect 5533 -644 5567 -610
rect 5533 -712 5567 -678
rect 5533 -780 5567 -746
rect 5533 -848 5567 -814
rect 5533 -916 5567 -882
rect 5533 -984 5567 -950
<< psubdiff >>
rect -5681 1149 -5559 1183
rect -5525 1149 -5491 1183
rect -5457 1149 -5423 1183
rect -5389 1149 -5355 1183
rect -5321 1149 -5287 1183
rect -5253 1149 -5219 1183
rect -5185 1149 -5151 1183
rect -5117 1149 -5083 1183
rect -5049 1149 -5015 1183
rect -4981 1149 -4947 1183
rect -4913 1149 -4879 1183
rect -4845 1149 -4811 1183
rect -4777 1149 -4743 1183
rect -4709 1149 -4675 1183
rect -4641 1149 -4607 1183
rect -4573 1149 -4539 1183
rect -4505 1149 -4471 1183
rect -4437 1149 -4403 1183
rect -4369 1149 -4335 1183
rect -4301 1149 -4267 1183
rect -4233 1149 -4199 1183
rect -4165 1149 -4131 1183
rect -4097 1149 -4063 1183
rect -4029 1149 -3995 1183
rect -3961 1149 -3927 1183
rect -3893 1149 -3859 1183
rect -3825 1149 -3791 1183
rect -3757 1149 -3723 1183
rect -3689 1149 -3655 1183
rect -3621 1149 -3587 1183
rect -3553 1149 -3519 1183
rect -3485 1149 -3451 1183
rect -3417 1149 -3383 1183
rect -3349 1149 -3315 1183
rect -3281 1149 -3247 1183
rect -3213 1149 -3179 1183
rect -3145 1149 -3111 1183
rect -3077 1149 -3043 1183
rect -3009 1149 -2975 1183
rect -2941 1149 -2907 1183
rect -2873 1149 -2839 1183
rect -2805 1149 -2771 1183
rect -2737 1149 -2703 1183
rect -2669 1149 -2635 1183
rect -2601 1149 -2567 1183
rect -2533 1149 -2499 1183
rect -2465 1149 -2431 1183
rect -2397 1149 -2363 1183
rect -2329 1149 -2295 1183
rect -2261 1149 -2227 1183
rect -2193 1149 -2159 1183
rect -2125 1149 -2091 1183
rect -2057 1149 -2023 1183
rect -1989 1149 -1955 1183
rect -1921 1149 -1887 1183
rect -1853 1149 -1819 1183
rect -1785 1149 -1751 1183
rect -1717 1149 -1683 1183
rect -1649 1149 -1615 1183
rect -1581 1149 -1547 1183
rect -1513 1149 -1479 1183
rect -1445 1149 -1411 1183
rect -1377 1149 -1343 1183
rect -1309 1149 -1275 1183
rect -1241 1149 -1207 1183
rect -1173 1149 -1139 1183
rect -1105 1149 -1071 1183
rect -1037 1149 -1003 1183
rect -969 1149 -935 1183
rect -901 1149 -867 1183
rect -833 1149 -799 1183
rect -765 1149 -731 1183
rect -697 1149 -663 1183
rect -629 1149 -595 1183
rect -561 1149 -527 1183
rect -493 1149 -459 1183
rect -425 1149 -391 1183
rect -357 1149 -323 1183
rect -289 1149 -255 1183
rect -221 1149 -187 1183
rect -153 1149 -119 1183
rect -85 1149 -51 1183
rect -17 1149 17 1183
rect 51 1149 85 1183
rect 119 1149 153 1183
rect 187 1149 221 1183
rect 255 1149 289 1183
rect 323 1149 357 1183
rect 391 1149 425 1183
rect 459 1149 493 1183
rect 527 1149 561 1183
rect 595 1149 629 1183
rect 663 1149 697 1183
rect 731 1149 765 1183
rect 799 1149 833 1183
rect 867 1149 901 1183
rect 935 1149 969 1183
rect 1003 1149 1037 1183
rect 1071 1149 1105 1183
rect 1139 1149 1173 1183
rect 1207 1149 1241 1183
rect 1275 1149 1309 1183
rect 1343 1149 1377 1183
rect 1411 1149 1445 1183
rect 1479 1149 1513 1183
rect 1547 1149 1581 1183
rect 1615 1149 1649 1183
rect 1683 1149 1717 1183
rect 1751 1149 1785 1183
rect 1819 1149 1853 1183
rect 1887 1149 1921 1183
rect 1955 1149 1989 1183
rect 2023 1149 2057 1183
rect 2091 1149 2125 1183
rect 2159 1149 2193 1183
rect 2227 1149 2261 1183
rect 2295 1149 2329 1183
rect 2363 1149 2397 1183
rect 2431 1149 2465 1183
rect 2499 1149 2533 1183
rect 2567 1149 2601 1183
rect 2635 1149 2669 1183
rect 2703 1149 2737 1183
rect 2771 1149 2805 1183
rect 2839 1149 2873 1183
rect 2907 1149 2941 1183
rect 2975 1149 3009 1183
rect 3043 1149 3077 1183
rect 3111 1149 3145 1183
rect 3179 1149 3213 1183
rect 3247 1149 3281 1183
rect 3315 1149 3349 1183
rect 3383 1149 3417 1183
rect 3451 1149 3485 1183
rect 3519 1149 3553 1183
rect 3587 1149 3621 1183
rect 3655 1149 3689 1183
rect 3723 1149 3757 1183
rect 3791 1149 3825 1183
rect 3859 1149 3893 1183
rect 3927 1149 3961 1183
rect 3995 1149 4029 1183
rect 4063 1149 4097 1183
rect 4131 1149 4165 1183
rect 4199 1149 4233 1183
rect 4267 1149 4301 1183
rect 4335 1149 4369 1183
rect 4403 1149 4437 1183
rect 4471 1149 4505 1183
rect 4539 1149 4573 1183
rect 4607 1149 4641 1183
rect 4675 1149 4709 1183
rect 4743 1149 4777 1183
rect 4811 1149 4845 1183
rect 4879 1149 4913 1183
rect 4947 1149 4981 1183
rect 5015 1149 5049 1183
rect 5083 1149 5117 1183
rect 5151 1149 5185 1183
rect 5219 1149 5253 1183
rect 5287 1149 5321 1183
rect 5355 1149 5389 1183
rect 5423 1149 5457 1183
rect 5491 1149 5525 1183
rect 5559 1149 5681 1183
rect -5681 1071 -5647 1149
rect -5681 1003 -5647 1037
rect 5647 1071 5681 1149
rect -5681 935 -5647 969
rect -5681 867 -5647 901
rect -5681 799 -5647 833
rect -5681 731 -5647 765
rect -5681 663 -5647 697
rect -5681 595 -5647 629
rect -5681 527 -5647 561
rect -5681 459 -5647 493
rect -5681 391 -5647 425
rect -5681 323 -5647 357
rect -5681 255 -5647 289
rect -5681 187 -5647 221
rect -5681 119 -5647 153
rect 5647 1003 5681 1037
rect 5647 935 5681 969
rect 5647 867 5681 901
rect 5647 799 5681 833
rect 5647 731 5681 765
rect 5647 663 5681 697
rect 5647 595 5681 629
rect 5647 527 5681 561
rect 5647 459 5681 493
rect 5647 391 5681 425
rect 5647 323 5681 357
rect 5647 255 5681 289
rect 5647 187 5681 221
rect 5647 119 5681 153
rect -5681 51 -5647 85
rect 5647 51 5681 85
rect -5681 -17 -5647 17
rect 5647 -17 5681 17
rect -5681 -85 -5647 -51
rect 5647 -85 5681 -51
rect -5681 -153 -5647 -119
rect -5681 -221 -5647 -187
rect -5681 -289 -5647 -255
rect -5681 -357 -5647 -323
rect -5681 -425 -5647 -391
rect -5681 -493 -5647 -459
rect -5681 -561 -5647 -527
rect -5681 -629 -5647 -595
rect -5681 -697 -5647 -663
rect -5681 -765 -5647 -731
rect -5681 -833 -5647 -799
rect -5681 -901 -5647 -867
rect -5681 -969 -5647 -935
rect -5681 -1037 -5647 -1003
rect 5647 -153 5681 -119
rect 5647 -221 5681 -187
rect 5647 -289 5681 -255
rect 5647 -357 5681 -323
rect 5647 -425 5681 -391
rect 5647 -493 5681 -459
rect 5647 -561 5681 -527
rect 5647 -629 5681 -595
rect 5647 -697 5681 -663
rect 5647 -765 5681 -731
rect 5647 -833 5681 -799
rect 5647 -901 5681 -867
rect 5647 -969 5681 -935
rect -5681 -1149 -5647 -1071
rect 5647 -1037 5681 -1003
rect 5647 -1149 5681 -1071
rect -5681 -1183 -5559 -1149
rect -5525 -1183 -5491 -1149
rect -5457 -1183 -5423 -1149
rect -5389 -1183 -5355 -1149
rect -5321 -1183 -5287 -1149
rect -5253 -1183 -5219 -1149
rect -5185 -1183 -5151 -1149
rect -5117 -1183 -5083 -1149
rect -5049 -1183 -5015 -1149
rect -4981 -1183 -4947 -1149
rect -4913 -1183 -4879 -1149
rect -4845 -1183 -4811 -1149
rect -4777 -1183 -4743 -1149
rect -4709 -1183 -4675 -1149
rect -4641 -1183 -4607 -1149
rect -4573 -1183 -4539 -1149
rect -4505 -1183 -4471 -1149
rect -4437 -1183 -4403 -1149
rect -4369 -1183 -4335 -1149
rect -4301 -1183 -4267 -1149
rect -4233 -1183 -4199 -1149
rect -4165 -1183 -4131 -1149
rect -4097 -1183 -4063 -1149
rect -4029 -1183 -3995 -1149
rect -3961 -1183 -3927 -1149
rect -3893 -1183 -3859 -1149
rect -3825 -1183 -3791 -1149
rect -3757 -1183 -3723 -1149
rect -3689 -1183 -3655 -1149
rect -3621 -1183 -3587 -1149
rect -3553 -1183 -3519 -1149
rect -3485 -1183 -3451 -1149
rect -3417 -1183 -3383 -1149
rect -3349 -1183 -3315 -1149
rect -3281 -1183 -3247 -1149
rect -3213 -1183 -3179 -1149
rect -3145 -1183 -3111 -1149
rect -3077 -1183 -3043 -1149
rect -3009 -1183 -2975 -1149
rect -2941 -1183 -2907 -1149
rect -2873 -1183 -2839 -1149
rect -2805 -1183 -2771 -1149
rect -2737 -1183 -2703 -1149
rect -2669 -1183 -2635 -1149
rect -2601 -1183 -2567 -1149
rect -2533 -1183 -2499 -1149
rect -2465 -1183 -2431 -1149
rect -2397 -1183 -2363 -1149
rect -2329 -1183 -2295 -1149
rect -2261 -1183 -2227 -1149
rect -2193 -1183 -2159 -1149
rect -2125 -1183 -2091 -1149
rect -2057 -1183 -2023 -1149
rect -1989 -1183 -1955 -1149
rect -1921 -1183 -1887 -1149
rect -1853 -1183 -1819 -1149
rect -1785 -1183 -1751 -1149
rect -1717 -1183 -1683 -1149
rect -1649 -1183 -1615 -1149
rect -1581 -1183 -1547 -1149
rect -1513 -1183 -1479 -1149
rect -1445 -1183 -1411 -1149
rect -1377 -1183 -1343 -1149
rect -1309 -1183 -1275 -1149
rect -1241 -1183 -1207 -1149
rect -1173 -1183 -1139 -1149
rect -1105 -1183 -1071 -1149
rect -1037 -1183 -1003 -1149
rect -969 -1183 -935 -1149
rect -901 -1183 -867 -1149
rect -833 -1183 -799 -1149
rect -765 -1183 -731 -1149
rect -697 -1183 -663 -1149
rect -629 -1183 -595 -1149
rect -561 -1183 -527 -1149
rect -493 -1183 -459 -1149
rect -425 -1183 -391 -1149
rect -357 -1183 -323 -1149
rect -289 -1183 -255 -1149
rect -221 -1183 -187 -1149
rect -153 -1183 -119 -1149
rect -85 -1183 -51 -1149
rect -17 -1183 17 -1149
rect 51 -1183 85 -1149
rect 119 -1183 153 -1149
rect 187 -1183 221 -1149
rect 255 -1183 289 -1149
rect 323 -1183 357 -1149
rect 391 -1183 425 -1149
rect 459 -1183 493 -1149
rect 527 -1183 561 -1149
rect 595 -1183 629 -1149
rect 663 -1183 697 -1149
rect 731 -1183 765 -1149
rect 799 -1183 833 -1149
rect 867 -1183 901 -1149
rect 935 -1183 969 -1149
rect 1003 -1183 1037 -1149
rect 1071 -1183 1105 -1149
rect 1139 -1183 1173 -1149
rect 1207 -1183 1241 -1149
rect 1275 -1183 1309 -1149
rect 1343 -1183 1377 -1149
rect 1411 -1183 1445 -1149
rect 1479 -1183 1513 -1149
rect 1547 -1183 1581 -1149
rect 1615 -1183 1649 -1149
rect 1683 -1183 1717 -1149
rect 1751 -1183 1785 -1149
rect 1819 -1183 1853 -1149
rect 1887 -1183 1921 -1149
rect 1955 -1183 1989 -1149
rect 2023 -1183 2057 -1149
rect 2091 -1183 2125 -1149
rect 2159 -1183 2193 -1149
rect 2227 -1183 2261 -1149
rect 2295 -1183 2329 -1149
rect 2363 -1183 2397 -1149
rect 2431 -1183 2465 -1149
rect 2499 -1183 2533 -1149
rect 2567 -1183 2601 -1149
rect 2635 -1183 2669 -1149
rect 2703 -1183 2737 -1149
rect 2771 -1183 2805 -1149
rect 2839 -1183 2873 -1149
rect 2907 -1183 2941 -1149
rect 2975 -1183 3009 -1149
rect 3043 -1183 3077 -1149
rect 3111 -1183 3145 -1149
rect 3179 -1183 3213 -1149
rect 3247 -1183 3281 -1149
rect 3315 -1183 3349 -1149
rect 3383 -1183 3417 -1149
rect 3451 -1183 3485 -1149
rect 3519 -1183 3553 -1149
rect 3587 -1183 3621 -1149
rect 3655 -1183 3689 -1149
rect 3723 -1183 3757 -1149
rect 3791 -1183 3825 -1149
rect 3859 -1183 3893 -1149
rect 3927 -1183 3961 -1149
rect 3995 -1183 4029 -1149
rect 4063 -1183 4097 -1149
rect 4131 -1183 4165 -1149
rect 4199 -1183 4233 -1149
rect 4267 -1183 4301 -1149
rect 4335 -1183 4369 -1149
rect 4403 -1183 4437 -1149
rect 4471 -1183 4505 -1149
rect 4539 -1183 4573 -1149
rect 4607 -1183 4641 -1149
rect 4675 -1183 4709 -1149
rect 4743 -1183 4777 -1149
rect 4811 -1183 4845 -1149
rect 4879 -1183 4913 -1149
rect 4947 -1183 4981 -1149
rect 5015 -1183 5049 -1149
rect 5083 -1183 5117 -1149
rect 5151 -1183 5185 -1149
rect 5219 -1183 5253 -1149
rect 5287 -1183 5321 -1149
rect 5355 -1183 5389 -1149
rect 5423 -1183 5457 -1149
rect 5491 -1183 5525 -1149
rect 5559 -1183 5681 -1149
<< psubdiffcont >>
rect -5559 1149 -5525 1183
rect -5491 1149 -5457 1183
rect -5423 1149 -5389 1183
rect -5355 1149 -5321 1183
rect -5287 1149 -5253 1183
rect -5219 1149 -5185 1183
rect -5151 1149 -5117 1183
rect -5083 1149 -5049 1183
rect -5015 1149 -4981 1183
rect -4947 1149 -4913 1183
rect -4879 1149 -4845 1183
rect -4811 1149 -4777 1183
rect -4743 1149 -4709 1183
rect -4675 1149 -4641 1183
rect -4607 1149 -4573 1183
rect -4539 1149 -4505 1183
rect -4471 1149 -4437 1183
rect -4403 1149 -4369 1183
rect -4335 1149 -4301 1183
rect -4267 1149 -4233 1183
rect -4199 1149 -4165 1183
rect -4131 1149 -4097 1183
rect -4063 1149 -4029 1183
rect -3995 1149 -3961 1183
rect -3927 1149 -3893 1183
rect -3859 1149 -3825 1183
rect -3791 1149 -3757 1183
rect -3723 1149 -3689 1183
rect -3655 1149 -3621 1183
rect -3587 1149 -3553 1183
rect -3519 1149 -3485 1183
rect -3451 1149 -3417 1183
rect -3383 1149 -3349 1183
rect -3315 1149 -3281 1183
rect -3247 1149 -3213 1183
rect -3179 1149 -3145 1183
rect -3111 1149 -3077 1183
rect -3043 1149 -3009 1183
rect -2975 1149 -2941 1183
rect -2907 1149 -2873 1183
rect -2839 1149 -2805 1183
rect -2771 1149 -2737 1183
rect -2703 1149 -2669 1183
rect -2635 1149 -2601 1183
rect -2567 1149 -2533 1183
rect -2499 1149 -2465 1183
rect -2431 1149 -2397 1183
rect -2363 1149 -2329 1183
rect -2295 1149 -2261 1183
rect -2227 1149 -2193 1183
rect -2159 1149 -2125 1183
rect -2091 1149 -2057 1183
rect -2023 1149 -1989 1183
rect -1955 1149 -1921 1183
rect -1887 1149 -1853 1183
rect -1819 1149 -1785 1183
rect -1751 1149 -1717 1183
rect -1683 1149 -1649 1183
rect -1615 1149 -1581 1183
rect -1547 1149 -1513 1183
rect -1479 1149 -1445 1183
rect -1411 1149 -1377 1183
rect -1343 1149 -1309 1183
rect -1275 1149 -1241 1183
rect -1207 1149 -1173 1183
rect -1139 1149 -1105 1183
rect -1071 1149 -1037 1183
rect -1003 1149 -969 1183
rect -935 1149 -901 1183
rect -867 1149 -833 1183
rect -799 1149 -765 1183
rect -731 1149 -697 1183
rect -663 1149 -629 1183
rect -595 1149 -561 1183
rect -527 1149 -493 1183
rect -459 1149 -425 1183
rect -391 1149 -357 1183
rect -323 1149 -289 1183
rect -255 1149 -221 1183
rect -187 1149 -153 1183
rect -119 1149 -85 1183
rect -51 1149 -17 1183
rect 17 1149 51 1183
rect 85 1149 119 1183
rect 153 1149 187 1183
rect 221 1149 255 1183
rect 289 1149 323 1183
rect 357 1149 391 1183
rect 425 1149 459 1183
rect 493 1149 527 1183
rect 561 1149 595 1183
rect 629 1149 663 1183
rect 697 1149 731 1183
rect 765 1149 799 1183
rect 833 1149 867 1183
rect 901 1149 935 1183
rect 969 1149 1003 1183
rect 1037 1149 1071 1183
rect 1105 1149 1139 1183
rect 1173 1149 1207 1183
rect 1241 1149 1275 1183
rect 1309 1149 1343 1183
rect 1377 1149 1411 1183
rect 1445 1149 1479 1183
rect 1513 1149 1547 1183
rect 1581 1149 1615 1183
rect 1649 1149 1683 1183
rect 1717 1149 1751 1183
rect 1785 1149 1819 1183
rect 1853 1149 1887 1183
rect 1921 1149 1955 1183
rect 1989 1149 2023 1183
rect 2057 1149 2091 1183
rect 2125 1149 2159 1183
rect 2193 1149 2227 1183
rect 2261 1149 2295 1183
rect 2329 1149 2363 1183
rect 2397 1149 2431 1183
rect 2465 1149 2499 1183
rect 2533 1149 2567 1183
rect 2601 1149 2635 1183
rect 2669 1149 2703 1183
rect 2737 1149 2771 1183
rect 2805 1149 2839 1183
rect 2873 1149 2907 1183
rect 2941 1149 2975 1183
rect 3009 1149 3043 1183
rect 3077 1149 3111 1183
rect 3145 1149 3179 1183
rect 3213 1149 3247 1183
rect 3281 1149 3315 1183
rect 3349 1149 3383 1183
rect 3417 1149 3451 1183
rect 3485 1149 3519 1183
rect 3553 1149 3587 1183
rect 3621 1149 3655 1183
rect 3689 1149 3723 1183
rect 3757 1149 3791 1183
rect 3825 1149 3859 1183
rect 3893 1149 3927 1183
rect 3961 1149 3995 1183
rect 4029 1149 4063 1183
rect 4097 1149 4131 1183
rect 4165 1149 4199 1183
rect 4233 1149 4267 1183
rect 4301 1149 4335 1183
rect 4369 1149 4403 1183
rect 4437 1149 4471 1183
rect 4505 1149 4539 1183
rect 4573 1149 4607 1183
rect 4641 1149 4675 1183
rect 4709 1149 4743 1183
rect 4777 1149 4811 1183
rect 4845 1149 4879 1183
rect 4913 1149 4947 1183
rect 4981 1149 5015 1183
rect 5049 1149 5083 1183
rect 5117 1149 5151 1183
rect 5185 1149 5219 1183
rect 5253 1149 5287 1183
rect 5321 1149 5355 1183
rect 5389 1149 5423 1183
rect 5457 1149 5491 1183
rect 5525 1149 5559 1183
rect -5681 1037 -5647 1071
rect 5647 1037 5681 1071
rect -5681 969 -5647 1003
rect -5681 901 -5647 935
rect -5681 833 -5647 867
rect -5681 765 -5647 799
rect -5681 697 -5647 731
rect -5681 629 -5647 663
rect -5681 561 -5647 595
rect -5681 493 -5647 527
rect -5681 425 -5647 459
rect -5681 357 -5647 391
rect -5681 289 -5647 323
rect -5681 221 -5647 255
rect -5681 153 -5647 187
rect -5681 85 -5647 119
rect 5647 969 5681 1003
rect 5647 901 5681 935
rect 5647 833 5681 867
rect 5647 765 5681 799
rect 5647 697 5681 731
rect 5647 629 5681 663
rect 5647 561 5681 595
rect 5647 493 5681 527
rect 5647 425 5681 459
rect 5647 357 5681 391
rect 5647 289 5681 323
rect 5647 221 5681 255
rect 5647 153 5681 187
rect -5681 17 -5647 51
rect 5647 85 5681 119
rect -5681 -51 -5647 -17
rect 5647 17 5681 51
rect -5681 -119 -5647 -85
rect 5647 -51 5681 -17
rect -5681 -187 -5647 -153
rect -5681 -255 -5647 -221
rect -5681 -323 -5647 -289
rect -5681 -391 -5647 -357
rect -5681 -459 -5647 -425
rect -5681 -527 -5647 -493
rect -5681 -595 -5647 -561
rect -5681 -663 -5647 -629
rect -5681 -731 -5647 -697
rect -5681 -799 -5647 -765
rect -5681 -867 -5647 -833
rect -5681 -935 -5647 -901
rect -5681 -1003 -5647 -969
rect 5647 -119 5681 -85
rect 5647 -187 5681 -153
rect 5647 -255 5681 -221
rect 5647 -323 5681 -289
rect 5647 -391 5681 -357
rect 5647 -459 5681 -425
rect 5647 -527 5681 -493
rect 5647 -595 5681 -561
rect 5647 -663 5681 -629
rect 5647 -731 5681 -697
rect 5647 -799 5681 -765
rect 5647 -867 5681 -833
rect 5647 -935 5681 -901
rect 5647 -1003 5681 -969
rect -5681 -1071 -5647 -1037
rect 5647 -1071 5681 -1037
rect -5559 -1183 -5525 -1149
rect -5491 -1183 -5457 -1149
rect -5423 -1183 -5389 -1149
rect -5355 -1183 -5321 -1149
rect -5287 -1183 -5253 -1149
rect -5219 -1183 -5185 -1149
rect -5151 -1183 -5117 -1149
rect -5083 -1183 -5049 -1149
rect -5015 -1183 -4981 -1149
rect -4947 -1183 -4913 -1149
rect -4879 -1183 -4845 -1149
rect -4811 -1183 -4777 -1149
rect -4743 -1183 -4709 -1149
rect -4675 -1183 -4641 -1149
rect -4607 -1183 -4573 -1149
rect -4539 -1183 -4505 -1149
rect -4471 -1183 -4437 -1149
rect -4403 -1183 -4369 -1149
rect -4335 -1183 -4301 -1149
rect -4267 -1183 -4233 -1149
rect -4199 -1183 -4165 -1149
rect -4131 -1183 -4097 -1149
rect -4063 -1183 -4029 -1149
rect -3995 -1183 -3961 -1149
rect -3927 -1183 -3893 -1149
rect -3859 -1183 -3825 -1149
rect -3791 -1183 -3757 -1149
rect -3723 -1183 -3689 -1149
rect -3655 -1183 -3621 -1149
rect -3587 -1183 -3553 -1149
rect -3519 -1183 -3485 -1149
rect -3451 -1183 -3417 -1149
rect -3383 -1183 -3349 -1149
rect -3315 -1183 -3281 -1149
rect -3247 -1183 -3213 -1149
rect -3179 -1183 -3145 -1149
rect -3111 -1183 -3077 -1149
rect -3043 -1183 -3009 -1149
rect -2975 -1183 -2941 -1149
rect -2907 -1183 -2873 -1149
rect -2839 -1183 -2805 -1149
rect -2771 -1183 -2737 -1149
rect -2703 -1183 -2669 -1149
rect -2635 -1183 -2601 -1149
rect -2567 -1183 -2533 -1149
rect -2499 -1183 -2465 -1149
rect -2431 -1183 -2397 -1149
rect -2363 -1183 -2329 -1149
rect -2295 -1183 -2261 -1149
rect -2227 -1183 -2193 -1149
rect -2159 -1183 -2125 -1149
rect -2091 -1183 -2057 -1149
rect -2023 -1183 -1989 -1149
rect -1955 -1183 -1921 -1149
rect -1887 -1183 -1853 -1149
rect -1819 -1183 -1785 -1149
rect -1751 -1183 -1717 -1149
rect -1683 -1183 -1649 -1149
rect -1615 -1183 -1581 -1149
rect -1547 -1183 -1513 -1149
rect -1479 -1183 -1445 -1149
rect -1411 -1183 -1377 -1149
rect -1343 -1183 -1309 -1149
rect -1275 -1183 -1241 -1149
rect -1207 -1183 -1173 -1149
rect -1139 -1183 -1105 -1149
rect -1071 -1183 -1037 -1149
rect -1003 -1183 -969 -1149
rect -935 -1183 -901 -1149
rect -867 -1183 -833 -1149
rect -799 -1183 -765 -1149
rect -731 -1183 -697 -1149
rect -663 -1183 -629 -1149
rect -595 -1183 -561 -1149
rect -527 -1183 -493 -1149
rect -459 -1183 -425 -1149
rect -391 -1183 -357 -1149
rect -323 -1183 -289 -1149
rect -255 -1183 -221 -1149
rect -187 -1183 -153 -1149
rect -119 -1183 -85 -1149
rect -51 -1183 -17 -1149
rect 17 -1183 51 -1149
rect 85 -1183 119 -1149
rect 153 -1183 187 -1149
rect 221 -1183 255 -1149
rect 289 -1183 323 -1149
rect 357 -1183 391 -1149
rect 425 -1183 459 -1149
rect 493 -1183 527 -1149
rect 561 -1183 595 -1149
rect 629 -1183 663 -1149
rect 697 -1183 731 -1149
rect 765 -1183 799 -1149
rect 833 -1183 867 -1149
rect 901 -1183 935 -1149
rect 969 -1183 1003 -1149
rect 1037 -1183 1071 -1149
rect 1105 -1183 1139 -1149
rect 1173 -1183 1207 -1149
rect 1241 -1183 1275 -1149
rect 1309 -1183 1343 -1149
rect 1377 -1183 1411 -1149
rect 1445 -1183 1479 -1149
rect 1513 -1183 1547 -1149
rect 1581 -1183 1615 -1149
rect 1649 -1183 1683 -1149
rect 1717 -1183 1751 -1149
rect 1785 -1183 1819 -1149
rect 1853 -1183 1887 -1149
rect 1921 -1183 1955 -1149
rect 1989 -1183 2023 -1149
rect 2057 -1183 2091 -1149
rect 2125 -1183 2159 -1149
rect 2193 -1183 2227 -1149
rect 2261 -1183 2295 -1149
rect 2329 -1183 2363 -1149
rect 2397 -1183 2431 -1149
rect 2465 -1183 2499 -1149
rect 2533 -1183 2567 -1149
rect 2601 -1183 2635 -1149
rect 2669 -1183 2703 -1149
rect 2737 -1183 2771 -1149
rect 2805 -1183 2839 -1149
rect 2873 -1183 2907 -1149
rect 2941 -1183 2975 -1149
rect 3009 -1183 3043 -1149
rect 3077 -1183 3111 -1149
rect 3145 -1183 3179 -1149
rect 3213 -1183 3247 -1149
rect 3281 -1183 3315 -1149
rect 3349 -1183 3383 -1149
rect 3417 -1183 3451 -1149
rect 3485 -1183 3519 -1149
rect 3553 -1183 3587 -1149
rect 3621 -1183 3655 -1149
rect 3689 -1183 3723 -1149
rect 3757 -1183 3791 -1149
rect 3825 -1183 3859 -1149
rect 3893 -1183 3927 -1149
rect 3961 -1183 3995 -1149
rect 4029 -1183 4063 -1149
rect 4097 -1183 4131 -1149
rect 4165 -1183 4199 -1149
rect 4233 -1183 4267 -1149
rect 4301 -1183 4335 -1149
rect 4369 -1183 4403 -1149
rect 4437 -1183 4471 -1149
rect 4505 -1183 4539 -1149
rect 4573 -1183 4607 -1149
rect 4641 -1183 4675 -1149
rect 4709 -1183 4743 -1149
rect 4777 -1183 4811 -1149
rect 4845 -1183 4879 -1149
rect 4913 -1183 4947 -1149
rect 4981 -1183 5015 -1149
rect 5049 -1183 5083 -1149
rect 5117 -1183 5151 -1149
rect 5185 -1183 5219 -1149
rect 5253 -1183 5287 -1149
rect 5321 -1183 5355 -1149
rect 5389 -1183 5423 -1149
rect 5457 -1183 5491 -1149
rect 5525 -1183 5559 -1149
<< poly >>
rect -5521 1081 -5431 1097
rect -5521 1047 -5493 1081
rect -5459 1047 -5431 1081
rect -5521 1009 -5431 1047
rect -5373 1081 -5283 1097
rect -5373 1047 -5345 1081
rect -5311 1047 -5283 1081
rect -5373 1009 -5283 1047
rect -5225 1081 -5135 1097
rect -5225 1047 -5197 1081
rect -5163 1047 -5135 1081
rect -5225 1009 -5135 1047
rect -5077 1081 -4987 1097
rect -5077 1047 -5049 1081
rect -5015 1047 -4987 1081
rect -5077 1009 -4987 1047
rect -4929 1081 -4839 1097
rect -4929 1047 -4901 1081
rect -4867 1047 -4839 1081
rect -4929 1009 -4839 1047
rect -4781 1081 -4691 1097
rect -4781 1047 -4753 1081
rect -4719 1047 -4691 1081
rect -4781 1009 -4691 1047
rect -4633 1081 -4543 1097
rect -4633 1047 -4605 1081
rect -4571 1047 -4543 1081
rect -4633 1009 -4543 1047
rect -4485 1081 -4395 1097
rect -4485 1047 -4457 1081
rect -4423 1047 -4395 1081
rect -4485 1009 -4395 1047
rect -4337 1081 -4247 1097
rect -4337 1047 -4309 1081
rect -4275 1047 -4247 1081
rect -4337 1009 -4247 1047
rect -4189 1081 -4099 1097
rect -4189 1047 -4161 1081
rect -4127 1047 -4099 1081
rect -4189 1009 -4099 1047
rect -4041 1081 -3951 1097
rect -4041 1047 -4013 1081
rect -3979 1047 -3951 1081
rect -4041 1009 -3951 1047
rect -3893 1081 -3803 1097
rect -3893 1047 -3865 1081
rect -3831 1047 -3803 1081
rect -3893 1009 -3803 1047
rect -3745 1081 -3655 1097
rect -3745 1047 -3717 1081
rect -3683 1047 -3655 1081
rect -3745 1009 -3655 1047
rect -3597 1081 -3507 1097
rect -3597 1047 -3569 1081
rect -3535 1047 -3507 1081
rect -3597 1009 -3507 1047
rect -3449 1081 -3359 1097
rect -3449 1047 -3421 1081
rect -3387 1047 -3359 1081
rect -3449 1009 -3359 1047
rect -3301 1081 -3211 1097
rect -3301 1047 -3273 1081
rect -3239 1047 -3211 1081
rect -3301 1009 -3211 1047
rect -3153 1081 -3063 1097
rect -3153 1047 -3125 1081
rect -3091 1047 -3063 1081
rect -3153 1009 -3063 1047
rect -3005 1081 -2915 1097
rect -3005 1047 -2977 1081
rect -2943 1047 -2915 1081
rect -3005 1009 -2915 1047
rect -2857 1081 -2767 1097
rect -2857 1047 -2829 1081
rect -2795 1047 -2767 1081
rect -2857 1009 -2767 1047
rect -2709 1081 -2619 1097
rect -2709 1047 -2681 1081
rect -2647 1047 -2619 1081
rect -2709 1009 -2619 1047
rect -2561 1081 -2471 1097
rect -2561 1047 -2533 1081
rect -2499 1047 -2471 1081
rect -2561 1009 -2471 1047
rect -2413 1081 -2323 1097
rect -2413 1047 -2385 1081
rect -2351 1047 -2323 1081
rect -2413 1009 -2323 1047
rect -2265 1081 -2175 1097
rect -2265 1047 -2237 1081
rect -2203 1047 -2175 1081
rect -2265 1009 -2175 1047
rect -2117 1081 -2027 1097
rect -2117 1047 -2089 1081
rect -2055 1047 -2027 1081
rect -2117 1009 -2027 1047
rect -1969 1081 -1879 1097
rect -1969 1047 -1941 1081
rect -1907 1047 -1879 1081
rect -1969 1009 -1879 1047
rect -1821 1081 -1731 1097
rect -1821 1047 -1793 1081
rect -1759 1047 -1731 1081
rect -1821 1009 -1731 1047
rect -1673 1081 -1583 1097
rect -1673 1047 -1645 1081
rect -1611 1047 -1583 1081
rect -1673 1009 -1583 1047
rect -1525 1081 -1435 1097
rect -1525 1047 -1497 1081
rect -1463 1047 -1435 1081
rect -1525 1009 -1435 1047
rect -1377 1081 -1287 1097
rect -1377 1047 -1349 1081
rect -1315 1047 -1287 1081
rect -1377 1009 -1287 1047
rect -1229 1081 -1139 1097
rect -1229 1047 -1201 1081
rect -1167 1047 -1139 1081
rect -1229 1009 -1139 1047
rect -1081 1081 -991 1097
rect -1081 1047 -1053 1081
rect -1019 1047 -991 1081
rect -1081 1009 -991 1047
rect -933 1081 -843 1097
rect -933 1047 -905 1081
rect -871 1047 -843 1081
rect -933 1009 -843 1047
rect -785 1081 -695 1097
rect -785 1047 -757 1081
rect -723 1047 -695 1081
rect -785 1009 -695 1047
rect -637 1081 -547 1097
rect -637 1047 -609 1081
rect -575 1047 -547 1081
rect -637 1009 -547 1047
rect -489 1081 -399 1097
rect -489 1047 -461 1081
rect -427 1047 -399 1081
rect -489 1009 -399 1047
rect -341 1081 -251 1097
rect -341 1047 -313 1081
rect -279 1047 -251 1081
rect -341 1009 -251 1047
rect -193 1081 -103 1097
rect -193 1047 -165 1081
rect -131 1047 -103 1081
rect -193 1009 -103 1047
rect -45 1081 45 1097
rect -45 1047 -17 1081
rect 17 1047 45 1081
rect -45 1009 45 1047
rect 103 1081 193 1097
rect 103 1047 131 1081
rect 165 1047 193 1081
rect 103 1009 193 1047
rect 251 1081 341 1097
rect 251 1047 279 1081
rect 313 1047 341 1081
rect 251 1009 341 1047
rect 399 1081 489 1097
rect 399 1047 427 1081
rect 461 1047 489 1081
rect 399 1009 489 1047
rect 547 1081 637 1097
rect 547 1047 575 1081
rect 609 1047 637 1081
rect 547 1009 637 1047
rect 695 1081 785 1097
rect 695 1047 723 1081
rect 757 1047 785 1081
rect 695 1009 785 1047
rect 843 1081 933 1097
rect 843 1047 871 1081
rect 905 1047 933 1081
rect 843 1009 933 1047
rect 991 1081 1081 1097
rect 991 1047 1019 1081
rect 1053 1047 1081 1081
rect 991 1009 1081 1047
rect 1139 1081 1229 1097
rect 1139 1047 1167 1081
rect 1201 1047 1229 1081
rect 1139 1009 1229 1047
rect 1287 1081 1377 1097
rect 1287 1047 1315 1081
rect 1349 1047 1377 1081
rect 1287 1009 1377 1047
rect 1435 1081 1525 1097
rect 1435 1047 1463 1081
rect 1497 1047 1525 1081
rect 1435 1009 1525 1047
rect 1583 1081 1673 1097
rect 1583 1047 1611 1081
rect 1645 1047 1673 1081
rect 1583 1009 1673 1047
rect 1731 1081 1821 1097
rect 1731 1047 1759 1081
rect 1793 1047 1821 1081
rect 1731 1009 1821 1047
rect 1879 1081 1969 1097
rect 1879 1047 1907 1081
rect 1941 1047 1969 1081
rect 1879 1009 1969 1047
rect 2027 1081 2117 1097
rect 2027 1047 2055 1081
rect 2089 1047 2117 1081
rect 2027 1009 2117 1047
rect 2175 1081 2265 1097
rect 2175 1047 2203 1081
rect 2237 1047 2265 1081
rect 2175 1009 2265 1047
rect 2323 1081 2413 1097
rect 2323 1047 2351 1081
rect 2385 1047 2413 1081
rect 2323 1009 2413 1047
rect 2471 1081 2561 1097
rect 2471 1047 2499 1081
rect 2533 1047 2561 1081
rect 2471 1009 2561 1047
rect 2619 1081 2709 1097
rect 2619 1047 2647 1081
rect 2681 1047 2709 1081
rect 2619 1009 2709 1047
rect 2767 1081 2857 1097
rect 2767 1047 2795 1081
rect 2829 1047 2857 1081
rect 2767 1009 2857 1047
rect 2915 1081 3005 1097
rect 2915 1047 2943 1081
rect 2977 1047 3005 1081
rect 2915 1009 3005 1047
rect 3063 1081 3153 1097
rect 3063 1047 3091 1081
rect 3125 1047 3153 1081
rect 3063 1009 3153 1047
rect 3211 1081 3301 1097
rect 3211 1047 3239 1081
rect 3273 1047 3301 1081
rect 3211 1009 3301 1047
rect 3359 1081 3449 1097
rect 3359 1047 3387 1081
rect 3421 1047 3449 1081
rect 3359 1009 3449 1047
rect 3507 1081 3597 1097
rect 3507 1047 3535 1081
rect 3569 1047 3597 1081
rect 3507 1009 3597 1047
rect 3655 1081 3745 1097
rect 3655 1047 3683 1081
rect 3717 1047 3745 1081
rect 3655 1009 3745 1047
rect 3803 1081 3893 1097
rect 3803 1047 3831 1081
rect 3865 1047 3893 1081
rect 3803 1009 3893 1047
rect 3951 1081 4041 1097
rect 3951 1047 3979 1081
rect 4013 1047 4041 1081
rect 3951 1009 4041 1047
rect 4099 1081 4189 1097
rect 4099 1047 4127 1081
rect 4161 1047 4189 1081
rect 4099 1009 4189 1047
rect 4247 1081 4337 1097
rect 4247 1047 4275 1081
rect 4309 1047 4337 1081
rect 4247 1009 4337 1047
rect 4395 1081 4485 1097
rect 4395 1047 4423 1081
rect 4457 1047 4485 1081
rect 4395 1009 4485 1047
rect 4543 1081 4633 1097
rect 4543 1047 4571 1081
rect 4605 1047 4633 1081
rect 4543 1009 4633 1047
rect 4691 1081 4781 1097
rect 4691 1047 4719 1081
rect 4753 1047 4781 1081
rect 4691 1009 4781 1047
rect 4839 1081 4929 1097
rect 4839 1047 4867 1081
rect 4901 1047 4929 1081
rect 4839 1009 4929 1047
rect 4987 1081 5077 1097
rect 4987 1047 5015 1081
rect 5049 1047 5077 1081
rect 4987 1009 5077 1047
rect 5135 1081 5225 1097
rect 5135 1047 5163 1081
rect 5197 1047 5225 1081
rect 5135 1009 5225 1047
rect 5283 1081 5373 1097
rect 5283 1047 5311 1081
rect 5345 1047 5373 1081
rect 5283 1009 5373 1047
rect 5431 1081 5521 1097
rect 5431 1047 5459 1081
rect 5493 1047 5521 1081
rect 5431 1009 5521 1047
rect -5521 71 -5431 109
rect -5521 37 -5493 71
rect -5459 37 -5431 71
rect -5521 21 -5431 37
rect -5373 71 -5283 109
rect -5373 37 -5345 71
rect -5311 37 -5283 71
rect -5373 21 -5283 37
rect -5225 71 -5135 109
rect -5225 37 -5197 71
rect -5163 37 -5135 71
rect -5225 21 -5135 37
rect -5077 71 -4987 109
rect -5077 37 -5049 71
rect -5015 37 -4987 71
rect -5077 21 -4987 37
rect -4929 71 -4839 109
rect -4929 37 -4901 71
rect -4867 37 -4839 71
rect -4929 21 -4839 37
rect -4781 71 -4691 109
rect -4781 37 -4753 71
rect -4719 37 -4691 71
rect -4781 21 -4691 37
rect -4633 71 -4543 109
rect -4633 37 -4605 71
rect -4571 37 -4543 71
rect -4633 21 -4543 37
rect -4485 71 -4395 109
rect -4485 37 -4457 71
rect -4423 37 -4395 71
rect -4485 21 -4395 37
rect -4337 71 -4247 109
rect -4337 37 -4309 71
rect -4275 37 -4247 71
rect -4337 21 -4247 37
rect -4189 71 -4099 109
rect -4189 37 -4161 71
rect -4127 37 -4099 71
rect -4189 21 -4099 37
rect -4041 71 -3951 109
rect -4041 37 -4013 71
rect -3979 37 -3951 71
rect -4041 21 -3951 37
rect -3893 71 -3803 109
rect -3893 37 -3865 71
rect -3831 37 -3803 71
rect -3893 21 -3803 37
rect -3745 71 -3655 109
rect -3745 37 -3717 71
rect -3683 37 -3655 71
rect -3745 21 -3655 37
rect -3597 71 -3507 109
rect -3597 37 -3569 71
rect -3535 37 -3507 71
rect -3597 21 -3507 37
rect -3449 71 -3359 109
rect -3449 37 -3421 71
rect -3387 37 -3359 71
rect -3449 21 -3359 37
rect -3301 71 -3211 109
rect -3301 37 -3273 71
rect -3239 37 -3211 71
rect -3301 21 -3211 37
rect -3153 71 -3063 109
rect -3153 37 -3125 71
rect -3091 37 -3063 71
rect -3153 21 -3063 37
rect -3005 71 -2915 109
rect -3005 37 -2977 71
rect -2943 37 -2915 71
rect -3005 21 -2915 37
rect -2857 71 -2767 109
rect -2857 37 -2829 71
rect -2795 37 -2767 71
rect -2857 21 -2767 37
rect -2709 71 -2619 109
rect -2709 37 -2681 71
rect -2647 37 -2619 71
rect -2709 21 -2619 37
rect -2561 71 -2471 109
rect -2561 37 -2533 71
rect -2499 37 -2471 71
rect -2561 21 -2471 37
rect -2413 71 -2323 109
rect -2413 37 -2385 71
rect -2351 37 -2323 71
rect -2413 21 -2323 37
rect -2265 71 -2175 109
rect -2265 37 -2237 71
rect -2203 37 -2175 71
rect -2265 21 -2175 37
rect -2117 71 -2027 109
rect -2117 37 -2089 71
rect -2055 37 -2027 71
rect -2117 21 -2027 37
rect -1969 71 -1879 109
rect -1969 37 -1941 71
rect -1907 37 -1879 71
rect -1969 21 -1879 37
rect -1821 71 -1731 109
rect -1821 37 -1793 71
rect -1759 37 -1731 71
rect -1821 21 -1731 37
rect -1673 71 -1583 109
rect -1673 37 -1645 71
rect -1611 37 -1583 71
rect -1673 21 -1583 37
rect -1525 71 -1435 109
rect -1525 37 -1497 71
rect -1463 37 -1435 71
rect -1525 21 -1435 37
rect -1377 71 -1287 109
rect -1377 37 -1349 71
rect -1315 37 -1287 71
rect -1377 21 -1287 37
rect -1229 71 -1139 109
rect -1229 37 -1201 71
rect -1167 37 -1139 71
rect -1229 21 -1139 37
rect -1081 71 -991 109
rect -1081 37 -1053 71
rect -1019 37 -991 71
rect -1081 21 -991 37
rect -933 71 -843 109
rect -933 37 -905 71
rect -871 37 -843 71
rect -933 21 -843 37
rect -785 71 -695 109
rect -785 37 -757 71
rect -723 37 -695 71
rect -785 21 -695 37
rect -637 71 -547 109
rect -637 37 -609 71
rect -575 37 -547 71
rect -637 21 -547 37
rect -489 71 -399 109
rect -489 37 -461 71
rect -427 37 -399 71
rect -489 21 -399 37
rect -341 71 -251 109
rect -341 37 -313 71
rect -279 37 -251 71
rect -341 21 -251 37
rect -193 71 -103 109
rect -193 37 -165 71
rect -131 37 -103 71
rect -193 21 -103 37
rect -45 71 45 109
rect -45 37 -17 71
rect 17 37 45 71
rect -45 21 45 37
rect 103 71 193 109
rect 103 37 131 71
rect 165 37 193 71
rect 103 21 193 37
rect 251 71 341 109
rect 251 37 279 71
rect 313 37 341 71
rect 251 21 341 37
rect 399 71 489 109
rect 399 37 427 71
rect 461 37 489 71
rect 399 21 489 37
rect 547 71 637 109
rect 547 37 575 71
rect 609 37 637 71
rect 547 21 637 37
rect 695 71 785 109
rect 695 37 723 71
rect 757 37 785 71
rect 695 21 785 37
rect 843 71 933 109
rect 843 37 871 71
rect 905 37 933 71
rect 843 21 933 37
rect 991 71 1081 109
rect 991 37 1019 71
rect 1053 37 1081 71
rect 991 21 1081 37
rect 1139 71 1229 109
rect 1139 37 1167 71
rect 1201 37 1229 71
rect 1139 21 1229 37
rect 1287 71 1377 109
rect 1287 37 1315 71
rect 1349 37 1377 71
rect 1287 21 1377 37
rect 1435 71 1525 109
rect 1435 37 1463 71
rect 1497 37 1525 71
rect 1435 21 1525 37
rect 1583 71 1673 109
rect 1583 37 1611 71
rect 1645 37 1673 71
rect 1583 21 1673 37
rect 1731 71 1821 109
rect 1731 37 1759 71
rect 1793 37 1821 71
rect 1731 21 1821 37
rect 1879 71 1969 109
rect 1879 37 1907 71
rect 1941 37 1969 71
rect 1879 21 1969 37
rect 2027 71 2117 109
rect 2027 37 2055 71
rect 2089 37 2117 71
rect 2027 21 2117 37
rect 2175 71 2265 109
rect 2175 37 2203 71
rect 2237 37 2265 71
rect 2175 21 2265 37
rect 2323 71 2413 109
rect 2323 37 2351 71
rect 2385 37 2413 71
rect 2323 21 2413 37
rect 2471 71 2561 109
rect 2471 37 2499 71
rect 2533 37 2561 71
rect 2471 21 2561 37
rect 2619 71 2709 109
rect 2619 37 2647 71
rect 2681 37 2709 71
rect 2619 21 2709 37
rect 2767 71 2857 109
rect 2767 37 2795 71
rect 2829 37 2857 71
rect 2767 21 2857 37
rect 2915 71 3005 109
rect 2915 37 2943 71
rect 2977 37 3005 71
rect 2915 21 3005 37
rect 3063 71 3153 109
rect 3063 37 3091 71
rect 3125 37 3153 71
rect 3063 21 3153 37
rect 3211 71 3301 109
rect 3211 37 3239 71
rect 3273 37 3301 71
rect 3211 21 3301 37
rect 3359 71 3449 109
rect 3359 37 3387 71
rect 3421 37 3449 71
rect 3359 21 3449 37
rect 3507 71 3597 109
rect 3507 37 3535 71
rect 3569 37 3597 71
rect 3507 21 3597 37
rect 3655 71 3745 109
rect 3655 37 3683 71
rect 3717 37 3745 71
rect 3655 21 3745 37
rect 3803 71 3893 109
rect 3803 37 3831 71
rect 3865 37 3893 71
rect 3803 21 3893 37
rect 3951 71 4041 109
rect 3951 37 3979 71
rect 4013 37 4041 71
rect 3951 21 4041 37
rect 4099 71 4189 109
rect 4099 37 4127 71
rect 4161 37 4189 71
rect 4099 21 4189 37
rect 4247 71 4337 109
rect 4247 37 4275 71
rect 4309 37 4337 71
rect 4247 21 4337 37
rect 4395 71 4485 109
rect 4395 37 4423 71
rect 4457 37 4485 71
rect 4395 21 4485 37
rect 4543 71 4633 109
rect 4543 37 4571 71
rect 4605 37 4633 71
rect 4543 21 4633 37
rect 4691 71 4781 109
rect 4691 37 4719 71
rect 4753 37 4781 71
rect 4691 21 4781 37
rect 4839 71 4929 109
rect 4839 37 4867 71
rect 4901 37 4929 71
rect 4839 21 4929 37
rect 4987 71 5077 109
rect 4987 37 5015 71
rect 5049 37 5077 71
rect 4987 21 5077 37
rect 5135 71 5225 109
rect 5135 37 5163 71
rect 5197 37 5225 71
rect 5135 21 5225 37
rect 5283 71 5373 109
rect 5283 37 5311 71
rect 5345 37 5373 71
rect 5283 21 5373 37
rect 5431 71 5521 109
rect 5431 37 5459 71
rect 5493 37 5521 71
rect 5431 21 5521 37
rect -5521 -37 -5431 -21
rect -5521 -71 -5493 -37
rect -5459 -71 -5431 -37
rect -5521 -109 -5431 -71
rect -5373 -37 -5283 -21
rect -5373 -71 -5345 -37
rect -5311 -71 -5283 -37
rect -5373 -109 -5283 -71
rect -5225 -37 -5135 -21
rect -5225 -71 -5197 -37
rect -5163 -71 -5135 -37
rect -5225 -109 -5135 -71
rect -5077 -37 -4987 -21
rect -5077 -71 -5049 -37
rect -5015 -71 -4987 -37
rect -5077 -109 -4987 -71
rect -4929 -37 -4839 -21
rect -4929 -71 -4901 -37
rect -4867 -71 -4839 -37
rect -4929 -109 -4839 -71
rect -4781 -37 -4691 -21
rect -4781 -71 -4753 -37
rect -4719 -71 -4691 -37
rect -4781 -109 -4691 -71
rect -4633 -37 -4543 -21
rect -4633 -71 -4605 -37
rect -4571 -71 -4543 -37
rect -4633 -109 -4543 -71
rect -4485 -37 -4395 -21
rect -4485 -71 -4457 -37
rect -4423 -71 -4395 -37
rect -4485 -109 -4395 -71
rect -4337 -37 -4247 -21
rect -4337 -71 -4309 -37
rect -4275 -71 -4247 -37
rect -4337 -109 -4247 -71
rect -4189 -37 -4099 -21
rect -4189 -71 -4161 -37
rect -4127 -71 -4099 -37
rect -4189 -109 -4099 -71
rect -4041 -37 -3951 -21
rect -4041 -71 -4013 -37
rect -3979 -71 -3951 -37
rect -4041 -109 -3951 -71
rect -3893 -37 -3803 -21
rect -3893 -71 -3865 -37
rect -3831 -71 -3803 -37
rect -3893 -109 -3803 -71
rect -3745 -37 -3655 -21
rect -3745 -71 -3717 -37
rect -3683 -71 -3655 -37
rect -3745 -109 -3655 -71
rect -3597 -37 -3507 -21
rect -3597 -71 -3569 -37
rect -3535 -71 -3507 -37
rect -3597 -109 -3507 -71
rect -3449 -37 -3359 -21
rect -3449 -71 -3421 -37
rect -3387 -71 -3359 -37
rect -3449 -109 -3359 -71
rect -3301 -37 -3211 -21
rect -3301 -71 -3273 -37
rect -3239 -71 -3211 -37
rect -3301 -109 -3211 -71
rect -3153 -37 -3063 -21
rect -3153 -71 -3125 -37
rect -3091 -71 -3063 -37
rect -3153 -109 -3063 -71
rect -3005 -37 -2915 -21
rect -3005 -71 -2977 -37
rect -2943 -71 -2915 -37
rect -3005 -109 -2915 -71
rect -2857 -37 -2767 -21
rect -2857 -71 -2829 -37
rect -2795 -71 -2767 -37
rect -2857 -109 -2767 -71
rect -2709 -37 -2619 -21
rect -2709 -71 -2681 -37
rect -2647 -71 -2619 -37
rect -2709 -109 -2619 -71
rect -2561 -37 -2471 -21
rect -2561 -71 -2533 -37
rect -2499 -71 -2471 -37
rect -2561 -109 -2471 -71
rect -2413 -37 -2323 -21
rect -2413 -71 -2385 -37
rect -2351 -71 -2323 -37
rect -2413 -109 -2323 -71
rect -2265 -37 -2175 -21
rect -2265 -71 -2237 -37
rect -2203 -71 -2175 -37
rect -2265 -109 -2175 -71
rect -2117 -37 -2027 -21
rect -2117 -71 -2089 -37
rect -2055 -71 -2027 -37
rect -2117 -109 -2027 -71
rect -1969 -37 -1879 -21
rect -1969 -71 -1941 -37
rect -1907 -71 -1879 -37
rect -1969 -109 -1879 -71
rect -1821 -37 -1731 -21
rect -1821 -71 -1793 -37
rect -1759 -71 -1731 -37
rect -1821 -109 -1731 -71
rect -1673 -37 -1583 -21
rect -1673 -71 -1645 -37
rect -1611 -71 -1583 -37
rect -1673 -109 -1583 -71
rect -1525 -37 -1435 -21
rect -1525 -71 -1497 -37
rect -1463 -71 -1435 -37
rect -1525 -109 -1435 -71
rect -1377 -37 -1287 -21
rect -1377 -71 -1349 -37
rect -1315 -71 -1287 -37
rect -1377 -109 -1287 -71
rect -1229 -37 -1139 -21
rect -1229 -71 -1201 -37
rect -1167 -71 -1139 -37
rect -1229 -109 -1139 -71
rect -1081 -37 -991 -21
rect -1081 -71 -1053 -37
rect -1019 -71 -991 -37
rect -1081 -109 -991 -71
rect -933 -37 -843 -21
rect -933 -71 -905 -37
rect -871 -71 -843 -37
rect -933 -109 -843 -71
rect -785 -37 -695 -21
rect -785 -71 -757 -37
rect -723 -71 -695 -37
rect -785 -109 -695 -71
rect -637 -37 -547 -21
rect -637 -71 -609 -37
rect -575 -71 -547 -37
rect -637 -109 -547 -71
rect -489 -37 -399 -21
rect -489 -71 -461 -37
rect -427 -71 -399 -37
rect -489 -109 -399 -71
rect -341 -37 -251 -21
rect -341 -71 -313 -37
rect -279 -71 -251 -37
rect -341 -109 -251 -71
rect -193 -37 -103 -21
rect -193 -71 -165 -37
rect -131 -71 -103 -37
rect -193 -109 -103 -71
rect -45 -37 45 -21
rect -45 -71 -17 -37
rect 17 -71 45 -37
rect -45 -109 45 -71
rect 103 -37 193 -21
rect 103 -71 131 -37
rect 165 -71 193 -37
rect 103 -109 193 -71
rect 251 -37 341 -21
rect 251 -71 279 -37
rect 313 -71 341 -37
rect 251 -109 341 -71
rect 399 -37 489 -21
rect 399 -71 427 -37
rect 461 -71 489 -37
rect 399 -109 489 -71
rect 547 -37 637 -21
rect 547 -71 575 -37
rect 609 -71 637 -37
rect 547 -109 637 -71
rect 695 -37 785 -21
rect 695 -71 723 -37
rect 757 -71 785 -37
rect 695 -109 785 -71
rect 843 -37 933 -21
rect 843 -71 871 -37
rect 905 -71 933 -37
rect 843 -109 933 -71
rect 991 -37 1081 -21
rect 991 -71 1019 -37
rect 1053 -71 1081 -37
rect 991 -109 1081 -71
rect 1139 -37 1229 -21
rect 1139 -71 1167 -37
rect 1201 -71 1229 -37
rect 1139 -109 1229 -71
rect 1287 -37 1377 -21
rect 1287 -71 1315 -37
rect 1349 -71 1377 -37
rect 1287 -109 1377 -71
rect 1435 -37 1525 -21
rect 1435 -71 1463 -37
rect 1497 -71 1525 -37
rect 1435 -109 1525 -71
rect 1583 -37 1673 -21
rect 1583 -71 1611 -37
rect 1645 -71 1673 -37
rect 1583 -109 1673 -71
rect 1731 -37 1821 -21
rect 1731 -71 1759 -37
rect 1793 -71 1821 -37
rect 1731 -109 1821 -71
rect 1879 -37 1969 -21
rect 1879 -71 1907 -37
rect 1941 -71 1969 -37
rect 1879 -109 1969 -71
rect 2027 -37 2117 -21
rect 2027 -71 2055 -37
rect 2089 -71 2117 -37
rect 2027 -109 2117 -71
rect 2175 -37 2265 -21
rect 2175 -71 2203 -37
rect 2237 -71 2265 -37
rect 2175 -109 2265 -71
rect 2323 -37 2413 -21
rect 2323 -71 2351 -37
rect 2385 -71 2413 -37
rect 2323 -109 2413 -71
rect 2471 -37 2561 -21
rect 2471 -71 2499 -37
rect 2533 -71 2561 -37
rect 2471 -109 2561 -71
rect 2619 -37 2709 -21
rect 2619 -71 2647 -37
rect 2681 -71 2709 -37
rect 2619 -109 2709 -71
rect 2767 -37 2857 -21
rect 2767 -71 2795 -37
rect 2829 -71 2857 -37
rect 2767 -109 2857 -71
rect 2915 -37 3005 -21
rect 2915 -71 2943 -37
rect 2977 -71 3005 -37
rect 2915 -109 3005 -71
rect 3063 -37 3153 -21
rect 3063 -71 3091 -37
rect 3125 -71 3153 -37
rect 3063 -109 3153 -71
rect 3211 -37 3301 -21
rect 3211 -71 3239 -37
rect 3273 -71 3301 -37
rect 3211 -109 3301 -71
rect 3359 -37 3449 -21
rect 3359 -71 3387 -37
rect 3421 -71 3449 -37
rect 3359 -109 3449 -71
rect 3507 -37 3597 -21
rect 3507 -71 3535 -37
rect 3569 -71 3597 -37
rect 3507 -109 3597 -71
rect 3655 -37 3745 -21
rect 3655 -71 3683 -37
rect 3717 -71 3745 -37
rect 3655 -109 3745 -71
rect 3803 -37 3893 -21
rect 3803 -71 3831 -37
rect 3865 -71 3893 -37
rect 3803 -109 3893 -71
rect 3951 -37 4041 -21
rect 3951 -71 3979 -37
rect 4013 -71 4041 -37
rect 3951 -109 4041 -71
rect 4099 -37 4189 -21
rect 4099 -71 4127 -37
rect 4161 -71 4189 -37
rect 4099 -109 4189 -71
rect 4247 -37 4337 -21
rect 4247 -71 4275 -37
rect 4309 -71 4337 -37
rect 4247 -109 4337 -71
rect 4395 -37 4485 -21
rect 4395 -71 4423 -37
rect 4457 -71 4485 -37
rect 4395 -109 4485 -71
rect 4543 -37 4633 -21
rect 4543 -71 4571 -37
rect 4605 -71 4633 -37
rect 4543 -109 4633 -71
rect 4691 -37 4781 -21
rect 4691 -71 4719 -37
rect 4753 -71 4781 -37
rect 4691 -109 4781 -71
rect 4839 -37 4929 -21
rect 4839 -71 4867 -37
rect 4901 -71 4929 -37
rect 4839 -109 4929 -71
rect 4987 -37 5077 -21
rect 4987 -71 5015 -37
rect 5049 -71 5077 -37
rect 4987 -109 5077 -71
rect 5135 -37 5225 -21
rect 5135 -71 5163 -37
rect 5197 -71 5225 -37
rect 5135 -109 5225 -71
rect 5283 -37 5373 -21
rect 5283 -71 5311 -37
rect 5345 -71 5373 -37
rect 5283 -109 5373 -71
rect 5431 -37 5521 -21
rect 5431 -71 5459 -37
rect 5493 -71 5521 -37
rect 5431 -109 5521 -71
rect -5521 -1047 -5431 -1009
rect -5521 -1081 -5493 -1047
rect -5459 -1081 -5431 -1047
rect -5521 -1097 -5431 -1081
rect -5373 -1047 -5283 -1009
rect -5373 -1081 -5345 -1047
rect -5311 -1081 -5283 -1047
rect -5373 -1097 -5283 -1081
rect -5225 -1047 -5135 -1009
rect -5225 -1081 -5197 -1047
rect -5163 -1081 -5135 -1047
rect -5225 -1097 -5135 -1081
rect -5077 -1047 -4987 -1009
rect -5077 -1081 -5049 -1047
rect -5015 -1081 -4987 -1047
rect -5077 -1097 -4987 -1081
rect -4929 -1047 -4839 -1009
rect -4929 -1081 -4901 -1047
rect -4867 -1081 -4839 -1047
rect -4929 -1097 -4839 -1081
rect -4781 -1047 -4691 -1009
rect -4781 -1081 -4753 -1047
rect -4719 -1081 -4691 -1047
rect -4781 -1097 -4691 -1081
rect -4633 -1047 -4543 -1009
rect -4633 -1081 -4605 -1047
rect -4571 -1081 -4543 -1047
rect -4633 -1097 -4543 -1081
rect -4485 -1047 -4395 -1009
rect -4485 -1081 -4457 -1047
rect -4423 -1081 -4395 -1047
rect -4485 -1097 -4395 -1081
rect -4337 -1047 -4247 -1009
rect -4337 -1081 -4309 -1047
rect -4275 -1081 -4247 -1047
rect -4337 -1097 -4247 -1081
rect -4189 -1047 -4099 -1009
rect -4189 -1081 -4161 -1047
rect -4127 -1081 -4099 -1047
rect -4189 -1097 -4099 -1081
rect -4041 -1047 -3951 -1009
rect -4041 -1081 -4013 -1047
rect -3979 -1081 -3951 -1047
rect -4041 -1097 -3951 -1081
rect -3893 -1047 -3803 -1009
rect -3893 -1081 -3865 -1047
rect -3831 -1081 -3803 -1047
rect -3893 -1097 -3803 -1081
rect -3745 -1047 -3655 -1009
rect -3745 -1081 -3717 -1047
rect -3683 -1081 -3655 -1047
rect -3745 -1097 -3655 -1081
rect -3597 -1047 -3507 -1009
rect -3597 -1081 -3569 -1047
rect -3535 -1081 -3507 -1047
rect -3597 -1097 -3507 -1081
rect -3449 -1047 -3359 -1009
rect -3449 -1081 -3421 -1047
rect -3387 -1081 -3359 -1047
rect -3449 -1097 -3359 -1081
rect -3301 -1047 -3211 -1009
rect -3301 -1081 -3273 -1047
rect -3239 -1081 -3211 -1047
rect -3301 -1097 -3211 -1081
rect -3153 -1047 -3063 -1009
rect -3153 -1081 -3125 -1047
rect -3091 -1081 -3063 -1047
rect -3153 -1097 -3063 -1081
rect -3005 -1047 -2915 -1009
rect -3005 -1081 -2977 -1047
rect -2943 -1081 -2915 -1047
rect -3005 -1097 -2915 -1081
rect -2857 -1047 -2767 -1009
rect -2857 -1081 -2829 -1047
rect -2795 -1081 -2767 -1047
rect -2857 -1097 -2767 -1081
rect -2709 -1047 -2619 -1009
rect -2709 -1081 -2681 -1047
rect -2647 -1081 -2619 -1047
rect -2709 -1097 -2619 -1081
rect -2561 -1047 -2471 -1009
rect -2561 -1081 -2533 -1047
rect -2499 -1081 -2471 -1047
rect -2561 -1097 -2471 -1081
rect -2413 -1047 -2323 -1009
rect -2413 -1081 -2385 -1047
rect -2351 -1081 -2323 -1047
rect -2413 -1097 -2323 -1081
rect -2265 -1047 -2175 -1009
rect -2265 -1081 -2237 -1047
rect -2203 -1081 -2175 -1047
rect -2265 -1097 -2175 -1081
rect -2117 -1047 -2027 -1009
rect -2117 -1081 -2089 -1047
rect -2055 -1081 -2027 -1047
rect -2117 -1097 -2027 -1081
rect -1969 -1047 -1879 -1009
rect -1969 -1081 -1941 -1047
rect -1907 -1081 -1879 -1047
rect -1969 -1097 -1879 -1081
rect -1821 -1047 -1731 -1009
rect -1821 -1081 -1793 -1047
rect -1759 -1081 -1731 -1047
rect -1821 -1097 -1731 -1081
rect -1673 -1047 -1583 -1009
rect -1673 -1081 -1645 -1047
rect -1611 -1081 -1583 -1047
rect -1673 -1097 -1583 -1081
rect -1525 -1047 -1435 -1009
rect -1525 -1081 -1497 -1047
rect -1463 -1081 -1435 -1047
rect -1525 -1097 -1435 -1081
rect -1377 -1047 -1287 -1009
rect -1377 -1081 -1349 -1047
rect -1315 -1081 -1287 -1047
rect -1377 -1097 -1287 -1081
rect -1229 -1047 -1139 -1009
rect -1229 -1081 -1201 -1047
rect -1167 -1081 -1139 -1047
rect -1229 -1097 -1139 -1081
rect -1081 -1047 -991 -1009
rect -1081 -1081 -1053 -1047
rect -1019 -1081 -991 -1047
rect -1081 -1097 -991 -1081
rect -933 -1047 -843 -1009
rect -933 -1081 -905 -1047
rect -871 -1081 -843 -1047
rect -933 -1097 -843 -1081
rect -785 -1047 -695 -1009
rect -785 -1081 -757 -1047
rect -723 -1081 -695 -1047
rect -785 -1097 -695 -1081
rect -637 -1047 -547 -1009
rect -637 -1081 -609 -1047
rect -575 -1081 -547 -1047
rect -637 -1097 -547 -1081
rect -489 -1047 -399 -1009
rect -489 -1081 -461 -1047
rect -427 -1081 -399 -1047
rect -489 -1097 -399 -1081
rect -341 -1047 -251 -1009
rect -341 -1081 -313 -1047
rect -279 -1081 -251 -1047
rect -341 -1097 -251 -1081
rect -193 -1047 -103 -1009
rect -193 -1081 -165 -1047
rect -131 -1081 -103 -1047
rect -193 -1097 -103 -1081
rect -45 -1047 45 -1009
rect -45 -1081 -17 -1047
rect 17 -1081 45 -1047
rect -45 -1097 45 -1081
rect 103 -1047 193 -1009
rect 103 -1081 131 -1047
rect 165 -1081 193 -1047
rect 103 -1097 193 -1081
rect 251 -1047 341 -1009
rect 251 -1081 279 -1047
rect 313 -1081 341 -1047
rect 251 -1097 341 -1081
rect 399 -1047 489 -1009
rect 399 -1081 427 -1047
rect 461 -1081 489 -1047
rect 399 -1097 489 -1081
rect 547 -1047 637 -1009
rect 547 -1081 575 -1047
rect 609 -1081 637 -1047
rect 547 -1097 637 -1081
rect 695 -1047 785 -1009
rect 695 -1081 723 -1047
rect 757 -1081 785 -1047
rect 695 -1097 785 -1081
rect 843 -1047 933 -1009
rect 843 -1081 871 -1047
rect 905 -1081 933 -1047
rect 843 -1097 933 -1081
rect 991 -1047 1081 -1009
rect 991 -1081 1019 -1047
rect 1053 -1081 1081 -1047
rect 991 -1097 1081 -1081
rect 1139 -1047 1229 -1009
rect 1139 -1081 1167 -1047
rect 1201 -1081 1229 -1047
rect 1139 -1097 1229 -1081
rect 1287 -1047 1377 -1009
rect 1287 -1081 1315 -1047
rect 1349 -1081 1377 -1047
rect 1287 -1097 1377 -1081
rect 1435 -1047 1525 -1009
rect 1435 -1081 1463 -1047
rect 1497 -1081 1525 -1047
rect 1435 -1097 1525 -1081
rect 1583 -1047 1673 -1009
rect 1583 -1081 1611 -1047
rect 1645 -1081 1673 -1047
rect 1583 -1097 1673 -1081
rect 1731 -1047 1821 -1009
rect 1731 -1081 1759 -1047
rect 1793 -1081 1821 -1047
rect 1731 -1097 1821 -1081
rect 1879 -1047 1969 -1009
rect 1879 -1081 1907 -1047
rect 1941 -1081 1969 -1047
rect 1879 -1097 1969 -1081
rect 2027 -1047 2117 -1009
rect 2027 -1081 2055 -1047
rect 2089 -1081 2117 -1047
rect 2027 -1097 2117 -1081
rect 2175 -1047 2265 -1009
rect 2175 -1081 2203 -1047
rect 2237 -1081 2265 -1047
rect 2175 -1097 2265 -1081
rect 2323 -1047 2413 -1009
rect 2323 -1081 2351 -1047
rect 2385 -1081 2413 -1047
rect 2323 -1097 2413 -1081
rect 2471 -1047 2561 -1009
rect 2471 -1081 2499 -1047
rect 2533 -1081 2561 -1047
rect 2471 -1097 2561 -1081
rect 2619 -1047 2709 -1009
rect 2619 -1081 2647 -1047
rect 2681 -1081 2709 -1047
rect 2619 -1097 2709 -1081
rect 2767 -1047 2857 -1009
rect 2767 -1081 2795 -1047
rect 2829 -1081 2857 -1047
rect 2767 -1097 2857 -1081
rect 2915 -1047 3005 -1009
rect 2915 -1081 2943 -1047
rect 2977 -1081 3005 -1047
rect 2915 -1097 3005 -1081
rect 3063 -1047 3153 -1009
rect 3063 -1081 3091 -1047
rect 3125 -1081 3153 -1047
rect 3063 -1097 3153 -1081
rect 3211 -1047 3301 -1009
rect 3211 -1081 3239 -1047
rect 3273 -1081 3301 -1047
rect 3211 -1097 3301 -1081
rect 3359 -1047 3449 -1009
rect 3359 -1081 3387 -1047
rect 3421 -1081 3449 -1047
rect 3359 -1097 3449 -1081
rect 3507 -1047 3597 -1009
rect 3507 -1081 3535 -1047
rect 3569 -1081 3597 -1047
rect 3507 -1097 3597 -1081
rect 3655 -1047 3745 -1009
rect 3655 -1081 3683 -1047
rect 3717 -1081 3745 -1047
rect 3655 -1097 3745 -1081
rect 3803 -1047 3893 -1009
rect 3803 -1081 3831 -1047
rect 3865 -1081 3893 -1047
rect 3803 -1097 3893 -1081
rect 3951 -1047 4041 -1009
rect 3951 -1081 3979 -1047
rect 4013 -1081 4041 -1047
rect 3951 -1097 4041 -1081
rect 4099 -1047 4189 -1009
rect 4099 -1081 4127 -1047
rect 4161 -1081 4189 -1047
rect 4099 -1097 4189 -1081
rect 4247 -1047 4337 -1009
rect 4247 -1081 4275 -1047
rect 4309 -1081 4337 -1047
rect 4247 -1097 4337 -1081
rect 4395 -1047 4485 -1009
rect 4395 -1081 4423 -1047
rect 4457 -1081 4485 -1047
rect 4395 -1097 4485 -1081
rect 4543 -1047 4633 -1009
rect 4543 -1081 4571 -1047
rect 4605 -1081 4633 -1047
rect 4543 -1097 4633 -1081
rect 4691 -1047 4781 -1009
rect 4691 -1081 4719 -1047
rect 4753 -1081 4781 -1047
rect 4691 -1097 4781 -1081
rect 4839 -1047 4929 -1009
rect 4839 -1081 4867 -1047
rect 4901 -1081 4929 -1047
rect 4839 -1097 4929 -1081
rect 4987 -1047 5077 -1009
rect 4987 -1081 5015 -1047
rect 5049 -1081 5077 -1047
rect 4987 -1097 5077 -1081
rect 5135 -1047 5225 -1009
rect 5135 -1081 5163 -1047
rect 5197 -1081 5225 -1047
rect 5135 -1097 5225 -1081
rect 5283 -1047 5373 -1009
rect 5283 -1081 5311 -1047
rect 5345 -1081 5373 -1047
rect 5283 -1097 5373 -1081
rect 5431 -1047 5521 -1009
rect 5431 -1081 5459 -1047
rect 5493 -1081 5521 -1047
rect 5431 -1097 5521 -1081
<< polycont >>
rect -5493 1047 -5459 1081
rect -5345 1047 -5311 1081
rect -5197 1047 -5163 1081
rect -5049 1047 -5015 1081
rect -4901 1047 -4867 1081
rect -4753 1047 -4719 1081
rect -4605 1047 -4571 1081
rect -4457 1047 -4423 1081
rect -4309 1047 -4275 1081
rect -4161 1047 -4127 1081
rect -4013 1047 -3979 1081
rect -3865 1047 -3831 1081
rect -3717 1047 -3683 1081
rect -3569 1047 -3535 1081
rect -3421 1047 -3387 1081
rect -3273 1047 -3239 1081
rect -3125 1047 -3091 1081
rect -2977 1047 -2943 1081
rect -2829 1047 -2795 1081
rect -2681 1047 -2647 1081
rect -2533 1047 -2499 1081
rect -2385 1047 -2351 1081
rect -2237 1047 -2203 1081
rect -2089 1047 -2055 1081
rect -1941 1047 -1907 1081
rect -1793 1047 -1759 1081
rect -1645 1047 -1611 1081
rect -1497 1047 -1463 1081
rect -1349 1047 -1315 1081
rect -1201 1047 -1167 1081
rect -1053 1047 -1019 1081
rect -905 1047 -871 1081
rect -757 1047 -723 1081
rect -609 1047 -575 1081
rect -461 1047 -427 1081
rect -313 1047 -279 1081
rect -165 1047 -131 1081
rect -17 1047 17 1081
rect 131 1047 165 1081
rect 279 1047 313 1081
rect 427 1047 461 1081
rect 575 1047 609 1081
rect 723 1047 757 1081
rect 871 1047 905 1081
rect 1019 1047 1053 1081
rect 1167 1047 1201 1081
rect 1315 1047 1349 1081
rect 1463 1047 1497 1081
rect 1611 1047 1645 1081
rect 1759 1047 1793 1081
rect 1907 1047 1941 1081
rect 2055 1047 2089 1081
rect 2203 1047 2237 1081
rect 2351 1047 2385 1081
rect 2499 1047 2533 1081
rect 2647 1047 2681 1081
rect 2795 1047 2829 1081
rect 2943 1047 2977 1081
rect 3091 1047 3125 1081
rect 3239 1047 3273 1081
rect 3387 1047 3421 1081
rect 3535 1047 3569 1081
rect 3683 1047 3717 1081
rect 3831 1047 3865 1081
rect 3979 1047 4013 1081
rect 4127 1047 4161 1081
rect 4275 1047 4309 1081
rect 4423 1047 4457 1081
rect 4571 1047 4605 1081
rect 4719 1047 4753 1081
rect 4867 1047 4901 1081
rect 5015 1047 5049 1081
rect 5163 1047 5197 1081
rect 5311 1047 5345 1081
rect 5459 1047 5493 1081
rect -5493 37 -5459 71
rect -5345 37 -5311 71
rect -5197 37 -5163 71
rect -5049 37 -5015 71
rect -4901 37 -4867 71
rect -4753 37 -4719 71
rect -4605 37 -4571 71
rect -4457 37 -4423 71
rect -4309 37 -4275 71
rect -4161 37 -4127 71
rect -4013 37 -3979 71
rect -3865 37 -3831 71
rect -3717 37 -3683 71
rect -3569 37 -3535 71
rect -3421 37 -3387 71
rect -3273 37 -3239 71
rect -3125 37 -3091 71
rect -2977 37 -2943 71
rect -2829 37 -2795 71
rect -2681 37 -2647 71
rect -2533 37 -2499 71
rect -2385 37 -2351 71
rect -2237 37 -2203 71
rect -2089 37 -2055 71
rect -1941 37 -1907 71
rect -1793 37 -1759 71
rect -1645 37 -1611 71
rect -1497 37 -1463 71
rect -1349 37 -1315 71
rect -1201 37 -1167 71
rect -1053 37 -1019 71
rect -905 37 -871 71
rect -757 37 -723 71
rect -609 37 -575 71
rect -461 37 -427 71
rect -313 37 -279 71
rect -165 37 -131 71
rect -17 37 17 71
rect 131 37 165 71
rect 279 37 313 71
rect 427 37 461 71
rect 575 37 609 71
rect 723 37 757 71
rect 871 37 905 71
rect 1019 37 1053 71
rect 1167 37 1201 71
rect 1315 37 1349 71
rect 1463 37 1497 71
rect 1611 37 1645 71
rect 1759 37 1793 71
rect 1907 37 1941 71
rect 2055 37 2089 71
rect 2203 37 2237 71
rect 2351 37 2385 71
rect 2499 37 2533 71
rect 2647 37 2681 71
rect 2795 37 2829 71
rect 2943 37 2977 71
rect 3091 37 3125 71
rect 3239 37 3273 71
rect 3387 37 3421 71
rect 3535 37 3569 71
rect 3683 37 3717 71
rect 3831 37 3865 71
rect 3979 37 4013 71
rect 4127 37 4161 71
rect 4275 37 4309 71
rect 4423 37 4457 71
rect 4571 37 4605 71
rect 4719 37 4753 71
rect 4867 37 4901 71
rect 5015 37 5049 71
rect 5163 37 5197 71
rect 5311 37 5345 71
rect 5459 37 5493 71
rect -5493 -71 -5459 -37
rect -5345 -71 -5311 -37
rect -5197 -71 -5163 -37
rect -5049 -71 -5015 -37
rect -4901 -71 -4867 -37
rect -4753 -71 -4719 -37
rect -4605 -71 -4571 -37
rect -4457 -71 -4423 -37
rect -4309 -71 -4275 -37
rect -4161 -71 -4127 -37
rect -4013 -71 -3979 -37
rect -3865 -71 -3831 -37
rect -3717 -71 -3683 -37
rect -3569 -71 -3535 -37
rect -3421 -71 -3387 -37
rect -3273 -71 -3239 -37
rect -3125 -71 -3091 -37
rect -2977 -71 -2943 -37
rect -2829 -71 -2795 -37
rect -2681 -71 -2647 -37
rect -2533 -71 -2499 -37
rect -2385 -71 -2351 -37
rect -2237 -71 -2203 -37
rect -2089 -71 -2055 -37
rect -1941 -71 -1907 -37
rect -1793 -71 -1759 -37
rect -1645 -71 -1611 -37
rect -1497 -71 -1463 -37
rect -1349 -71 -1315 -37
rect -1201 -71 -1167 -37
rect -1053 -71 -1019 -37
rect -905 -71 -871 -37
rect -757 -71 -723 -37
rect -609 -71 -575 -37
rect -461 -71 -427 -37
rect -313 -71 -279 -37
rect -165 -71 -131 -37
rect -17 -71 17 -37
rect 131 -71 165 -37
rect 279 -71 313 -37
rect 427 -71 461 -37
rect 575 -71 609 -37
rect 723 -71 757 -37
rect 871 -71 905 -37
rect 1019 -71 1053 -37
rect 1167 -71 1201 -37
rect 1315 -71 1349 -37
rect 1463 -71 1497 -37
rect 1611 -71 1645 -37
rect 1759 -71 1793 -37
rect 1907 -71 1941 -37
rect 2055 -71 2089 -37
rect 2203 -71 2237 -37
rect 2351 -71 2385 -37
rect 2499 -71 2533 -37
rect 2647 -71 2681 -37
rect 2795 -71 2829 -37
rect 2943 -71 2977 -37
rect 3091 -71 3125 -37
rect 3239 -71 3273 -37
rect 3387 -71 3421 -37
rect 3535 -71 3569 -37
rect 3683 -71 3717 -37
rect 3831 -71 3865 -37
rect 3979 -71 4013 -37
rect 4127 -71 4161 -37
rect 4275 -71 4309 -37
rect 4423 -71 4457 -37
rect 4571 -71 4605 -37
rect 4719 -71 4753 -37
rect 4867 -71 4901 -37
rect 5015 -71 5049 -37
rect 5163 -71 5197 -37
rect 5311 -71 5345 -37
rect 5459 -71 5493 -37
rect -5493 -1081 -5459 -1047
rect -5345 -1081 -5311 -1047
rect -5197 -1081 -5163 -1047
rect -5049 -1081 -5015 -1047
rect -4901 -1081 -4867 -1047
rect -4753 -1081 -4719 -1047
rect -4605 -1081 -4571 -1047
rect -4457 -1081 -4423 -1047
rect -4309 -1081 -4275 -1047
rect -4161 -1081 -4127 -1047
rect -4013 -1081 -3979 -1047
rect -3865 -1081 -3831 -1047
rect -3717 -1081 -3683 -1047
rect -3569 -1081 -3535 -1047
rect -3421 -1081 -3387 -1047
rect -3273 -1081 -3239 -1047
rect -3125 -1081 -3091 -1047
rect -2977 -1081 -2943 -1047
rect -2829 -1081 -2795 -1047
rect -2681 -1081 -2647 -1047
rect -2533 -1081 -2499 -1047
rect -2385 -1081 -2351 -1047
rect -2237 -1081 -2203 -1047
rect -2089 -1081 -2055 -1047
rect -1941 -1081 -1907 -1047
rect -1793 -1081 -1759 -1047
rect -1645 -1081 -1611 -1047
rect -1497 -1081 -1463 -1047
rect -1349 -1081 -1315 -1047
rect -1201 -1081 -1167 -1047
rect -1053 -1081 -1019 -1047
rect -905 -1081 -871 -1047
rect -757 -1081 -723 -1047
rect -609 -1081 -575 -1047
rect -461 -1081 -427 -1047
rect -313 -1081 -279 -1047
rect -165 -1081 -131 -1047
rect -17 -1081 17 -1047
rect 131 -1081 165 -1047
rect 279 -1081 313 -1047
rect 427 -1081 461 -1047
rect 575 -1081 609 -1047
rect 723 -1081 757 -1047
rect 871 -1081 905 -1047
rect 1019 -1081 1053 -1047
rect 1167 -1081 1201 -1047
rect 1315 -1081 1349 -1047
rect 1463 -1081 1497 -1047
rect 1611 -1081 1645 -1047
rect 1759 -1081 1793 -1047
rect 1907 -1081 1941 -1047
rect 2055 -1081 2089 -1047
rect 2203 -1081 2237 -1047
rect 2351 -1081 2385 -1047
rect 2499 -1081 2533 -1047
rect 2647 -1081 2681 -1047
rect 2795 -1081 2829 -1047
rect 2943 -1081 2977 -1047
rect 3091 -1081 3125 -1047
rect 3239 -1081 3273 -1047
rect 3387 -1081 3421 -1047
rect 3535 -1081 3569 -1047
rect 3683 -1081 3717 -1047
rect 3831 -1081 3865 -1047
rect 3979 -1081 4013 -1047
rect 4127 -1081 4161 -1047
rect 4275 -1081 4309 -1047
rect 4423 -1081 4457 -1047
rect 4571 -1081 4605 -1047
rect 4719 -1081 4753 -1047
rect 4867 -1081 4901 -1047
rect 5015 -1081 5049 -1047
rect 5163 -1081 5197 -1047
rect 5311 -1081 5345 -1047
rect 5459 -1081 5493 -1047
<< locali >>
rect -5681 1149 -5559 1183
rect -5525 1149 -5491 1183
rect -5457 1149 -5423 1183
rect -5389 1149 -5355 1183
rect -5321 1149 -5287 1183
rect -5253 1149 -5219 1183
rect -5185 1149 -5151 1183
rect -5117 1149 -5083 1183
rect -5049 1149 -5015 1183
rect -4981 1149 -4947 1183
rect -4913 1149 -4879 1183
rect -4845 1149 -4811 1183
rect -4777 1149 -4743 1183
rect -4709 1149 -4675 1183
rect -4641 1149 -4607 1183
rect -4573 1149 -4539 1183
rect -4505 1149 -4471 1183
rect -4437 1149 -4403 1183
rect -4369 1149 -4335 1183
rect -4301 1149 -4267 1183
rect -4233 1149 -4199 1183
rect -4165 1149 -4131 1183
rect -4097 1149 -4063 1183
rect -4029 1149 -3995 1183
rect -3961 1149 -3927 1183
rect -3893 1149 -3859 1183
rect -3825 1149 -3791 1183
rect -3757 1149 -3723 1183
rect -3689 1149 -3655 1183
rect -3621 1149 -3587 1183
rect -3553 1149 -3519 1183
rect -3485 1149 -3451 1183
rect -3417 1149 -3383 1183
rect -3349 1149 -3315 1183
rect -3281 1149 -3247 1183
rect -3213 1149 -3179 1183
rect -3145 1149 -3111 1183
rect -3077 1149 -3043 1183
rect -3009 1149 -2975 1183
rect -2941 1149 -2907 1183
rect -2873 1149 -2839 1183
rect -2805 1149 -2771 1183
rect -2737 1149 -2703 1183
rect -2669 1149 -2635 1183
rect -2601 1149 -2567 1183
rect -2533 1149 -2499 1183
rect -2465 1149 -2431 1183
rect -2397 1149 -2363 1183
rect -2329 1149 -2295 1183
rect -2261 1149 -2227 1183
rect -2193 1149 -2159 1183
rect -2125 1149 -2091 1183
rect -2057 1149 -2023 1183
rect -1989 1149 -1955 1183
rect -1921 1149 -1887 1183
rect -1853 1149 -1819 1183
rect -1785 1149 -1751 1183
rect -1717 1149 -1683 1183
rect -1649 1149 -1615 1183
rect -1581 1149 -1547 1183
rect -1513 1149 -1479 1183
rect -1445 1149 -1411 1183
rect -1377 1149 -1343 1183
rect -1309 1149 -1275 1183
rect -1241 1149 -1207 1183
rect -1173 1149 -1139 1183
rect -1105 1149 -1071 1183
rect -1037 1149 -1003 1183
rect -969 1149 -935 1183
rect -901 1149 -867 1183
rect -833 1149 -799 1183
rect -765 1149 -731 1183
rect -697 1149 -663 1183
rect -629 1149 -595 1183
rect -561 1149 -527 1183
rect -493 1149 -459 1183
rect -425 1149 -391 1183
rect -357 1149 -323 1183
rect -289 1149 -255 1183
rect -221 1149 -187 1183
rect -153 1149 -119 1183
rect -85 1149 -51 1183
rect -17 1149 17 1183
rect 51 1149 85 1183
rect 119 1149 153 1183
rect 187 1149 221 1183
rect 255 1149 289 1183
rect 323 1149 357 1183
rect 391 1149 425 1183
rect 459 1149 493 1183
rect 527 1149 561 1183
rect 595 1149 629 1183
rect 663 1149 697 1183
rect 731 1149 765 1183
rect 799 1149 833 1183
rect 867 1149 901 1183
rect 935 1149 969 1183
rect 1003 1149 1037 1183
rect 1071 1149 1105 1183
rect 1139 1149 1173 1183
rect 1207 1149 1241 1183
rect 1275 1149 1309 1183
rect 1343 1149 1377 1183
rect 1411 1149 1445 1183
rect 1479 1149 1513 1183
rect 1547 1149 1581 1183
rect 1615 1149 1649 1183
rect 1683 1149 1717 1183
rect 1751 1149 1785 1183
rect 1819 1149 1853 1183
rect 1887 1149 1921 1183
rect 1955 1149 1989 1183
rect 2023 1149 2057 1183
rect 2091 1149 2125 1183
rect 2159 1149 2193 1183
rect 2227 1149 2261 1183
rect 2295 1149 2329 1183
rect 2363 1149 2397 1183
rect 2431 1149 2465 1183
rect 2499 1149 2533 1183
rect 2567 1149 2601 1183
rect 2635 1149 2669 1183
rect 2703 1149 2737 1183
rect 2771 1149 2805 1183
rect 2839 1149 2873 1183
rect 2907 1149 2941 1183
rect 2975 1149 3009 1183
rect 3043 1149 3077 1183
rect 3111 1149 3145 1183
rect 3179 1149 3213 1183
rect 3247 1149 3281 1183
rect 3315 1149 3349 1183
rect 3383 1149 3417 1183
rect 3451 1149 3485 1183
rect 3519 1149 3553 1183
rect 3587 1149 3621 1183
rect 3655 1149 3689 1183
rect 3723 1149 3757 1183
rect 3791 1149 3825 1183
rect 3859 1149 3893 1183
rect 3927 1149 3961 1183
rect 3995 1149 4029 1183
rect 4063 1149 4097 1183
rect 4131 1149 4165 1183
rect 4199 1149 4233 1183
rect 4267 1149 4301 1183
rect 4335 1149 4369 1183
rect 4403 1149 4437 1183
rect 4471 1149 4505 1183
rect 4539 1149 4573 1183
rect 4607 1149 4641 1183
rect 4675 1149 4709 1183
rect 4743 1149 4777 1183
rect 4811 1149 4845 1183
rect 4879 1149 4913 1183
rect 4947 1149 4981 1183
rect 5015 1149 5049 1183
rect 5083 1149 5117 1183
rect 5151 1149 5185 1183
rect 5219 1149 5253 1183
rect 5287 1149 5321 1183
rect 5355 1149 5389 1183
rect 5423 1149 5457 1183
rect 5491 1149 5525 1183
rect 5559 1149 5681 1183
rect -5681 1071 -5647 1149
rect -5521 1047 -5493 1081
rect -5459 1047 -5431 1081
rect -5373 1047 -5345 1081
rect -5311 1047 -5283 1081
rect -5225 1047 -5197 1081
rect -5163 1047 -5135 1081
rect -5077 1047 -5049 1081
rect -5015 1047 -4987 1081
rect -4929 1047 -4901 1081
rect -4867 1047 -4839 1081
rect -4781 1047 -4753 1081
rect -4719 1047 -4691 1081
rect -4633 1047 -4605 1081
rect -4571 1047 -4543 1081
rect -4485 1047 -4457 1081
rect -4423 1047 -4395 1081
rect -4337 1047 -4309 1081
rect -4275 1047 -4247 1081
rect -4189 1047 -4161 1081
rect -4127 1047 -4099 1081
rect -4041 1047 -4013 1081
rect -3979 1047 -3951 1081
rect -3893 1047 -3865 1081
rect -3831 1047 -3803 1081
rect -3745 1047 -3717 1081
rect -3683 1047 -3655 1081
rect -3597 1047 -3569 1081
rect -3535 1047 -3507 1081
rect -3449 1047 -3421 1081
rect -3387 1047 -3359 1081
rect -3301 1047 -3273 1081
rect -3239 1047 -3211 1081
rect -3153 1047 -3125 1081
rect -3091 1047 -3063 1081
rect -3005 1047 -2977 1081
rect -2943 1047 -2915 1081
rect -2857 1047 -2829 1081
rect -2795 1047 -2767 1081
rect -2709 1047 -2681 1081
rect -2647 1047 -2619 1081
rect -2561 1047 -2533 1081
rect -2499 1047 -2471 1081
rect -2413 1047 -2385 1081
rect -2351 1047 -2323 1081
rect -2265 1047 -2237 1081
rect -2203 1047 -2175 1081
rect -2117 1047 -2089 1081
rect -2055 1047 -2027 1081
rect -1969 1047 -1941 1081
rect -1907 1047 -1879 1081
rect -1821 1047 -1793 1081
rect -1759 1047 -1731 1081
rect -1673 1047 -1645 1081
rect -1611 1047 -1583 1081
rect -1525 1047 -1497 1081
rect -1463 1047 -1435 1081
rect -1377 1047 -1349 1081
rect -1315 1047 -1287 1081
rect -1229 1047 -1201 1081
rect -1167 1047 -1139 1081
rect -1081 1047 -1053 1081
rect -1019 1047 -991 1081
rect -933 1047 -905 1081
rect -871 1047 -843 1081
rect -785 1047 -757 1081
rect -723 1047 -695 1081
rect -637 1047 -609 1081
rect -575 1047 -547 1081
rect -489 1047 -461 1081
rect -427 1047 -399 1081
rect -341 1047 -313 1081
rect -279 1047 -251 1081
rect -193 1047 -165 1081
rect -131 1047 -103 1081
rect -45 1047 -17 1081
rect 17 1047 45 1081
rect 103 1047 131 1081
rect 165 1047 193 1081
rect 251 1047 279 1081
rect 313 1047 341 1081
rect 399 1047 427 1081
rect 461 1047 489 1081
rect 547 1047 575 1081
rect 609 1047 637 1081
rect 695 1047 723 1081
rect 757 1047 785 1081
rect 843 1047 871 1081
rect 905 1047 933 1081
rect 991 1047 1019 1081
rect 1053 1047 1081 1081
rect 1139 1047 1167 1081
rect 1201 1047 1229 1081
rect 1287 1047 1315 1081
rect 1349 1047 1377 1081
rect 1435 1047 1463 1081
rect 1497 1047 1525 1081
rect 1583 1047 1611 1081
rect 1645 1047 1673 1081
rect 1731 1047 1759 1081
rect 1793 1047 1821 1081
rect 1879 1047 1907 1081
rect 1941 1047 1969 1081
rect 2027 1047 2055 1081
rect 2089 1047 2117 1081
rect 2175 1047 2203 1081
rect 2237 1047 2265 1081
rect 2323 1047 2351 1081
rect 2385 1047 2413 1081
rect 2471 1047 2499 1081
rect 2533 1047 2561 1081
rect 2619 1047 2647 1081
rect 2681 1047 2709 1081
rect 2767 1047 2795 1081
rect 2829 1047 2857 1081
rect 2915 1047 2943 1081
rect 2977 1047 3005 1081
rect 3063 1047 3091 1081
rect 3125 1047 3153 1081
rect 3211 1047 3239 1081
rect 3273 1047 3301 1081
rect 3359 1047 3387 1081
rect 3421 1047 3449 1081
rect 3507 1047 3535 1081
rect 3569 1047 3597 1081
rect 3655 1047 3683 1081
rect 3717 1047 3745 1081
rect 3803 1047 3831 1081
rect 3865 1047 3893 1081
rect 3951 1047 3979 1081
rect 4013 1047 4041 1081
rect 4099 1047 4127 1081
rect 4161 1047 4189 1081
rect 4247 1047 4275 1081
rect 4309 1047 4337 1081
rect 4395 1047 4423 1081
rect 4457 1047 4485 1081
rect 4543 1047 4571 1081
rect 4605 1047 4633 1081
rect 4691 1047 4719 1081
rect 4753 1047 4781 1081
rect 4839 1047 4867 1081
rect 4901 1047 4929 1081
rect 4987 1047 5015 1081
rect 5049 1047 5077 1081
rect 5135 1047 5163 1081
rect 5197 1047 5225 1081
rect 5283 1047 5311 1081
rect 5345 1047 5373 1081
rect 5431 1047 5459 1081
rect 5493 1047 5521 1081
rect 5647 1071 5681 1149
rect -5681 1003 -5647 1037
rect -5681 935 -5647 969
rect -5681 867 -5647 901
rect -5681 799 -5647 833
rect -5681 731 -5647 765
rect -5681 663 -5647 697
rect -5681 595 -5647 629
rect -5681 527 -5647 561
rect -5681 459 -5647 493
rect -5681 391 -5647 425
rect -5681 323 -5647 357
rect -5681 255 -5647 289
rect -5681 187 -5647 221
rect -5681 119 -5647 153
rect -5567 984 -5533 1013
rect -5567 916 -5533 938
rect -5567 848 -5533 866
rect -5567 780 -5533 794
rect -5567 712 -5533 722
rect -5567 644 -5533 650
rect -5567 576 -5533 578
rect -5567 540 -5533 542
rect -5567 468 -5533 474
rect -5567 396 -5533 406
rect -5567 324 -5533 338
rect -5567 252 -5533 270
rect -5567 180 -5533 202
rect -5567 105 -5533 134
rect -5419 984 -5385 1013
rect -5419 916 -5385 938
rect -5419 848 -5385 866
rect -5419 780 -5385 794
rect -5419 712 -5385 722
rect -5419 644 -5385 650
rect -5419 576 -5385 578
rect -5419 540 -5385 542
rect -5419 468 -5385 474
rect -5419 396 -5385 406
rect -5419 324 -5385 338
rect -5419 252 -5385 270
rect -5419 180 -5385 202
rect -5419 105 -5385 134
rect -5271 984 -5237 1013
rect -5271 916 -5237 938
rect -5271 848 -5237 866
rect -5271 780 -5237 794
rect -5271 712 -5237 722
rect -5271 644 -5237 650
rect -5271 576 -5237 578
rect -5271 540 -5237 542
rect -5271 468 -5237 474
rect -5271 396 -5237 406
rect -5271 324 -5237 338
rect -5271 252 -5237 270
rect -5271 180 -5237 202
rect -5271 105 -5237 134
rect -5123 984 -5089 1013
rect -5123 916 -5089 938
rect -5123 848 -5089 866
rect -5123 780 -5089 794
rect -5123 712 -5089 722
rect -5123 644 -5089 650
rect -5123 576 -5089 578
rect -5123 540 -5089 542
rect -5123 468 -5089 474
rect -5123 396 -5089 406
rect -5123 324 -5089 338
rect -5123 252 -5089 270
rect -5123 180 -5089 202
rect -5123 105 -5089 134
rect -4975 984 -4941 1013
rect -4975 916 -4941 938
rect -4975 848 -4941 866
rect -4975 780 -4941 794
rect -4975 712 -4941 722
rect -4975 644 -4941 650
rect -4975 576 -4941 578
rect -4975 540 -4941 542
rect -4975 468 -4941 474
rect -4975 396 -4941 406
rect -4975 324 -4941 338
rect -4975 252 -4941 270
rect -4975 180 -4941 202
rect -4975 105 -4941 134
rect -4827 984 -4793 1013
rect -4827 916 -4793 938
rect -4827 848 -4793 866
rect -4827 780 -4793 794
rect -4827 712 -4793 722
rect -4827 644 -4793 650
rect -4827 576 -4793 578
rect -4827 540 -4793 542
rect -4827 468 -4793 474
rect -4827 396 -4793 406
rect -4827 324 -4793 338
rect -4827 252 -4793 270
rect -4827 180 -4793 202
rect -4827 105 -4793 134
rect -4679 984 -4645 1013
rect -4679 916 -4645 938
rect -4679 848 -4645 866
rect -4679 780 -4645 794
rect -4679 712 -4645 722
rect -4679 644 -4645 650
rect -4679 576 -4645 578
rect -4679 540 -4645 542
rect -4679 468 -4645 474
rect -4679 396 -4645 406
rect -4679 324 -4645 338
rect -4679 252 -4645 270
rect -4679 180 -4645 202
rect -4679 105 -4645 134
rect -4531 984 -4497 1013
rect -4531 916 -4497 938
rect -4531 848 -4497 866
rect -4531 780 -4497 794
rect -4531 712 -4497 722
rect -4531 644 -4497 650
rect -4531 576 -4497 578
rect -4531 540 -4497 542
rect -4531 468 -4497 474
rect -4531 396 -4497 406
rect -4531 324 -4497 338
rect -4531 252 -4497 270
rect -4531 180 -4497 202
rect -4531 105 -4497 134
rect -4383 984 -4349 1013
rect -4383 916 -4349 938
rect -4383 848 -4349 866
rect -4383 780 -4349 794
rect -4383 712 -4349 722
rect -4383 644 -4349 650
rect -4383 576 -4349 578
rect -4383 540 -4349 542
rect -4383 468 -4349 474
rect -4383 396 -4349 406
rect -4383 324 -4349 338
rect -4383 252 -4349 270
rect -4383 180 -4349 202
rect -4383 105 -4349 134
rect -4235 984 -4201 1013
rect -4235 916 -4201 938
rect -4235 848 -4201 866
rect -4235 780 -4201 794
rect -4235 712 -4201 722
rect -4235 644 -4201 650
rect -4235 576 -4201 578
rect -4235 540 -4201 542
rect -4235 468 -4201 474
rect -4235 396 -4201 406
rect -4235 324 -4201 338
rect -4235 252 -4201 270
rect -4235 180 -4201 202
rect -4235 105 -4201 134
rect -4087 984 -4053 1013
rect -4087 916 -4053 938
rect -4087 848 -4053 866
rect -4087 780 -4053 794
rect -4087 712 -4053 722
rect -4087 644 -4053 650
rect -4087 576 -4053 578
rect -4087 540 -4053 542
rect -4087 468 -4053 474
rect -4087 396 -4053 406
rect -4087 324 -4053 338
rect -4087 252 -4053 270
rect -4087 180 -4053 202
rect -4087 105 -4053 134
rect -3939 984 -3905 1013
rect -3939 916 -3905 938
rect -3939 848 -3905 866
rect -3939 780 -3905 794
rect -3939 712 -3905 722
rect -3939 644 -3905 650
rect -3939 576 -3905 578
rect -3939 540 -3905 542
rect -3939 468 -3905 474
rect -3939 396 -3905 406
rect -3939 324 -3905 338
rect -3939 252 -3905 270
rect -3939 180 -3905 202
rect -3939 105 -3905 134
rect -3791 984 -3757 1013
rect -3791 916 -3757 938
rect -3791 848 -3757 866
rect -3791 780 -3757 794
rect -3791 712 -3757 722
rect -3791 644 -3757 650
rect -3791 576 -3757 578
rect -3791 540 -3757 542
rect -3791 468 -3757 474
rect -3791 396 -3757 406
rect -3791 324 -3757 338
rect -3791 252 -3757 270
rect -3791 180 -3757 202
rect -3791 105 -3757 134
rect -3643 984 -3609 1013
rect -3643 916 -3609 938
rect -3643 848 -3609 866
rect -3643 780 -3609 794
rect -3643 712 -3609 722
rect -3643 644 -3609 650
rect -3643 576 -3609 578
rect -3643 540 -3609 542
rect -3643 468 -3609 474
rect -3643 396 -3609 406
rect -3643 324 -3609 338
rect -3643 252 -3609 270
rect -3643 180 -3609 202
rect -3643 105 -3609 134
rect -3495 984 -3461 1013
rect -3495 916 -3461 938
rect -3495 848 -3461 866
rect -3495 780 -3461 794
rect -3495 712 -3461 722
rect -3495 644 -3461 650
rect -3495 576 -3461 578
rect -3495 540 -3461 542
rect -3495 468 -3461 474
rect -3495 396 -3461 406
rect -3495 324 -3461 338
rect -3495 252 -3461 270
rect -3495 180 -3461 202
rect -3495 105 -3461 134
rect -3347 984 -3313 1013
rect -3347 916 -3313 938
rect -3347 848 -3313 866
rect -3347 780 -3313 794
rect -3347 712 -3313 722
rect -3347 644 -3313 650
rect -3347 576 -3313 578
rect -3347 540 -3313 542
rect -3347 468 -3313 474
rect -3347 396 -3313 406
rect -3347 324 -3313 338
rect -3347 252 -3313 270
rect -3347 180 -3313 202
rect -3347 105 -3313 134
rect -3199 984 -3165 1013
rect -3199 916 -3165 938
rect -3199 848 -3165 866
rect -3199 780 -3165 794
rect -3199 712 -3165 722
rect -3199 644 -3165 650
rect -3199 576 -3165 578
rect -3199 540 -3165 542
rect -3199 468 -3165 474
rect -3199 396 -3165 406
rect -3199 324 -3165 338
rect -3199 252 -3165 270
rect -3199 180 -3165 202
rect -3199 105 -3165 134
rect -3051 984 -3017 1013
rect -3051 916 -3017 938
rect -3051 848 -3017 866
rect -3051 780 -3017 794
rect -3051 712 -3017 722
rect -3051 644 -3017 650
rect -3051 576 -3017 578
rect -3051 540 -3017 542
rect -3051 468 -3017 474
rect -3051 396 -3017 406
rect -3051 324 -3017 338
rect -3051 252 -3017 270
rect -3051 180 -3017 202
rect -3051 105 -3017 134
rect -2903 984 -2869 1013
rect -2903 916 -2869 938
rect -2903 848 -2869 866
rect -2903 780 -2869 794
rect -2903 712 -2869 722
rect -2903 644 -2869 650
rect -2903 576 -2869 578
rect -2903 540 -2869 542
rect -2903 468 -2869 474
rect -2903 396 -2869 406
rect -2903 324 -2869 338
rect -2903 252 -2869 270
rect -2903 180 -2869 202
rect -2903 105 -2869 134
rect -2755 984 -2721 1013
rect -2755 916 -2721 938
rect -2755 848 -2721 866
rect -2755 780 -2721 794
rect -2755 712 -2721 722
rect -2755 644 -2721 650
rect -2755 576 -2721 578
rect -2755 540 -2721 542
rect -2755 468 -2721 474
rect -2755 396 -2721 406
rect -2755 324 -2721 338
rect -2755 252 -2721 270
rect -2755 180 -2721 202
rect -2755 105 -2721 134
rect -2607 984 -2573 1013
rect -2607 916 -2573 938
rect -2607 848 -2573 866
rect -2607 780 -2573 794
rect -2607 712 -2573 722
rect -2607 644 -2573 650
rect -2607 576 -2573 578
rect -2607 540 -2573 542
rect -2607 468 -2573 474
rect -2607 396 -2573 406
rect -2607 324 -2573 338
rect -2607 252 -2573 270
rect -2607 180 -2573 202
rect -2607 105 -2573 134
rect -2459 984 -2425 1013
rect -2459 916 -2425 938
rect -2459 848 -2425 866
rect -2459 780 -2425 794
rect -2459 712 -2425 722
rect -2459 644 -2425 650
rect -2459 576 -2425 578
rect -2459 540 -2425 542
rect -2459 468 -2425 474
rect -2459 396 -2425 406
rect -2459 324 -2425 338
rect -2459 252 -2425 270
rect -2459 180 -2425 202
rect -2459 105 -2425 134
rect -2311 984 -2277 1013
rect -2311 916 -2277 938
rect -2311 848 -2277 866
rect -2311 780 -2277 794
rect -2311 712 -2277 722
rect -2311 644 -2277 650
rect -2311 576 -2277 578
rect -2311 540 -2277 542
rect -2311 468 -2277 474
rect -2311 396 -2277 406
rect -2311 324 -2277 338
rect -2311 252 -2277 270
rect -2311 180 -2277 202
rect -2311 105 -2277 134
rect -2163 984 -2129 1013
rect -2163 916 -2129 938
rect -2163 848 -2129 866
rect -2163 780 -2129 794
rect -2163 712 -2129 722
rect -2163 644 -2129 650
rect -2163 576 -2129 578
rect -2163 540 -2129 542
rect -2163 468 -2129 474
rect -2163 396 -2129 406
rect -2163 324 -2129 338
rect -2163 252 -2129 270
rect -2163 180 -2129 202
rect -2163 105 -2129 134
rect -2015 984 -1981 1013
rect -2015 916 -1981 938
rect -2015 848 -1981 866
rect -2015 780 -1981 794
rect -2015 712 -1981 722
rect -2015 644 -1981 650
rect -2015 576 -1981 578
rect -2015 540 -1981 542
rect -2015 468 -1981 474
rect -2015 396 -1981 406
rect -2015 324 -1981 338
rect -2015 252 -1981 270
rect -2015 180 -1981 202
rect -2015 105 -1981 134
rect -1867 984 -1833 1013
rect -1867 916 -1833 938
rect -1867 848 -1833 866
rect -1867 780 -1833 794
rect -1867 712 -1833 722
rect -1867 644 -1833 650
rect -1867 576 -1833 578
rect -1867 540 -1833 542
rect -1867 468 -1833 474
rect -1867 396 -1833 406
rect -1867 324 -1833 338
rect -1867 252 -1833 270
rect -1867 180 -1833 202
rect -1867 105 -1833 134
rect -1719 984 -1685 1013
rect -1719 916 -1685 938
rect -1719 848 -1685 866
rect -1719 780 -1685 794
rect -1719 712 -1685 722
rect -1719 644 -1685 650
rect -1719 576 -1685 578
rect -1719 540 -1685 542
rect -1719 468 -1685 474
rect -1719 396 -1685 406
rect -1719 324 -1685 338
rect -1719 252 -1685 270
rect -1719 180 -1685 202
rect -1719 105 -1685 134
rect -1571 984 -1537 1013
rect -1571 916 -1537 938
rect -1571 848 -1537 866
rect -1571 780 -1537 794
rect -1571 712 -1537 722
rect -1571 644 -1537 650
rect -1571 576 -1537 578
rect -1571 540 -1537 542
rect -1571 468 -1537 474
rect -1571 396 -1537 406
rect -1571 324 -1537 338
rect -1571 252 -1537 270
rect -1571 180 -1537 202
rect -1571 105 -1537 134
rect -1423 984 -1389 1013
rect -1423 916 -1389 938
rect -1423 848 -1389 866
rect -1423 780 -1389 794
rect -1423 712 -1389 722
rect -1423 644 -1389 650
rect -1423 576 -1389 578
rect -1423 540 -1389 542
rect -1423 468 -1389 474
rect -1423 396 -1389 406
rect -1423 324 -1389 338
rect -1423 252 -1389 270
rect -1423 180 -1389 202
rect -1423 105 -1389 134
rect -1275 984 -1241 1013
rect -1275 916 -1241 938
rect -1275 848 -1241 866
rect -1275 780 -1241 794
rect -1275 712 -1241 722
rect -1275 644 -1241 650
rect -1275 576 -1241 578
rect -1275 540 -1241 542
rect -1275 468 -1241 474
rect -1275 396 -1241 406
rect -1275 324 -1241 338
rect -1275 252 -1241 270
rect -1275 180 -1241 202
rect -1275 105 -1241 134
rect -1127 984 -1093 1013
rect -1127 916 -1093 938
rect -1127 848 -1093 866
rect -1127 780 -1093 794
rect -1127 712 -1093 722
rect -1127 644 -1093 650
rect -1127 576 -1093 578
rect -1127 540 -1093 542
rect -1127 468 -1093 474
rect -1127 396 -1093 406
rect -1127 324 -1093 338
rect -1127 252 -1093 270
rect -1127 180 -1093 202
rect -1127 105 -1093 134
rect -979 984 -945 1013
rect -979 916 -945 938
rect -979 848 -945 866
rect -979 780 -945 794
rect -979 712 -945 722
rect -979 644 -945 650
rect -979 576 -945 578
rect -979 540 -945 542
rect -979 468 -945 474
rect -979 396 -945 406
rect -979 324 -945 338
rect -979 252 -945 270
rect -979 180 -945 202
rect -979 105 -945 134
rect -831 984 -797 1013
rect -831 916 -797 938
rect -831 848 -797 866
rect -831 780 -797 794
rect -831 712 -797 722
rect -831 644 -797 650
rect -831 576 -797 578
rect -831 540 -797 542
rect -831 468 -797 474
rect -831 396 -797 406
rect -831 324 -797 338
rect -831 252 -797 270
rect -831 180 -797 202
rect -831 105 -797 134
rect -683 984 -649 1013
rect -683 916 -649 938
rect -683 848 -649 866
rect -683 780 -649 794
rect -683 712 -649 722
rect -683 644 -649 650
rect -683 576 -649 578
rect -683 540 -649 542
rect -683 468 -649 474
rect -683 396 -649 406
rect -683 324 -649 338
rect -683 252 -649 270
rect -683 180 -649 202
rect -683 105 -649 134
rect -535 984 -501 1013
rect -535 916 -501 938
rect -535 848 -501 866
rect -535 780 -501 794
rect -535 712 -501 722
rect -535 644 -501 650
rect -535 576 -501 578
rect -535 540 -501 542
rect -535 468 -501 474
rect -535 396 -501 406
rect -535 324 -501 338
rect -535 252 -501 270
rect -535 180 -501 202
rect -535 105 -501 134
rect -387 984 -353 1013
rect -387 916 -353 938
rect -387 848 -353 866
rect -387 780 -353 794
rect -387 712 -353 722
rect -387 644 -353 650
rect -387 576 -353 578
rect -387 540 -353 542
rect -387 468 -353 474
rect -387 396 -353 406
rect -387 324 -353 338
rect -387 252 -353 270
rect -387 180 -353 202
rect -387 105 -353 134
rect -239 984 -205 1013
rect -239 916 -205 938
rect -239 848 -205 866
rect -239 780 -205 794
rect -239 712 -205 722
rect -239 644 -205 650
rect -239 576 -205 578
rect -239 540 -205 542
rect -239 468 -205 474
rect -239 396 -205 406
rect -239 324 -205 338
rect -239 252 -205 270
rect -239 180 -205 202
rect -239 105 -205 134
rect -91 984 -57 1013
rect -91 916 -57 938
rect -91 848 -57 866
rect -91 780 -57 794
rect -91 712 -57 722
rect -91 644 -57 650
rect -91 576 -57 578
rect -91 540 -57 542
rect -91 468 -57 474
rect -91 396 -57 406
rect -91 324 -57 338
rect -91 252 -57 270
rect -91 180 -57 202
rect -91 105 -57 134
rect 57 984 91 1013
rect 57 916 91 938
rect 57 848 91 866
rect 57 780 91 794
rect 57 712 91 722
rect 57 644 91 650
rect 57 576 91 578
rect 57 540 91 542
rect 57 468 91 474
rect 57 396 91 406
rect 57 324 91 338
rect 57 252 91 270
rect 57 180 91 202
rect 57 105 91 134
rect 205 984 239 1013
rect 205 916 239 938
rect 205 848 239 866
rect 205 780 239 794
rect 205 712 239 722
rect 205 644 239 650
rect 205 576 239 578
rect 205 540 239 542
rect 205 468 239 474
rect 205 396 239 406
rect 205 324 239 338
rect 205 252 239 270
rect 205 180 239 202
rect 205 105 239 134
rect 353 984 387 1013
rect 353 916 387 938
rect 353 848 387 866
rect 353 780 387 794
rect 353 712 387 722
rect 353 644 387 650
rect 353 576 387 578
rect 353 540 387 542
rect 353 468 387 474
rect 353 396 387 406
rect 353 324 387 338
rect 353 252 387 270
rect 353 180 387 202
rect 353 105 387 134
rect 501 984 535 1013
rect 501 916 535 938
rect 501 848 535 866
rect 501 780 535 794
rect 501 712 535 722
rect 501 644 535 650
rect 501 576 535 578
rect 501 540 535 542
rect 501 468 535 474
rect 501 396 535 406
rect 501 324 535 338
rect 501 252 535 270
rect 501 180 535 202
rect 501 105 535 134
rect 649 984 683 1013
rect 649 916 683 938
rect 649 848 683 866
rect 649 780 683 794
rect 649 712 683 722
rect 649 644 683 650
rect 649 576 683 578
rect 649 540 683 542
rect 649 468 683 474
rect 649 396 683 406
rect 649 324 683 338
rect 649 252 683 270
rect 649 180 683 202
rect 649 105 683 134
rect 797 984 831 1013
rect 797 916 831 938
rect 797 848 831 866
rect 797 780 831 794
rect 797 712 831 722
rect 797 644 831 650
rect 797 576 831 578
rect 797 540 831 542
rect 797 468 831 474
rect 797 396 831 406
rect 797 324 831 338
rect 797 252 831 270
rect 797 180 831 202
rect 797 105 831 134
rect 945 984 979 1013
rect 945 916 979 938
rect 945 848 979 866
rect 945 780 979 794
rect 945 712 979 722
rect 945 644 979 650
rect 945 576 979 578
rect 945 540 979 542
rect 945 468 979 474
rect 945 396 979 406
rect 945 324 979 338
rect 945 252 979 270
rect 945 180 979 202
rect 945 105 979 134
rect 1093 984 1127 1013
rect 1093 916 1127 938
rect 1093 848 1127 866
rect 1093 780 1127 794
rect 1093 712 1127 722
rect 1093 644 1127 650
rect 1093 576 1127 578
rect 1093 540 1127 542
rect 1093 468 1127 474
rect 1093 396 1127 406
rect 1093 324 1127 338
rect 1093 252 1127 270
rect 1093 180 1127 202
rect 1093 105 1127 134
rect 1241 984 1275 1013
rect 1241 916 1275 938
rect 1241 848 1275 866
rect 1241 780 1275 794
rect 1241 712 1275 722
rect 1241 644 1275 650
rect 1241 576 1275 578
rect 1241 540 1275 542
rect 1241 468 1275 474
rect 1241 396 1275 406
rect 1241 324 1275 338
rect 1241 252 1275 270
rect 1241 180 1275 202
rect 1241 105 1275 134
rect 1389 984 1423 1013
rect 1389 916 1423 938
rect 1389 848 1423 866
rect 1389 780 1423 794
rect 1389 712 1423 722
rect 1389 644 1423 650
rect 1389 576 1423 578
rect 1389 540 1423 542
rect 1389 468 1423 474
rect 1389 396 1423 406
rect 1389 324 1423 338
rect 1389 252 1423 270
rect 1389 180 1423 202
rect 1389 105 1423 134
rect 1537 984 1571 1013
rect 1537 916 1571 938
rect 1537 848 1571 866
rect 1537 780 1571 794
rect 1537 712 1571 722
rect 1537 644 1571 650
rect 1537 576 1571 578
rect 1537 540 1571 542
rect 1537 468 1571 474
rect 1537 396 1571 406
rect 1537 324 1571 338
rect 1537 252 1571 270
rect 1537 180 1571 202
rect 1537 105 1571 134
rect 1685 984 1719 1013
rect 1685 916 1719 938
rect 1685 848 1719 866
rect 1685 780 1719 794
rect 1685 712 1719 722
rect 1685 644 1719 650
rect 1685 576 1719 578
rect 1685 540 1719 542
rect 1685 468 1719 474
rect 1685 396 1719 406
rect 1685 324 1719 338
rect 1685 252 1719 270
rect 1685 180 1719 202
rect 1685 105 1719 134
rect 1833 984 1867 1013
rect 1833 916 1867 938
rect 1833 848 1867 866
rect 1833 780 1867 794
rect 1833 712 1867 722
rect 1833 644 1867 650
rect 1833 576 1867 578
rect 1833 540 1867 542
rect 1833 468 1867 474
rect 1833 396 1867 406
rect 1833 324 1867 338
rect 1833 252 1867 270
rect 1833 180 1867 202
rect 1833 105 1867 134
rect 1981 984 2015 1013
rect 1981 916 2015 938
rect 1981 848 2015 866
rect 1981 780 2015 794
rect 1981 712 2015 722
rect 1981 644 2015 650
rect 1981 576 2015 578
rect 1981 540 2015 542
rect 1981 468 2015 474
rect 1981 396 2015 406
rect 1981 324 2015 338
rect 1981 252 2015 270
rect 1981 180 2015 202
rect 1981 105 2015 134
rect 2129 984 2163 1013
rect 2129 916 2163 938
rect 2129 848 2163 866
rect 2129 780 2163 794
rect 2129 712 2163 722
rect 2129 644 2163 650
rect 2129 576 2163 578
rect 2129 540 2163 542
rect 2129 468 2163 474
rect 2129 396 2163 406
rect 2129 324 2163 338
rect 2129 252 2163 270
rect 2129 180 2163 202
rect 2129 105 2163 134
rect 2277 984 2311 1013
rect 2277 916 2311 938
rect 2277 848 2311 866
rect 2277 780 2311 794
rect 2277 712 2311 722
rect 2277 644 2311 650
rect 2277 576 2311 578
rect 2277 540 2311 542
rect 2277 468 2311 474
rect 2277 396 2311 406
rect 2277 324 2311 338
rect 2277 252 2311 270
rect 2277 180 2311 202
rect 2277 105 2311 134
rect 2425 984 2459 1013
rect 2425 916 2459 938
rect 2425 848 2459 866
rect 2425 780 2459 794
rect 2425 712 2459 722
rect 2425 644 2459 650
rect 2425 576 2459 578
rect 2425 540 2459 542
rect 2425 468 2459 474
rect 2425 396 2459 406
rect 2425 324 2459 338
rect 2425 252 2459 270
rect 2425 180 2459 202
rect 2425 105 2459 134
rect 2573 984 2607 1013
rect 2573 916 2607 938
rect 2573 848 2607 866
rect 2573 780 2607 794
rect 2573 712 2607 722
rect 2573 644 2607 650
rect 2573 576 2607 578
rect 2573 540 2607 542
rect 2573 468 2607 474
rect 2573 396 2607 406
rect 2573 324 2607 338
rect 2573 252 2607 270
rect 2573 180 2607 202
rect 2573 105 2607 134
rect 2721 984 2755 1013
rect 2721 916 2755 938
rect 2721 848 2755 866
rect 2721 780 2755 794
rect 2721 712 2755 722
rect 2721 644 2755 650
rect 2721 576 2755 578
rect 2721 540 2755 542
rect 2721 468 2755 474
rect 2721 396 2755 406
rect 2721 324 2755 338
rect 2721 252 2755 270
rect 2721 180 2755 202
rect 2721 105 2755 134
rect 2869 984 2903 1013
rect 2869 916 2903 938
rect 2869 848 2903 866
rect 2869 780 2903 794
rect 2869 712 2903 722
rect 2869 644 2903 650
rect 2869 576 2903 578
rect 2869 540 2903 542
rect 2869 468 2903 474
rect 2869 396 2903 406
rect 2869 324 2903 338
rect 2869 252 2903 270
rect 2869 180 2903 202
rect 2869 105 2903 134
rect 3017 984 3051 1013
rect 3017 916 3051 938
rect 3017 848 3051 866
rect 3017 780 3051 794
rect 3017 712 3051 722
rect 3017 644 3051 650
rect 3017 576 3051 578
rect 3017 540 3051 542
rect 3017 468 3051 474
rect 3017 396 3051 406
rect 3017 324 3051 338
rect 3017 252 3051 270
rect 3017 180 3051 202
rect 3017 105 3051 134
rect 3165 984 3199 1013
rect 3165 916 3199 938
rect 3165 848 3199 866
rect 3165 780 3199 794
rect 3165 712 3199 722
rect 3165 644 3199 650
rect 3165 576 3199 578
rect 3165 540 3199 542
rect 3165 468 3199 474
rect 3165 396 3199 406
rect 3165 324 3199 338
rect 3165 252 3199 270
rect 3165 180 3199 202
rect 3165 105 3199 134
rect 3313 984 3347 1013
rect 3313 916 3347 938
rect 3313 848 3347 866
rect 3313 780 3347 794
rect 3313 712 3347 722
rect 3313 644 3347 650
rect 3313 576 3347 578
rect 3313 540 3347 542
rect 3313 468 3347 474
rect 3313 396 3347 406
rect 3313 324 3347 338
rect 3313 252 3347 270
rect 3313 180 3347 202
rect 3313 105 3347 134
rect 3461 984 3495 1013
rect 3461 916 3495 938
rect 3461 848 3495 866
rect 3461 780 3495 794
rect 3461 712 3495 722
rect 3461 644 3495 650
rect 3461 576 3495 578
rect 3461 540 3495 542
rect 3461 468 3495 474
rect 3461 396 3495 406
rect 3461 324 3495 338
rect 3461 252 3495 270
rect 3461 180 3495 202
rect 3461 105 3495 134
rect 3609 984 3643 1013
rect 3609 916 3643 938
rect 3609 848 3643 866
rect 3609 780 3643 794
rect 3609 712 3643 722
rect 3609 644 3643 650
rect 3609 576 3643 578
rect 3609 540 3643 542
rect 3609 468 3643 474
rect 3609 396 3643 406
rect 3609 324 3643 338
rect 3609 252 3643 270
rect 3609 180 3643 202
rect 3609 105 3643 134
rect 3757 984 3791 1013
rect 3757 916 3791 938
rect 3757 848 3791 866
rect 3757 780 3791 794
rect 3757 712 3791 722
rect 3757 644 3791 650
rect 3757 576 3791 578
rect 3757 540 3791 542
rect 3757 468 3791 474
rect 3757 396 3791 406
rect 3757 324 3791 338
rect 3757 252 3791 270
rect 3757 180 3791 202
rect 3757 105 3791 134
rect 3905 984 3939 1013
rect 3905 916 3939 938
rect 3905 848 3939 866
rect 3905 780 3939 794
rect 3905 712 3939 722
rect 3905 644 3939 650
rect 3905 576 3939 578
rect 3905 540 3939 542
rect 3905 468 3939 474
rect 3905 396 3939 406
rect 3905 324 3939 338
rect 3905 252 3939 270
rect 3905 180 3939 202
rect 3905 105 3939 134
rect 4053 984 4087 1013
rect 4053 916 4087 938
rect 4053 848 4087 866
rect 4053 780 4087 794
rect 4053 712 4087 722
rect 4053 644 4087 650
rect 4053 576 4087 578
rect 4053 540 4087 542
rect 4053 468 4087 474
rect 4053 396 4087 406
rect 4053 324 4087 338
rect 4053 252 4087 270
rect 4053 180 4087 202
rect 4053 105 4087 134
rect 4201 984 4235 1013
rect 4201 916 4235 938
rect 4201 848 4235 866
rect 4201 780 4235 794
rect 4201 712 4235 722
rect 4201 644 4235 650
rect 4201 576 4235 578
rect 4201 540 4235 542
rect 4201 468 4235 474
rect 4201 396 4235 406
rect 4201 324 4235 338
rect 4201 252 4235 270
rect 4201 180 4235 202
rect 4201 105 4235 134
rect 4349 984 4383 1013
rect 4349 916 4383 938
rect 4349 848 4383 866
rect 4349 780 4383 794
rect 4349 712 4383 722
rect 4349 644 4383 650
rect 4349 576 4383 578
rect 4349 540 4383 542
rect 4349 468 4383 474
rect 4349 396 4383 406
rect 4349 324 4383 338
rect 4349 252 4383 270
rect 4349 180 4383 202
rect 4349 105 4383 134
rect 4497 984 4531 1013
rect 4497 916 4531 938
rect 4497 848 4531 866
rect 4497 780 4531 794
rect 4497 712 4531 722
rect 4497 644 4531 650
rect 4497 576 4531 578
rect 4497 540 4531 542
rect 4497 468 4531 474
rect 4497 396 4531 406
rect 4497 324 4531 338
rect 4497 252 4531 270
rect 4497 180 4531 202
rect 4497 105 4531 134
rect 4645 984 4679 1013
rect 4645 916 4679 938
rect 4645 848 4679 866
rect 4645 780 4679 794
rect 4645 712 4679 722
rect 4645 644 4679 650
rect 4645 576 4679 578
rect 4645 540 4679 542
rect 4645 468 4679 474
rect 4645 396 4679 406
rect 4645 324 4679 338
rect 4645 252 4679 270
rect 4645 180 4679 202
rect 4645 105 4679 134
rect 4793 984 4827 1013
rect 4793 916 4827 938
rect 4793 848 4827 866
rect 4793 780 4827 794
rect 4793 712 4827 722
rect 4793 644 4827 650
rect 4793 576 4827 578
rect 4793 540 4827 542
rect 4793 468 4827 474
rect 4793 396 4827 406
rect 4793 324 4827 338
rect 4793 252 4827 270
rect 4793 180 4827 202
rect 4793 105 4827 134
rect 4941 984 4975 1013
rect 4941 916 4975 938
rect 4941 848 4975 866
rect 4941 780 4975 794
rect 4941 712 4975 722
rect 4941 644 4975 650
rect 4941 576 4975 578
rect 4941 540 4975 542
rect 4941 468 4975 474
rect 4941 396 4975 406
rect 4941 324 4975 338
rect 4941 252 4975 270
rect 4941 180 4975 202
rect 4941 105 4975 134
rect 5089 984 5123 1013
rect 5089 916 5123 938
rect 5089 848 5123 866
rect 5089 780 5123 794
rect 5089 712 5123 722
rect 5089 644 5123 650
rect 5089 576 5123 578
rect 5089 540 5123 542
rect 5089 468 5123 474
rect 5089 396 5123 406
rect 5089 324 5123 338
rect 5089 252 5123 270
rect 5089 180 5123 202
rect 5089 105 5123 134
rect 5237 984 5271 1013
rect 5237 916 5271 938
rect 5237 848 5271 866
rect 5237 780 5271 794
rect 5237 712 5271 722
rect 5237 644 5271 650
rect 5237 576 5271 578
rect 5237 540 5271 542
rect 5237 468 5271 474
rect 5237 396 5271 406
rect 5237 324 5271 338
rect 5237 252 5271 270
rect 5237 180 5271 202
rect 5237 105 5271 134
rect 5385 984 5419 1013
rect 5385 916 5419 938
rect 5385 848 5419 866
rect 5385 780 5419 794
rect 5385 712 5419 722
rect 5385 644 5419 650
rect 5385 576 5419 578
rect 5385 540 5419 542
rect 5385 468 5419 474
rect 5385 396 5419 406
rect 5385 324 5419 338
rect 5385 252 5419 270
rect 5385 180 5419 202
rect 5385 105 5419 134
rect 5533 984 5567 1013
rect 5533 916 5567 938
rect 5533 848 5567 866
rect 5533 780 5567 794
rect 5533 712 5567 722
rect 5533 644 5567 650
rect 5533 576 5567 578
rect 5533 540 5567 542
rect 5533 468 5567 474
rect 5533 396 5567 406
rect 5533 324 5567 338
rect 5533 252 5567 270
rect 5533 180 5567 202
rect 5533 105 5567 134
rect 5647 1003 5681 1037
rect 5647 935 5681 969
rect 5647 867 5681 901
rect 5647 799 5681 833
rect 5647 731 5681 765
rect 5647 663 5681 697
rect 5647 595 5681 629
rect 5647 527 5681 561
rect 5647 459 5681 493
rect 5647 391 5681 425
rect 5647 323 5681 357
rect 5647 255 5681 289
rect 5647 187 5681 221
rect 5647 119 5681 153
rect -5681 51 -5647 85
rect -5521 37 -5493 71
rect -5459 37 -5431 71
rect -5373 37 -5345 71
rect -5311 37 -5283 71
rect -5225 37 -5197 71
rect -5163 37 -5135 71
rect -5077 37 -5049 71
rect -5015 37 -4987 71
rect -4929 37 -4901 71
rect -4867 37 -4839 71
rect -4781 37 -4753 71
rect -4719 37 -4691 71
rect -4633 37 -4605 71
rect -4571 37 -4543 71
rect -4485 37 -4457 71
rect -4423 37 -4395 71
rect -4337 37 -4309 71
rect -4275 37 -4247 71
rect -4189 37 -4161 71
rect -4127 37 -4099 71
rect -4041 37 -4013 71
rect -3979 37 -3951 71
rect -3893 37 -3865 71
rect -3831 37 -3803 71
rect -3745 37 -3717 71
rect -3683 37 -3655 71
rect -3597 37 -3569 71
rect -3535 37 -3507 71
rect -3449 37 -3421 71
rect -3387 37 -3359 71
rect -3301 37 -3273 71
rect -3239 37 -3211 71
rect -3153 37 -3125 71
rect -3091 37 -3063 71
rect -3005 37 -2977 71
rect -2943 37 -2915 71
rect -2857 37 -2829 71
rect -2795 37 -2767 71
rect -2709 37 -2681 71
rect -2647 37 -2619 71
rect -2561 37 -2533 71
rect -2499 37 -2471 71
rect -2413 37 -2385 71
rect -2351 37 -2323 71
rect -2265 37 -2237 71
rect -2203 37 -2175 71
rect -2117 37 -2089 71
rect -2055 37 -2027 71
rect -1969 37 -1941 71
rect -1907 37 -1879 71
rect -1821 37 -1793 71
rect -1759 37 -1731 71
rect -1673 37 -1645 71
rect -1611 37 -1583 71
rect -1525 37 -1497 71
rect -1463 37 -1435 71
rect -1377 37 -1349 71
rect -1315 37 -1287 71
rect -1229 37 -1201 71
rect -1167 37 -1139 71
rect -1081 37 -1053 71
rect -1019 37 -991 71
rect -933 37 -905 71
rect -871 37 -843 71
rect -785 37 -757 71
rect -723 37 -695 71
rect -637 37 -609 71
rect -575 37 -547 71
rect -489 37 -461 71
rect -427 37 -399 71
rect -341 37 -313 71
rect -279 37 -251 71
rect -193 37 -165 71
rect -131 37 -103 71
rect -45 37 -17 71
rect 17 37 45 71
rect 103 37 131 71
rect 165 37 193 71
rect 251 37 279 71
rect 313 37 341 71
rect 399 37 427 71
rect 461 37 489 71
rect 547 37 575 71
rect 609 37 637 71
rect 695 37 723 71
rect 757 37 785 71
rect 843 37 871 71
rect 905 37 933 71
rect 991 37 1019 71
rect 1053 37 1081 71
rect 1139 37 1167 71
rect 1201 37 1229 71
rect 1287 37 1315 71
rect 1349 37 1377 71
rect 1435 37 1463 71
rect 1497 37 1525 71
rect 1583 37 1611 71
rect 1645 37 1673 71
rect 1731 37 1759 71
rect 1793 37 1821 71
rect 1879 37 1907 71
rect 1941 37 1969 71
rect 2027 37 2055 71
rect 2089 37 2117 71
rect 2175 37 2203 71
rect 2237 37 2265 71
rect 2323 37 2351 71
rect 2385 37 2413 71
rect 2471 37 2499 71
rect 2533 37 2561 71
rect 2619 37 2647 71
rect 2681 37 2709 71
rect 2767 37 2795 71
rect 2829 37 2857 71
rect 2915 37 2943 71
rect 2977 37 3005 71
rect 3063 37 3091 71
rect 3125 37 3153 71
rect 3211 37 3239 71
rect 3273 37 3301 71
rect 3359 37 3387 71
rect 3421 37 3449 71
rect 3507 37 3535 71
rect 3569 37 3597 71
rect 3655 37 3683 71
rect 3717 37 3745 71
rect 3803 37 3831 71
rect 3865 37 3893 71
rect 3951 37 3979 71
rect 4013 37 4041 71
rect 4099 37 4127 71
rect 4161 37 4189 71
rect 4247 37 4275 71
rect 4309 37 4337 71
rect 4395 37 4423 71
rect 4457 37 4485 71
rect 4543 37 4571 71
rect 4605 37 4633 71
rect 4691 37 4719 71
rect 4753 37 4781 71
rect 4839 37 4867 71
rect 4901 37 4929 71
rect 4987 37 5015 71
rect 5049 37 5077 71
rect 5135 37 5163 71
rect 5197 37 5225 71
rect 5283 37 5311 71
rect 5345 37 5373 71
rect 5431 37 5459 71
rect 5493 37 5521 71
rect 5647 51 5681 85
rect -5681 -17 -5647 17
rect 5647 -17 5681 17
rect -5681 -85 -5647 -51
rect -5521 -71 -5493 -37
rect -5459 -71 -5431 -37
rect -5373 -71 -5345 -37
rect -5311 -71 -5283 -37
rect -5225 -71 -5197 -37
rect -5163 -71 -5135 -37
rect -5077 -71 -5049 -37
rect -5015 -71 -4987 -37
rect -4929 -71 -4901 -37
rect -4867 -71 -4839 -37
rect -4781 -71 -4753 -37
rect -4719 -71 -4691 -37
rect -4633 -71 -4605 -37
rect -4571 -71 -4543 -37
rect -4485 -71 -4457 -37
rect -4423 -71 -4395 -37
rect -4337 -71 -4309 -37
rect -4275 -71 -4247 -37
rect -4189 -71 -4161 -37
rect -4127 -71 -4099 -37
rect -4041 -71 -4013 -37
rect -3979 -71 -3951 -37
rect -3893 -71 -3865 -37
rect -3831 -71 -3803 -37
rect -3745 -71 -3717 -37
rect -3683 -71 -3655 -37
rect -3597 -71 -3569 -37
rect -3535 -71 -3507 -37
rect -3449 -71 -3421 -37
rect -3387 -71 -3359 -37
rect -3301 -71 -3273 -37
rect -3239 -71 -3211 -37
rect -3153 -71 -3125 -37
rect -3091 -71 -3063 -37
rect -3005 -71 -2977 -37
rect -2943 -71 -2915 -37
rect -2857 -71 -2829 -37
rect -2795 -71 -2767 -37
rect -2709 -71 -2681 -37
rect -2647 -71 -2619 -37
rect -2561 -71 -2533 -37
rect -2499 -71 -2471 -37
rect -2413 -71 -2385 -37
rect -2351 -71 -2323 -37
rect -2265 -71 -2237 -37
rect -2203 -71 -2175 -37
rect -2117 -71 -2089 -37
rect -2055 -71 -2027 -37
rect -1969 -71 -1941 -37
rect -1907 -71 -1879 -37
rect -1821 -71 -1793 -37
rect -1759 -71 -1731 -37
rect -1673 -71 -1645 -37
rect -1611 -71 -1583 -37
rect -1525 -71 -1497 -37
rect -1463 -71 -1435 -37
rect -1377 -71 -1349 -37
rect -1315 -71 -1287 -37
rect -1229 -71 -1201 -37
rect -1167 -71 -1139 -37
rect -1081 -71 -1053 -37
rect -1019 -71 -991 -37
rect -933 -71 -905 -37
rect -871 -71 -843 -37
rect -785 -71 -757 -37
rect -723 -71 -695 -37
rect -637 -71 -609 -37
rect -575 -71 -547 -37
rect -489 -71 -461 -37
rect -427 -71 -399 -37
rect -341 -71 -313 -37
rect -279 -71 -251 -37
rect -193 -71 -165 -37
rect -131 -71 -103 -37
rect -45 -71 -17 -37
rect 17 -71 45 -37
rect 103 -71 131 -37
rect 165 -71 193 -37
rect 251 -71 279 -37
rect 313 -71 341 -37
rect 399 -71 427 -37
rect 461 -71 489 -37
rect 547 -71 575 -37
rect 609 -71 637 -37
rect 695 -71 723 -37
rect 757 -71 785 -37
rect 843 -71 871 -37
rect 905 -71 933 -37
rect 991 -71 1019 -37
rect 1053 -71 1081 -37
rect 1139 -71 1167 -37
rect 1201 -71 1229 -37
rect 1287 -71 1315 -37
rect 1349 -71 1377 -37
rect 1435 -71 1463 -37
rect 1497 -71 1525 -37
rect 1583 -71 1611 -37
rect 1645 -71 1673 -37
rect 1731 -71 1759 -37
rect 1793 -71 1821 -37
rect 1879 -71 1907 -37
rect 1941 -71 1969 -37
rect 2027 -71 2055 -37
rect 2089 -71 2117 -37
rect 2175 -71 2203 -37
rect 2237 -71 2265 -37
rect 2323 -71 2351 -37
rect 2385 -71 2413 -37
rect 2471 -71 2499 -37
rect 2533 -71 2561 -37
rect 2619 -71 2647 -37
rect 2681 -71 2709 -37
rect 2767 -71 2795 -37
rect 2829 -71 2857 -37
rect 2915 -71 2943 -37
rect 2977 -71 3005 -37
rect 3063 -71 3091 -37
rect 3125 -71 3153 -37
rect 3211 -71 3239 -37
rect 3273 -71 3301 -37
rect 3359 -71 3387 -37
rect 3421 -71 3449 -37
rect 3507 -71 3535 -37
rect 3569 -71 3597 -37
rect 3655 -71 3683 -37
rect 3717 -71 3745 -37
rect 3803 -71 3831 -37
rect 3865 -71 3893 -37
rect 3951 -71 3979 -37
rect 4013 -71 4041 -37
rect 4099 -71 4127 -37
rect 4161 -71 4189 -37
rect 4247 -71 4275 -37
rect 4309 -71 4337 -37
rect 4395 -71 4423 -37
rect 4457 -71 4485 -37
rect 4543 -71 4571 -37
rect 4605 -71 4633 -37
rect 4691 -71 4719 -37
rect 4753 -71 4781 -37
rect 4839 -71 4867 -37
rect 4901 -71 4929 -37
rect 4987 -71 5015 -37
rect 5049 -71 5077 -37
rect 5135 -71 5163 -37
rect 5197 -71 5225 -37
rect 5283 -71 5311 -37
rect 5345 -71 5373 -37
rect 5431 -71 5459 -37
rect 5493 -71 5521 -37
rect 5647 -85 5681 -51
rect -5681 -153 -5647 -119
rect -5681 -221 -5647 -187
rect -5681 -289 -5647 -255
rect -5681 -357 -5647 -323
rect -5681 -425 -5647 -391
rect -5681 -493 -5647 -459
rect -5681 -561 -5647 -527
rect -5681 -629 -5647 -595
rect -5681 -697 -5647 -663
rect -5681 -765 -5647 -731
rect -5681 -833 -5647 -799
rect -5681 -901 -5647 -867
rect -5681 -969 -5647 -935
rect -5681 -1037 -5647 -1003
rect -5567 -134 -5533 -105
rect -5567 -202 -5533 -180
rect -5567 -270 -5533 -252
rect -5567 -338 -5533 -324
rect -5567 -406 -5533 -396
rect -5567 -474 -5533 -468
rect -5567 -542 -5533 -540
rect -5567 -578 -5533 -576
rect -5567 -650 -5533 -644
rect -5567 -722 -5533 -712
rect -5567 -794 -5533 -780
rect -5567 -866 -5533 -848
rect -5567 -938 -5533 -916
rect -5567 -1013 -5533 -984
rect -5419 -134 -5385 -105
rect -5419 -202 -5385 -180
rect -5419 -270 -5385 -252
rect -5419 -338 -5385 -324
rect -5419 -406 -5385 -396
rect -5419 -474 -5385 -468
rect -5419 -542 -5385 -540
rect -5419 -578 -5385 -576
rect -5419 -650 -5385 -644
rect -5419 -722 -5385 -712
rect -5419 -794 -5385 -780
rect -5419 -866 -5385 -848
rect -5419 -938 -5385 -916
rect -5419 -1013 -5385 -984
rect -5271 -134 -5237 -105
rect -5271 -202 -5237 -180
rect -5271 -270 -5237 -252
rect -5271 -338 -5237 -324
rect -5271 -406 -5237 -396
rect -5271 -474 -5237 -468
rect -5271 -542 -5237 -540
rect -5271 -578 -5237 -576
rect -5271 -650 -5237 -644
rect -5271 -722 -5237 -712
rect -5271 -794 -5237 -780
rect -5271 -866 -5237 -848
rect -5271 -938 -5237 -916
rect -5271 -1013 -5237 -984
rect -5123 -134 -5089 -105
rect -5123 -202 -5089 -180
rect -5123 -270 -5089 -252
rect -5123 -338 -5089 -324
rect -5123 -406 -5089 -396
rect -5123 -474 -5089 -468
rect -5123 -542 -5089 -540
rect -5123 -578 -5089 -576
rect -5123 -650 -5089 -644
rect -5123 -722 -5089 -712
rect -5123 -794 -5089 -780
rect -5123 -866 -5089 -848
rect -5123 -938 -5089 -916
rect -5123 -1013 -5089 -984
rect -4975 -134 -4941 -105
rect -4975 -202 -4941 -180
rect -4975 -270 -4941 -252
rect -4975 -338 -4941 -324
rect -4975 -406 -4941 -396
rect -4975 -474 -4941 -468
rect -4975 -542 -4941 -540
rect -4975 -578 -4941 -576
rect -4975 -650 -4941 -644
rect -4975 -722 -4941 -712
rect -4975 -794 -4941 -780
rect -4975 -866 -4941 -848
rect -4975 -938 -4941 -916
rect -4975 -1013 -4941 -984
rect -4827 -134 -4793 -105
rect -4827 -202 -4793 -180
rect -4827 -270 -4793 -252
rect -4827 -338 -4793 -324
rect -4827 -406 -4793 -396
rect -4827 -474 -4793 -468
rect -4827 -542 -4793 -540
rect -4827 -578 -4793 -576
rect -4827 -650 -4793 -644
rect -4827 -722 -4793 -712
rect -4827 -794 -4793 -780
rect -4827 -866 -4793 -848
rect -4827 -938 -4793 -916
rect -4827 -1013 -4793 -984
rect -4679 -134 -4645 -105
rect -4679 -202 -4645 -180
rect -4679 -270 -4645 -252
rect -4679 -338 -4645 -324
rect -4679 -406 -4645 -396
rect -4679 -474 -4645 -468
rect -4679 -542 -4645 -540
rect -4679 -578 -4645 -576
rect -4679 -650 -4645 -644
rect -4679 -722 -4645 -712
rect -4679 -794 -4645 -780
rect -4679 -866 -4645 -848
rect -4679 -938 -4645 -916
rect -4679 -1013 -4645 -984
rect -4531 -134 -4497 -105
rect -4531 -202 -4497 -180
rect -4531 -270 -4497 -252
rect -4531 -338 -4497 -324
rect -4531 -406 -4497 -396
rect -4531 -474 -4497 -468
rect -4531 -542 -4497 -540
rect -4531 -578 -4497 -576
rect -4531 -650 -4497 -644
rect -4531 -722 -4497 -712
rect -4531 -794 -4497 -780
rect -4531 -866 -4497 -848
rect -4531 -938 -4497 -916
rect -4531 -1013 -4497 -984
rect -4383 -134 -4349 -105
rect -4383 -202 -4349 -180
rect -4383 -270 -4349 -252
rect -4383 -338 -4349 -324
rect -4383 -406 -4349 -396
rect -4383 -474 -4349 -468
rect -4383 -542 -4349 -540
rect -4383 -578 -4349 -576
rect -4383 -650 -4349 -644
rect -4383 -722 -4349 -712
rect -4383 -794 -4349 -780
rect -4383 -866 -4349 -848
rect -4383 -938 -4349 -916
rect -4383 -1013 -4349 -984
rect -4235 -134 -4201 -105
rect -4235 -202 -4201 -180
rect -4235 -270 -4201 -252
rect -4235 -338 -4201 -324
rect -4235 -406 -4201 -396
rect -4235 -474 -4201 -468
rect -4235 -542 -4201 -540
rect -4235 -578 -4201 -576
rect -4235 -650 -4201 -644
rect -4235 -722 -4201 -712
rect -4235 -794 -4201 -780
rect -4235 -866 -4201 -848
rect -4235 -938 -4201 -916
rect -4235 -1013 -4201 -984
rect -4087 -134 -4053 -105
rect -4087 -202 -4053 -180
rect -4087 -270 -4053 -252
rect -4087 -338 -4053 -324
rect -4087 -406 -4053 -396
rect -4087 -474 -4053 -468
rect -4087 -542 -4053 -540
rect -4087 -578 -4053 -576
rect -4087 -650 -4053 -644
rect -4087 -722 -4053 -712
rect -4087 -794 -4053 -780
rect -4087 -866 -4053 -848
rect -4087 -938 -4053 -916
rect -4087 -1013 -4053 -984
rect -3939 -134 -3905 -105
rect -3939 -202 -3905 -180
rect -3939 -270 -3905 -252
rect -3939 -338 -3905 -324
rect -3939 -406 -3905 -396
rect -3939 -474 -3905 -468
rect -3939 -542 -3905 -540
rect -3939 -578 -3905 -576
rect -3939 -650 -3905 -644
rect -3939 -722 -3905 -712
rect -3939 -794 -3905 -780
rect -3939 -866 -3905 -848
rect -3939 -938 -3905 -916
rect -3939 -1013 -3905 -984
rect -3791 -134 -3757 -105
rect -3791 -202 -3757 -180
rect -3791 -270 -3757 -252
rect -3791 -338 -3757 -324
rect -3791 -406 -3757 -396
rect -3791 -474 -3757 -468
rect -3791 -542 -3757 -540
rect -3791 -578 -3757 -576
rect -3791 -650 -3757 -644
rect -3791 -722 -3757 -712
rect -3791 -794 -3757 -780
rect -3791 -866 -3757 -848
rect -3791 -938 -3757 -916
rect -3791 -1013 -3757 -984
rect -3643 -134 -3609 -105
rect -3643 -202 -3609 -180
rect -3643 -270 -3609 -252
rect -3643 -338 -3609 -324
rect -3643 -406 -3609 -396
rect -3643 -474 -3609 -468
rect -3643 -542 -3609 -540
rect -3643 -578 -3609 -576
rect -3643 -650 -3609 -644
rect -3643 -722 -3609 -712
rect -3643 -794 -3609 -780
rect -3643 -866 -3609 -848
rect -3643 -938 -3609 -916
rect -3643 -1013 -3609 -984
rect -3495 -134 -3461 -105
rect -3495 -202 -3461 -180
rect -3495 -270 -3461 -252
rect -3495 -338 -3461 -324
rect -3495 -406 -3461 -396
rect -3495 -474 -3461 -468
rect -3495 -542 -3461 -540
rect -3495 -578 -3461 -576
rect -3495 -650 -3461 -644
rect -3495 -722 -3461 -712
rect -3495 -794 -3461 -780
rect -3495 -866 -3461 -848
rect -3495 -938 -3461 -916
rect -3495 -1013 -3461 -984
rect -3347 -134 -3313 -105
rect -3347 -202 -3313 -180
rect -3347 -270 -3313 -252
rect -3347 -338 -3313 -324
rect -3347 -406 -3313 -396
rect -3347 -474 -3313 -468
rect -3347 -542 -3313 -540
rect -3347 -578 -3313 -576
rect -3347 -650 -3313 -644
rect -3347 -722 -3313 -712
rect -3347 -794 -3313 -780
rect -3347 -866 -3313 -848
rect -3347 -938 -3313 -916
rect -3347 -1013 -3313 -984
rect -3199 -134 -3165 -105
rect -3199 -202 -3165 -180
rect -3199 -270 -3165 -252
rect -3199 -338 -3165 -324
rect -3199 -406 -3165 -396
rect -3199 -474 -3165 -468
rect -3199 -542 -3165 -540
rect -3199 -578 -3165 -576
rect -3199 -650 -3165 -644
rect -3199 -722 -3165 -712
rect -3199 -794 -3165 -780
rect -3199 -866 -3165 -848
rect -3199 -938 -3165 -916
rect -3199 -1013 -3165 -984
rect -3051 -134 -3017 -105
rect -3051 -202 -3017 -180
rect -3051 -270 -3017 -252
rect -3051 -338 -3017 -324
rect -3051 -406 -3017 -396
rect -3051 -474 -3017 -468
rect -3051 -542 -3017 -540
rect -3051 -578 -3017 -576
rect -3051 -650 -3017 -644
rect -3051 -722 -3017 -712
rect -3051 -794 -3017 -780
rect -3051 -866 -3017 -848
rect -3051 -938 -3017 -916
rect -3051 -1013 -3017 -984
rect -2903 -134 -2869 -105
rect -2903 -202 -2869 -180
rect -2903 -270 -2869 -252
rect -2903 -338 -2869 -324
rect -2903 -406 -2869 -396
rect -2903 -474 -2869 -468
rect -2903 -542 -2869 -540
rect -2903 -578 -2869 -576
rect -2903 -650 -2869 -644
rect -2903 -722 -2869 -712
rect -2903 -794 -2869 -780
rect -2903 -866 -2869 -848
rect -2903 -938 -2869 -916
rect -2903 -1013 -2869 -984
rect -2755 -134 -2721 -105
rect -2755 -202 -2721 -180
rect -2755 -270 -2721 -252
rect -2755 -338 -2721 -324
rect -2755 -406 -2721 -396
rect -2755 -474 -2721 -468
rect -2755 -542 -2721 -540
rect -2755 -578 -2721 -576
rect -2755 -650 -2721 -644
rect -2755 -722 -2721 -712
rect -2755 -794 -2721 -780
rect -2755 -866 -2721 -848
rect -2755 -938 -2721 -916
rect -2755 -1013 -2721 -984
rect -2607 -134 -2573 -105
rect -2607 -202 -2573 -180
rect -2607 -270 -2573 -252
rect -2607 -338 -2573 -324
rect -2607 -406 -2573 -396
rect -2607 -474 -2573 -468
rect -2607 -542 -2573 -540
rect -2607 -578 -2573 -576
rect -2607 -650 -2573 -644
rect -2607 -722 -2573 -712
rect -2607 -794 -2573 -780
rect -2607 -866 -2573 -848
rect -2607 -938 -2573 -916
rect -2607 -1013 -2573 -984
rect -2459 -134 -2425 -105
rect -2459 -202 -2425 -180
rect -2459 -270 -2425 -252
rect -2459 -338 -2425 -324
rect -2459 -406 -2425 -396
rect -2459 -474 -2425 -468
rect -2459 -542 -2425 -540
rect -2459 -578 -2425 -576
rect -2459 -650 -2425 -644
rect -2459 -722 -2425 -712
rect -2459 -794 -2425 -780
rect -2459 -866 -2425 -848
rect -2459 -938 -2425 -916
rect -2459 -1013 -2425 -984
rect -2311 -134 -2277 -105
rect -2311 -202 -2277 -180
rect -2311 -270 -2277 -252
rect -2311 -338 -2277 -324
rect -2311 -406 -2277 -396
rect -2311 -474 -2277 -468
rect -2311 -542 -2277 -540
rect -2311 -578 -2277 -576
rect -2311 -650 -2277 -644
rect -2311 -722 -2277 -712
rect -2311 -794 -2277 -780
rect -2311 -866 -2277 -848
rect -2311 -938 -2277 -916
rect -2311 -1013 -2277 -984
rect -2163 -134 -2129 -105
rect -2163 -202 -2129 -180
rect -2163 -270 -2129 -252
rect -2163 -338 -2129 -324
rect -2163 -406 -2129 -396
rect -2163 -474 -2129 -468
rect -2163 -542 -2129 -540
rect -2163 -578 -2129 -576
rect -2163 -650 -2129 -644
rect -2163 -722 -2129 -712
rect -2163 -794 -2129 -780
rect -2163 -866 -2129 -848
rect -2163 -938 -2129 -916
rect -2163 -1013 -2129 -984
rect -2015 -134 -1981 -105
rect -2015 -202 -1981 -180
rect -2015 -270 -1981 -252
rect -2015 -338 -1981 -324
rect -2015 -406 -1981 -396
rect -2015 -474 -1981 -468
rect -2015 -542 -1981 -540
rect -2015 -578 -1981 -576
rect -2015 -650 -1981 -644
rect -2015 -722 -1981 -712
rect -2015 -794 -1981 -780
rect -2015 -866 -1981 -848
rect -2015 -938 -1981 -916
rect -2015 -1013 -1981 -984
rect -1867 -134 -1833 -105
rect -1867 -202 -1833 -180
rect -1867 -270 -1833 -252
rect -1867 -338 -1833 -324
rect -1867 -406 -1833 -396
rect -1867 -474 -1833 -468
rect -1867 -542 -1833 -540
rect -1867 -578 -1833 -576
rect -1867 -650 -1833 -644
rect -1867 -722 -1833 -712
rect -1867 -794 -1833 -780
rect -1867 -866 -1833 -848
rect -1867 -938 -1833 -916
rect -1867 -1013 -1833 -984
rect -1719 -134 -1685 -105
rect -1719 -202 -1685 -180
rect -1719 -270 -1685 -252
rect -1719 -338 -1685 -324
rect -1719 -406 -1685 -396
rect -1719 -474 -1685 -468
rect -1719 -542 -1685 -540
rect -1719 -578 -1685 -576
rect -1719 -650 -1685 -644
rect -1719 -722 -1685 -712
rect -1719 -794 -1685 -780
rect -1719 -866 -1685 -848
rect -1719 -938 -1685 -916
rect -1719 -1013 -1685 -984
rect -1571 -134 -1537 -105
rect -1571 -202 -1537 -180
rect -1571 -270 -1537 -252
rect -1571 -338 -1537 -324
rect -1571 -406 -1537 -396
rect -1571 -474 -1537 -468
rect -1571 -542 -1537 -540
rect -1571 -578 -1537 -576
rect -1571 -650 -1537 -644
rect -1571 -722 -1537 -712
rect -1571 -794 -1537 -780
rect -1571 -866 -1537 -848
rect -1571 -938 -1537 -916
rect -1571 -1013 -1537 -984
rect -1423 -134 -1389 -105
rect -1423 -202 -1389 -180
rect -1423 -270 -1389 -252
rect -1423 -338 -1389 -324
rect -1423 -406 -1389 -396
rect -1423 -474 -1389 -468
rect -1423 -542 -1389 -540
rect -1423 -578 -1389 -576
rect -1423 -650 -1389 -644
rect -1423 -722 -1389 -712
rect -1423 -794 -1389 -780
rect -1423 -866 -1389 -848
rect -1423 -938 -1389 -916
rect -1423 -1013 -1389 -984
rect -1275 -134 -1241 -105
rect -1275 -202 -1241 -180
rect -1275 -270 -1241 -252
rect -1275 -338 -1241 -324
rect -1275 -406 -1241 -396
rect -1275 -474 -1241 -468
rect -1275 -542 -1241 -540
rect -1275 -578 -1241 -576
rect -1275 -650 -1241 -644
rect -1275 -722 -1241 -712
rect -1275 -794 -1241 -780
rect -1275 -866 -1241 -848
rect -1275 -938 -1241 -916
rect -1275 -1013 -1241 -984
rect -1127 -134 -1093 -105
rect -1127 -202 -1093 -180
rect -1127 -270 -1093 -252
rect -1127 -338 -1093 -324
rect -1127 -406 -1093 -396
rect -1127 -474 -1093 -468
rect -1127 -542 -1093 -540
rect -1127 -578 -1093 -576
rect -1127 -650 -1093 -644
rect -1127 -722 -1093 -712
rect -1127 -794 -1093 -780
rect -1127 -866 -1093 -848
rect -1127 -938 -1093 -916
rect -1127 -1013 -1093 -984
rect -979 -134 -945 -105
rect -979 -202 -945 -180
rect -979 -270 -945 -252
rect -979 -338 -945 -324
rect -979 -406 -945 -396
rect -979 -474 -945 -468
rect -979 -542 -945 -540
rect -979 -578 -945 -576
rect -979 -650 -945 -644
rect -979 -722 -945 -712
rect -979 -794 -945 -780
rect -979 -866 -945 -848
rect -979 -938 -945 -916
rect -979 -1013 -945 -984
rect -831 -134 -797 -105
rect -831 -202 -797 -180
rect -831 -270 -797 -252
rect -831 -338 -797 -324
rect -831 -406 -797 -396
rect -831 -474 -797 -468
rect -831 -542 -797 -540
rect -831 -578 -797 -576
rect -831 -650 -797 -644
rect -831 -722 -797 -712
rect -831 -794 -797 -780
rect -831 -866 -797 -848
rect -831 -938 -797 -916
rect -831 -1013 -797 -984
rect -683 -134 -649 -105
rect -683 -202 -649 -180
rect -683 -270 -649 -252
rect -683 -338 -649 -324
rect -683 -406 -649 -396
rect -683 -474 -649 -468
rect -683 -542 -649 -540
rect -683 -578 -649 -576
rect -683 -650 -649 -644
rect -683 -722 -649 -712
rect -683 -794 -649 -780
rect -683 -866 -649 -848
rect -683 -938 -649 -916
rect -683 -1013 -649 -984
rect -535 -134 -501 -105
rect -535 -202 -501 -180
rect -535 -270 -501 -252
rect -535 -338 -501 -324
rect -535 -406 -501 -396
rect -535 -474 -501 -468
rect -535 -542 -501 -540
rect -535 -578 -501 -576
rect -535 -650 -501 -644
rect -535 -722 -501 -712
rect -535 -794 -501 -780
rect -535 -866 -501 -848
rect -535 -938 -501 -916
rect -535 -1013 -501 -984
rect -387 -134 -353 -105
rect -387 -202 -353 -180
rect -387 -270 -353 -252
rect -387 -338 -353 -324
rect -387 -406 -353 -396
rect -387 -474 -353 -468
rect -387 -542 -353 -540
rect -387 -578 -353 -576
rect -387 -650 -353 -644
rect -387 -722 -353 -712
rect -387 -794 -353 -780
rect -387 -866 -353 -848
rect -387 -938 -353 -916
rect -387 -1013 -353 -984
rect -239 -134 -205 -105
rect -239 -202 -205 -180
rect -239 -270 -205 -252
rect -239 -338 -205 -324
rect -239 -406 -205 -396
rect -239 -474 -205 -468
rect -239 -542 -205 -540
rect -239 -578 -205 -576
rect -239 -650 -205 -644
rect -239 -722 -205 -712
rect -239 -794 -205 -780
rect -239 -866 -205 -848
rect -239 -938 -205 -916
rect -239 -1013 -205 -984
rect -91 -134 -57 -105
rect -91 -202 -57 -180
rect -91 -270 -57 -252
rect -91 -338 -57 -324
rect -91 -406 -57 -396
rect -91 -474 -57 -468
rect -91 -542 -57 -540
rect -91 -578 -57 -576
rect -91 -650 -57 -644
rect -91 -722 -57 -712
rect -91 -794 -57 -780
rect -91 -866 -57 -848
rect -91 -938 -57 -916
rect -91 -1013 -57 -984
rect 57 -134 91 -105
rect 57 -202 91 -180
rect 57 -270 91 -252
rect 57 -338 91 -324
rect 57 -406 91 -396
rect 57 -474 91 -468
rect 57 -542 91 -540
rect 57 -578 91 -576
rect 57 -650 91 -644
rect 57 -722 91 -712
rect 57 -794 91 -780
rect 57 -866 91 -848
rect 57 -938 91 -916
rect 57 -1013 91 -984
rect 205 -134 239 -105
rect 205 -202 239 -180
rect 205 -270 239 -252
rect 205 -338 239 -324
rect 205 -406 239 -396
rect 205 -474 239 -468
rect 205 -542 239 -540
rect 205 -578 239 -576
rect 205 -650 239 -644
rect 205 -722 239 -712
rect 205 -794 239 -780
rect 205 -866 239 -848
rect 205 -938 239 -916
rect 205 -1013 239 -984
rect 353 -134 387 -105
rect 353 -202 387 -180
rect 353 -270 387 -252
rect 353 -338 387 -324
rect 353 -406 387 -396
rect 353 -474 387 -468
rect 353 -542 387 -540
rect 353 -578 387 -576
rect 353 -650 387 -644
rect 353 -722 387 -712
rect 353 -794 387 -780
rect 353 -866 387 -848
rect 353 -938 387 -916
rect 353 -1013 387 -984
rect 501 -134 535 -105
rect 501 -202 535 -180
rect 501 -270 535 -252
rect 501 -338 535 -324
rect 501 -406 535 -396
rect 501 -474 535 -468
rect 501 -542 535 -540
rect 501 -578 535 -576
rect 501 -650 535 -644
rect 501 -722 535 -712
rect 501 -794 535 -780
rect 501 -866 535 -848
rect 501 -938 535 -916
rect 501 -1013 535 -984
rect 649 -134 683 -105
rect 649 -202 683 -180
rect 649 -270 683 -252
rect 649 -338 683 -324
rect 649 -406 683 -396
rect 649 -474 683 -468
rect 649 -542 683 -540
rect 649 -578 683 -576
rect 649 -650 683 -644
rect 649 -722 683 -712
rect 649 -794 683 -780
rect 649 -866 683 -848
rect 649 -938 683 -916
rect 649 -1013 683 -984
rect 797 -134 831 -105
rect 797 -202 831 -180
rect 797 -270 831 -252
rect 797 -338 831 -324
rect 797 -406 831 -396
rect 797 -474 831 -468
rect 797 -542 831 -540
rect 797 -578 831 -576
rect 797 -650 831 -644
rect 797 -722 831 -712
rect 797 -794 831 -780
rect 797 -866 831 -848
rect 797 -938 831 -916
rect 797 -1013 831 -984
rect 945 -134 979 -105
rect 945 -202 979 -180
rect 945 -270 979 -252
rect 945 -338 979 -324
rect 945 -406 979 -396
rect 945 -474 979 -468
rect 945 -542 979 -540
rect 945 -578 979 -576
rect 945 -650 979 -644
rect 945 -722 979 -712
rect 945 -794 979 -780
rect 945 -866 979 -848
rect 945 -938 979 -916
rect 945 -1013 979 -984
rect 1093 -134 1127 -105
rect 1093 -202 1127 -180
rect 1093 -270 1127 -252
rect 1093 -338 1127 -324
rect 1093 -406 1127 -396
rect 1093 -474 1127 -468
rect 1093 -542 1127 -540
rect 1093 -578 1127 -576
rect 1093 -650 1127 -644
rect 1093 -722 1127 -712
rect 1093 -794 1127 -780
rect 1093 -866 1127 -848
rect 1093 -938 1127 -916
rect 1093 -1013 1127 -984
rect 1241 -134 1275 -105
rect 1241 -202 1275 -180
rect 1241 -270 1275 -252
rect 1241 -338 1275 -324
rect 1241 -406 1275 -396
rect 1241 -474 1275 -468
rect 1241 -542 1275 -540
rect 1241 -578 1275 -576
rect 1241 -650 1275 -644
rect 1241 -722 1275 -712
rect 1241 -794 1275 -780
rect 1241 -866 1275 -848
rect 1241 -938 1275 -916
rect 1241 -1013 1275 -984
rect 1389 -134 1423 -105
rect 1389 -202 1423 -180
rect 1389 -270 1423 -252
rect 1389 -338 1423 -324
rect 1389 -406 1423 -396
rect 1389 -474 1423 -468
rect 1389 -542 1423 -540
rect 1389 -578 1423 -576
rect 1389 -650 1423 -644
rect 1389 -722 1423 -712
rect 1389 -794 1423 -780
rect 1389 -866 1423 -848
rect 1389 -938 1423 -916
rect 1389 -1013 1423 -984
rect 1537 -134 1571 -105
rect 1537 -202 1571 -180
rect 1537 -270 1571 -252
rect 1537 -338 1571 -324
rect 1537 -406 1571 -396
rect 1537 -474 1571 -468
rect 1537 -542 1571 -540
rect 1537 -578 1571 -576
rect 1537 -650 1571 -644
rect 1537 -722 1571 -712
rect 1537 -794 1571 -780
rect 1537 -866 1571 -848
rect 1537 -938 1571 -916
rect 1537 -1013 1571 -984
rect 1685 -134 1719 -105
rect 1685 -202 1719 -180
rect 1685 -270 1719 -252
rect 1685 -338 1719 -324
rect 1685 -406 1719 -396
rect 1685 -474 1719 -468
rect 1685 -542 1719 -540
rect 1685 -578 1719 -576
rect 1685 -650 1719 -644
rect 1685 -722 1719 -712
rect 1685 -794 1719 -780
rect 1685 -866 1719 -848
rect 1685 -938 1719 -916
rect 1685 -1013 1719 -984
rect 1833 -134 1867 -105
rect 1833 -202 1867 -180
rect 1833 -270 1867 -252
rect 1833 -338 1867 -324
rect 1833 -406 1867 -396
rect 1833 -474 1867 -468
rect 1833 -542 1867 -540
rect 1833 -578 1867 -576
rect 1833 -650 1867 -644
rect 1833 -722 1867 -712
rect 1833 -794 1867 -780
rect 1833 -866 1867 -848
rect 1833 -938 1867 -916
rect 1833 -1013 1867 -984
rect 1981 -134 2015 -105
rect 1981 -202 2015 -180
rect 1981 -270 2015 -252
rect 1981 -338 2015 -324
rect 1981 -406 2015 -396
rect 1981 -474 2015 -468
rect 1981 -542 2015 -540
rect 1981 -578 2015 -576
rect 1981 -650 2015 -644
rect 1981 -722 2015 -712
rect 1981 -794 2015 -780
rect 1981 -866 2015 -848
rect 1981 -938 2015 -916
rect 1981 -1013 2015 -984
rect 2129 -134 2163 -105
rect 2129 -202 2163 -180
rect 2129 -270 2163 -252
rect 2129 -338 2163 -324
rect 2129 -406 2163 -396
rect 2129 -474 2163 -468
rect 2129 -542 2163 -540
rect 2129 -578 2163 -576
rect 2129 -650 2163 -644
rect 2129 -722 2163 -712
rect 2129 -794 2163 -780
rect 2129 -866 2163 -848
rect 2129 -938 2163 -916
rect 2129 -1013 2163 -984
rect 2277 -134 2311 -105
rect 2277 -202 2311 -180
rect 2277 -270 2311 -252
rect 2277 -338 2311 -324
rect 2277 -406 2311 -396
rect 2277 -474 2311 -468
rect 2277 -542 2311 -540
rect 2277 -578 2311 -576
rect 2277 -650 2311 -644
rect 2277 -722 2311 -712
rect 2277 -794 2311 -780
rect 2277 -866 2311 -848
rect 2277 -938 2311 -916
rect 2277 -1013 2311 -984
rect 2425 -134 2459 -105
rect 2425 -202 2459 -180
rect 2425 -270 2459 -252
rect 2425 -338 2459 -324
rect 2425 -406 2459 -396
rect 2425 -474 2459 -468
rect 2425 -542 2459 -540
rect 2425 -578 2459 -576
rect 2425 -650 2459 -644
rect 2425 -722 2459 -712
rect 2425 -794 2459 -780
rect 2425 -866 2459 -848
rect 2425 -938 2459 -916
rect 2425 -1013 2459 -984
rect 2573 -134 2607 -105
rect 2573 -202 2607 -180
rect 2573 -270 2607 -252
rect 2573 -338 2607 -324
rect 2573 -406 2607 -396
rect 2573 -474 2607 -468
rect 2573 -542 2607 -540
rect 2573 -578 2607 -576
rect 2573 -650 2607 -644
rect 2573 -722 2607 -712
rect 2573 -794 2607 -780
rect 2573 -866 2607 -848
rect 2573 -938 2607 -916
rect 2573 -1013 2607 -984
rect 2721 -134 2755 -105
rect 2721 -202 2755 -180
rect 2721 -270 2755 -252
rect 2721 -338 2755 -324
rect 2721 -406 2755 -396
rect 2721 -474 2755 -468
rect 2721 -542 2755 -540
rect 2721 -578 2755 -576
rect 2721 -650 2755 -644
rect 2721 -722 2755 -712
rect 2721 -794 2755 -780
rect 2721 -866 2755 -848
rect 2721 -938 2755 -916
rect 2721 -1013 2755 -984
rect 2869 -134 2903 -105
rect 2869 -202 2903 -180
rect 2869 -270 2903 -252
rect 2869 -338 2903 -324
rect 2869 -406 2903 -396
rect 2869 -474 2903 -468
rect 2869 -542 2903 -540
rect 2869 -578 2903 -576
rect 2869 -650 2903 -644
rect 2869 -722 2903 -712
rect 2869 -794 2903 -780
rect 2869 -866 2903 -848
rect 2869 -938 2903 -916
rect 2869 -1013 2903 -984
rect 3017 -134 3051 -105
rect 3017 -202 3051 -180
rect 3017 -270 3051 -252
rect 3017 -338 3051 -324
rect 3017 -406 3051 -396
rect 3017 -474 3051 -468
rect 3017 -542 3051 -540
rect 3017 -578 3051 -576
rect 3017 -650 3051 -644
rect 3017 -722 3051 -712
rect 3017 -794 3051 -780
rect 3017 -866 3051 -848
rect 3017 -938 3051 -916
rect 3017 -1013 3051 -984
rect 3165 -134 3199 -105
rect 3165 -202 3199 -180
rect 3165 -270 3199 -252
rect 3165 -338 3199 -324
rect 3165 -406 3199 -396
rect 3165 -474 3199 -468
rect 3165 -542 3199 -540
rect 3165 -578 3199 -576
rect 3165 -650 3199 -644
rect 3165 -722 3199 -712
rect 3165 -794 3199 -780
rect 3165 -866 3199 -848
rect 3165 -938 3199 -916
rect 3165 -1013 3199 -984
rect 3313 -134 3347 -105
rect 3313 -202 3347 -180
rect 3313 -270 3347 -252
rect 3313 -338 3347 -324
rect 3313 -406 3347 -396
rect 3313 -474 3347 -468
rect 3313 -542 3347 -540
rect 3313 -578 3347 -576
rect 3313 -650 3347 -644
rect 3313 -722 3347 -712
rect 3313 -794 3347 -780
rect 3313 -866 3347 -848
rect 3313 -938 3347 -916
rect 3313 -1013 3347 -984
rect 3461 -134 3495 -105
rect 3461 -202 3495 -180
rect 3461 -270 3495 -252
rect 3461 -338 3495 -324
rect 3461 -406 3495 -396
rect 3461 -474 3495 -468
rect 3461 -542 3495 -540
rect 3461 -578 3495 -576
rect 3461 -650 3495 -644
rect 3461 -722 3495 -712
rect 3461 -794 3495 -780
rect 3461 -866 3495 -848
rect 3461 -938 3495 -916
rect 3461 -1013 3495 -984
rect 3609 -134 3643 -105
rect 3609 -202 3643 -180
rect 3609 -270 3643 -252
rect 3609 -338 3643 -324
rect 3609 -406 3643 -396
rect 3609 -474 3643 -468
rect 3609 -542 3643 -540
rect 3609 -578 3643 -576
rect 3609 -650 3643 -644
rect 3609 -722 3643 -712
rect 3609 -794 3643 -780
rect 3609 -866 3643 -848
rect 3609 -938 3643 -916
rect 3609 -1013 3643 -984
rect 3757 -134 3791 -105
rect 3757 -202 3791 -180
rect 3757 -270 3791 -252
rect 3757 -338 3791 -324
rect 3757 -406 3791 -396
rect 3757 -474 3791 -468
rect 3757 -542 3791 -540
rect 3757 -578 3791 -576
rect 3757 -650 3791 -644
rect 3757 -722 3791 -712
rect 3757 -794 3791 -780
rect 3757 -866 3791 -848
rect 3757 -938 3791 -916
rect 3757 -1013 3791 -984
rect 3905 -134 3939 -105
rect 3905 -202 3939 -180
rect 3905 -270 3939 -252
rect 3905 -338 3939 -324
rect 3905 -406 3939 -396
rect 3905 -474 3939 -468
rect 3905 -542 3939 -540
rect 3905 -578 3939 -576
rect 3905 -650 3939 -644
rect 3905 -722 3939 -712
rect 3905 -794 3939 -780
rect 3905 -866 3939 -848
rect 3905 -938 3939 -916
rect 3905 -1013 3939 -984
rect 4053 -134 4087 -105
rect 4053 -202 4087 -180
rect 4053 -270 4087 -252
rect 4053 -338 4087 -324
rect 4053 -406 4087 -396
rect 4053 -474 4087 -468
rect 4053 -542 4087 -540
rect 4053 -578 4087 -576
rect 4053 -650 4087 -644
rect 4053 -722 4087 -712
rect 4053 -794 4087 -780
rect 4053 -866 4087 -848
rect 4053 -938 4087 -916
rect 4053 -1013 4087 -984
rect 4201 -134 4235 -105
rect 4201 -202 4235 -180
rect 4201 -270 4235 -252
rect 4201 -338 4235 -324
rect 4201 -406 4235 -396
rect 4201 -474 4235 -468
rect 4201 -542 4235 -540
rect 4201 -578 4235 -576
rect 4201 -650 4235 -644
rect 4201 -722 4235 -712
rect 4201 -794 4235 -780
rect 4201 -866 4235 -848
rect 4201 -938 4235 -916
rect 4201 -1013 4235 -984
rect 4349 -134 4383 -105
rect 4349 -202 4383 -180
rect 4349 -270 4383 -252
rect 4349 -338 4383 -324
rect 4349 -406 4383 -396
rect 4349 -474 4383 -468
rect 4349 -542 4383 -540
rect 4349 -578 4383 -576
rect 4349 -650 4383 -644
rect 4349 -722 4383 -712
rect 4349 -794 4383 -780
rect 4349 -866 4383 -848
rect 4349 -938 4383 -916
rect 4349 -1013 4383 -984
rect 4497 -134 4531 -105
rect 4497 -202 4531 -180
rect 4497 -270 4531 -252
rect 4497 -338 4531 -324
rect 4497 -406 4531 -396
rect 4497 -474 4531 -468
rect 4497 -542 4531 -540
rect 4497 -578 4531 -576
rect 4497 -650 4531 -644
rect 4497 -722 4531 -712
rect 4497 -794 4531 -780
rect 4497 -866 4531 -848
rect 4497 -938 4531 -916
rect 4497 -1013 4531 -984
rect 4645 -134 4679 -105
rect 4645 -202 4679 -180
rect 4645 -270 4679 -252
rect 4645 -338 4679 -324
rect 4645 -406 4679 -396
rect 4645 -474 4679 -468
rect 4645 -542 4679 -540
rect 4645 -578 4679 -576
rect 4645 -650 4679 -644
rect 4645 -722 4679 -712
rect 4645 -794 4679 -780
rect 4645 -866 4679 -848
rect 4645 -938 4679 -916
rect 4645 -1013 4679 -984
rect 4793 -134 4827 -105
rect 4793 -202 4827 -180
rect 4793 -270 4827 -252
rect 4793 -338 4827 -324
rect 4793 -406 4827 -396
rect 4793 -474 4827 -468
rect 4793 -542 4827 -540
rect 4793 -578 4827 -576
rect 4793 -650 4827 -644
rect 4793 -722 4827 -712
rect 4793 -794 4827 -780
rect 4793 -866 4827 -848
rect 4793 -938 4827 -916
rect 4793 -1013 4827 -984
rect 4941 -134 4975 -105
rect 4941 -202 4975 -180
rect 4941 -270 4975 -252
rect 4941 -338 4975 -324
rect 4941 -406 4975 -396
rect 4941 -474 4975 -468
rect 4941 -542 4975 -540
rect 4941 -578 4975 -576
rect 4941 -650 4975 -644
rect 4941 -722 4975 -712
rect 4941 -794 4975 -780
rect 4941 -866 4975 -848
rect 4941 -938 4975 -916
rect 4941 -1013 4975 -984
rect 5089 -134 5123 -105
rect 5089 -202 5123 -180
rect 5089 -270 5123 -252
rect 5089 -338 5123 -324
rect 5089 -406 5123 -396
rect 5089 -474 5123 -468
rect 5089 -542 5123 -540
rect 5089 -578 5123 -576
rect 5089 -650 5123 -644
rect 5089 -722 5123 -712
rect 5089 -794 5123 -780
rect 5089 -866 5123 -848
rect 5089 -938 5123 -916
rect 5089 -1013 5123 -984
rect 5237 -134 5271 -105
rect 5237 -202 5271 -180
rect 5237 -270 5271 -252
rect 5237 -338 5271 -324
rect 5237 -406 5271 -396
rect 5237 -474 5271 -468
rect 5237 -542 5271 -540
rect 5237 -578 5271 -576
rect 5237 -650 5271 -644
rect 5237 -722 5271 -712
rect 5237 -794 5271 -780
rect 5237 -866 5271 -848
rect 5237 -938 5271 -916
rect 5237 -1013 5271 -984
rect 5385 -134 5419 -105
rect 5385 -202 5419 -180
rect 5385 -270 5419 -252
rect 5385 -338 5419 -324
rect 5385 -406 5419 -396
rect 5385 -474 5419 -468
rect 5385 -542 5419 -540
rect 5385 -578 5419 -576
rect 5385 -650 5419 -644
rect 5385 -722 5419 -712
rect 5385 -794 5419 -780
rect 5385 -866 5419 -848
rect 5385 -938 5419 -916
rect 5385 -1013 5419 -984
rect 5533 -134 5567 -105
rect 5533 -202 5567 -180
rect 5533 -270 5567 -252
rect 5533 -338 5567 -324
rect 5533 -406 5567 -396
rect 5533 -474 5567 -468
rect 5533 -542 5567 -540
rect 5533 -578 5567 -576
rect 5533 -650 5567 -644
rect 5533 -722 5567 -712
rect 5533 -794 5567 -780
rect 5533 -866 5567 -848
rect 5533 -938 5567 -916
rect 5533 -1013 5567 -984
rect 5647 -153 5681 -119
rect 5647 -221 5681 -187
rect 5647 -289 5681 -255
rect 5647 -357 5681 -323
rect 5647 -425 5681 -391
rect 5647 -493 5681 -459
rect 5647 -561 5681 -527
rect 5647 -629 5681 -595
rect 5647 -697 5681 -663
rect 5647 -765 5681 -731
rect 5647 -833 5681 -799
rect 5647 -901 5681 -867
rect 5647 -969 5681 -935
rect 5647 -1037 5681 -1003
rect -5681 -1149 -5647 -1071
rect -5521 -1081 -5493 -1047
rect -5459 -1081 -5431 -1047
rect -5373 -1081 -5345 -1047
rect -5311 -1081 -5283 -1047
rect -5225 -1081 -5197 -1047
rect -5163 -1081 -5135 -1047
rect -5077 -1081 -5049 -1047
rect -5015 -1081 -4987 -1047
rect -4929 -1081 -4901 -1047
rect -4867 -1081 -4839 -1047
rect -4781 -1081 -4753 -1047
rect -4719 -1081 -4691 -1047
rect -4633 -1081 -4605 -1047
rect -4571 -1081 -4543 -1047
rect -4485 -1081 -4457 -1047
rect -4423 -1081 -4395 -1047
rect -4337 -1081 -4309 -1047
rect -4275 -1081 -4247 -1047
rect -4189 -1081 -4161 -1047
rect -4127 -1081 -4099 -1047
rect -4041 -1081 -4013 -1047
rect -3979 -1081 -3951 -1047
rect -3893 -1081 -3865 -1047
rect -3831 -1081 -3803 -1047
rect -3745 -1081 -3717 -1047
rect -3683 -1081 -3655 -1047
rect -3597 -1081 -3569 -1047
rect -3535 -1081 -3507 -1047
rect -3449 -1081 -3421 -1047
rect -3387 -1081 -3359 -1047
rect -3301 -1081 -3273 -1047
rect -3239 -1081 -3211 -1047
rect -3153 -1081 -3125 -1047
rect -3091 -1081 -3063 -1047
rect -3005 -1081 -2977 -1047
rect -2943 -1081 -2915 -1047
rect -2857 -1081 -2829 -1047
rect -2795 -1081 -2767 -1047
rect -2709 -1081 -2681 -1047
rect -2647 -1081 -2619 -1047
rect -2561 -1081 -2533 -1047
rect -2499 -1081 -2471 -1047
rect -2413 -1081 -2385 -1047
rect -2351 -1081 -2323 -1047
rect -2265 -1081 -2237 -1047
rect -2203 -1081 -2175 -1047
rect -2117 -1081 -2089 -1047
rect -2055 -1081 -2027 -1047
rect -1969 -1081 -1941 -1047
rect -1907 -1081 -1879 -1047
rect -1821 -1081 -1793 -1047
rect -1759 -1081 -1731 -1047
rect -1673 -1081 -1645 -1047
rect -1611 -1081 -1583 -1047
rect -1525 -1081 -1497 -1047
rect -1463 -1081 -1435 -1047
rect -1377 -1081 -1349 -1047
rect -1315 -1081 -1287 -1047
rect -1229 -1081 -1201 -1047
rect -1167 -1081 -1139 -1047
rect -1081 -1081 -1053 -1047
rect -1019 -1081 -991 -1047
rect -933 -1081 -905 -1047
rect -871 -1081 -843 -1047
rect -785 -1081 -757 -1047
rect -723 -1081 -695 -1047
rect -637 -1081 -609 -1047
rect -575 -1081 -547 -1047
rect -489 -1081 -461 -1047
rect -427 -1081 -399 -1047
rect -341 -1081 -313 -1047
rect -279 -1081 -251 -1047
rect -193 -1081 -165 -1047
rect -131 -1081 -103 -1047
rect -45 -1081 -17 -1047
rect 17 -1081 45 -1047
rect 103 -1081 131 -1047
rect 165 -1081 193 -1047
rect 251 -1081 279 -1047
rect 313 -1081 341 -1047
rect 399 -1081 427 -1047
rect 461 -1081 489 -1047
rect 547 -1081 575 -1047
rect 609 -1081 637 -1047
rect 695 -1081 723 -1047
rect 757 -1081 785 -1047
rect 843 -1081 871 -1047
rect 905 -1081 933 -1047
rect 991 -1081 1019 -1047
rect 1053 -1081 1081 -1047
rect 1139 -1081 1167 -1047
rect 1201 -1081 1229 -1047
rect 1287 -1081 1315 -1047
rect 1349 -1081 1377 -1047
rect 1435 -1081 1463 -1047
rect 1497 -1081 1525 -1047
rect 1583 -1081 1611 -1047
rect 1645 -1081 1673 -1047
rect 1731 -1081 1759 -1047
rect 1793 -1081 1821 -1047
rect 1879 -1081 1907 -1047
rect 1941 -1081 1969 -1047
rect 2027 -1081 2055 -1047
rect 2089 -1081 2117 -1047
rect 2175 -1081 2203 -1047
rect 2237 -1081 2265 -1047
rect 2323 -1081 2351 -1047
rect 2385 -1081 2413 -1047
rect 2471 -1081 2499 -1047
rect 2533 -1081 2561 -1047
rect 2619 -1081 2647 -1047
rect 2681 -1081 2709 -1047
rect 2767 -1081 2795 -1047
rect 2829 -1081 2857 -1047
rect 2915 -1081 2943 -1047
rect 2977 -1081 3005 -1047
rect 3063 -1081 3091 -1047
rect 3125 -1081 3153 -1047
rect 3211 -1081 3239 -1047
rect 3273 -1081 3301 -1047
rect 3359 -1081 3387 -1047
rect 3421 -1081 3449 -1047
rect 3507 -1081 3535 -1047
rect 3569 -1081 3597 -1047
rect 3655 -1081 3683 -1047
rect 3717 -1081 3745 -1047
rect 3803 -1081 3831 -1047
rect 3865 -1081 3893 -1047
rect 3951 -1081 3979 -1047
rect 4013 -1081 4041 -1047
rect 4099 -1081 4127 -1047
rect 4161 -1081 4189 -1047
rect 4247 -1081 4275 -1047
rect 4309 -1081 4337 -1047
rect 4395 -1081 4423 -1047
rect 4457 -1081 4485 -1047
rect 4543 -1081 4571 -1047
rect 4605 -1081 4633 -1047
rect 4691 -1081 4719 -1047
rect 4753 -1081 4781 -1047
rect 4839 -1081 4867 -1047
rect 4901 -1081 4929 -1047
rect 4987 -1081 5015 -1047
rect 5049 -1081 5077 -1047
rect 5135 -1081 5163 -1047
rect 5197 -1081 5225 -1047
rect 5283 -1081 5311 -1047
rect 5345 -1081 5373 -1047
rect 5431 -1081 5459 -1047
rect 5493 -1081 5521 -1047
rect 5647 -1149 5681 -1071
rect -5681 -1183 -5559 -1149
rect -5525 -1183 -5491 -1149
rect -5457 -1183 -5423 -1149
rect -5389 -1183 -5355 -1149
rect -5321 -1183 -5287 -1149
rect -5253 -1183 -5219 -1149
rect -5185 -1183 -5151 -1149
rect -5117 -1183 -5083 -1149
rect -5049 -1183 -5015 -1149
rect -4981 -1183 -4947 -1149
rect -4913 -1183 -4879 -1149
rect -4845 -1183 -4811 -1149
rect -4777 -1183 -4743 -1149
rect -4709 -1183 -4675 -1149
rect -4641 -1183 -4607 -1149
rect -4573 -1183 -4539 -1149
rect -4505 -1183 -4471 -1149
rect -4437 -1183 -4403 -1149
rect -4369 -1183 -4335 -1149
rect -4301 -1183 -4267 -1149
rect -4233 -1183 -4199 -1149
rect -4165 -1183 -4131 -1149
rect -4097 -1183 -4063 -1149
rect -4029 -1183 -3995 -1149
rect -3961 -1183 -3927 -1149
rect -3893 -1183 -3859 -1149
rect -3825 -1183 -3791 -1149
rect -3757 -1183 -3723 -1149
rect -3689 -1183 -3655 -1149
rect -3621 -1183 -3587 -1149
rect -3553 -1183 -3519 -1149
rect -3485 -1183 -3451 -1149
rect -3417 -1183 -3383 -1149
rect -3349 -1183 -3315 -1149
rect -3281 -1183 -3247 -1149
rect -3213 -1183 -3179 -1149
rect -3145 -1183 -3111 -1149
rect -3077 -1183 -3043 -1149
rect -3009 -1183 -2975 -1149
rect -2941 -1183 -2907 -1149
rect -2873 -1183 -2839 -1149
rect -2805 -1183 -2771 -1149
rect -2737 -1183 -2703 -1149
rect -2669 -1183 -2635 -1149
rect -2601 -1183 -2567 -1149
rect -2533 -1183 -2499 -1149
rect -2465 -1183 -2431 -1149
rect -2397 -1183 -2363 -1149
rect -2329 -1183 -2295 -1149
rect -2261 -1183 -2227 -1149
rect -2193 -1183 -2159 -1149
rect -2125 -1183 -2091 -1149
rect -2057 -1183 -2023 -1149
rect -1989 -1183 -1955 -1149
rect -1921 -1183 -1887 -1149
rect -1853 -1183 -1819 -1149
rect -1785 -1183 -1751 -1149
rect -1717 -1183 -1683 -1149
rect -1649 -1183 -1615 -1149
rect -1581 -1183 -1547 -1149
rect -1513 -1183 -1479 -1149
rect -1445 -1183 -1411 -1149
rect -1377 -1183 -1343 -1149
rect -1309 -1183 -1275 -1149
rect -1241 -1183 -1207 -1149
rect -1173 -1183 -1139 -1149
rect -1105 -1183 -1071 -1149
rect -1037 -1183 -1003 -1149
rect -969 -1183 -935 -1149
rect -901 -1183 -867 -1149
rect -833 -1183 -799 -1149
rect -765 -1183 -731 -1149
rect -697 -1183 -663 -1149
rect -629 -1183 -595 -1149
rect -561 -1183 -527 -1149
rect -493 -1183 -459 -1149
rect -425 -1183 -391 -1149
rect -357 -1183 -323 -1149
rect -289 -1183 -255 -1149
rect -221 -1183 -187 -1149
rect -153 -1183 -119 -1149
rect -85 -1183 -51 -1149
rect -17 -1183 17 -1149
rect 51 -1183 85 -1149
rect 119 -1183 153 -1149
rect 187 -1183 221 -1149
rect 255 -1183 289 -1149
rect 323 -1183 357 -1149
rect 391 -1183 425 -1149
rect 459 -1183 493 -1149
rect 527 -1183 561 -1149
rect 595 -1183 629 -1149
rect 663 -1183 697 -1149
rect 731 -1183 765 -1149
rect 799 -1183 833 -1149
rect 867 -1183 901 -1149
rect 935 -1183 969 -1149
rect 1003 -1183 1037 -1149
rect 1071 -1183 1105 -1149
rect 1139 -1183 1173 -1149
rect 1207 -1183 1241 -1149
rect 1275 -1183 1309 -1149
rect 1343 -1183 1377 -1149
rect 1411 -1183 1445 -1149
rect 1479 -1183 1513 -1149
rect 1547 -1183 1581 -1149
rect 1615 -1183 1649 -1149
rect 1683 -1183 1717 -1149
rect 1751 -1183 1785 -1149
rect 1819 -1183 1853 -1149
rect 1887 -1183 1921 -1149
rect 1955 -1183 1989 -1149
rect 2023 -1183 2057 -1149
rect 2091 -1183 2125 -1149
rect 2159 -1183 2193 -1149
rect 2227 -1183 2261 -1149
rect 2295 -1183 2329 -1149
rect 2363 -1183 2397 -1149
rect 2431 -1183 2465 -1149
rect 2499 -1183 2533 -1149
rect 2567 -1183 2601 -1149
rect 2635 -1183 2669 -1149
rect 2703 -1183 2737 -1149
rect 2771 -1183 2805 -1149
rect 2839 -1183 2873 -1149
rect 2907 -1183 2941 -1149
rect 2975 -1183 3009 -1149
rect 3043 -1183 3077 -1149
rect 3111 -1183 3145 -1149
rect 3179 -1183 3213 -1149
rect 3247 -1183 3281 -1149
rect 3315 -1183 3349 -1149
rect 3383 -1183 3417 -1149
rect 3451 -1183 3485 -1149
rect 3519 -1183 3553 -1149
rect 3587 -1183 3621 -1149
rect 3655 -1183 3689 -1149
rect 3723 -1183 3757 -1149
rect 3791 -1183 3825 -1149
rect 3859 -1183 3893 -1149
rect 3927 -1183 3961 -1149
rect 3995 -1183 4029 -1149
rect 4063 -1183 4097 -1149
rect 4131 -1183 4165 -1149
rect 4199 -1183 4233 -1149
rect 4267 -1183 4301 -1149
rect 4335 -1183 4369 -1149
rect 4403 -1183 4437 -1149
rect 4471 -1183 4505 -1149
rect 4539 -1183 4573 -1149
rect 4607 -1183 4641 -1149
rect 4675 -1183 4709 -1149
rect 4743 -1183 4777 -1149
rect 4811 -1183 4845 -1149
rect 4879 -1183 4913 -1149
rect 4947 -1183 4981 -1149
rect 5015 -1183 5049 -1149
rect 5083 -1183 5117 -1149
rect 5151 -1183 5185 -1149
rect 5219 -1183 5253 -1149
rect 5287 -1183 5321 -1149
rect 5355 -1183 5389 -1149
rect 5423 -1183 5457 -1149
rect 5491 -1183 5525 -1149
rect 5559 -1183 5681 -1149
<< viali >>
rect -5493 1047 -5459 1081
rect -5345 1047 -5311 1081
rect -5197 1047 -5163 1081
rect -5049 1047 -5015 1081
rect -4901 1047 -4867 1081
rect -4753 1047 -4719 1081
rect -4605 1047 -4571 1081
rect -4457 1047 -4423 1081
rect -4309 1047 -4275 1081
rect -4161 1047 -4127 1081
rect -4013 1047 -3979 1081
rect -3865 1047 -3831 1081
rect -3717 1047 -3683 1081
rect -3569 1047 -3535 1081
rect -3421 1047 -3387 1081
rect -3273 1047 -3239 1081
rect -3125 1047 -3091 1081
rect -2977 1047 -2943 1081
rect -2829 1047 -2795 1081
rect -2681 1047 -2647 1081
rect -2533 1047 -2499 1081
rect -2385 1047 -2351 1081
rect -2237 1047 -2203 1081
rect -2089 1047 -2055 1081
rect -1941 1047 -1907 1081
rect -1793 1047 -1759 1081
rect -1645 1047 -1611 1081
rect -1497 1047 -1463 1081
rect -1349 1047 -1315 1081
rect -1201 1047 -1167 1081
rect -1053 1047 -1019 1081
rect -905 1047 -871 1081
rect -757 1047 -723 1081
rect -609 1047 -575 1081
rect -461 1047 -427 1081
rect -313 1047 -279 1081
rect -165 1047 -131 1081
rect -17 1047 17 1081
rect 131 1047 165 1081
rect 279 1047 313 1081
rect 427 1047 461 1081
rect 575 1047 609 1081
rect 723 1047 757 1081
rect 871 1047 905 1081
rect 1019 1047 1053 1081
rect 1167 1047 1201 1081
rect 1315 1047 1349 1081
rect 1463 1047 1497 1081
rect 1611 1047 1645 1081
rect 1759 1047 1793 1081
rect 1907 1047 1941 1081
rect 2055 1047 2089 1081
rect 2203 1047 2237 1081
rect 2351 1047 2385 1081
rect 2499 1047 2533 1081
rect 2647 1047 2681 1081
rect 2795 1047 2829 1081
rect 2943 1047 2977 1081
rect 3091 1047 3125 1081
rect 3239 1047 3273 1081
rect 3387 1047 3421 1081
rect 3535 1047 3569 1081
rect 3683 1047 3717 1081
rect 3831 1047 3865 1081
rect 3979 1047 4013 1081
rect 4127 1047 4161 1081
rect 4275 1047 4309 1081
rect 4423 1047 4457 1081
rect 4571 1047 4605 1081
rect 4719 1047 4753 1081
rect 4867 1047 4901 1081
rect 5015 1047 5049 1081
rect 5163 1047 5197 1081
rect 5311 1047 5345 1081
rect 5459 1047 5493 1081
rect -5567 950 -5533 972
rect -5567 938 -5533 950
rect -5567 882 -5533 900
rect -5567 866 -5533 882
rect -5567 814 -5533 828
rect -5567 794 -5533 814
rect -5567 746 -5533 756
rect -5567 722 -5533 746
rect -5567 678 -5533 684
rect -5567 650 -5533 678
rect -5567 610 -5533 612
rect -5567 578 -5533 610
rect -5567 508 -5533 540
rect -5567 506 -5533 508
rect -5567 440 -5533 468
rect -5567 434 -5533 440
rect -5567 372 -5533 396
rect -5567 362 -5533 372
rect -5567 304 -5533 324
rect -5567 290 -5533 304
rect -5567 236 -5533 252
rect -5567 218 -5533 236
rect -5567 168 -5533 180
rect -5567 146 -5533 168
rect -5419 950 -5385 972
rect -5419 938 -5385 950
rect -5419 882 -5385 900
rect -5419 866 -5385 882
rect -5419 814 -5385 828
rect -5419 794 -5385 814
rect -5419 746 -5385 756
rect -5419 722 -5385 746
rect -5419 678 -5385 684
rect -5419 650 -5385 678
rect -5419 610 -5385 612
rect -5419 578 -5385 610
rect -5419 508 -5385 540
rect -5419 506 -5385 508
rect -5419 440 -5385 468
rect -5419 434 -5385 440
rect -5419 372 -5385 396
rect -5419 362 -5385 372
rect -5419 304 -5385 324
rect -5419 290 -5385 304
rect -5419 236 -5385 252
rect -5419 218 -5385 236
rect -5419 168 -5385 180
rect -5419 146 -5385 168
rect -5271 950 -5237 972
rect -5271 938 -5237 950
rect -5271 882 -5237 900
rect -5271 866 -5237 882
rect -5271 814 -5237 828
rect -5271 794 -5237 814
rect -5271 746 -5237 756
rect -5271 722 -5237 746
rect -5271 678 -5237 684
rect -5271 650 -5237 678
rect -5271 610 -5237 612
rect -5271 578 -5237 610
rect -5271 508 -5237 540
rect -5271 506 -5237 508
rect -5271 440 -5237 468
rect -5271 434 -5237 440
rect -5271 372 -5237 396
rect -5271 362 -5237 372
rect -5271 304 -5237 324
rect -5271 290 -5237 304
rect -5271 236 -5237 252
rect -5271 218 -5237 236
rect -5271 168 -5237 180
rect -5271 146 -5237 168
rect -5123 950 -5089 972
rect -5123 938 -5089 950
rect -5123 882 -5089 900
rect -5123 866 -5089 882
rect -5123 814 -5089 828
rect -5123 794 -5089 814
rect -5123 746 -5089 756
rect -5123 722 -5089 746
rect -5123 678 -5089 684
rect -5123 650 -5089 678
rect -5123 610 -5089 612
rect -5123 578 -5089 610
rect -5123 508 -5089 540
rect -5123 506 -5089 508
rect -5123 440 -5089 468
rect -5123 434 -5089 440
rect -5123 372 -5089 396
rect -5123 362 -5089 372
rect -5123 304 -5089 324
rect -5123 290 -5089 304
rect -5123 236 -5089 252
rect -5123 218 -5089 236
rect -5123 168 -5089 180
rect -5123 146 -5089 168
rect -4975 950 -4941 972
rect -4975 938 -4941 950
rect -4975 882 -4941 900
rect -4975 866 -4941 882
rect -4975 814 -4941 828
rect -4975 794 -4941 814
rect -4975 746 -4941 756
rect -4975 722 -4941 746
rect -4975 678 -4941 684
rect -4975 650 -4941 678
rect -4975 610 -4941 612
rect -4975 578 -4941 610
rect -4975 508 -4941 540
rect -4975 506 -4941 508
rect -4975 440 -4941 468
rect -4975 434 -4941 440
rect -4975 372 -4941 396
rect -4975 362 -4941 372
rect -4975 304 -4941 324
rect -4975 290 -4941 304
rect -4975 236 -4941 252
rect -4975 218 -4941 236
rect -4975 168 -4941 180
rect -4975 146 -4941 168
rect -4827 950 -4793 972
rect -4827 938 -4793 950
rect -4827 882 -4793 900
rect -4827 866 -4793 882
rect -4827 814 -4793 828
rect -4827 794 -4793 814
rect -4827 746 -4793 756
rect -4827 722 -4793 746
rect -4827 678 -4793 684
rect -4827 650 -4793 678
rect -4827 610 -4793 612
rect -4827 578 -4793 610
rect -4827 508 -4793 540
rect -4827 506 -4793 508
rect -4827 440 -4793 468
rect -4827 434 -4793 440
rect -4827 372 -4793 396
rect -4827 362 -4793 372
rect -4827 304 -4793 324
rect -4827 290 -4793 304
rect -4827 236 -4793 252
rect -4827 218 -4793 236
rect -4827 168 -4793 180
rect -4827 146 -4793 168
rect -4679 950 -4645 972
rect -4679 938 -4645 950
rect -4679 882 -4645 900
rect -4679 866 -4645 882
rect -4679 814 -4645 828
rect -4679 794 -4645 814
rect -4679 746 -4645 756
rect -4679 722 -4645 746
rect -4679 678 -4645 684
rect -4679 650 -4645 678
rect -4679 610 -4645 612
rect -4679 578 -4645 610
rect -4679 508 -4645 540
rect -4679 506 -4645 508
rect -4679 440 -4645 468
rect -4679 434 -4645 440
rect -4679 372 -4645 396
rect -4679 362 -4645 372
rect -4679 304 -4645 324
rect -4679 290 -4645 304
rect -4679 236 -4645 252
rect -4679 218 -4645 236
rect -4679 168 -4645 180
rect -4679 146 -4645 168
rect -4531 950 -4497 972
rect -4531 938 -4497 950
rect -4531 882 -4497 900
rect -4531 866 -4497 882
rect -4531 814 -4497 828
rect -4531 794 -4497 814
rect -4531 746 -4497 756
rect -4531 722 -4497 746
rect -4531 678 -4497 684
rect -4531 650 -4497 678
rect -4531 610 -4497 612
rect -4531 578 -4497 610
rect -4531 508 -4497 540
rect -4531 506 -4497 508
rect -4531 440 -4497 468
rect -4531 434 -4497 440
rect -4531 372 -4497 396
rect -4531 362 -4497 372
rect -4531 304 -4497 324
rect -4531 290 -4497 304
rect -4531 236 -4497 252
rect -4531 218 -4497 236
rect -4531 168 -4497 180
rect -4531 146 -4497 168
rect -4383 950 -4349 972
rect -4383 938 -4349 950
rect -4383 882 -4349 900
rect -4383 866 -4349 882
rect -4383 814 -4349 828
rect -4383 794 -4349 814
rect -4383 746 -4349 756
rect -4383 722 -4349 746
rect -4383 678 -4349 684
rect -4383 650 -4349 678
rect -4383 610 -4349 612
rect -4383 578 -4349 610
rect -4383 508 -4349 540
rect -4383 506 -4349 508
rect -4383 440 -4349 468
rect -4383 434 -4349 440
rect -4383 372 -4349 396
rect -4383 362 -4349 372
rect -4383 304 -4349 324
rect -4383 290 -4349 304
rect -4383 236 -4349 252
rect -4383 218 -4349 236
rect -4383 168 -4349 180
rect -4383 146 -4349 168
rect -4235 950 -4201 972
rect -4235 938 -4201 950
rect -4235 882 -4201 900
rect -4235 866 -4201 882
rect -4235 814 -4201 828
rect -4235 794 -4201 814
rect -4235 746 -4201 756
rect -4235 722 -4201 746
rect -4235 678 -4201 684
rect -4235 650 -4201 678
rect -4235 610 -4201 612
rect -4235 578 -4201 610
rect -4235 508 -4201 540
rect -4235 506 -4201 508
rect -4235 440 -4201 468
rect -4235 434 -4201 440
rect -4235 372 -4201 396
rect -4235 362 -4201 372
rect -4235 304 -4201 324
rect -4235 290 -4201 304
rect -4235 236 -4201 252
rect -4235 218 -4201 236
rect -4235 168 -4201 180
rect -4235 146 -4201 168
rect -4087 950 -4053 972
rect -4087 938 -4053 950
rect -4087 882 -4053 900
rect -4087 866 -4053 882
rect -4087 814 -4053 828
rect -4087 794 -4053 814
rect -4087 746 -4053 756
rect -4087 722 -4053 746
rect -4087 678 -4053 684
rect -4087 650 -4053 678
rect -4087 610 -4053 612
rect -4087 578 -4053 610
rect -4087 508 -4053 540
rect -4087 506 -4053 508
rect -4087 440 -4053 468
rect -4087 434 -4053 440
rect -4087 372 -4053 396
rect -4087 362 -4053 372
rect -4087 304 -4053 324
rect -4087 290 -4053 304
rect -4087 236 -4053 252
rect -4087 218 -4053 236
rect -4087 168 -4053 180
rect -4087 146 -4053 168
rect -3939 950 -3905 972
rect -3939 938 -3905 950
rect -3939 882 -3905 900
rect -3939 866 -3905 882
rect -3939 814 -3905 828
rect -3939 794 -3905 814
rect -3939 746 -3905 756
rect -3939 722 -3905 746
rect -3939 678 -3905 684
rect -3939 650 -3905 678
rect -3939 610 -3905 612
rect -3939 578 -3905 610
rect -3939 508 -3905 540
rect -3939 506 -3905 508
rect -3939 440 -3905 468
rect -3939 434 -3905 440
rect -3939 372 -3905 396
rect -3939 362 -3905 372
rect -3939 304 -3905 324
rect -3939 290 -3905 304
rect -3939 236 -3905 252
rect -3939 218 -3905 236
rect -3939 168 -3905 180
rect -3939 146 -3905 168
rect -3791 950 -3757 972
rect -3791 938 -3757 950
rect -3791 882 -3757 900
rect -3791 866 -3757 882
rect -3791 814 -3757 828
rect -3791 794 -3757 814
rect -3791 746 -3757 756
rect -3791 722 -3757 746
rect -3791 678 -3757 684
rect -3791 650 -3757 678
rect -3791 610 -3757 612
rect -3791 578 -3757 610
rect -3791 508 -3757 540
rect -3791 506 -3757 508
rect -3791 440 -3757 468
rect -3791 434 -3757 440
rect -3791 372 -3757 396
rect -3791 362 -3757 372
rect -3791 304 -3757 324
rect -3791 290 -3757 304
rect -3791 236 -3757 252
rect -3791 218 -3757 236
rect -3791 168 -3757 180
rect -3791 146 -3757 168
rect -3643 950 -3609 972
rect -3643 938 -3609 950
rect -3643 882 -3609 900
rect -3643 866 -3609 882
rect -3643 814 -3609 828
rect -3643 794 -3609 814
rect -3643 746 -3609 756
rect -3643 722 -3609 746
rect -3643 678 -3609 684
rect -3643 650 -3609 678
rect -3643 610 -3609 612
rect -3643 578 -3609 610
rect -3643 508 -3609 540
rect -3643 506 -3609 508
rect -3643 440 -3609 468
rect -3643 434 -3609 440
rect -3643 372 -3609 396
rect -3643 362 -3609 372
rect -3643 304 -3609 324
rect -3643 290 -3609 304
rect -3643 236 -3609 252
rect -3643 218 -3609 236
rect -3643 168 -3609 180
rect -3643 146 -3609 168
rect -3495 950 -3461 972
rect -3495 938 -3461 950
rect -3495 882 -3461 900
rect -3495 866 -3461 882
rect -3495 814 -3461 828
rect -3495 794 -3461 814
rect -3495 746 -3461 756
rect -3495 722 -3461 746
rect -3495 678 -3461 684
rect -3495 650 -3461 678
rect -3495 610 -3461 612
rect -3495 578 -3461 610
rect -3495 508 -3461 540
rect -3495 506 -3461 508
rect -3495 440 -3461 468
rect -3495 434 -3461 440
rect -3495 372 -3461 396
rect -3495 362 -3461 372
rect -3495 304 -3461 324
rect -3495 290 -3461 304
rect -3495 236 -3461 252
rect -3495 218 -3461 236
rect -3495 168 -3461 180
rect -3495 146 -3461 168
rect -3347 950 -3313 972
rect -3347 938 -3313 950
rect -3347 882 -3313 900
rect -3347 866 -3313 882
rect -3347 814 -3313 828
rect -3347 794 -3313 814
rect -3347 746 -3313 756
rect -3347 722 -3313 746
rect -3347 678 -3313 684
rect -3347 650 -3313 678
rect -3347 610 -3313 612
rect -3347 578 -3313 610
rect -3347 508 -3313 540
rect -3347 506 -3313 508
rect -3347 440 -3313 468
rect -3347 434 -3313 440
rect -3347 372 -3313 396
rect -3347 362 -3313 372
rect -3347 304 -3313 324
rect -3347 290 -3313 304
rect -3347 236 -3313 252
rect -3347 218 -3313 236
rect -3347 168 -3313 180
rect -3347 146 -3313 168
rect -3199 950 -3165 972
rect -3199 938 -3165 950
rect -3199 882 -3165 900
rect -3199 866 -3165 882
rect -3199 814 -3165 828
rect -3199 794 -3165 814
rect -3199 746 -3165 756
rect -3199 722 -3165 746
rect -3199 678 -3165 684
rect -3199 650 -3165 678
rect -3199 610 -3165 612
rect -3199 578 -3165 610
rect -3199 508 -3165 540
rect -3199 506 -3165 508
rect -3199 440 -3165 468
rect -3199 434 -3165 440
rect -3199 372 -3165 396
rect -3199 362 -3165 372
rect -3199 304 -3165 324
rect -3199 290 -3165 304
rect -3199 236 -3165 252
rect -3199 218 -3165 236
rect -3199 168 -3165 180
rect -3199 146 -3165 168
rect -3051 950 -3017 972
rect -3051 938 -3017 950
rect -3051 882 -3017 900
rect -3051 866 -3017 882
rect -3051 814 -3017 828
rect -3051 794 -3017 814
rect -3051 746 -3017 756
rect -3051 722 -3017 746
rect -3051 678 -3017 684
rect -3051 650 -3017 678
rect -3051 610 -3017 612
rect -3051 578 -3017 610
rect -3051 508 -3017 540
rect -3051 506 -3017 508
rect -3051 440 -3017 468
rect -3051 434 -3017 440
rect -3051 372 -3017 396
rect -3051 362 -3017 372
rect -3051 304 -3017 324
rect -3051 290 -3017 304
rect -3051 236 -3017 252
rect -3051 218 -3017 236
rect -3051 168 -3017 180
rect -3051 146 -3017 168
rect -2903 950 -2869 972
rect -2903 938 -2869 950
rect -2903 882 -2869 900
rect -2903 866 -2869 882
rect -2903 814 -2869 828
rect -2903 794 -2869 814
rect -2903 746 -2869 756
rect -2903 722 -2869 746
rect -2903 678 -2869 684
rect -2903 650 -2869 678
rect -2903 610 -2869 612
rect -2903 578 -2869 610
rect -2903 508 -2869 540
rect -2903 506 -2869 508
rect -2903 440 -2869 468
rect -2903 434 -2869 440
rect -2903 372 -2869 396
rect -2903 362 -2869 372
rect -2903 304 -2869 324
rect -2903 290 -2869 304
rect -2903 236 -2869 252
rect -2903 218 -2869 236
rect -2903 168 -2869 180
rect -2903 146 -2869 168
rect -2755 950 -2721 972
rect -2755 938 -2721 950
rect -2755 882 -2721 900
rect -2755 866 -2721 882
rect -2755 814 -2721 828
rect -2755 794 -2721 814
rect -2755 746 -2721 756
rect -2755 722 -2721 746
rect -2755 678 -2721 684
rect -2755 650 -2721 678
rect -2755 610 -2721 612
rect -2755 578 -2721 610
rect -2755 508 -2721 540
rect -2755 506 -2721 508
rect -2755 440 -2721 468
rect -2755 434 -2721 440
rect -2755 372 -2721 396
rect -2755 362 -2721 372
rect -2755 304 -2721 324
rect -2755 290 -2721 304
rect -2755 236 -2721 252
rect -2755 218 -2721 236
rect -2755 168 -2721 180
rect -2755 146 -2721 168
rect -2607 950 -2573 972
rect -2607 938 -2573 950
rect -2607 882 -2573 900
rect -2607 866 -2573 882
rect -2607 814 -2573 828
rect -2607 794 -2573 814
rect -2607 746 -2573 756
rect -2607 722 -2573 746
rect -2607 678 -2573 684
rect -2607 650 -2573 678
rect -2607 610 -2573 612
rect -2607 578 -2573 610
rect -2607 508 -2573 540
rect -2607 506 -2573 508
rect -2607 440 -2573 468
rect -2607 434 -2573 440
rect -2607 372 -2573 396
rect -2607 362 -2573 372
rect -2607 304 -2573 324
rect -2607 290 -2573 304
rect -2607 236 -2573 252
rect -2607 218 -2573 236
rect -2607 168 -2573 180
rect -2607 146 -2573 168
rect -2459 950 -2425 972
rect -2459 938 -2425 950
rect -2459 882 -2425 900
rect -2459 866 -2425 882
rect -2459 814 -2425 828
rect -2459 794 -2425 814
rect -2459 746 -2425 756
rect -2459 722 -2425 746
rect -2459 678 -2425 684
rect -2459 650 -2425 678
rect -2459 610 -2425 612
rect -2459 578 -2425 610
rect -2459 508 -2425 540
rect -2459 506 -2425 508
rect -2459 440 -2425 468
rect -2459 434 -2425 440
rect -2459 372 -2425 396
rect -2459 362 -2425 372
rect -2459 304 -2425 324
rect -2459 290 -2425 304
rect -2459 236 -2425 252
rect -2459 218 -2425 236
rect -2459 168 -2425 180
rect -2459 146 -2425 168
rect -2311 950 -2277 972
rect -2311 938 -2277 950
rect -2311 882 -2277 900
rect -2311 866 -2277 882
rect -2311 814 -2277 828
rect -2311 794 -2277 814
rect -2311 746 -2277 756
rect -2311 722 -2277 746
rect -2311 678 -2277 684
rect -2311 650 -2277 678
rect -2311 610 -2277 612
rect -2311 578 -2277 610
rect -2311 508 -2277 540
rect -2311 506 -2277 508
rect -2311 440 -2277 468
rect -2311 434 -2277 440
rect -2311 372 -2277 396
rect -2311 362 -2277 372
rect -2311 304 -2277 324
rect -2311 290 -2277 304
rect -2311 236 -2277 252
rect -2311 218 -2277 236
rect -2311 168 -2277 180
rect -2311 146 -2277 168
rect -2163 950 -2129 972
rect -2163 938 -2129 950
rect -2163 882 -2129 900
rect -2163 866 -2129 882
rect -2163 814 -2129 828
rect -2163 794 -2129 814
rect -2163 746 -2129 756
rect -2163 722 -2129 746
rect -2163 678 -2129 684
rect -2163 650 -2129 678
rect -2163 610 -2129 612
rect -2163 578 -2129 610
rect -2163 508 -2129 540
rect -2163 506 -2129 508
rect -2163 440 -2129 468
rect -2163 434 -2129 440
rect -2163 372 -2129 396
rect -2163 362 -2129 372
rect -2163 304 -2129 324
rect -2163 290 -2129 304
rect -2163 236 -2129 252
rect -2163 218 -2129 236
rect -2163 168 -2129 180
rect -2163 146 -2129 168
rect -2015 950 -1981 972
rect -2015 938 -1981 950
rect -2015 882 -1981 900
rect -2015 866 -1981 882
rect -2015 814 -1981 828
rect -2015 794 -1981 814
rect -2015 746 -1981 756
rect -2015 722 -1981 746
rect -2015 678 -1981 684
rect -2015 650 -1981 678
rect -2015 610 -1981 612
rect -2015 578 -1981 610
rect -2015 508 -1981 540
rect -2015 506 -1981 508
rect -2015 440 -1981 468
rect -2015 434 -1981 440
rect -2015 372 -1981 396
rect -2015 362 -1981 372
rect -2015 304 -1981 324
rect -2015 290 -1981 304
rect -2015 236 -1981 252
rect -2015 218 -1981 236
rect -2015 168 -1981 180
rect -2015 146 -1981 168
rect -1867 950 -1833 972
rect -1867 938 -1833 950
rect -1867 882 -1833 900
rect -1867 866 -1833 882
rect -1867 814 -1833 828
rect -1867 794 -1833 814
rect -1867 746 -1833 756
rect -1867 722 -1833 746
rect -1867 678 -1833 684
rect -1867 650 -1833 678
rect -1867 610 -1833 612
rect -1867 578 -1833 610
rect -1867 508 -1833 540
rect -1867 506 -1833 508
rect -1867 440 -1833 468
rect -1867 434 -1833 440
rect -1867 372 -1833 396
rect -1867 362 -1833 372
rect -1867 304 -1833 324
rect -1867 290 -1833 304
rect -1867 236 -1833 252
rect -1867 218 -1833 236
rect -1867 168 -1833 180
rect -1867 146 -1833 168
rect -1719 950 -1685 972
rect -1719 938 -1685 950
rect -1719 882 -1685 900
rect -1719 866 -1685 882
rect -1719 814 -1685 828
rect -1719 794 -1685 814
rect -1719 746 -1685 756
rect -1719 722 -1685 746
rect -1719 678 -1685 684
rect -1719 650 -1685 678
rect -1719 610 -1685 612
rect -1719 578 -1685 610
rect -1719 508 -1685 540
rect -1719 506 -1685 508
rect -1719 440 -1685 468
rect -1719 434 -1685 440
rect -1719 372 -1685 396
rect -1719 362 -1685 372
rect -1719 304 -1685 324
rect -1719 290 -1685 304
rect -1719 236 -1685 252
rect -1719 218 -1685 236
rect -1719 168 -1685 180
rect -1719 146 -1685 168
rect -1571 950 -1537 972
rect -1571 938 -1537 950
rect -1571 882 -1537 900
rect -1571 866 -1537 882
rect -1571 814 -1537 828
rect -1571 794 -1537 814
rect -1571 746 -1537 756
rect -1571 722 -1537 746
rect -1571 678 -1537 684
rect -1571 650 -1537 678
rect -1571 610 -1537 612
rect -1571 578 -1537 610
rect -1571 508 -1537 540
rect -1571 506 -1537 508
rect -1571 440 -1537 468
rect -1571 434 -1537 440
rect -1571 372 -1537 396
rect -1571 362 -1537 372
rect -1571 304 -1537 324
rect -1571 290 -1537 304
rect -1571 236 -1537 252
rect -1571 218 -1537 236
rect -1571 168 -1537 180
rect -1571 146 -1537 168
rect -1423 950 -1389 972
rect -1423 938 -1389 950
rect -1423 882 -1389 900
rect -1423 866 -1389 882
rect -1423 814 -1389 828
rect -1423 794 -1389 814
rect -1423 746 -1389 756
rect -1423 722 -1389 746
rect -1423 678 -1389 684
rect -1423 650 -1389 678
rect -1423 610 -1389 612
rect -1423 578 -1389 610
rect -1423 508 -1389 540
rect -1423 506 -1389 508
rect -1423 440 -1389 468
rect -1423 434 -1389 440
rect -1423 372 -1389 396
rect -1423 362 -1389 372
rect -1423 304 -1389 324
rect -1423 290 -1389 304
rect -1423 236 -1389 252
rect -1423 218 -1389 236
rect -1423 168 -1389 180
rect -1423 146 -1389 168
rect -1275 950 -1241 972
rect -1275 938 -1241 950
rect -1275 882 -1241 900
rect -1275 866 -1241 882
rect -1275 814 -1241 828
rect -1275 794 -1241 814
rect -1275 746 -1241 756
rect -1275 722 -1241 746
rect -1275 678 -1241 684
rect -1275 650 -1241 678
rect -1275 610 -1241 612
rect -1275 578 -1241 610
rect -1275 508 -1241 540
rect -1275 506 -1241 508
rect -1275 440 -1241 468
rect -1275 434 -1241 440
rect -1275 372 -1241 396
rect -1275 362 -1241 372
rect -1275 304 -1241 324
rect -1275 290 -1241 304
rect -1275 236 -1241 252
rect -1275 218 -1241 236
rect -1275 168 -1241 180
rect -1275 146 -1241 168
rect -1127 950 -1093 972
rect -1127 938 -1093 950
rect -1127 882 -1093 900
rect -1127 866 -1093 882
rect -1127 814 -1093 828
rect -1127 794 -1093 814
rect -1127 746 -1093 756
rect -1127 722 -1093 746
rect -1127 678 -1093 684
rect -1127 650 -1093 678
rect -1127 610 -1093 612
rect -1127 578 -1093 610
rect -1127 508 -1093 540
rect -1127 506 -1093 508
rect -1127 440 -1093 468
rect -1127 434 -1093 440
rect -1127 372 -1093 396
rect -1127 362 -1093 372
rect -1127 304 -1093 324
rect -1127 290 -1093 304
rect -1127 236 -1093 252
rect -1127 218 -1093 236
rect -1127 168 -1093 180
rect -1127 146 -1093 168
rect -979 950 -945 972
rect -979 938 -945 950
rect -979 882 -945 900
rect -979 866 -945 882
rect -979 814 -945 828
rect -979 794 -945 814
rect -979 746 -945 756
rect -979 722 -945 746
rect -979 678 -945 684
rect -979 650 -945 678
rect -979 610 -945 612
rect -979 578 -945 610
rect -979 508 -945 540
rect -979 506 -945 508
rect -979 440 -945 468
rect -979 434 -945 440
rect -979 372 -945 396
rect -979 362 -945 372
rect -979 304 -945 324
rect -979 290 -945 304
rect -979 236 -945 252
rect -979 218 -945 236
rect -979 168 -945 180
rect -979 146 -945 168
rect -831 950 -797 972
rect -831 938 -797 950
rect -831 882 -797 900
rect -831 866 -797 882
rect -831 814 -797 828
rect -831 794 -797 814
rect -831 746 -797 756
rect -831 722 -797 746
rect -831 678 -797 684
rect -831 650 -797 678
rect -831 610 -797 612
rect -831 578 -797 610
rect -831 508 -797 540
rect -831 506 -797 508
rect -831 440 -797 468
rect -831 434 -797 440
rect -831 372 -797 396
rect -831 362 -797 372
rect -831 304 -797 324
rect -831 290 -797 304
rect -831 236 -797 252
rect -831 218 -797 236
rect -831 168 -797 180
rect -831 146 -797 168
rect -683 950 -649 972
rect -683 938 -649 950
rect -683 882 -649 900
rect -683 866 -649 882
rect -683 814 -649 828
rect -683 794 -649 814
rect -683 746 -649 756
rect -683 722 -649 746
rect -683 678 -649 684
rect -683 650 -649 678
rect -683 610 -649 612
rect -683 578 -649 610
rect -683 508 -649 540
rect -683 506 -649 508
rect -683 440 -649 468
rect -683 434 -649 440
rect -683 372 -649 396
rect -683 362 -649 372
rect -683 304 -649 324
rect -683 290 -649 304
rect -683 236 -649 252
rect -683 218 -649 236
rect -683 168 -649 180
rect -683 146 -649 168
rect -535 950 -501 972
rect -535 938 -501 950
rect -535 882 -501 900
rect -535 866 -501 882
rect -535 814 -501 828
rect -535 794 -501 814
rect -535 746 -501 756
rect -535 722 -501 746
rect -535 678 -501 684
rect -535 650 -501 678
rect -535 610 -501 612
rect -535 578 -501 610
rect -535 508 -501 540
rect -535 506 -501 508
rect -535 440 -501 468
rect -535 434 -501 440
rect -535 372 -501 396
rect -535 362 -501 372
rect -535 304 -501 324
rect -535 290 -501 304
rect -535 236 -501 252
rect -535 218 -501 236
rect -535 168 -501 180
rect -535 146 -501 168
rect -387 950 -353 972
rect -387 938 -353 950
rect -387 882 -353 900
rect -387 866 -353 882
rect -387 814 -353 828
rect -387 794 -353 814
rect -387 746 -353 756
rect -387 722 -353 746
rect -387 678 -353 684
rect -387 650 -353 678
rect -387 610 -353 612
rect -387 578 -353 610
rect -387 508 -353 540
rect -387 506 -353 508
rect -387 440 -353 468
rect -387 434 -353 440
rect -387 372 -353 396
rect -387 362 -353 372
rect -387 304 -353 324
rect -387 290 -353 304
rect -387 236 -353 252
rect -387 218 -353 236
rect -387 168 -353 180
rect -387 146 -353 168
rect -239 950 -205 972
rect -239 938 -205 950
rect -239 882 -205 900
rect -239 866 -205 882
rect -239 814 -205 828
rect -239 794 -205 814
rect -239 746 -205 756
rect -239 722 -205 746
rect -239 678 -205 684
rect -239 650 -205 678
rect -239 610 -205 612
rect -239 578 -205 610
rect -239 508 -205 540
rect -239 506 -205 508
rect -239 440 -205 468
rect -239 434 -205 440
rect -239 372 -205 396
rect -239 362 -205 372
rect -239 304 -205 324
rect -239 290 -205 304
rect -239 236 -205 252
rect -239 218 -205 236
rect -239 168 -205 180
rect -239 146 -205 168
rect -91 950 -57 972
rect -91 938 -57 950
rect -91 882 -57 900
rect -91 866 -57 882
rect -91 814 -57 828
rect -91 794 -57 814
rect -91 746 -57 756
rect -91 722 -57 746
rect -91 678 -57 684
rect -91 650 -57 678
rect -91 610 -57 612
rect -91 578 -57 610
rect -91 508 -57 540
rect -91 506 -57 508
rect -91 440 -57 468
rect -91 434 -57 440
rect -91 372 -57 396
rect -91 362 -57 372
rect -91 304 -57 324
rect -91 290 -57 304
rect -91 236 -57 252
rect -91 218 -57 236
rect -91 168 -57 180
rect -91 146 -57 168
rect 57 950 91 972
rect 57 938 91 950
rect 57 882 91 900
rect 57 866 91 882
rect 57 814 91 828
rect 57 794 91 814
rect 57 746 91 756
rect 57 722 91 746
rect 57 678 91 684
rect 57 650 91 678
rect 57 610 91 612
rect 57 578 91 610
rect 57 508 91 540
rect 57 506 91 508
rect 57 440 91 468
rect 57 434 91 440
rect 57 372 91 396
rect 57 362 91 372
rect 57 304 91 324
rect 57 290 91 304
rect 57 236 91 252
rect 57 218 91 236
rect 57 168 91 180
rect 57 146 91 168
rect 205 950 239 972
rect 205 938 239 950
rect 205 882 239 900
rect 205 866 239 882
rect 205 814 239 828
rect 205 794 239 814
rect 205 746 239 756
rect 205 722 239 746
rect 205 678 239 684
rect 205 650 239 678
rect 205 610 239 612
rect 205 578 239 610
rect 205 508 239 540
rect 205 506 239 508
rect 205 440 239 468
rect 205 434 239 440
rect 205 372 239 396
rect 205 362 239 372
rect 205 304 239 324
rect 205 290 239 304
rect 205 236 239 252
rect 205 218 239 236
rect 205 168 239 180
rect 205 146 239 168
rect 353 950 387 972
rect 353 938 387 950
rect 353 882 387 900
rect 353 866 387 882
rect 353 814 387 828
rect 353 794 387 814
rect 353 746 387 756
rect 353 722 387 746
rect 353 678 387 684
rect 353 650 387 678
rect 353 610 387 612
rect 353 578 387 610
rect 353 508 387 540
rect 353 506 387 508
rect 353 440 387 468
rect 353 434 387 440
rect 353 372 387 396
rect 353 362 387 372
rect 353 304 387 324
rect 353 290 387 304
rect 353 236 387 252
rect 353 218 387 236
rect 353 168 387 180
rect 353 146 387 168
rect 501 950 535 972
rect 501 938 535 950
rect 501 882 535 900
rect 501 866 535 882
rect 501 814 535 828
rect 501 794 535 814
rect 501 746 535 756
rect 501 722 535 746
rect 501 678 535 684
rect 501 650 535 678
rect 501 610 535 612
rect 501 578 535 610
rect 501 508 535 540
rect 501 506 535 508
rect 501 440 535 468
rect 501 434 535 440
rect 501 372 535 396
rect 501 362 535 372
rect 501 304 535 324
rect 501 290 535 304
rect 501 236 535 252
rect 501 218 535 236
rect 501 168 535 180
rect 501 146 535 168
rect 649 950 683 972
rect 649 938 683 950
rect 649 882 683 900
rect 649 866 683 882
rect 649 814 683 828
rect 649 794 683 814
rect 649 746 683 756
rect 649 722 683 746
rect 649 678 683 684
rect 649 650 683 678
rect 649 610 683 612
rect 649 578 683 610
rect 649 508 683 540
rect 649 506 683 508
rect 649 440 683 468
rect 649 434 683 440
rect 649 372 683 396
rect 649 362 683 372
rect 649 304 683 324
rect 649 290 683 304
rect 649 236 683 252
rect 649 218 683 236
rect 649 168 683 180
rect 649 146 683 168
rect 797 950 831 972
rect 797 938 831 950
rect 797 882 831 900
rect 797 866 831 882
rect 797 814 831 828
rect 797 794 831 814
rect 797 746 831 756
rect 797 722 831 746
rect 797 678 831 684
rect 797 650 831 678
rect 797 610 831 612
rect 797 578 831 610
rect 797 508 831 540
rect 797 506 831 508
rect 797 440 831 468
rect 797 434 831 440
rect 797 372 831 396
rect 797 362 831 372
rect 797 304 831 324
rect 797 290 831 304
rect 797 236 831 252
rect 797 218 831 236
rect 797 168 831 180
rect 797 146 831 168
rect 945 950 979 972
rect 945 938 979 950
rect 945 882 979 900
rect 945 866 979 882
rect 945 814 979 828
rect 945 794 979 814
rect 945 746 979 756
rect 945 722 979 746
rect 945 678 979 684
rect 945 650 979 678
rect 945 610 979 612
rect 945 578 979 610
rect 945 508 979 540
rect 945 506 979 508
rect 945 440 979 468
rect 945 434 979 440
rect 945 372 979 396
rect 945 362 979 372
rect 945 304 979 324
rect 945 290 979 304
rect 945 236 979 252
rect 945 218 979 236
rect 945 168 979 180
rect 945 146 979 168
rect 1093 950 1127 972
rect 1093 938 1127 950
rect 1093 882 1127 900
rect 1093 866 1127 882
rect 1093 814 1127 828
rect 1093 794 1127 814
rect 1093 746 1127 756
rect 1093 722 1127 746
rect 1093 678 1127 684
rect 1093 650 1127 678
rect 1093 610 1127 612
rect 1093 578 1127 610
rect 1093 508 1127 540
rect 1093 506 1127 508
rect 1093 440 1127 468
rect 1093 434 1127 440
rect 1093 372 1127 396
rect 1093 362 1127 372
rect 1093 304 1127 324
rect 1093 290 1127 304
rect 1093 236 1127 252
rect 1093 218 1127 236
rect 1093 168 1127 180
rect 1093 146 1127 168
rect 1241 950 1275 972
rect 1241 938 1275 950
rect 1241 882 1275 900
rect 1241 866 1275 882
rect 1241 814 1275 828
rect 1241 794 1275 814
rect 1241 746 1275 756
rect 1241 722 1275 746
rect 1241 678 1275 684
rect 1241 650 1275 678
rect 1241 610 1275 612
rect 1241 578 1275 610
rect 1241 508 1275 540
rect 1241 506 1275 508
rect 1241 440 1275 468
rect 1241 434 1275 440
rect 1241 372 1275 396
rect 1241 362 1275 372
rect 1241 304 1275 324
rect 1241 290 1275 304
rect 1241 236 1275 252
rect 1241 218 1275 236
rect 1241 168 1275 180
rect 1241 146 1275 168
rect 1389 950 1423 972
rect 1389 938 1423 950
rect 1389 882 1423 900
rect 1389 866 1423 882
rect 1389 814 1423 828
rect 1389 794 1423 814
rect 1389 746 1423 756
rect 1389 722 1423 746
rect 1389 678 1423 684
rect 1389 650 1423 678
rect 1389 610 1423 612
rect 1389 578 1423 610
rect 1389 508 1423 540
rect 1389 506 1423 508
rect 1389 440 1423 468
rect 1389 434 1423 440
rect 1389 372 1423 396
rect 1389 362 1423 372
rect 1389 304 1423 324
rect 1389 290 1423 304
rect 1389 236 1423 252
rect 1389 218 1423 236
rect 1389 168 1423 180
rect 1389 146 1423 168
rect 1537 950 1571 972
rect 1537 938 1571 950
rect 1537 882 1571 900
rect 1537 866 1571 882
rect 1537 814 1571 828
rect 1537 794 1571 814
rect 1537 746 1571 756
rect 1537 722 1571 746
rect 1537 678 1571 684
rect 1537 650 1571 678
rect 1537 610 1571 612
rect 1537 578 1571 610
rect 1537 508 1571 540
rect 1537 506 1571 508
rect 1537 440 1571 468
rect 1537 434 1571 440
rect 1537 372 1571 396
rect 1537 362 1571 372
rect 1537 304 1571 324
rect 1537 290 1571 304
rect 1537 236 1571 252
rect 1537 218 1571 236
rect 1537 168 1571 180
rect 1537 146 1571 168
rect 1685 950 1719 972
rect 1685 938 1719 950
rect 1685 882 1719 900
rect 1685 866 1719 882
rect 1685 814 1719 828
rect 1685 794 1719 814
rect 1685 746 1719 756
rect 1685 722 1719 746
rect 1685 678 1719 684
rect 1685 650 1719 678
rect 1685 610 1719 612
rect 1685 578 1719 610
rect 1685 508 1719 540
rect 1685 506 1719 508
rect 1685 440 1719 468
rect 1685 434 1719 440
rect 1685 372 1719 396
rect 1685 362 1719 372
rect 1685 304 1719 324
rect 1685 290 1719 304
rect 1685 236 1719 252
rect 1685 218 1719 236
rect 1685 168 1719 180
rect 1685 146 1719 168
rect 1833 950 1867 972
rect 1833 938 1867 950
rect 1833 882 1867 900
rect 1833 866 1867 882
rect 1833 814 1867 828
rect 1833 794 1867 814
rect 1833 746 1867 756
rect 1833 722 1867 746
rect 1833 678 1867 684
rect 1833 650 1867 678
rect 1833 610 1867 612
rect 1833 578 1867 610
rect 1833 508 1867 540
rect 1833 506 1867 508
rect 1833 440 1867 468
rect 1833 434 1867 440
rect 1833 372 1867 396
rect 1833 362 1867 372
rect 1833 304 1867 324
rect 1833 290 1867 304
rect 1833 236 1867 252
rect 1833 218 1867 236
rect 1833 168 1867 180
rect 1833 146 1867 168
rect 1981 950 2015 972
rect 1981 938 2015 950
rect 1981 882 2015 900
rect 1981 866 2015 882
rect 1981 814 2015 828
rect 1981 794 2015 814
rect 1981 746 2015 756
rect 1981 722 2015 746
rect 1981 678 2015 684
rect 1981 650 2015 678
rect 1981 610 2015 612
rect 1981 578 2015 610
rect 1981 508 2015 540
rect 1981 506 2015 508
rect 1981 440 2015 468
rect 1981 434 2015 440
rect 1981 372 2015 396
rect 1981 362 2015 372
rect 1981 304 2015 324
rect 1981 290 2015 304
rect 1981 236 2015 252
rect 1981 218 2015 236
rect 1981 168 2015 180
rect 1981 146 2015 168
rect 2129 950 2163 972
rect 2129 938 2163 950
rect 2129 882 2163 900
rect 2129 866 2163 882
rect 2129 814 2163 828
rect 2129 794 2163 814
rect 2129 746 2163 756
rect 2129 722 2163 746
rect 2129 678 2163 684
rect 2129 650 2163 678
rect 2129 610 2163 612
rect 2129 578 2163 610
rect 2129 508 2163 540
rect 2129 506 2163 508
rect 2129 440 2163 468
rect 2129 434 2163 440
rect 2129 372 2163 396
rect 2129 362 2163 372
rect 2129 304 2163 324
rect 2129 290 2163 304
rect 2129 236 2163 252
rect 2129 218 2163 236
rect 2129 168 2163 180
rect 2129 146 2163 168
rect 2277 950 2311 972
rect 2277 938 2311 950
rect 2277 882 2311 900
rect 2277 866 2311 882
rect 2277 814 2311 828
rect 2277 794 2311 814
rect 2277 746 2311 756
rect 2277 722 2311 746
rect 2277 678 2311 684
rect 2277 650 2311 678
rect 2277 610 2311 612
rect 2277 578 2311 610
rect 2277 508 2311 540
rect 2277 506 2311 508
rect 2277 440 2311 468
rect 2277 434 2311 440
rect 2277 372 2311 396
rect 2277 362 2311 372
rect 2277 304 2311 324
rect 2277 290 2311 304
rect 2277 236 2311 252
rect 2277 218 2311 236
rect 2277 168 2311 180
rect 2277 146 2311 168
rect 2425 950 2459 972
rect 2425 938 2459 950
rect 2425 882 2459 900
rect 2425 866 2459 882
rect 2425 814 2459 828
rect 2425 794 2459 814
rect 2425 746 2459 756
rect 2425 722 2459 746
rect 2425 678 2459 684
rect 2425 650 2459 678
rect 2425 610 2459 612
rect 2425 578 2459 610
rect 2425 508 2459 540
rect 2425 506 2459 508
rect 2425 440 2459 468
rect 2425 434 2459 440
rect 2425 372 2459 396
rect 2425 362 2459 372
rect 2425 304 2459 324
rect 2425 290 2459 304
rect 2425 236 2459 252
rect 2425 218 2459 236
rect 2425 168 2459 180
rect 2425 146 2459 168
rect 2573 950 2607 972
rect 2573 938 2607 950
rect 2573 882 2607 900
rect 2573 866 2607 882
rect 2573 814 2607 828
rect 2573 794 2607 814
rect 2573 746 2607 756
rect 2573 722 2607 746
rect 2573 678 2607 684
rect 2573 650 2607 678
rect 2573 610 2607 612
rect 2573 578 2607 610
rect 2573 508 2607 540
rect 2573 506 2607 508
rect 2573 440 2607 468
rect 2573 434 2607 440
rect 2573 372 2607 396
rect 2573 362 2607 372
rect 2573 304 2607 324
rect 2573 290 2607 304
rect 2573 236 2607 252
rect 2573 218 2607 236
rect 2573 168 2607 180
rect 2573 146 2607 168
rect 2721 950 2755 972
rect 2721 938 2755 950
rect 2721 882 2755 900
rect 2721 866 2755 882
rect 2721 814 2755 828
rect 2721 794 2755 814
rect 2721 746 2755 756
rect 2721 722 2755 746
rect 2721 678 2755 684
rect 2721 650 2755 678
rect 2721 610 2755 612
rect 2721 578 2755 610
rect 2721 508 2755 540
rect 2721 506 2755 508
rect 2721 440 2755 468
rect 2721 434 2755 440
rect 2721 372 2755 396
rect 2721 362 2755 372
rect 2721 304 2755 324
rect 2721 290 2755 304
rect 2721 236 2755 252
rect 2721 218 2755 236
rect 2721 168 2755 180
rect 2721 146 2755 168
rect 2869 950 2903 972
rect 2869 938 2903 950
rect 2869 882 2903 900
rect 2869 866 2903 882
rect 2869 814 2903 828
rect 2869 794 2903 814
rect 2869 746 2903 756
rect 2869 722 2903 746
rect 2869 678 2903 684
rect 2869 650 2903 678
rect 2869 610 2903 612
rect 2869 578 2903 610
rect 2869 508 2903 540
rect 2869 506 2903 508
rect 2869 440 2903 468
rect 2869 434 2903 440
rect 2869 372 2903 396
rect 2869 362 2903 372
rect 2869 304 2903 324
rect 2869 290 2903 304
rect 2869 236 2903 252
rect 2869 218 2903 236
rect 2869 168 2903 180
rect 2869 146 2903 168
rect 3017 950 3051 972
rect 3017 938 3051 950
rect 3017 882 3051 900
rect 3017 866 3051 882
rect 3017 814 3051 828
rect 3017 794 3051 814
rect 3017 746 3051 756
rect 3017 722 3051 746
rect 3017 678 3051 684
rect 3017 650 3051 678
rect 3017 610 3051 612
rect 3017 578 3051 610
rect 3017 508 3051 540
rect 3017 506 3051 508
rect 3017 440 3051 468
rect 3017 434 3051 440
rect 3017 372 3051 396
rect 3017 362 3051 372
rect 3017 304 3051 324
rect 3017 290 3051 304
rect 3017 236 3051 252
rect 3017 218 3051 236
rect 3017 168 3051 180
rect 3017 146 3051 168
rect 3165 950 3199 972
rect 3165 938 3199 950
rect 3165 882 3199 900
rect 3165 866 3199 882
rect 3165 814 3199 828
rect 3165 794 3199 814
rect 3165 746 3199 756
rect 3165 722 3199 746
rect 3165 678 3199 684
rect 3165 650 3199 678
rect 3165 610 3199 612
rect 3165 578 3199 610
rect 3165 508 3199 540
rect 3165 506 3199 508
rect 3165 440 3199 468
rect 3165 434 3199 440
rect 3165 372 3199 396
rect 3165 362 3199 372
rect 3165 304 3199 324
rect 3165 290 3199 304
rect 3165 236 3199 252
rect 3165 218 3199 236
rect 3165 168 3199 180
rect 3165 146 3199 168
rect 3313 950 3347 972
rect 3313 938 3347 950
rect 3313 882 3347 900
rect 3313 866 3347 882
rect 3313 814 3347 828
rect 3313 794 3347 814
rect 3313 746 3347 756
rect 3313 722 3347 746
rect 3313 678 3347 684
rect 3313 650 3347 678
rect 3313 610 3347 612
rect 3313 578 3347 610
rect 3313 508 3347 540
rect 3313 506 3347 508
rect 3313 440 3347 468
rect 3313 434 3347 440
rect 3313 372 3347 396
rect 3313 362 3347 372
rect 3313 304 3347 324
rect 3313 290 3347 304
rect 3313 236 3347 252
rect 3313 218 3347 236
rect 3313 168 3347 180
rect 3313 146 3347 168
rect 3461 950 3495 972
rect 3461 938 3495 950
rect 3461 882 3495 900
rect 3461 866 3495 882
rect 3461 814 3495 828
rect 3461 794 3495 814
rect 3461 746 3495 756
rect 3461 722 3495 746
rect 3461 678 3495 684
rect 3461 650 3495 678
rect 3461 610 3495 612
rect 3461 578 3495 610
rect 3461 508 3495 540
rect 3461 506 3495 508
rect 3461 440 3495 468
rect 3461 434 3495 440
rect 3461 372 3495 396
rect 3461 362 3495 372
rect 3461 304 3495 324
rect 3461 290 3495 304
rect 3461 236 3495 252
rect 3461 218 3495 236
rect 3461 168 3495 180
rect 3461 146 3495 168
rect 3609 950 3643 972
rect 3609 938 3643 950
rect 3609 882 3643 900
rect 3609 866 3643 882
rect 3609 814 3643 828
rect 3609 794 3643 814
rect 3609 746 3643 756
rect 3609 722 3643 746
rect 3609 678 3643 684
rect 3609 650 3643 678
rect 3609 610 3643 612
rect 3609 578 3643 610
rect 3609 508 3643 540
rect 3609 506 3643 508
rect 3609 440 3643 468
rect 3609 434 3643 440
rect 3609 372 3643 396
rect 3609 362 3643 372
rect 3609 304 3643 324
rect 3609 290 3643 304
rect 3609 236 3643 252
rect 3609 218 3643 236
rect 3609 168 3643 180
rect 3609 146 3643 168
rect 3757 950 3791 972
rect 3757 938 3791 950
rect 3757 882 3791 900
rect 3757 866 3791 882
rect 3757 814 3791 828
rect 3757 794 3791 814
rect 3757 746 3791 756
rect 3757 722 3791 746
rect 3757 678 3791 684
rect 3757 650 3791 678
rect 3757 610 3791 612
rect 3757 578 3791 610
rect 3757 508 3791 540
rect 3757 506 3791 508
rect 3757 440 3791 468
rect 3757 434 3791 440
rect 3757 372 3791 396
rect 3757 362 3791 372
rect 3757 304 3791 324
rect 3757 290 3791 304
rect 3757 236 3791 252
rect 3757 218 3791 236
rect 3757 168 3791 180
rect 3757 146 3791 168
rect 3905 950 3939 972
rect 3905 938 3939 950
rect 3905 882 3939 900
rect 3905 866 3939 882
rect 3905 814 3939 828
rect 3905 794 3939 814
rect 3905 746 3939 756
rect 3905 722 3939 746
rect 3905 678 3939 684
rect 3905 650 3939 678
rect 3905 610 3939 612
rect 3905 578 3939 610
rect 3905 508 3939 540
rect 3905 506 3939 508
rect 3905 440 3939 468
rect 3905 434 3939 440
rect 3905 372 3939 396
rect 3905 362 3939 372
rect 3905 304 3939 324
rect 3905 290 3939 304
rect 3905 236 3939 252
rect 3905 218 3939 236
rect 3905 168 3939 180
rect 3905 146 3939 168
rect 4053 950 4087 972
rect 4053 938 4087 950
rect 4053 882 4087 900
rect 4053 866 4087 882
rect 4053 814 4087 828
rect 4053 794 4087 814
rect 4053 746 4087 756
rect 4053 722 4087 746
rect 4053 678 4087 684
rect 4053 650 4087 678
rect 4053 610 4087 612
rect 4053 578 4087 610
rect 4053 508 4087 540
rect 4053 506 4087 508
rect 4053 440 4087 468
rect 4053 434 4087 440
rect 4053 372 4087 396
rect 4053 362 4087 372
rect 4053 304 4087 324
rect 4053 290 4087 304
rect 4053 236 4087 252
rect 4053 218 4087 236
rect 4053 168 4087 180
rect 4053 146 4087 168
rect 4201 950 4235 972
rect 4201 938 4235 950
rect 4201 882 4235 900
rect 4201 866 4235 882
rect 4201 814 4235 828
rect 4201 794 4235 814
rect 4201 746 4235 756
rect 4201 722 4235 746
rect 4201 678 4235 684
rect 4201 650 4235 678
rect 4201 610 4235 612
rect 4201 578 4235 610
rect 4201 508 4235 540
rect 4201 506 4235 508
rect 4201 440 4235 468
rect 4201 434 4235 440
rect 4201 372 4235 396
rect 4201 362 4235 372
rect 4201 304 4235 324
rect 4201 290 4235 304
rect 4201 236 4235 252
rect 4201 218 4235 236
rect 4201 168 4235 180
rect 4201 146 4235 168
rect 4349 950 4383 972
rect 4349 938 4383 950
rect 4349 882 4383 900
rect 4349 866 4383 882
rect 4349 814 4383 828
rect 4349 794 4383 814
rect 4349 746 4383 756
rect 4349 722 4383 746
rect 4349 678 4383 684
rect 4349 650 4383 678
rect 4349 610 4383 612
rect 4349 578 4383 610
rect 4349 508 4383 540
rect 4349 506 4383 508
rect 4349 440 4383 468
rect 4349 434 4383 440
rect 4349 372 4383 396
rect 4349 362 4383 372
rect 4349 304 4383 324
rect 4349 290 4383 304
rect 4349 236 4383 252
rect 4349 218 4383 236
rect 4349 168 4383 180
rect 4349 146 4383 168
rect 4497 950 4531 972
rect 4497 938 4531 950
rect 4497 882 4531 900
rect 4497 866 4531 882
rect 4497 814 4531 828
rect 4497 794 4531 814
rect 4497 746 4531 756
rect 4497 722 4531 746
rect 4497 678 4531 684
rect 4497 650 4531 678
rect 4497 610 4531 612
rect 4497 578 4531 610
rect 4497 508 4531 540
rect 4497 506 4531 508
rect 4497 440 4531 468
rect 4497 434 4531 440
rect 4497 372 4531 396
rect 4497 362 4531 372
rect 4497 304 4531 324
rect 4497 290 4531 304
rect 4497 236 4531 252
rect 4497 218 4531 236
rect 4497 168 4531 180
rect 4497 146 4531 168
rect 4645 950 4679 972
rect 4645 938 4679 950
rect 4645 882 4679 900
rect 4645 866 4679 882
rect 4645 814 4679 828
rect 4645 794 4679 814
rect 4645 746 4679 756
rect 4645 722 4679 746
rect 4645 678 4679 684
rect 4645 650 4679 678
rect 4645 610 4679 612
rect 4645 578 4679 610
rect 4645 508 4679 540
rect 4645 506 4679 508
rect 4645 440 4679 468
rect 4645 434 4679 440
rect 4645 372 4679 396
rect 4645 362 4679 372
rect 4645 304 4679 324
rect 4645 290 4679 304
rect 4645 236 4679 252
rect 4645 218 4679 236
rect 4645 168 4679 180
rect 4645 146 4679 168
rect 4793 950 4827 972
rect 4793 938 4827 950
rect 4793 882 4827 900
rect 4793 866 4827 882
rect 4793 814 4827 828
rect 4793 794 4827 814
rect 4793 746 4827 756
rect 4793 722 4827 746
rect 4793 678 4827 684
rect 4793 650 4827 678
rect 4793 610 4827 612
rect 4793 578 4827 610
rect 4793 508 4827 540
rect 4793 506 4827 508
rect 4793 440 4827 468
rect 4793 434 4827 440
rect 4793 372 4827 396
rect 4793 362 4827 372
rect 4793 304 4827 324
rect 4793 290 4827 304
rect 4793 236 4827 252
rect 4793 218 4827 236
rect 4793 168 4827 180
rect 4793 146 4827 168
rect 4941 950 4975 972
rect 4941 938 4975 950
rect 4941 882 4975 900
rect 4941 866 4975 882
rect 4941 814 4975 828
rect 4941 794 4975 814
rect 4941 746 4975 756
rect 4941 722 4975 746
rect 4941 678 4975 684
rect 4941 650 4975 678
rect 4941 610 4975 612
rect 4941 578 4975 610
rect 4941 508 4975 540
rect 4941 506 4975 508
rect 4941 440 4975 468
rect 4941 434 4975 440
rect 4941 372 4975 396
rect 4941 362 4975 372
rect 4941 304 4975 324
rect 4941 290 4975 304
rect 4941 236 4975 252
rect 4941 218 4975 236
rect 4941 168 4975 180
rect 4941 146 4975 168
rect 5089 950 5123 972
rect 5089 938 5123 950
rect 5089 882 5123 900
rect 5089 866 5123 882
rect 5089 814 5123 828
rect 5089 794 5123 814
rect 5089 746 5123 756
rect 5089 722 5123 746
rect 5089 678 5123 684
rect 5089 650 5123 678
rect 5089 610 5123 612
rect 5089 578 5123 610
rect 5089 508 5123 540
rect 5089 506 5123 508
rect 5089 440 5123 468
rect 5089 434 5123 440
rect 5089 372 5123 396
rect 5089 362 5123 372
rect 5089 304 5123 324
rect 5089 290 5123 304
rect 5089 236 5123 252
rect 5089 218 5123 236
rect 5089 168 5123 180
rect 5089 146 5123 168
rect 5237 950 5271 972
rect 5237 938 5271 950
rect 5237 882 5271 900
rect 5237 866 5271 882
rect 5237 814 5271 828
rect 5237 794 5271 814
rect 5237 746 5271 756
rect 5237 722 5271 746
rect 5237 678 5271 684
rect 5237 650 5271 678
rect 5237 610 5271 612
rect 5237 578 5271 610
rect 5237 508 5271 540
rect 5237 506 5271 508
rect 5237 440 5271 468
rect 5237 434 5271 440
rect 5237 372 5271 396
rect 5237 362 5271 372
rect 5237 304 5271 324
rect 5237 290 5271 304
rect 5237 236 5271 252
rect 5237 218 5271 236
rect 5237 168 5271 180
rect 5237 146 5271 168
rect 5385 950 5419 972
rect 5385 938 5419 950
rect 5385 882 5419 900
rect 5385 866 5419 882
rect 5385 814 5419 828
rect 5385 794 5419 814
rect 5385 746 5419 756
rect 5385 722 5419 746
rect 5385 678 5419 684
rect 5385 650 5419 678
rect 5385 610 5419 612
rect 5385 578 5419 610
rect 5385 508 5419 540
rect 5385 506 5419 508
rect 5385 440 5419 468
rect 5385 434 5419 440
rect 5385 372 5419 396
rect 5385 362 5419 372
rect 5385 304 5419 324
rect 5385 290 5419 304
rect 5385 236 5419 252
rect 5385 218 5419 236
rect 5385 168 5419 180
rect 5385 146 5419 168
rect 5533 950 5567 972
rect 5533 938 5567 950
rect 5533 882 5567 900
rect 5533 866 5567 882
rect 5533 814 5567 828
rect 5533 794 5567 814
rect 5533 746 5567 756
rect 5533 722 5567 746
rect 5533 678 5567 684
rect 5533 650 5567 678
rect 5533 610 5567 612
rect 5533 578 5567 610
rect 5533 508 5567 540
rect 5533 506 5567 508
rect 5533 440 5567 468
rect 5533 434 5567 440
rect 5533 372 5567 396
rect 5533 362 5567 372
rect 5533 304 5567 324
rect 5533 290 5567 304
rect 5533 236 5567 252
rect 5533 218 5567 236
rect 5533 168 5567 180
rect 5533 146 5567 168
rect -5493 37 -5459 71
rect -5345 37 -5311 71
rect -5197 37 -5163 71
rect -5049 37 -5015 71
rect -4901 37 -4867 71
rect -4753 37 -4719 71
rect -4605 37 -4571 71
rect -4457 37 -4423 71
rect -4309 37 -4275 71
rect -4161 37 -4127 71
rect -4013 37 -3979 71
rect -3865 37 -3831 71
rect -3717 37 -3683 71
rect -3569 37 -3535 71
rect -3421 37 -3387 71
rect -3273 37 -3239 71
rect -3125 37 -3091 71
rect -2977 37 -2943 71
rect -2829 37 -2795 71
rect -2681 37 -2647 71
rect -2533 37 -2499 71
rect -2385 37 -2351 71
rect -2237 37 -2203 71
rect -2089 37 -2055 71
rect -1941 37 -1907 71
rect -1793 37 -1759 71
rect -1645 37 -1611 71
rect -1497 37 -1463 71
rect -1349 37 -1315 71
rect -1201 37 -1167 71
rect -1053 37 -1019 71
rect -905 37 -871 71
rect -757 37 -723 71
rect -609 37 -575 71
rect -461 37 -427 71
rect -313 37 -279 71
rect -165 37 -131 71
rect -17 37 17 71
rect 131 37 165 71
rect 279 37 313 71
rect 427 37 461 71
rect 575 37 609 71
rect 723 37 757 71
rect 871 37 905 71
rect 1019 37 1053 71
rect 1167 37 1201 71
rect 1315 37 1349 71
rect 1463 37 1497 71
rect 1611 37 1645 71
rect 1759 37 1793 71
rect 1907 37 1941 71
rect 2055 37 2089 71
rect 2203 37 2237 71
rect 2351 37 2385 71
rect 2499 37 2533 71
rect 2647 37 2681 71
rect 2795 37 2829 71
rect 2943 37 2977 71
rect 3091 37 3125 71
rect 3239 37 3273 71
rect 3387 37 3421 71
rect 3535 37 3569 71
rect 3683 37 3717 71
rect 3831 37 3865 71
rect 3979 37 4013 71
rect 4127 37 4161 71
rect 4275 37 4309 71
rect 4423 37 4457 71
rect 4571 37 4605 71
rect 4719 37 4753 71
rect 4867 37 4901 71
rect 5015 37 5049 71
rect 5163 37 5197 71
rect 5311 37 5345 71
rect 5459 37 5493 71
rect -5493 -71 -5459 -37
rect -5345 -71 -5311 -37
rect -5197 -71 -5163 -37
rect -5049 -71 -5015 -37
rect -4901 -71 -4867 -37
rect -4753 -71 -4719 -37
rect -4605 -71 -4571 -37
rect -4457 -71 -4423 -37
rect -4309 -71 -4275 -37
rect -4161 -71 -4127 -37
rect -4013 -71 -3979 -37
rect -3865 -71 -3831 -37
rect -3717 -71 -3683 -37
rect -3569 -71 -3535 -37
rect -3421 -71 -3387 -37
rect -3273 -71 -3239 -37
rect -3125 -71 -3091 -37
rect -2977 -71 -2943 -37
rect -2829 -71 -2795 -37
rect -2681 -71 -2647 -37
rect -2533 -71 -2499 -37
rect -2385 -71 -2351 -37
rect -2237 -71 -2203 -37
rect -2089 -71 -2055 -37
rect -1941 -71 -1907 -37
rect -1793 -71 -1759 -37
rect -1645 -71 -1611 -37
rect -1497 -71 -1463 -37
rect -1349 -71 -1315 -37
rect -1201 -71 -1167 -37
rect -1053 -71 -1019 -37
rect -905 -71 -871 -37
rect -757 -71 -723 -37
rect -609 -71 -575 -37
rect -461 -71 -427 -37
rect -313 -71 -279 -37
rect -165 -71 -131 -37
rect -17 -71 17 -37
rect 131 -71 165 -37
rect 279 -71 313 -37
rect 427 -71 461 -37
rect 575 -71 609 -37
rect 723 -71 757 -37
rect 871 -71 905 -37
rect 1019 -71 1053 -37
rect 1167 -71 1201 -37
rect 1315 -71 1349 -37
rect 1463 -71 1497 -37
rect 1611 -71 1645 -37
rect 1759 -71 1793 -37
rect 1907 -71 1941 -37
rect 2055 -71 2089 -37
rect 2203 -71 2237 -37
rect 2351 -71 2385 -37
rect 2499 -71 2533 -37
rect 2647 -71 2681 -37
rect 2795 -71 2829 -37
rect 2943 -71 2977 -37
rect 3091 -71 3125 -37
rect 3239 -71 3273 -37
rect 3387 -71 3421 -37
rect 3535 -71 3569 -37
rect 3683 -71 3717 -37
rect 3831 -71 3865 -37
rect 3979 -71 4013 -37
rect 4127 -71 4161 -37
rect 4275 -71 4309 -37
rect 4423 -71 4457 -37
rect 4571 -71 4605 -37
rect 4719 -71 4753 -37
rect 4867 -71 4901 -37
rect 5015 -71 5049 -37
rect 5163 -71 5197 -37
rect 5311 -71 5345 -37
rect 5459 -71 5493 -37
rect -5567 -168 -5533 -146
rect -5567 -180 -5533 -168
rect -5567 -236 -5533 -218
rect -5567 -252 -5533 -236
rect -5567 -304 -5533 -290
rect -5567 -324 -5533 -304
rect -5567 -372 -5533 -362
rect -5567 -396 -5533 -372
rect -5567 -440 -5533 -434
rect -5567 -468 -5533 -440
rect -5567 -508 -5533 -506
rect -5567 -540 -5533 -508
rect -5567 -610 -5533 -578
rect -5567 -612 -5533 -610
rect -5567 -678 -5533 -650
rect -5567 -684 -5533 -678
rect -5567 -746 -5533 -722
rect -5567 -756 -5533 -746
rect -5567 -814 -5533 -794
rect -5567 -828 -5533 -814
rect -5567 -882 -5533 -866
rect -5567 -900 -5533 -882
rect -5567 -950 -5533 -938
rect -5567 -972 -5533 -950
rect -5419 -168 -5385 -146
rect -5419 -180 -5385 -168
rect -5419 -236 -5385 -218
rect -5419 -252 -5385 -236
rect -5419 -304 -5385 -290
rect -5419 -324 -5385 -304
rect -5419 -372 -5385 -362
rect -5419 -396 -5385 -372
rect -5419 -440 -5385 -434
rect -5419 -468 -5385 -440
rect -5419 -508 -5385 -506
rect -5419 -540 -5385 -508
rect -5419 -610 -5385 -578
rect -5419 -612 -5385 -610
rect -5419 -678 -5385 -650
rect -5419 -684 -5385 -678
rect -5419 -746 -5385 -722
rect -5419 -756 -5385 -746
rect -5419 -814 -5385 -794
rect -5419 -828 -5385 -814
rect -5419 -882 -5385 -866
rect -5419 -900 -5385 -882
rect -5419 -950 -5385 -938
rect -5419 -972 -5385 -950
rect -5271 -168 -5237 -146
rect -5271 -180 -5237 -168
rect -5271 -236 -5237 -218
rect -5271 -252 -5237 -236
rect -5271 -304 -5237 -290
rect -5271 -324 -5237 -304
rect -5271 -372 -5237 -362
rect -5271 -396 -5237 -372
rect -5271 -440 -5237 -434
rect -5271 -468 -5237 -440
rect -5271 -508 -5237 -506
rect -5271 -540 -5237 -508
rect -5271 -610 -5237 -578
rect -5271 -612 -5237 -610
rect -5271 -678 -5237 -650
rect -5271 -684 -5237 -678
rect -5271 -746 -5237 -722
rect -5271 -756 -5237 -746
rect -5271 -814 -5237 -794
rect -5271 -828 -5237 -814
rect -5271 -882 -5237 -866
rect -5271 -900 -5237 -882
rect -5271 -950 -5237 -938
rect -5271 -972 -5237 -950
rect -5123 -168 -5089 -146
rect -5123 -180 -5089 -168
rect -5123 -236 -5089 -218
rect -5123 -252 -5089 -236
rect -5123 -304 -5089 -290
rect -5123 -324 -5089 -304
rect -5123 -372 -5089 -362
rect -5123 -396 -5089 -372
rect -5123 -440 -5089 -434
rect -5123 -468 -5089 -440
rect -5123 -508 -5089 -506
rect -5123 -540 -5089 -508
rect -5123 -610 -5089 -578
rect -5123 -612 -5089 -610
rect -5123 -678 -5089 -650
rect -5123 -684 -5089 -678
rect -5123 -746 -5089 -722
rect -5123 -756 -5089 -746
rect -5123 -814 -5089 -794
rect -5123 -828 -5089 -814
rect -5123 -882 -5089 -866
rect -5123 -900 -5089 -882
rect -5123 -950 -5089 -938
rect -5123 -972 -5089 -950
rect -4975 -168 -4941 -146
rect -4975 -180 -4941 -168
rect -4975 -236 -4941 -218
rect -4975 -252 -4941 -236
rect -4975 -304 -4941 -290
rect -4975 -324 -4941 -304
rect -4975 -372 -4941 -362
rect -4975 -396 -4941 -372
rect -4975 -440 -4941 -434
rect -4975 -468 -4941 -440
rect -4975 -508 -4941 -506
rect -4975 -540 -4941 -508
rect -4975 -610 -4941 -578
rect -4975 -612 -4941 -610
rect -4975 -678 -4941 -650
rect -4975 -684 -4941 -678
rect -4975 -746 -4941 -722
rect -4975 -756 -4941 -746
rect -4975 -814 -4941 -794
rect -4975 -828 -4941 -814
rect -4975 -882 -4941 -866
rect -4975 -900 -4941 -882
rect -4975 -950 -4941 -938
rect -4975 -972 -4941 -950
rect -4827 -168 -4793 -146
rect -4827 -180 -4793 -168
rect -4827 -236 -4793 -218
rect -4827 -252 -4793 -236
rect -4827 -304 -4793 -290
rect -4827 -324 -4793 -304
rect -4827 -372 -4793 -362
rect -4827 -396 -4793 -372
rect -4827 -440 -4793 -434
rect -4827 -468 -4793 -440
rect -4827 -508 -4793 -506
rect -4827 -540 -4793 -508
rect -4827 -610 -4793 -578
rect -4827 -612 -4793 -610
rect -4827 -678 -4793 -650
rect -4827 -684 -4793 -678
rect -4827 -746 -4793 -722
rect -4827 -756 -4793 -746
rect -4827 -814 -4793 -794
rect -4827 -828 -4793 -814
rect -4827 -882 -4793 -866
rect -4827 -900 -4793 -882
rect -4827 -950 -4793 -938
rect -4827 -972 -4793 -950
rect -4679 -168 -4645 -146
rect -4679 -180 -4645 -168
rect -4679 -236 -4645 -218
rect -4679 -252 -4645 -236
rect -4679 -304 -4645 -290
rect -4679 -324 -4645 -304
rect -4679 -372 -4645 -362
rect -4679 -396 -4645 -372
rect -4679 -440 -4645 -434
rect -4679 -468 -4645 -440
rect -4679 -508 -4645 -506
rect -4679 -540 -4645 -508
rect -4679 -610 -4645 -578
rect -4679 -612 -4645 -610
rect -4679 -678 -4645 -650
rect -4679 -684 -4645 -678
rect -4679 -746 -4645 -722
rect -4679 -756 -4645 -746
rect -4679 -814 -4645 -794
rect -4679 -828 -4645 -814
rect -4679 -882 -4645 -866
rect -4679 -900 -4645 -882
rect -4679 -950 -4645 -938
rect -4679 -972 -4645 -950
rect -4531 -168 -4497 -146
rect -4531 -180 -4497 -168
rect -4531 -236 -4497 -218
rect -4531 -252 -4497 -236
rect -4531 -304 -4497 -290
rect -4531 -324 -4497 -304
rect -4531 -372 -4497 -362
rect -4531 -396 -4497 -372
rect -4531 -440 -4497 -434
rect -4531 -468 -4497 -440
rect -4531 -508 -4497 -506
rect -4531 -540 -4497 -508
rect -4531 -610 -4497 -578
rect -4531 -612 -4497 -610
rect -4531 -678 -4497 -650
rect -4531 -684 -4497 -678
rect -4531 -746 -4497 -722
rect -4531 -756 -4497 -746
rect -4531 -814 -4497 -794
rect -4531 -828 -4497 -814
rect -4531 -882 -4497 -866
rect -4531 -900 -4497 -882
rect -4531 -950 -4497 -938
rect -4531 -972 -4497 -950
rect -4383 -168 -4349 -146
rect -4383 -180 -4349 -168
rect -4383 -236 -4349 -218
rect -4383 -252 -4349 -236
rect -4383 -304 -4349 -290
rect -4383 -324 -4349 -304
rect -4383 -372 -4349 -362
rect -4383 -396 -4349 -372
rect -4383 -440 -4349 -434
rect -4383 -468 -4349 -440
rect -4383 -508 -4349 -506
rect -4383 -540 -4349 -508
rect -4383 -610 -4349 -578
rect -4383 -612 -4349 -610
rect -4383 -678 -4349 -650
rect -4383 -684 -4349 -678
rect -4383 -746 -4349 -722
rect -4383 -756 -4349 -746
rect -4383 -814 -4349 -794
rect -4383 -828 -4349 -814
rect -4383 -882 -4349 -866
rect -4383 -900 -4349 -882
rect -4383 -950 -4349 -938
rect -4383 -972 -4349 -950
rect -4235 -168 -4201 -146
rect -4235 -180 -4201 -168
rect -4235 -236 -4201 -218
rect -4235 -252 -4201 -236
rect -4235 -304 -4201 -290
rect -4235 -324 -4201 -304
rect -4235 -372 -4201 -362
rect -4235 -396 -4201 -372
rect -4235 -440 -4201 -434
rect -4235 -468 -4201 -440
rect -4235 -508 -4201 -506
rect -4235 -540 -4201 -508
rect -4235 -610 -4201 -578
rect -4235 -612 -4201 -610
rect -4235 -678 -4201 -650
rect -4235 -684 -4201 -678
rect -4235 -746 -4201 -722
rect -4235 -756 -4201 -746
rect -4235 -814 -4201 -794
rect -4235 -828 -4201 -814
rect -4235 -882 -4201 -866
rect -4235 -900 -4201 -882
rect -4235 -950 -4201 -938
rect -4235 -972 -4201 -950
rect -4087 -168 -4053 -146
rect -4087 -180 -4053 -168
rect -4087 -236 -4053 -218
rect -4087 -252 -4053 -236
rect -4087 -304 -4053 -290
rect -4087 -324 -4053 -304
rect -4087 -372 -4053 -362
rect -4087 -396 -4053 -372
rect -4087 -440 -4053 -434
rect -4087 -468 -4053 -440
rect -4087 -508 -4053 -506
rect -4087 -540 -4053 -508
rect -4087 -610 -4053 -578
rect -4087 -612 -4053 -610
rect -4087 -678 -4053 -650
rect -4087 -684 -4053 -678
rect -4087 -746 -4053 -722
rect -4087 -756 -4053 -746
rect -4087 -814 -4053 -794
rect -4087 -828 -4053 -814
rect -4087 -882 -4053 -866
rect -4087 -900 -4053 -882
rect -4087 -950 -4053 -938
rect -4087 -972 -4053 -950
rect -3939 -168 -3905 -146
rect -3939 -180 -3905 -168
rect -3939 -236 -3905 -218
rect -3939 -252 -3905 -236
rect -3939 -304 -3905 -290
rect -3939 -324 -3905 -304
rect -3939 -372 -3905 -362
rect -3939 -396 -3905 -372
rect -3939 -440 -3905 -434
rect -3939 -468 -3905 -440
rect -3939 -508 -3905 -506
rect -3939 -540 -3905 -508
rect -3939 -610 -3905 -578
rect -3939 -612 -3905 -610
rect -3939 -678 -3905 -650
rect -3939 -684 -3905 -678
rect -3939 -746 -3905 -722
rect -3939 -756 -3905 -746
rect -3939 -814 -3905 -794
rect -3939 -828 -3905 -814
rect -3939 -882 -3905 -866
rect -3939 -900 -3905 -882
rect -3939 -950 -3905 -938
rect -3939 -972 -3905 -950
rect -3791 -168 -3757 -146
rect -3791 -180 -3757 -168
rect -3791 -236 -3757 -218
rect -3791 -252 -3757 -236
rect -3791 -304 -3757 -290
rect -3791 -324 -3757 -304
rect -3791 -372 -3757 -362
rect -3791 -396 -3757 -372
rect -3791 -440 -3757 -434
rect -3791 -468 -3757 -440
rect -3791 -508 -3757 -506
rect -3791 -540 -3757 -508
rect -3791 -610 -3757 -578
rect -3791 -612 -3757 -610
rect -3791 -678 -3757 -650
rect -3791 -684 -3757 -678
rect -3791 -746 -3757 -722
rect -3791 -756 -3757 -746
rect -3791 -814 -3757 -794
rect -3791 -828 -3757 -814
rect -3791 -882 -3757 -866
rect -3791 -900 -3757 -882
rect -3791 -950 -3757 -938
rect -3791 -972 -3757 -950
rect -3643 -168 -3609 -146
rect -3643 -180 -3609 -168
rect -3643 -236 -3609 -218
rect -3643 -252 -3609 -236
rect -3643 -304 -3609 -290
rect -3643 -324 -3609 -304
rect -3643 -372 -3609 -362
rect -3643 -396 -3609 -372
rect -3643 -440 -3609 -434
rect -3643 -468 -3609 -440
rect -3643 -508 -3609 -506
rect -3643 -540 -3609 -508
rect -3643 -610 -3609 -578
rect -3643 -612 -3609 -610
rect -3643 -678 -3609 -650
rect -3643 -684 -3609 -678
rect -3643 -746 -3609 -722
rect -3643 -756 -3609 -746
rect -3643 -814 -3609 -794
rect -3643 -828 -3609 -814
rect -3643 -882 -3609 -866
rect -3643 -900 -3609 -882
rect -3643 -950 -3609 -938
rect -3643 -972 -3609 -950
rect -3495 -168 -3461 -146
rect -3495 -180 -3461 -168
rect -3495 -236 -3461 -218
rect -3495 -252 -3461 -236
rect -3495 -304 -3461 -290
rect -3495 -324 -3461 -304
rect -3495 -372 -3461 -362
rect -3495 -396 -3461 -372
rect -3495 -440 -3461 -434
rect -3495 -468 -3461 -440
rect -3495 -508 -3461 -506
rect -3495 -540 -3461 -508
rect -3495 -610 -3461 -578
rect -3495 -612 -3461 -610
rect -3495 -678 -3461 -650
rect -3495 -684 -3461 -678
rect -3495 -746 -3461 -722
rect -3495 -756 -3461 -746
rect -3495 -814 -3461 -794
rect -3495 -828 -3461 -814
rect -3495 -882 -3461 -866
rect -3495 -900 -3461 -882
rect -3495 -950 -3461 -938
rect -3495 -972 -3461 -950
rect -3347 -168 -3313 -146
rect -3347 -180 -3313 -168
rect -3347 -236 -3313 -218
rect -3347 -252 -3313 -236
rect -3347 -304 -3313 -290
rect -3347 -324 -3313 -304
rect -3347 -372 -3313 -362
rect -3347 -396 -3313 -372
rect -3347 -440 -3313 -434
rect -3347 -468 -3313 -440
rect -3347 -508 -3313 -506
rect -3347 -540 -3313 -508
rect -3347 -610 -3313 -578
rect -3347 -612 -3313 -610
rect -3347 -678 -3313 -650
rect -3347 -684 -3313 -678
rect -3347 -746 -3313 -722
rect -3347 -756 -3313 -746
rect -3347 -814 -3313 -794
rect -3347 -828 -3313 -814
rect -3347 -882 -3313 -866
rect -3347 -900 -3313 -882
rect -3347 -950 -3313 -938
rect -3347 -972 -3313 -950
rect -3199 -168 -3165 -146
rect -3199 -180 -3165 -168
rect -3199 -236 -3165 -218
rect -3199 -252 -3165 -236
rect -3199 -304 -3165 -290
rect -3199 -324 -3165 -304
rect -3199 -372 -3165 -362
rect -3199 -396 -3165 -372
rect -3199 -440 -3165 -434
rect -3199 -468 -3165 -440
rect -3199 -508 -3165 -506
rect -3199 -540 -3165 -508
rect -3199 -610 -3165 -578
rect -3199 -612 -3165 -610
rect -3199 -678 -3165 -650
rect -3199 -684 -3165 -678
rect -3199 -746 -3165 -722
rect -3199 -756 -3165 -746
rect -3199 -814 -3165 -794
rect -3199 -828 -3165 -814
rect -3199 -882 -3165 -866
rect -3199 -900 -3165 -882
rect -3199 -950 -3165 -938
rect -3199 -972 -3165 -950
rect -3051 -168 -3017 -146
rect -3051 -180 -3017 -168
rect -3051 -236 -3017 -218
rect -3051 -252 -3017 -236
rect -3051 -304 -3017 -290
rect -3051 -324 -3017 -304
rect -3051 -372 -3017 -362
rect -3051 -396 -3017 -372
rect -3051 -440 -3017 -434
rect -3051 -468 -3017 -440
rect -3051 -508 -3017 -506
rect -3051 -540 -3017 -508
rect -3051 -610 -3017 -578
rect -3051 -612 -3017 -610
rect -3051 -678 -3017 -650
rect -3051 -684 -3017 -678
rect -3051 -746 -3017 -722
rect -3051 -756 -3017 -746
rect -3051 -814 -3017 -794
rect -3051 -828 -3017 -814
rect -3051 -882 -3017 -866
rect -3051 -900 -3017 -882
rect -3051 -950 -3017 -938
rect -3051 -972 -3017 -950
rect -2903 -168 -2869 -146
rect -2903 -180 -2869 -168
rect -2903 -236 -2869 -218
rect -2903 -252 -2869 -236
rect -2903 -304 -2869 -290
rect -2903 -324 -2869 -304
rect -2903 -372 -2869 -362
rect -2903 -396 -2869 -372
rect -2903 -440 -2869 -434
rect -2903 -468 -2869 -440
rect -2903 -508 -2869 -506
rect -2903 -540 -2869 -508
rect -2903 -610 -2869 -578
rect -2903 -612 -2869 -610
rect -2903 -678 -2869 -650
rect -2903 -684 -2869 -678
rect -2903 -746 -2869 -722
rect -2903 -756 -2869 -746
rect -2903 -814 -2869 -794
rect -2903 -828 -2869 -814
rect -2903 -882 -2869 -866
rect -2903 -900 -2869 -882
rect -2903 -950 -2869 -938
rect -2903 -972 -2869 -950
rect -2755 -168 -2721 -146
rect -2755 -180 -2721 -168
rect -2755 -236 -2721 -218
rect -2755 -252 -2721 -236
rect -2755 -304 -2721 -290
rect -2755 -324 -2721 -304
rect -2755 -372 -2721 -362
rect -2755 -396 -2721 -372
rect -2755 -440 -2721 -434
rect -2755 -468 -2721 -440
rect -2755 -508 -2721 -506
rect -2755 -540 -2721 -508
rect -2755 -610 -2721 -578
rect -2755 -612 -2721 -610
rect -2755 -678 -2721 -650
rect -2755 -684 -2721 -678
rect -2755 -746 -2721 -722
rect -2755 -756 -2721 -746
rect -2755 -814 -2721 -794
rect -2755 -828 -2721 -814
rect -2755 -882 -2721 -866
rect -2755 -900 -2721 -882
rect -2755 -950 -2721 -938
rect -2755 -972 -2721 -950
rect -2607 -168 -2573 -146
rect -2607 -180 -2573 -168
rect -2607 -236 -2573 -218
rect -2607 -252 -2573 -236
rect -2607 -304 -2573 -290
rect -2607 -324 -2573 -304
rect -2607 -372 -2573 -362
rect -2607 -396 -2573 -372
rect -2607 -440 -2573 -434
rect -2607 -468 -2573 -440
rect -2607 -508 -2573 -506
rect -2607 -540 -2573 -508
rect -2607 -610 -2573 -578
rect -2607 -612 -2573 -610
rect -2607 -678 -2573 -650
rect -2607 -684 -2573 -678
rect -2607 -746 -2573 -722
rect -2607 -756 -2573 -746
rect -2607 -814 -2573 -794
rect -2607 -828 -2573 -814
rect -2607 -882 -2573 -866
rect -2607 -900 -2573 -882
rect -2607 -950 -2573 -938
rect -2607 -972 -2573 -950
rect -2459 -168 -2425 -146
rect -2459 -180 -2425 -168
rect -2459 -236 -2425 -218
rect -2459 -252 -2425 -236
rect -2459 -304 -2425 -290
rect -2459 -324 -2425 -304
rect -2459 -372 -2425 -362
rect -2459 -396 -2425 -372
rect -2459 -440 -2425 -434
rect -2459 -468 -2425 -440
rect -2459 -508 -2425 -506
rect -2459 -540 -2425 -508
rect -2459 -610 -2425 -578
rect -2459 -612 -2425 -610
rect -2459 -678 -2425 -650
rect -2459 -684 -2425 -678
rect -2459 -746 -2425 -722
rect -2459 -756 -2425 -746
rect -2459 -814 -2425 -794
rect -2459 -828 -2425 -814
rect -2459 -882 -2425 -866
rect -2459 -900 -2425 -882
rect -2459 -950 -2425 -938
rect -2459 -972 -2425 -950
rect -2311 -168 -2277 -146
rect -2311 -180 -2277 -168
rect -2311 -236 -2277 -218
rect -2311 -252 -2277 -236
rect -2311 -304 -2277 -290
rect -2311 -324 -2277 -304
rect -2311 -372 -2277 -362
rect -2311 -396 -2277 -372
rect -2311 -440 -2277 -434
rect -2311 -468 -2277 -440
rect -2311 -508 -2277 -506
rect -2311 -540 -2277 -508
rect -2311 -610 -2277 -578
rect -2311 -612 -2277 -610
rect -2311 -678 -2277 -650
rect -2311 -684 -2277 -678
rect -2311 -746 -2277 -722
rect -2311 -756 -2277 -746
rect -2311 -814 -2277 -794
rect -2311 -828 -2277 -814
rect -2311 -882 -2277 -866
rect -2311 -900 -2277 -882
rect -2311 -950 -2277 -938
rect -2311 -972 -2277 -950
rect -2163 -168 -2129 -146
rect -2163 -180 -2129 -168
rect -2163 -236 -2129 -218
rect -2163 -252 -2129 -236
rect -2163 -304 -2129 -290
rect -2163 -324 -2129 -304
rect -2163 -372 -2129 -362
rect -2163 -396 -2129 -372
rect -2163 -440 -2129 -434
rect -2163 -468 -2129 -440
rect -2163 -508 -2129 -506
rect -2163 -540 -2129 -508
rect -2163 -610 -2129 -578
rect -2163 -612 -2129 -610
rect -2163 -678 -2129 -650
rect -2163 -684 -2129 -678
rect -2163 -746 -2129 -722
rect -2163 -756 -2129 -746
rect -2163 -814 -2129 -794
rect -2163 -828 -2129 -814
rect -2163 -882 -2129 -866
rect -2163 -900 -2129 -882
rect -2163 -950 -2129 -938
rect -2163 -972 -2129 -950
rect -2015 -168 -1981 -146
rect -2015 -180 -1981 -168
rect -2015 -236 -1981 -218
rect -2015 -252 -1981 -236
rect -2015 -304 -1981 -290
rect -2015 -324 -1981 -304
rect -2015 -372 -1981 -362
rect -2015 -396 -1981 -372
rect -2015 -440 -1981 -434
rect -2015 -468 -1981 -440
rect -2015 -508 -1981 -506
rect -2015 -540 -1981 -508
rect -2015 -610 -1981 -578
rect -2015 -612 -1981 -610
rect -2015 -678 -1981 -650
rect -2015 -684 -1981 -678
rect -2015 -746 -1981 -722
rect -2015 -756 -1981 -746
rect -2015 -814 -1981 -794
rect -2015 -828 -1981 -814
rect -2015 -882 -1981 -866
rect -2015 -900 -1981 -882
rect -2015 -950 -1981 -938
rect -2015 -972 -1981 -950
rect -1867 -168 -1833 -146
rect -1867 -180 -1833 -168
rect -1867 -236 -1833 -218
rect -1867 -252 -1833 -236
rect -1867 -304 -1833 -290
rect -1867 -324 -1833 -304
rect -1867 -372 -1833 -362
rect -1867 -396 -1833 -372
rect -1867 -440 -1833 -434
rect -1867 -468 -1833 -440
rect -1867 -508 -1833 -506
rect -1867 -540 -1833 -508
rect -1867 -610 -1833 -578
rect -1867 -612 -1833 -610
rect -1867 -678 -1833 -650
rect -1867 -684 -1833 -678
rect -1867 -746 -1833 -722
rect -1867 -756 -1833 -746
rect -1867 -814 -1833 -794
rect -1867 -828 -1833 -814
rect -1867 -882 -1833 -866
rect -1867 -900 -1833 -882
rect -1867 -950 -1833 -938
rect -1867 -972 -1833 -950
rect -1719 -168 -1685 -146
rect -1719 -180 -1685 -168
rect -1719 -236 -1685 -218
rect -1719 -252 -1685 -236
rect -1719 -304 -1685 -290
rect -1719 -324 -1685 -304
rect -1719 -372 -1685 -362
rect -1719 -396 -1685 -372
rect -1719 -440 -1685 -434
rect -1719 -468 -1685 -440
rect -1719 -508 -1685 -506
rect -1719 -540 -1685 -508
rect -1719 -610 -1685 -578
rect -1719 -612 -1685 -610
rect -1719 -678 -1685 -650
rect -1719 -684 -1685 -678
rect -1719 -746 -1685 -722
rect -1719 -756 -1685 -746
rect -1719 -814 -1685 -794
rect -1719 -828 -1685 -814
rect -1719 -882 -1685 -866
rect -1719 -900 -1685 -882
rect -1719 -950 -1685 -938
rect -1719 -972 -1685 -950
rect -1571 -168 -1537 -146
rect -1571 -180 -1537 -168
rect -1571 -236 -1537 -218
rect -1571 -252 -1537 -236
rect -1571 -304 -1537 -290
rect -1571 -324 -1537 -304
rect -1571 -372 -1537 -362
rect -1571 -396 -1537 -372
rect -1571 -440 -1537 -434
rect -1571 -468 -1537 -440
rect -1571 -508 -1537 -506
rect -1571 -540 -1537 -508
rect -1571 -610 -1537 -578
rect -1571 -612 -1537 -610
rect -1571 -678 -1537 -650
rect -1571 -684 -1537 -678
rect -1571 -746 -1537 -722
rect -1571 -756 -1537 -746
rect -1571 -814 -1537 -794
rect -1571 -828 -1537 -814
rect -1571 -882 -1537 -866
rect -1571 -900 -1537 -882
rect -1571 -950 -1537 -938
rect -1571 -972 -1537 -950
rect -1423 -168 -1389 -146
rect -1423 -180 -1389 -168
rect -1423 -236 -1389 -218
rect -1423 -252 -1389 -236
rect -1423 -304 -1389 -290
rect -1423 -324 -1389 -304
rect -1423 -372 -1389 -362
rect -1423 -396 -1389 -372
rect -1423 -440 -1389 -434
rect -1423 -468 -1389 -440
rect -1423 -508 -1389 -506
rect -1423 -540 -1389 -508
rect -1423 -610 -1389 -578
rect -1423 -612 -1389 -610
rect -1423 -678 -1389 -650
rect -1423 -684 -1389 -678
rect -1423 -746 -1389 -722
rect -1423 -756 -1389 -746
rect -1423 -814 -1389 -794
rect -1423 -828 -1389 -814
rect -1423 -882 -1389 -866
rect -1423 -900 -1389 -882
rect -1423 -950 -1389 -938
rect -1423 -972 -1389 -950
rect -1275 -168 -1241 -146
rect -1275 -180 -1241 -168
rect -1275 -236 -1241 -218
rect -1275 -252 -1241 -236
rect -1275 -304 -1241 -290
rect -1275 -324 -1241 -304
rect -1275 -372 -1241 -362
rect -1275 -396 -1241 -372
rect -1275 -440 -1241 -434
rect -1275 -468 -1241 -440
rect -1275 -508 -1241 -506
rect -1275 -540 -1241 -508
rect -1275 -610 -1241 -578
rect -1275 -612 -1241 -610
rect -1275 -678 -1241 -650
rect -1275 -684 -1241 -678
rect -1275 -746 -1241 -722
rect -1275 -756 -1241 -746
rect -1275 -814 -1241 -794
rect -1275 -828 -1241 -814
rect -1275 -882 -1241 -866
rect -1275 -900 -1241 -882
rect -1275 -950 -1241 -938
rect -1275 -972 -1241 -950
rect -1127 -168 -1093 -146
rect -1127 -180 -1093 -168
rect -1127 -236 -1093 -218
rect -1127 -252 -1093 -236
rect -1127 -304 -1093 -290
rect -1127 -324 -1093 -304
rect -1127 -372 -1093 -362
rect -1127 -396 -1093 -372
rect -1127 -440 -1093 -434
rect -1127 -468 -1093 -440
rect -1127 -508 -1093 -506
rect -1127 -540 -1093 -508
rect -1127 -610 -1093 -578
rect -1127 -612 -1093 -610
rect -1127 -678 -1093 -650
rect -1127 -684 -1093 -678
rect -1127 -746 -1093 -722
rect -1127 -756 -1093 -746
rect -1127 -814 -1093 -794
rect -1127 -828 -1093 -814
rect -1127 -882 -1093 -866
rect -1127 -900 -1093 -882
rect -1127 -950 -1093 -938
rect -1127 -972 -1093 -950
rect -979 -168 -945 -146
rect -979 -180 -945 -168
rect -979 -236 -945 -218
rect -979 -252 -945 -236
rect -979 -304 -945 -290
rect -979 -324 -945 -304
rect -979 -372 -945 -362
rect -979 -396 -945 -372
rect -979 -440 -945 -434
rect -979 -468 -945 -440
rect -979 -508 -945 -506
rect -979 -540 -945 -508
rect -979 -610 -945 -578
rect -979 -612 -945 -610
rect -979 -678 -945 -650
rect -979 -684 -945 -678
rect -979 -746 -945 -722
rect -979 -756 -945 -746
rect -979 -814 -945 -794
rect -979 -828 -945 -814
rect -979 -882 -945 -866
rect -979 -900 -945 -882
rect -979 -950 -945 -938
rect -979 -972 -945 -950
rect -831 -168 -797 -146
rect -831 -180 -797 -168
rect -831 -236 -797 -218
rect -831 -252 -797 -236
rect -831 -304 -797 -290
rect -831 -324 -797 -304
rect -831 -372 -797 -362
rect -831 -396 -797 -372
rect -831 -440 -797 -434
rect -831 -468 -797 -440
rect -831 -508 -797 -506
rect -831 -540 -797 -508
rect -831 -610 -797 -578
rect -831 -612 -797 -610
rect -831 -678 -797 -650
rect -831 -684 -797 -678
rect -831 -746 -797 -722
rect -831 -756 -797 -746
rect -831 -814 -797 -794
rect -831 -828 -797 -814
rect -831 -882 -797 -866
rect -831 -900 -797 -882
rect -831 -950 -797 -938
rect -831 -972 -797 -950
rect -683 -168 -649 -146
rect -683 -180 -649 -168
rect -683 -236 -649 -218
rect -683 -252 -649 -236
rect -683 -304 -649 -290
rect -683 -324 -649 -304
rect -683 -372 -649 -362
rect -683 -396 -649 -372
rect -683 -440 -649 -434
rect -683 -468 -649 -440
rect -683 -508 -649 -506
rect -683 -540 -649 -508
rect -683 -610 -649 -578
rect -683 -612 -649 -610
rect -683 -678 -649 -650
rect -683 -684 -649 -678
rect -683 -746 -649 -722
rect -683 -756 -649 -746
rect -683 -814 -649 -794
rect -683 -828 -649 -814
rect -683 -882 -649 -866
rect -683 -900 -649 -882
rect -683 -950 -649 -938
rect -683 -972 -649 -950
rect -535 -168 -501 -146
rect -535 -180 -501 -168
rect -535 -236 -501 -218
rect -535 -252 -501 -236
rect -535 -304 -501 -290
rect -535 -324 -501 -304
rect -535 -372 -501 -362
rect -535 -396 -501 -372
rect -535 -440 -501 -434
rect -535 -468 -501 -440
rect -535 -508 -501 -506
rect -535 -540 -501 -508
rect -535 -610 -501 -578
rect -535 -612 -501 -610
rect -535 -678 -501 -650
rect -535 -684 -501 -678
rect -535 -746 -501 -722
rect -535 -756 -501 -746
rect -535 -814 -501 -794
rect -535 -828 -501 -814
rect -535 -882 -501 -866
rect -535 -900 -501 -882
rect -535 -950 -501 -938
rect -535 -972 -501 -950
rect -387 -168 -353 -146
rect -387 -180 -353 -168
rect -387 -236 -353 -218
rect -387 -252 -353 -236
rect -387 -304 -353 -290
rect -387 -324 -353 -304
rect -387 -372 -353 -362
rect -387 -396 -353 -372
rect -387 -440 -353 -434
rect -387 -468 -353 -440
rect -387 -508 -353 -506
rect -387 -540 -353 -508
rect -387 -610 -353 -578
rect -387 -612 -353 -610
rect -387 -678 -353 -650
rect -387 -684 -353 -678
rect -387 -746 -353 -722
rect -387 -756 -353 -746
rect -387 -814 -353 -794
rect -387 -828 -353 -814
rect -387 -882 -353 -866
rect -387 -900 -353 -882
rect -387 -950 -353 -938
rect -387 -972 -353 -950
rect -239 -168 -205 -146
rect -239 -180 -205 -168
rect -239 -236 -205 -218
rect -239 -252 -205 -236
rect -239 -304 -205 -290
rect -239 -324 -205 -304
rect -239 -372 -205 -362
rect -239 -396 -205 -372
rect -239 -440 -205 -434
rect -239 -468 -205 -440
rect -239 -508 -205 -506
rect -239 -540 -205 -508
rect -239 -610 -205 -578
rect -239 -612 -205 -610
rect -239 -678 -205 -650
rect -239 -684 -205 -678
rect -239 -746 -205 -722
rect -239 -756 -205 -746
rect -239 -814 -205 -794
rect -239 -828 -205 -814
rect -239 -882 -205 -866
rect -239 -900 -205 -882
rect -239 -950 -205 -938
rect -239 -972 -205 -950
rect -91 -168 -57 -146
rect -91 -180 -57 -168
rect -91 -236 -57 -218
rect -91 -252 -57 -236
rect -91 -304 -57 -290
rect -91 -324 -57 -304
rect -91 -372 -57 -362
rect -91 -396 -57 -372
rect -91 -440 -57 -434
rect -91 -468 -57 -440
rect -91 -508 -57 -506
rect -91 -540 -57 -508
rect -91 -610 -57 -578
rect -91 -612 -57 -610
rect -91 -678 -57 -650
rect -91 -684 -57 -678
rect -91 -746 -57 -722
rect -91 -756 -57 -746
rect -91 -814 -57 -794
rect -91 -828 -57 -814
rect -91 -882 -57 -866
rect -91 -900 -57 -882
rect -91 -950 -57 -938
rect -91 -972 -57 -950
rect 57 -168 91 -146
rect 57 -180 91 -168
rect 57 -236 91 -218
rect 57 -252 91 -236
rect 57 -304 91 -290
rect 57 -324 91 -304
rect 57 -372 91 -362
rect 57 -396 91 -372
rect 57 -440 91 -434
rect 57 -468 91 -440
rect 57 -508 91 -506
rect 57 -540 91 -508
rect 57 -610 91 -578
rect 57 -612 91 -610
rect 57 -678 91 -650
rect 57 -684 91 -678
rect 57 -746 91 -722
rect 57 -756 91 -746
rect 57 -814 91 -794
rect 57 -828 91 -814
rect 57 -882 91 -866
rect 57 -900 91 -882
rect 57 -950 91 -938
rect 57 -972 91 -950
rect 205 -168 239 -146
rect 205 -180 239 -168
rect 205 -236 239 -218
rect 205 -252 239 -236
rect 205 -304 239 -290
rect 205 -324 239 -304
rect 205 -372 239 -362
rect 205 -396 239 -372
rect 205 -440 239 -434
rect 205 -468 239 -440
rect 205 -508 239 -506
rect 205 -540 239 -508
rect 205 -610 239 -578
rect 205 -612 239 -610
rect 205 -678 239 -650
rect 205 -684 239 -678
rect 205 -746 239 -722
rect 205 -756 239 -746
rect 205 -814 239 -794
rect 205 -828 239 -814
rect 205 -882 239 -866
rect 205 -900 239 -882
rect 205 -950 239 -938
rect 205 -972 239 -950
rect 353 -168 387 -146
rect 353 -180 387 -168
rect 353 -236 387 -218
rect 353 -252 387 -236
rect 353 -304 387 -290
rect 353 -324 387 -304
rect 353 -372 387 -362
rect 353 -396 387 -372
rect 353 -440 387 -434
rect 353 -468 387 -440
rect 353 -508 387 -506
rect 353 -540 387 -508
rect 353 -610 387 -578
rect 353 -612 387 -610
rect 353 -678 387 -650
rect 353 -684 387 -678
rect 353 -746 387 -722
rect 353 -756 387 -746
rect 353 -814 387 -794
rect 353 -828 387 -814
rect 353 -882 387 -866
rect 353 -900 387 -882
rect 353 -950 387 -938
rect 353 -972 387 -950
rect 501 -168 535 -146
rect 501 -180 535 -168
rect 501 -236 535 -218
rect 501 -252 535 -236
rect 501 -304 535 -290
rect 501 -324 535 -304
rect 501 -372 535 -362
rect 501 -396 535 -372
rect 501 -440 535 -434
rect 501 -468 535 -440
rect 501 -508 535 -506
rect 501 -540 535 -508
rect 501 -610 535 -578
rect 501 -612 535 -610
rect 501 -678 535 -650
rect 501 -684 535 -678
rect 501 -746 535 -722
rect 501 -756 535 -746
rect 501 -814 535 -794
rect 501 -828 535 -814
rect 501 -882 535 -866
rect 501 -900 535 -882
rect 501 -950 535 -938
rect 501 -972 535 -950
rect 649 -168 683 -146
rect 649 -180 683 -168
rect 649 -236 683 -218
rect 649 -252 683 -236
rect 649 -304 683 -290
rect 649 -324 683 -304
rect 649 -372 683 -362
rect 649 -396 683 -372
rect 649 -440 683 -434
rect 649 -468 683 -440
rect 649 -508 683 -506
rect 649 -540 683 -508
rect 649 -610 683 -578
rect 649 -612 683 -610
rect 649 -678 683 -650
rect 649 -684 683 -678
rect 649 -746 683 -722
rect 649 -756 683 -746
rect 649 -814 683 -794
rect 649 -828 683 -814
rect 649 -882 683 -866
rect 649 -900 683 -882
rect 649 -950 683 -938
rect 649 -972 683 -950
rect 797 -168 831 -146
rect 797 -180 831 -168
rect 797 -236 831 -218
rect 797 -252 831 -236
rect 797 -304 831 -290
rect 797 -324 831 -304
rect 797 -372 831 -362
rect 797 -396 831 -372
rect 797 -440 831 -434
rect 797 -468 831 -440
rect 797 -508 831 -506
rect 797 -540 831 -508
rect 797 -610 831 -578
rect 797 -612 831 -610
rect 797 -678 831 -650
rect 797 -684 831 -678
rect 797 -746 831 -722
rect 797 -756 831 -746
rect 797 -814 831 -794
rect 797 -828 831 -814
rect 797 -882 831 -866
rect 797 -900 831 -882
rect 797 -950 831 -938
rect 797 -972 831 -950
rect 945 -168 979 -146
rect 945 -180 979 -168
rect 945 -236 979 -218
rect 945 -252 979 -236
rect 945 -304 979 -290
rect 945 -324 979 -304
rect 945 -372 979 -362
rect 945 -396 979 -372
rect 945 -440 979 -434
rect 945 -468 979 -440
rect 945 -508 979 -506
rect 945 -540 979 -508
rect 945 -610 979 -578
rect 945 -612 979 -610
rect 945 -678 979 -650
rect 945 -684 979 -678
rect 945 -746 979 -722
rect 945 -756 979 -746
rect 945 -814 979 -794
rect 945 -828 979 -814
rect 945 -882 979 -866
rect 945 -900 979 -882
rect 945 -950 979 -938
rect 945 -972 979 -950
rect 1093 -168 1127 -146
rect 1093 -180 1127 -168
rect 1093 -236 1127 -218
rect 1093 -252 1127 -236
rect 1093 -304 1127 -290
rect 1093 -324 1127 -304
rect 1093 -372 1127 -362
rect 1093 -396 1127 -372
rect 1093 -440 1127 -434
rect 1093 -468 1127 -440
rect 1093 -508 1127 -506
rect 1093 -540 1127 -508
rect 1093 -610 1127 -578
rect 1093 -612 1127 -610
rect 1093 -678 1127 -650
rect 1093 -684 1127 -678
rect 1093 -746 1127 -722
rect 1093 -756 1127 -746
rect 1093 -814 1127 -794
rect 1093 -828 1127 -814
rect 1093 -882 1127 -866
rect 1093 -900 1127 -882
rect 1093 -950 1127 -938
rect 1093 -972 1127 -950
rect 1241 -168 1275 -146
rect 1241 -180 1275 -168
rect 1241 -236 1275 -218
rect 1241 -252 1275 -236
rect 1241 -304 1275 -290
rect 1241 -324 1275 -304
rect 1241 -372 1275 -362
rect 1241 -396 1275 -372
rect 1241 -440 1275 -434
rect 1241 -468 1275 -440
rect 1241 -508 1275 -506
rect 1241 -540 1275 -508
rect 1241 -610 1275 -578
rect 1241 -612 1275 -610
rect 1241 -678 1275 -650
rect 1241 -684 1275 -678
rect 1241 -746 1275 -722
rect 1241 -756 1275 -746
rect 1241 -814 1275 -794
rect 1241 -828 1275 -814
rect 1241 -882 1275 -866
rect 1241 -900 1275 -882
rect 1241 -950 1275 -938
rect 1241 -972 1275 -950
rect 1389 -168 1423 -146
rect 1389 -180 1423 -168
rect 1389 -236 1423 -218
rect 1389 -252 1423 -236
rect 1389 -304 1423 -290
rect 1389 -324 1423 -304
rect 1389 -372 1423 -362
rect 1389 -396 1423 -372
rect 1389 -440 1423 -434
rect 1389 -468 1423 -440
rect 1389 -508 1423 -506
rect 1389 -540 1423 -508
rect 1389 -610 1423 -578
rect 1389 -612 1423 -610
rect 1389 -678 1423 -650
rect 1389 -684 1423 -678
rect 1389 -746 1423 -722
rect 1389 -756 1423 -746
rect 1389 -814 1423 -794
rect 1389 -828 1423 -814
rect 1389 -882 1423 -866
rect 1389 -900 1423 -882
rect 1389 -950 1423 -938
rect 1389 -972 1423 -950
rect 1537 -168 1571 -146
rect 1537 -180 1571 -168
rect 1537 -236 1571 -218
rect 1537 -252 1571 -236
rect 1537 -304 1571 -290
rect 1537 -324 1571 -304
rect 1537 -372 1571 -362
rect 1537 -396 1571 -372
rect 1537 -440 1571 -434
rect 1537 -468 1571 -440
rect 1537 -508 1571 -506
rect 1537 -540 1571 -508
rect 1537 -610 1571 -578
rect 1537 -612 1571 -610
rect 1537 -678 1571 -650
rect 1537 -684 1571 -678
rect 1537 -746 1571 -722
rect 1537 -756 1571 -746
rect 1537 -814 1571 -794
rect 1537 -828 1571 -814
rect 1537 -882 1571 -866
rect 1537 -900 1571 -882
rect 1537 -950 1571 -938
rect 1537 -972 1571 -950
rect 1685 -168 1719 -146
rect 1685 -180 1719 -168
rect 1685 -236 1719 -218
rect 1685 -252 1719 -236
rect 1685 -304 1719 -290
rect 1685 -324 1719 -304
rect 1685 -372 1719 -362
rect 1685 -396 1719 -372
rect 1685 -440 1719 -434
rect 1685 -468 1719 -440
rect 1685 -508 1719 -506
rect 1685 -540 1719 -508
rect 1685 -610 1719 -578
rect 1685 -612 1719 -610
rect 1685 -678 1719 -650
rect 1685 -684 1719 -678
rect 1685 -746 1719 -722
rect 1685 -756 1719 -746
rect 1685 -814 1719 -794
rect 1685 -828 1719 -814
rect 1685 -882 1719 -866
rect 1685 -900 1719 -882
rect 1685 -950 1719 -938
rect 1685 -972 1719 -950
rect 1833 -168 1867 -146
rect 1833 -180 1867 -168
rect 1833 -236 1867 -218
rect 1833 -252 1867 -236
rect 1833 -304 1867 -290
rect 1833 -324 1867 -304
rect 1833 -372 1867 -362
rect 1833 -396 1867 -372
rect 1833 -440 1867 -434
rect 1833 -468 1867 -440
rect 1833 -508 1867 -506
rect 1833 -540 1867 -508
rect 1833 -610 1867 -578
rect 1833 -612 1867 -610
rect 1833 -678 1867 -650
rect 1833 -684 1867 -678
rect 1833 -746 1867 -722
rect 1833 -756 1867 -746
rect 1833 -814 1867 -794
rect 1833 -828 1867 -814
rect 1833 -882 1867 -866
rect 1833 -900 1867 -882
rect 1833 -950 1867 -938
rect 1833 -972 1867 -950
rect 1981 -168 2015 -146
rect 1981 -180 2015 -168
rect 1981 -236 2015 -218
rect 1981 -252 2015 -236
rect 1981 -304 2015 -290
rect 1981 -324 2015 -304
rect 1981 -372 2015 -362
rect 1981 -396 2015 -372
rect 1981 -440 2015 -434
rect 1981 -468 2015 -440
rect 1981 -508 2015 -506
rect 1981 -540 2015 -508
rect 1981 -610 2015 -578
rect 1981 -612 2015 -610
rect 1981 -678 2015 -650
rect 1981 -684 2015 -678
rect 1981 -746 2015 -722
rect 1981 -756 2015 -746
rect 1981 -814 2015 -794
rect 1981 -828 2015 -814
rect 1981 -882 2015 -866
rect 1981 -900 2015 -882
rect 1981 -950 2015 -938
rect 1981 -972 2015 -950
rect 2129 -168 2163 -146
rect 2129 -180 2163 -168
rect 2129 -236 2163 -218
rect 2129 -252 2163 -236
rect 2129 -304 2163 -290
rect 2129 -324 2163 -304
rect 2129 -372 2163 -362
rect 2129 -396 2163 -372
rect 2129 -440 2163 -434
rect 2129 -468 2163 -440
rect 2129 -508 2163 -506
rect 2129 -540 2163 -508
rect 2129 -610 2163 -578
rect 2129 -612 2163 -610
rect 2129 -678 2163 -650
rect 2129 -684 2163 -678
rect 2129 -746 2163 -722
rect 2129 -756 2163 -746
rect 2129 -814 2163 -794
rect 2129 -828 2163 -814
rect 2129 -882 2163 -866
rect 2129 -900 2163 -882
rect 2129 -950 2163 -938
rect 2129 -972 2163 -950
rect 2277 -168 2311 -146
rect 2277 -180 2311 -168
rect 2277 -236 2311 -218
rect 2277 -252 2311 -236
rect 2277 -304 2311 -290
rect 2277 -324 2311 -304
rect 2277 -372 2311 -362
rect 2277 -396 2311 -372
rect 2277 -440 2311 -434
rect 2277 -468 2311 -440
rect 2277 -508 2311 -506
rect 2277 -540 2311 -508
rect 2277 -610 2311 -578
rect 2277 -612 2311 -610
rect 2277 -678 2311 -650
rect 2277 -684 2311 -678
rect 2277 -746 2311 -722
rect 2277 -756 2311 -746
rect 2277 -814 2311 -794
rect 2277 -828 2311 -814
rect 2277 -882 2311 -866
rect 2277 -900 2311 -882
rect 2277 -950 2311 -938
rect 2277 -972 2311 -950
rect 2425 -168 2459 -146
rect 2425 -180 2459 -168
rect 2425 -236 2459 -218
rect 2425 -252 2459 -236
rect 2425 -304 2459 -290
rect 2425 -324 2459 -304
rect 2425 -372 2459 -362
rect 2425 -396 2459 -372
rect 2425 -440 2459 -434
rect 2425 -468 2459 -440
rect 2425 -508 2459 -506
rect 2425 -540 2459 -508
rect 2425 -610 2459 -578
rect 2425 -612 2459 -610
rect 2425 -678 2459 -650
rect 2425 -684 2459 -678
rect 2425 -746 2459 -722
rect 2425 -756 2459 -746
rect 2425 -814 2459 -794
rect 2425 -828 2459 -814
rect 2425 -882 2459 -866
rect 2425 -900 2459 -882
rect 2425 -950 2459 -938
rect 2425 -972 2459 -950
rect 2573 -168 2607 -146
rect 2573 -180 2607 -168
rect 2573 -236 2607 -218
rect 2573 -252 2607 -236
rect 2573 -304 2607 -290
rect 2573 -324 2607 -304
rect 2573 -372 2607 -362
rect 2573 -396 2607 -372
rect 2573 -440 2607 -434
rect 2573 -468 2607 -440
rect 2573 -508 2607 -506
rect 2573 -540 2607 -508
rect 2573 -610 2607 -578
rect 2573 -612 2607 -610
rect 2573 -678 2607 -650
rect 2573 -684 2607 -678
rect 2573 -746 2607 -722
rect 2573 -756 2607 -746
rect 2573 -814 2607 -794
rect 2573 -828 2607 -814
rect 2573 -882 2607 -866
rect 2573 -900 2607 -882
rect 2573 -950 2607 -938
rect 2573 -972 2607 -950
rect 2721 -168 2755 -146
rect 2721 -180 2755 -168
rect 2721 -236 2755 -218
rect 2721 -252 2755 -236
rect 2721 -304 2755 -290
rect 2721 -324 2755 -304
rect 2721 -372 2755 -362
rect 2721 -396 2755 -372
rect 2721 -440 2755 -434
rect 2721 -468 2755 -440
rect 2721 -508 2755 -506
rect 2721 -540 2755 -508
rect 2721 -610 2755 -578
rect 2721 -612 2755 -610
rect 2721 -678 2755 -650
rect 2721 -684 2755 -678
rect 2721 -746 2755 -722
rect 2721 -756 2755 -746
rect 2721 -814 2755 -794
rect 2721 -828 2755 -814
rect 2721 -882 2755 -866
rect 2721 -900 2755 -882
rect 2721 -950 2755 -938
rect 2721 -972 2755 -950
rect 2869 -168 2903 -146
rect 2869 -180 2903 -168
rect 2869 -236 2903 -218
rect 2869 -252 2903 -236
rect 2869 -304 2903 -290
rect 2869 -324 2903 -304
rect 2869 -372 2903 -362
rect 2869 -396 2903 -372
rect 2869 -440 2903 -434
rect 2869 -468 2903 -440
rect 2869 -508 2903 -506
rect 2869 -540 2903 -508
rect 2869 -610 2903 -578
rect 2869 -612 2903 -610
rect 2869 -678 2903 -650
rect 2869 -684 2903 -678
rect 2869 -746 2903 -722
rect 2869 -756 2903 -746
rect 2869 -814 2903 -794
rect 2869 -828 2903 -814
rect 2869 -882 2903 -866
rect 2869 -900 2903 -882
rect 2869 -950 2903 -938
rect 2869 -972 2903 -950
rect 3017 -168 3051 -146
rect 3017 -180 3051 -168
rect 3017 -236 3051 -218
rect 3017 -252 3051 -236
rect 3017 -304 3051 -290
rect 3017 -324 3051 -304
rect 3017 -372 3051 -362
rect 3017 -396 3051 -372
rect 3017 -440 3051 -434
rect 3017 -468 3051 -440
rect 3017 -508 3051 -506
rect 3017 -540 3051 -508
rect 3017 -610 3051 -578
rect 3017 -612 3051 -610
rect 3017 -678 3051 -650
rect 3017 -684 3051 -678
rect 3017 -746 3051 -722
rect 3017 -756 3051 -746
rect 3017 -814 3051 -794
rect 3017 -828 3051 -814
rect 3017 -882 3051 -866
rect 3017 -900 3051 -882
rect 3017 -950 3051 -938
rect 3017 -972 3051 -950
rect 3165 -168 3199 -146
rect 3165 -180 3199 -168
rect 3165 -236 3199 -218
rect 3165 -252 3199 -236
rect 3165 -304 3199 -290
rect 3165 -324 3199 -304
rect 3165 -372 3199 -362
rect 3165 -396 3199 -372
rect 3165 -440 3199 -434
rect 3165 -468 3199 -440
rect 3165 -508 3199 -506
rect 3165 -540 3199 -508
rect 3165 -610 3199 -578
rect 3165 -612 3199 -610
rect 3165 -678 3199 -650
rect 3165 -684 3199 -678
rect 3165 -746 3199 -722
rect 3165 -756 3199 -746
rect 3165 -814 3199 -794
rect 3165 -828 3199 -814
rect 3165 -882 3199 -866
rect 3165 -900 3199 -882
rect 3165 -950 3199 -938
rect 3165 -972 3199 -950
rect 3313 -168 3347 -146
rect 3313 -180 3347 -168
rect 3313 -236 3347 -218
rect 3313 -252 3347 -236
rect 3313 -304 3347 -290
rect 3313 -324 3347 -304
rect 3313 -372 3347 -362
rect 3313 -396 3347 -372
rect 3313 -440 3347 -434
rect 3313 -468 3347 -440
rect 3313 -508 3347 -506
rect 3313 -540 3347 -508
rect 3313 -610 3347 -578
rect 3313 -612 3347 -610
rect 3313 -678 3347 -650
rect 3313 -684 3347 -678
rect 3313 -746 3347 -722
rect 3313 -756 3347 -746
rect 3313 -814 3347 -794
rect 3313 -828 3347 -814
rect 3313 -882 3347 -866
rect 3313 -900 3347 -882
rect 3313 -950 3347 -938
rect 3313 -972 3347 -950
rect 3461 -168 3495 -146
rect 3461 -180 3495 -168
rect 3461 -236 3495 -218
rect 3461 -252 3495 -236
rect 3461 -304 3495 -290
rect 3461 -324 3495 -304
rect 3461 -372 3495 -362
rect 3461 -396 3495 -372
rect 3461 -440 3495 -434
rect 3461 -468 3495 -440
rect 3461 -508 3495 -506
rect 3461 -540 3495 -508
rect 3461 -610 3495 -578
rect 3461 -612 3495 -610
rect 3461 -678 3495 -650
rect 3461 -684 3495 -678
rect 3461 -746 3495 -722
rect 3461 -756 3495 -746
rect 3461 -814 3495 -794
rect 3461 -828 3495 -814
rect 3461 -882 3495 -866
rect 3461 -900 3495 -882
rect 3461 -950 3495 -938
rect 3461 -972 3495 -950
rect 3609 -168 3643 -146
rect 3609 -180 3643 -168
rect 3609 -236 3643 -218
rect 3609 -252 3643 -236
rect 3609 -304 3643 -290
rect 3609 -324 3643 -304
rect 3609 -372 3643 -362
rect 3609 -396 3643 -372
rect 3609 -440 3643 -434
rect 3609 -468 3643 -440
rect 3609 -508 3643 -506
rect 3609 -540 3643 -508
rect 3609 -610 3643 -578
rect 3609 -612 3643 -610
rect 3609 -678 3643 -650
rect 3609 -684 3643 -678
rect 3609 -746 3643 -722
rect 3609 -756 3643 -746
rect 3609 -814 3643 -794
rect 3609 -828 3643 -814
rect 3609 -882 3643 -866
rect 3609 -900 3643 -882
rect 3609 -950 3643 -938
rect 3609 -972 3643 -950
rect 3757 -168 3791 -146
rect 3757 -180 3791 -168
rect 3757 -236 3791 -218
rect 3757 -252 3791 -236
rect 3757 -304 3791 -290
rect 3757 -324 3791 -304
rect 3757 -372 3791 -362
rect 3757 -396 3791 -372
rect 3757 -440 3791 -434
rect 3757 -468 3791 -440
rect 3757 -508 3791 -506
rect 3757 -540 3791 -508
rect 3757 -610 3791 -578
rect 3757 -612 3791 -610
rect 3757 -678 3791 -650
rect 3757 -684 3791 -678
rect 3757 -746 3791 -722
rect 3757 -756 3791 -746
rect 3757 -814 3791 -794
rect 3757 -828 3791 -814
rect 3757 -882 3791 -866
rect 3757 -900 3791 -882
rect 3757 -950 3791 -938
rect 3757 -972 3791 -950
rect 3905 -168 3939 -146
rect 3905 -180 3939 -168
rect 3905 -236 3939 -218
rect 3905 -252 3939 -236
rect 3905 -304 3939 -290
rect 3905 -324 3939 -304
rect 3905 -372 3939 -362
rect 3905 -396 3939 -372
rect 3905 -440 3939 -434
rect 3905 -468 3939 -440
rect 3905 -508 3939 -506
rect 3905 -540 3939 -508
rect 3905 -610 3939 -578
rect 3905 -612 3939 -610
rect 3905 -678 3939 -650
rect 3905 -684 3939 -678
rect 3905 -746 3939 -722
rect 3905 -756 3939 -746
rect 3905 -814 3939 -794
rect 3905 -828 3939 -814
rect 3905 -882 3939 -866
rect 3905 -900 3939 -882
rect 3905 -950 3939 -938
rect 3905 -972 3939 -950
rect 4053 -168 4087 -146
rect 4053 -180 4087 -168
rect 4053 -236 4087 -218
rect 4053 -252 4087 -236
rect 4053 -304 4087 -290
rect 4053 -324 4087 -304
rect 4053 -372 4087 -362
rect 4053 -396 4087 -372
rect 4053 -440 4087 -434
rect 4053 -468 4087 -440
rect 4053 -508 4087 -506
rect 4053 -540 4087 -508
rect 4053 -610 4087 -578
rect 4053 -612 4087 -610
rect 4053 -678 4087 -650
rect 4053 -684 4087 -678
rect 4053 -746 4087 -722
rect 4053 -756 4087 -746
rect 4053 -814 4087 -794
rect 4053 -828 4087 -814
rect 4053 -882 4087 -866
rect 4053 -900 4087 -882
rect 4053 -950 4087 -938
rect 4053 -972 4087 -950
rect 4201 -168 4235 -146
rect 4201 -180 4235 -168
rect 4201 -236 4235 -218
rect 4201 -252 4235 -236
rect 4201 -304 4235 -290
rect 4201 -324 4235 -304
rect 4201 -372 4235 -362
rect 4201 -396 4235 -372
rect 4201 -440 4235 -434
rect 4201 -468 4235 -440
rect 4201 -508 4235 -506
rect 4201 -540 4235 -508
rect 4201 -610 4235 -578
rect 4201 -612 4235 -610
rect 4201 -678 4235 -650
rect 4201 -684 4235 -678
rect 4201 -746 4235 -722
rect 4201 -756 4235 -746
rect 4201 -814 4235 -794
rect 4201 -828 4235 -814
rect 4201 -882 4235 -866
rect 4201 -900 4235 -882
rect 4201 -950 4235 -938
rect 4201 -972 4235 -950
rect 4349 -168 4383 -146
rect 4349 -180 4383 -168
rect 4349 -236 4383 -218
rect 4349 -252 4383 -236
rect 4349 -304 4383 -290
rect 4349 -324 4383 -304
rect 4349 -372 4383 -362
rect 4349 -396 4383 -372
rect 4349 -440 4383 -434
rect 4349 -468 4383 -440
rect 4349 -508 4383 -506
rect 4349 -540 4383 -508
rect 4349 -610 4383 -578
rect 4349 -612 4383 -610
rect 4349 -678 4383 -650
rect 4349 -684 4383 -678
rect 4349 -746 4383 -722
rect 4349 -756 4383 -746
rect 4349 -814 4383 -794
rect 4349 -828 4383 -814
rect 4349 -882 4383 -866
rect 4349 -900 4383 -882
rect 4349 -950 4383 -938
rect 4349 -972 4383 -950
rect 4497 -168 4531 -146
rect 4497 -180 4531 -168
rect 4497 -236 4531 -218
rect 4497 -252 4531 -236
rect 4497 -304 4531 -290
rect 4497 -324 4531 -304
rect 4497 -372 4531 -362
rect 4497 -396 4531 -372
rect 4497 -440 4531 -434
rect 4497 -468 4531 -440
rect 4497 -508 4531 -506
rect 4497 -540 4531 -508
rect 4497 -610 4531 -578
rect 4497 -612 4531 -610
rect 4497 -678 4531 -650
rect 4497 -684 4531 -678
rect 4497 -746 4531 -722
rect 4497 -756 4531 -746
rect 4497 -814 4531 -794
rect 4497 -828 4531 -814
rect 4497 -882 4531 -866
rect 4497 -900 4531 -882
rect 4497 -950 4531 -938
rect 4497 -972 4531 -950
rect 4645 -168 4679 -146
rect 4645 -180 4679 -168
rect 4645 -236 4679 -218
rect 4645 -252 4679 -236
rect 4645 -304 4679 -290
rect 4645 -324 4679 -304
rect 4645 -372 4679 -362
rect 4645 -396 4679 -372
rect 4645 -440 4679 -434
rect 4645 -468 4679 -440
rect 4645 -508 4679 -506
rect 4645 -540 4679 -508
rect 4645 -610 4679 -578
rect 4645 -612 4679 -610
rect 4645 -678 4679 -650
rect 4645 -684 4679 -678
rect 4645 -746 4679 -722
rect 4645 -756 4679 -746
rect 4645 -814 4679 -794
rect 4645 -828 4679 -814
rect 4645 -882 4679 -866
rect 4645 -900 4679 -882
rect 4645 -950 4679 -938
rect 4645 -972 4679 -950
rect 4793 -168 4827 -146
rect 4793 -180 4827 -168
rect 4793 -236 4827 -218
rect 4793 -252 4827 -236
rect 4793 -304 4827 -290
rect 4793 -324 4827 -304
rect 4793 -372 4827 -362
rect 4793 -396 4827 -372
rect 4793 -440 4827 -434
rect 4793 -468 4827 -440
rect 4793 -508 4827 -506
rect 4793 -540 4827 -508
rect 4793 -610 4827 -578
rect 4793 -612 4827 -610
rect 4793 -678 4827 -650
rect 4793 -684 4827 -678
rect 4793 -746 4827 -722
rect 4793 -756 4827 -746
rect 4793 -814 4827 -794
rect 4793 -828 4827 -814
rect 4793 -882 4827 -866
rect 4793 -900 4827 -882
rect 4793 -950 4827 -938
rect 4793 -972 4827 -950
rect 4941 -168 4975 -146
rect 4941 -180 4975 -168
rect 4941 -236 4975 -218
rect 4941 -252 4975 -236
rect 4941 -304 4975 -290
rect 4941 -324 4975 -304
rect 4941 -372 4975 -362
rect 4941 -396 4975 -372
rect 4941 -440 4975 -434
rect 4941 -468 4975 -440
rect 4941 -508 4975 -506
rect 4941 -540 4975 -508
rect 4941 -610 4975 -578
rect 4941 -612 4975 -610
rect 4941 -678 4975 -650
rect 4941 -684 4975 -678
rect 4941 -746 4975 -722
rect 4941 -756 4975 -746
rect 4941 -814 4975 -794
rect 4941 -828 4975 -814
rect 4941 -882 4975 -866
rect 4941 -900 4975 -882
rect 4941 -950 4975 -938
rect 4941 -972 4975 -950
rect 5089 -168 5123 -146
rect 5089 -180 5123 -168
rect 5089 -236 5123 -218
rect 5089 -252 5123 -236
rect 5089 -304 5123 -290
rect 5089 -324 5123 -304
rect 5089 -372 5123 -362
rect 5089 -396 5123 -372
rect 5089 -440 5123 -434
rect 5089 -468 5123 -440
rect 5089 -508 5123 -506
rect 5089 -540 5123 -508
rect 5089 -610 5123 -578
rect 5089 -612 5123 -610
rect 5089 -678 5123 -650
rect 5089 -684 5123 -678
rect 5089 -746 5123 -722
rect 5089 -756 5123 -746
rect 5089 -814 5123 -794
rect 5089 -828 5123 -814
rect 5089 -882 5123 -866
rect 5089 -900 5123 -882
rect 5089 -950 5123 -938
rect 5089 -972 5123 -950
rect 5237 -168 5271 -146
rect 5237 -180 5271 -168
rect 5237 -236 5271 -218
rect 5237 -252 5271 -236
rect 5237 -304 5271 -290
rect 5237 -324 5271 -304
rect 5237 -372 5271 -362
rect 5237 -396 5271 -372
rect 5237 -440 5271 -434
rect 5237 -468 5271 -440
rect 5237 -508 5271 -506
rect 5237 -540 5271 -508
rect 5237 -610 5271 -578
rect 5237 -612 5271 -610
rect 5237 -678 5271 -650
rect 5237 -684 5271 -678
rect 5237 -746 5271 -722
rect 5237 -756 5271 -746
rect 5237 -814 5271 -794
rect 5237 -828 5271 -814
rect 5237 -882 5271 -866
rect 5237 -900 5271 -882
rect 5237 -950 5271 -938
rect 5237 -972 5271 -950
rect 5385 -168 5419 -146
rect 5385 -180 5419 -168
rect 5385 -236 5419 -218
rect 5385 -252 5419 -236
rect 5385 -304 5419 -290
rect 5385 -324 5419 -304
rect 5385 -372 5419 -362
rect 5385 -396 5419 -372
rect 5385 -440 5419 -434
rect 5385 -468 5419 -440
rect 5385 -508 5419 -506
rect 5385 -540 5419 -508
rect 5385 -610 5419 -578
rect 5385 -612 5419 -610
rect 5385 -678 5419 -650
rect 5385 -684 5419 -678
rect 5385 -746 5419 -722
rect 5385 -756 5419 -746
rect 5385 -814 5419 -794
rect 5385 -828 5419 -814
rect 5385 -882 5419 -866
rect 5385 -900 5419 -882
rect 5385 -950 5419 -938
rect 5385 -972 5419 -950
rect 5533 -168 5567 -146
rect 5533 -180 5567 -168
rect 5533 -236 5567 -218
rect 5533 -252 5567 -236
rect 5533 -304 5567 -290
rect 5533 -324 5567 -304
rect 5533 -372 5567 -362
rect 5533 -396 5567 -372
rect 5533 -440 5567 -434
rect 5533 -468 5567 -440
rect 5533 -508 5567 -506
rect 5533 -540 5567 -508
rect 5533 -610 5567 -578
rect 5533 -612 5567 -610
rect 5533 -678 5567 -650
rect 5533 -684 5567 -678
rect 5533 -746 5567 -722
rect 5533 -756 5567 -746
rect 5533 -814 5567 -794
rect 5533 -828 5567 -814
rect 5533 -882 5567 -866
rect 5533 -900 5567 -882
rect 5533 -950 5567 -938
rect 5533 -972 5567 -950
rect -5493 -1081 -5459 -1047
rect -5345 -1081 -5311 -1047
rect -5197 -1081 -5163 -1047
rect -5049 -1081 -5015 -1047
rect -4901 -1081 -4867 -1047
rect -4753 -1081 -4719 -1047
rect -4605 -1081 -4571 -1047
rect -4457 -1081 -4423 -1047
rect -4309 -1081 -4275 -1047
rect -4161 -1081 -4127 -1047
rect -4013 -1081 -3979 -1047
rect -3865 -1081 -3831 -1047
rect -3717 -1081 -3683 -1047
rect -3569 -1081 -3535 -1047
rect -3421 -1081 -3387 -1047
rect -3273 -1081 -3239 -1047
rect -3125 -1081 -3091 -1047
rect -2977 -1081 -2943 -1047
rect -2829 -1081 -2795 -1047
rect -2681 -1081 -2647 -1047
rect -2533 -1081 -2499 -1047
rect -2385 -1081 -2351 -1047
rect -2237 -1081 -2203 -1047
rect -2089 -1081 -2055 -1047
rect -1941 -1081 -1907 -1047
rect -1793 -1081 -1759 -1047
rect -1645 -1081 -1611 -1047
rect -1497 -1081 -1463 -1047
rect -1349 -1081 -1315 -1047
rect -1201 -1081 -1167 -1047
rect -1053 -1081 -1019 -1047
rect -905 -1081 -871 -1047
rect -757 -1081 -723 -1047
rect -609 -1081 -575 -1047
rect -461 -1081 -427 -1047
rect -313 -1081 -279 -1047
rect -165 -1081 -131 -1047
rect -17 -1081 17 -1047
rect 131 -1081 165 -1047
rect 279 -1081 313 -1047
rect 427 -1081 461 -1047
rect 575 -1081 609 -1047
rect 723 -1081 757 -1047
rect 871 -1081 905 -1047
rect 1019 -1081 1053 -1047
rect 1167 -1081 1201 -1047
rect 1315 -1081 1349 -1047
rect 1463 -1081 1497 -1047
rect 1611 -1081 1645 -1047
rect 1759 -1081 1793 -1047
rect 1907 -1081 1941 -1047
rect 2055 -1081 2089 -1047
rect 2203 -1081 2237 -1047
rect 2351 -1081 2385 -1047
rect 2499 -1081 2533 -1047
rect 2647 -1081 2681 -1047
rect 2795 -1081 2829 -1047
rect 2943 -1081 2977 -1047
rect 3091 -1081 3125 -1047
rect 3239 -1081 3273 -1047
rect 3387 -1081 3421 -1047
rect 3535 -1081 3569 -1047
rect 3683 -1081 3717 -1047
rect 3831 -1081 3865 -1047
rect 3979 -1081 4013 -1047
rect 4127 -1081 4161 -1047
rect 4275 -1081 4309 -1047
rect 4423 -1081 4457 -1047
rect 4571 -1081 4605 -1047
rect 4719 -1081 4753 -1047
rect 4867 -1081 4901 -1047
rect 5015 -1081 5049 -1047
rect 5163 -1081 5197 -1047
rect 5311 -1081 5345 -1047
rect 5459 -1081 5493 -1047
<< metal1 >>
rect -5517 1081 -5435 1087
rect -5517 1047 -5493 1081
rect -5459 1047 -5435 1081
rect -5517 1041 -5435 1047
rect -5369 1081 -5287 1087
rect -5369 1047 -5345 1081
rect -5311 1047 -5287 1081
rect -5369 1041 -5287 1047
rect -5221 1081 -5139 1087
rect -5221 1047 -5197 1081
rect -5163 1047 -5139 1081
rect -5221 1041 -5139 1047
rect -5073 1081 -4991 1087
rect -5073 1047 -5049 1081
rect -5015 1047 -4991 1081
rect -5073 1041 -4991 1047
rect -4925 1081 -4843 1087
rect -4925 1047 -4901 1081
rect -4867 1047 -4843 1081
rect -4925 1041 -4843 1047
rect -4777 1081 -4695 1087
rect -4777 1047 -4753 1081
rect -4719 1047 -4695 1081
rect -4777 1041 -4695 1047
rect -4629 1081 -4547 1087
rect -4629 1047 -4605 1081
rect -4571 1047 -4547 1081
rect -4629 1041 -4547 1047
rect -4481 1081 -4399 1087
rect -4481 1047 -4457 1081
rect -4423 1047 -4399 1081
rect -4481 1041 -4399 1047
rect -4333 1081 -4251 1087
rect -4333 1047 -4309 1081
rect -4275 1047 -4251 1081
rect -4333 1041 -4251 1047
rect -4185 1081 -4103 1087
rect -4185 1047 -4161 1081
rect -4127 1047 -4103 1081
rect -4185 1041 -4103 1047
rect -4037 1081 -3955 1087
rect -4037 1047 -4013 1081
rect -3979 1047 -3955 1081
rect -4037 1041 -3955 1047
rect -3889 1081 -3807 1087
rect -3889 1047 -3865 1081
rect -3831 1047 -3807 1081
rect -3889 1041 -3807 1047
rect -3741 1081 -3659 1087
rect -3741 1047 -3717 1081
rect -3683 1047 -3659 1081
rect -3741 1041 -3659 1047
rect -3593 1081 -3511 1087
rect -3593 1047 -3569 1081
rect -3535 1047 -3511 1081
rect -3593 1041 -3511 1047
rect -3445 1081 -3363 1087
rect -3445 1047 -3421 1081
rect -3387 1047 -3363 1081
rect -3445 1041 -3363 1047
rect -3297 1081 -3215 1087
rect -3297 1047 -3273 1081
rect -3239 1047 -3215 1081
rect -3297 1041 -3215 1047
rect -3149 1081 -3067 1087
rect -3149 1047 -3125 1081
rect -3091 1047 -3067 1081
rect -3149 1041 -3067 1047
rect -3001 1081 -2919 1087
rect -3001 1047 -2977 1081
rect -2943 1047 -2919 1081
rect -3001 1041 -2919 1047
rect -2853 1081 -2771 1087
rect -2853 1047 -2829 1081
rect -2795 1047 -2771 1081
rect -2853 1041 -2771 1047
rect -2705 1081 -2623 1087
rect -2705 1047 -2681 1081
rect -2647 1047 -2623 1081
rect -2705 1041 -2623 1047
rect -2557 1081 -2475 1087
rect -2557 1047 -2533 1081
rect -2499 1047 -2475 1081
rect -2557 1041 -2475 1047
rect -2409 1081 -2327 1087
rect -2409 1047 -2385 1081
rect -2351 1047 -2327 1081
rect -2409 1041 -2327 1047
rect -2261 1081 -2179 1087
rect -2261 1047 -2237 1081
rect -2203 1047 -2179 1081
rect -2261 1041 -2179 1047
rect -2113 1081 -2031 1087
rect -2113 1047 -2089 1081
rect -2055 1047 -2031 1081
rect -2113 1041 -2031 1047
rect -1965 1081 -1883 1087
rect -1965 1047 -1941 1081
rect -1907 1047 -1883 1081
rect -1965 1041 -1883 1047
rect -1817 1081 -1735 1087
rect -1817 1047 -1793 1081
rect -1759 1047 -1735 1081
rect -1817 1041 -1735 1047
rect -1669 1081 -1587 1087
rect -1669 1047 -1645 1081
rect -1611 1047 -1587 1081
rect -1669 1041 -1587 1047
rect -1521 1081 -1439 1087
rect -1521 1047 -1497 1081
rect -1463 1047 -1439 1081
rect -1521 1041 -1439 1047
rect -1373 1081 -1291 1087
rect -1373 1047 -1349 1081
rect -1315 1047 -1291 1081
rect -1373 1041 -1291 1047
rect -1225 1081 -1143 1087
rect -1225 1047 -1201 1081
rect -1167 1047 -1143 1081
rect -1225 1041 -1143 1047
rect -1077 1081 -995 1087
rect -1077 1047 -1053 1081
rect -1019 1047 -995 1081
rect -1077 1041 -995 1047
rect -929 1081 -847 1087
rect -929 1047 -905 1081
rect -871 1047 -847 1081
rect -929 1041 -847 1047
rect -781 1081 -699 1087
rect -781 1047 -757 1081
rect -723 1047 -699 1081
rect -781 1041 -699 1047
rect -633 1081 -551 1087
rect -633 1047 -609 1081
rect -575 1047 -551 1081
rect -633 1041 -551 1047
rect -485 1081 -403 1087
rect -485 1047 -461 1081
rect -427 1047 -403 1081
rect -485 1041 -403 1047
rect -337 1081 -255 1087
rect -337 1047 -313 1081
rect -279 1047 -255 1081
rect -337 1041 -255 1047
rect -189 1081 -107 1087
rect -189 1047 -165 1081
rect -131 1047 -107 1081
rect -189 1041 -107 1047
rect -41 1081 41 1087
rect -41 1047 -17 1081
rect 17 1047 41 1081
rect -41 1041 41 1047
rect 107 1081 189 1087
rect 107 1047 131 1081
rect 165 1047 189 1081
rect 107 1041 189 1047
rect 255 1081 337 1087
rect 255 1047 279 1081
rect 313 1047 337 1081
rect 255 1041 337 1047
rect 403 1081 485 1087
rect 403 1047 427 1081
rect 461 1047 485 1081
rect 403 1041 485 1047
rect 551 1081 633 1087
rect 551 1047 575 1081
rect 609 1047 633 1081
rect 551 1041 633 1047
rect 699 1081 781 1087
rect 699 1047 723 1081
rect 757 1047 781 1081
rect 699 1041 781 1047
rect 847 1081 929 1087
rect 847 1047 871 1081
rect 905 1047 929 1081
rect 847 1041 929 1047
rect 995 1081 1077 1087
rect 995 1047 1019 1081
rect 1053 1047 1077 1081
rect 995 1041 1077 1047
rect 1143 1081 1225 1087
rect 1143 1047 1167 1081
rect 1201 1047 1225 1081
rect 1143 1041 1225 1047
rect 1291 1081 1373 1087
rect 1291 1047 1315 1081
rect 1349 1047 1373 1081
rect 1291 1041 1373 1047
rect 1439 1081 1521 1087
rect 1439 1047 1463 1081
rect 1497 1047 1521 1081
rect 1439 1041 1521 1047
rect 1587 1081 1669 1087
rect 1587 1047 1611 1081
rect 1645 1047 1669 1081
rect 1587 1041 1669 1047
rect 1735 1081 1817 1087
rect 1735 1047 1759 1081
rect 1793 1047 1817 1081
rect 1735 1041 1817 1047
rect 1883 1081 1965 1087
rect 1883 1047 1907 1081
rect 1941 1047 1965 1081
rect 1883 1041 1965 1047
rect 2031 1081 2113 1087
rect 2031 1047 2055 1081
rect 2089 1047 2113 1081
rect 2031 1041 2113 1047
rect 2179 1081 2261 1087
rect 2179 1047 2203 1081
rect 2237 1047 2261 1081
rect 2179 1041 2261 1047
rect 2327 1081 2409 1087
rect 2327 1047 2351 1081
rect 2385 1047 2409 1081
rect 2327 1041 2409 1047
rect 2475 1081 2557 1087
rect 2475 1047 2499 1081
rect 2533 1047 2557 1081
rect 2475 1041 2557 1047
rect 2623 1081 2705 1087
rect 2623 1047 2647 1081
rect 2681 1047 2705 1081
rect 2623 1041 2705 1047
rect 2771 1081 2853 1087
rect 2771 1047 2795 1081
rect 2829 1047 2853 1081
rect 2771 1041 2853 1047
rect 2919 1081 3001 1087
rect 2919 1047 2943 1081
rect 2977 1047 3001 1081
rect 2919 1041 3001 1047
rect 3067 1081 3149 1087
rect 3067 1047 3091 1081
rect 3125 1047 3149 1081
rect 3067 1041 3149 1047
rect 3215 1081 3297 1087
rect 3215 1047 3239 1081
rect 3273 1047 3297 1081
rect 3215 1041 3297 1047
rect 3363 1081 3445 1087
rect 3363 1047 3387 1081
rect 3421 1047 3445 1081
rect 3363 1041 3445 1047
rect 3511 1081 3593 1087
rect 3511 1047 3535 1081
rect 3569 1047 3593 1081
rect 3511 1041 3593 1047
rect 3659 1081 3741 1087
rect 3659 1047 3683 1081
rect 3717 1047 3741 1081
rect 3659 1041 3741 1047
rect 3807 1081 3889 1087
rect 3807 1047 3831 1081
rect 3865 1047 3889 1081
rect 3807 1041 3889 1047
rect 3955 1081 4037 1087
rect 3955 1047 3979 1081
rect 4013 1047 4037 1081
rect 3955 1041 4037 1047
rect 4103 1081 4185 1087
rect 4103 1047 4127 1081
rect 4161 1047 4185 1081
rect 4103 1041 4185 1047
rect 4251 1081 4333 1087
rect 4251 1047 4275 1081
rect 4309 1047 4333 1081
rect 4251 1041 4333 1047
rect 4399 1081 4481 1087
rect 4399 1047 4423 1081
rect 4457 1047 4481 1081
rect 4399 1041 4481 1047
rect 4547 1081 4629 1087
rect 4547 1047 4571 1081
rect 4605 1047 4629 1081
rect 4547 1041 4629 1047
rect 4695 1081 4777 1087
rect 4695 1047 4719 1081
rect 4753 1047 4777 1081
rect 4695 1041 4777 1047
rect 4843 1081 4925 1087
rect 4843 1047 4867 1081
rect 4901 1047 4925 1081
rect 4843 1041 4925 1047
rect 4991 1081 5073 1087
rect 4991 1047 5015 1081
rect 5049 1047 5073 1081
rect 4991 1041 5073 1047
rect 5139 1081 5221 1087
rect 5139 1047 5163 1081
rect 5197 1047 5221 1081
rect 5139 1041 5221 1047
rect 5287 1081 5369 1087
rect 5287 1047 5311 1081
rect 5345 1047 5369 1081
rect 5287 1041 5369 1047
rect 5435 1081 5517 1087
rect 5435 1047 5459 1081
rect 5493 1047 5517 1081
rect 5435 1041 5517 1047
rect -5573 972 -5527 1009
rect -5573 938 -5567 972
rect -5533 938 -5527 972
rect -5573 900 -5527 938
rect -5573 866 -5567 900
rect -5533 866 -5527 900
rect -5573 828 -5527 866
rect -5573 794 -5567 828
rect -5533 794 -5527 828
rect -5573 756 -5527 794
rect -5573 722 -5567 756
rect -5533 722 -5527 756
rect -5573 684 -5527 722
rect -5573 650 -5567 684
rect -5533 650 -5527 684
rect -5573 612 -5527 650
rect -5573 578 -5567 612
rect -5533 578 -5527 612
rect -5573 540 -5527 578
rect -5573 506 -5567 540
rect -5533 506 -5527 540
rect -5573 468 -5527 506
rect -5573 434 -5567 468
rect -5533 434 -5527 468
rect -5573 396 -5527 434
rect -5573 362 -5567 396
rect -5533 362 -5527 396
rect -5573 324 -5527 362
rect -5573 290 -5567 324
rect -5533 290 -5527 324
rect -5573 252 -5527 290
rect -5573 218 -5567 252
rect -5533 218 -5527 252
rect -5573 180 -5527 218
rect -5573 146 -5567 180
rect -5533 146 -5527 180
rect -5573 109 -5527 146
rect -5425 972 -5379 1009
rect -5425 938 -5419 972
rect -5385 938 -5379 972
rect -5425 900 -5379 938
rect -5425 866 -5419 900
rect -5385 866 -5379 900
rect -5425 828 -5379 866
rect -5425 794 -5419 828
rect -5385 794 -5379 828
rect -5425 756 -5379 794
rect -5425 722 -5419 756
rect -5385 722 -5379 756
rect -5425 684 -5379 722
rect -5425 650 -5419 684
rect -5385 650 -5379 684
rect -5425 612 -5379 650
rect -5425 578 -5419 612
rect -5385 578 -5379 612
rect -5425 540 -5379 578
rect -5425 506 -5419 540
rect -5385 506 -5379 540
rect -5425 468 -5379 506
rect -5425 434 -5419 468
rect -5385 434 -5379 468
rect -5425 396 -5379 434
rect -5425 362 -5419 396
rect -5385 362 -5379 396
rect -5425 324 -5379 362
rect -5425 290 -5419 324
rect -5385 290 -5379 324
rect -5425 252 -5379 290
rect -5425 218 -5419 252
rect -5385 218 -5379 252
rect -5425 180 -5379 218
rect -5425 146 -5419 180
rect -5385 146 -5379 180
rect -5425 109 -5379 146
rect -5277 972 -5231 1009
rect -5277 938 -5271 972
rect -5237 938 -5231 972
rect -5277 900 -5231 938
rect -5277 866 -5271 900
rect -5237 866 -5231 900
rect -5277 828 -5231 866
rect -5277 794 -5271 828
rect -5237 794 -5231 828
rect -5277 756 -5231 794
rect -5277 722 -5271 756
rect -5237 722 -5231 756
rect -5277 684 -5231 722
rect -5277 650 -5271 684
rect -5237 650 -5231 684
rect -5277 612 -5231 650
rect -5277 578 -5271 612
rect -5237 578 -5231 612
rect -5277 540 -5231 578
rect -5277 506 -5271 540
rect -5237 506 -5231 540
rect -5277 468 -5231 506
rect -5277 434 -5271 468
rect -5237 434 -5231 468
rect -5277 396 -5231 434
rect -5277 362 -5271 396
rect -5237 362 -5231 396
rect -5277 324 -5231 362
rect -5277 290 -5271 324
rect -5237 290 -5231 324
rect -5277 252 -5231 290
rect -5277 218 -5271 252
rect -5237 218 -5231 252
rect -5277 180 -5231 218
rect -5277 146 -5271 180
rect -5237 146 -5231 180
rect -5277 109 -5231 146
rect -5129 972 -5083 1009
rect -5129 938 -5123 972
rect -5089 938 -5083 972
rect -5129 900 -5083 938
rect -5129 866 -5123 900
rect -5089 866 -5083 900
rect -5129 828 -5083 866
rect -5129 794 -5123 828
rect -5089 794 -5083 828
rect -5129 756 -5083 794
rect -5129 722 -5123 756
rect -5089 722 -5083 756
rect -5129 684 -5083 722
rect -5129 650 -5123 684
rect -5089 650 -5083 684
rect -5129 612 -5083 650
rect -5129 578 -5123 612
rect -5089 578 -5083 612
rect -5129 540 -5083 578
rect -5129 506 -5123 540
rect -5089 506 -5083 540
rect -5129 468 -5083 506
rect -5129 434 -5123 468
rect -5089 434 -5083 468
rect -5129 396 -5083 434
rect -5129 362 -5123 396
rect -5089 362 -5083 396
rect -5129 324 -5083 362
rect -5129 290 -5123 324
rect -5089 290 -5083 324
rect -5129 252 -5083 290
rect -5129 218 -5123 252
rect -5089 218 -5083 252
rect -5129 180 -5083 218
rect -5129 146 -5123 180
rect -5089 146 -5083 180
rect -5129 109 -5083 146
rect -4981 972 -4935 1009
rect -4981 938 -4975 972
rect -4941 938 -4935 972
rect -4981 900 -4935 938
rect -4981 866 -4975 900
rect -4941 866 -4935 900
rect -4981 828 -4935 866
rect -4981 794 -4975 828
rect -4941 794 -4935 828
rect -4981 756 -4935 794
rect -4981 722 -4975 756
rect -4941 722 -4935 756
rect -4981 684 -4935 722
rect -4981 650 -4975 684
rect -4941 650 -4935 684
rect -4981 612 -4935 650
rect -4981 578 -4975 612
rect -4941 578 -4935 612
rect -4981 540 -4935 578
rect -4981 506 -4975 540
rect -4941 506 -4935 540
rect -4981 468 -4935 506
rect -4981 434 -4975 468
rect -4941 434 -4935 468
rect -4981 396 -4935 434
rect -4981 362 -4975 396
rect -4941 362 -4935 396
rect -4981 324 -4935 362
rect -4981 290 -4975 324
rect -4941 290 -4935 324
rect -4981 252 -4935 290
rect -4981 218 -4975 252
rect -4941 218 -4935 252
rect -4981 180 -4935 218
rect -4981 146 -4975 180
rect -4941 146 -4935 180
rect -4981 109 -4935 146
rect -4833 972 -4787 1009
rect -4833 938 -4827 972
rect -4793 938 -4787 972
rect -4833 900 -4787 938
rect -4833 866 -4827 900
rect -4793 866 -4787 900
rect -4833 828 -4787 866
rect -4833 794 -4827 828
rect -4793 794 -4787 828
rect -4833 756 -4787 794
rect -4833 722 -4827 756
rect -4793 722 -4787 756
rect -4833 684 -4787 722
rect -4833 650 -4827 684
rect -4793 650 -4787 684
rect -4833 612 -4787 650
rect -4833 578 -4827 612
rect -4793 578 -4787 612
rect -4833 540 -4787 578
rect -4833 506 -4827 540
rect -4793 506 -4787 540
rect -4833 468 -4787 506
rect -4833 434 -4827 468
rect -4793 434 -4787 468
rect -4833 396 -4787 434
rect -4833 362 -4827 396
rect -4793 362 -4787 396
rect -4833 324 -4787 362
rect -4833 290 -4827 324
rect -4793 290 -4787 324
rect -4833 252 -4787 290
rect -4833 218 -4827 252
rect -4793 218 -4787 252
rect -4833 180 -4787 218
rect -4833 146 -4827 180
rect -4793 146 -4787 180
rect -4833 109 -4787 146
rect -4685 972 -4639 1009
rect -4685 938 -4679 972
rect -4645 938 -4639 972
rect -4685 900 -4639 938
rect -4685 866 -4679 900
rect -4645 866 -4639 900
rect -4685 828 -4639 866
rect -4685 794 -4679 828
rect -4645 794 -4639 828
rect -4685 756 -4639 794
rect -4685 722 -4679 756
rect -4645 722 -4639 756
rect -4685 684 -4639 722
rect -4685 650 -4679 684
rect -4645 650 -4639 684
rect -4685 612 -4639 650
rect -4685 578 -4679 612
rect -4645 578 -4639 612
rect -4685 540 -4639 578
rect -4685 506 -4679 540
rect -4645 506 -4639 540
rect -4685 468 -4639 506
rect -4685 434 -4679 468
rect -4645 434 -4639 468
rect -4685 396 -4639 434
rect -4685 362 -4679 396
rect -4645 362 -4639 396
rect -4685 324 -4639 362
rect -4685 290 -4679 324
rect -4645 290 -4639 324
rect -4685 252 -4639 290
rect -4685 218 -4679 252
rect -4645 218 -4639 252
rect -4685 180 -4639 218
rect -4685 146 -4679 180
rect -4645 146 -4639 180
rect -4685 109 -4639 146
rect -4537 972 -4491 1009
rect -4537 938 -4531 972
rect -4497 938 -4491 972
rect -4537 900 -4491 938
rect -4537 866 -4531 900
rect -4497 866 -4491 900
rect -4537 828 -4491 866
rect -4537 794 -4531 828
rect -4497 794 -4491 828
rect -4537 756 -4491 794
rect -4537 722 -4531 756
rect -4497 722 -4491 756
rect -4537 684 -4491 722
rect -4537 650 -4531 684
rect -4497 650 -4491 684
rect -4537 612 -4491 650
rect -4537 578 -4531 612
rect -4497 578 -4491 612
rect -4537 540 -4491 578
rect -4537 506 -4531 540
rect -4497 506 -4491 540
rect -4537 468 -4491 506
rect -4537 434 -4531 468
rect -4497 434 -4491 468
rect -4537 396 -4491 434
rect -4537 362 -4531 396
rect -4497 362 -4491 396
rect -4537 324 -4491 362
rect -4537 290 -4531 324
rect -4497 290 -4491 324
rect -4537 252 -4491 290
rect -4537 218 -4531 252
rect -4497 218 -4491 252
rect -4537 180 -4491 218
rect -4537 146 -4531 180
rect -4497 146 -4491 180
rect -4537 109 -4491 146
rect -4389 972 -4343 1009
rect -4389 938 -4383 972
rect -4349 938 -4343 972
rect -4389 900 -4343 938
rect -4389 866 -4383 900
rect -4349 866 -4343 900
rect -4389 828 -4343 866
rect -4389 794 -4383 828
rect -4349 794 -4343 828
rect -4389 756 -4343 794
rect -4389 722 -4383 756
rect -4349 722 -4343 756
rect -4389 684 -4343 722
rect -4389 650 -4383 684
rect -4349 650 -4343 684
rect -4389 612 -4343 650
rect -4389 578 -4383 612
rect -4349 578 -4343 612
rect -4389 540 -4343 578
rect -4389 506 -4383 540
rect -4349 506 -4343 540
rect -4389 468 -4343 506
rect -4389 434 -4383 468
rect -4349 434 -4343 468
rect -4389 396 -4343 434
rect -4389 362 -4383 396
rect -4349 362 -4343 396
rect -4389 324 -4343 362
rect -4389 290 -4383 324
rect -4349 290 -4343 324
rect -4389 252 -4343 290
rect -4389 218 -4383 252
rect -4349 218 -4343 252
rect -4389 180 -4343 218
rect -4389 146 -4383 180
rect -4349 146 -4343 180
rect -4389 109 -4343 146
rect -4241 972 -4195 1009
rect -4241 938 -4235 972
rect -4201 938 -4195 972
rect -4241 900 -4195 938
rect -4241 866 -4235 900
rect -4201 866 -4195 900
rect -4241 828 -4195 866
rect -4241 794 -4235 828
rect -4201 794 -4195 828
rect -4241 756 -4195 794
rect -4241 722 -4235 756
rect -4201 722 -4195 756
rect -4241 684 -4195 722
rect -4241 650 -4235 684
rect -4201 650 -4195 684
rect -4241 612 -4195 650
rect -4241 578 -4235 612
rect -4201 578 -4195 612
rect -4241 540 -4195 578
rect -4241 506 -4235 540
rect -4201 506 -4195 540
rect -4241 468 -4195 506
rect -4241 434 -4235 468
rect -4201 434 -4195 468
rect -4241 396 -4195 434
rect -4241 362 -4235 396
rect -4201 362 -4195 396
rect -4241 324 -4195 362
rect -4241 290 -4235 324
rect -4201 290 -4195 324
rect -4241 252 -4195 290
rect -4241 218 -4235 252
rect -4201 218 -4195 252
rect -4241 180 -4195 218
rect -4241 146 -4235 180
rect -4201 146 -4195 180
rect -4241 109 -4195 146
rect -4093 972 -4047 1009
rect -4093 938 -4087 972
rect -4053 938 -4047 972
rect -4093 900 -4047 938
rect -4093 866 -4087 900
rect -4053 866 -4047 900
rect -4093 828 -4047 866
rect -4093 794 -4087 828
rect -4053 794 -4047 828
rect -4093 756 -4047 794
rect -4093 722 -4087 756
rect -4053 722 -4047 756
rect -4093 684 -4047 722
rect -4093 650 -4087 684
rect -4053 650 -4047 684
rect -4093 612 -4047 650
rect -4093 578 -4087 612
rect -4053 578 -4047 612
rect -4093 540 -4047 578
rect -4093 506 -4087 540
rect -4053 506 -4047 540
rect -4093 468 -4047 506
rect -4093 434 -4087 468
rect -4053 434 -4047 468
rect -4093 396 -4047 434
rect -4093 362 -4087 396
rect -4053 362 -4047 396
rect -4093 324 -4047 362
rect -4093 290 -4087 324
rect -4053 290 -4047 324
rect -4093 252 -4047 290
rect -4093 218 -4087 252
rect -4053 218 -4047 252
rect -4093 180 -4047 218
rect -4093 146 -4087 180
rect -4053 146 -4047 180
rect -4093 109 -4047 146
rect -3945 972 -3899 1009
rect -3945 938 -3939 972
rect -3905 938 -3899 972
rect -3945 900 -3899 938
rect -3945 866 -3939 900
rect -3905 866 -3899 900
rect -3945 828 -3899 866
rect -3945 794 -3939 828
rect -3905 794 -3899 828
rect -3945 756 -3899 794
rect -3945 722 -3939 756
rect -3905 722 -3899 756
rect -3945 684 -3899 722
rect -3945 650 -3939 684
rect -3905 650 -3899 684
rect -3945 612 -3899 650
rect -3945 578 -3939 612
rect -3905 578 -3899 612
rect -3945 540 -3899 578
rect -3945 506 -3939 540
rect -3905 506 -3899 540
rect -3945 468 -3899 506
rect -3945 434 -3939 468
rect -3905 434 -3899 468
rect -3945 396 -3899 434
rect -3945 362 -3939 396
rect -3905 362 -3899 396
rect -3945 324 -3899 362
rect -3945 290 -3939 324
rect -3905 290 -3899 324
rect -3945 252 -3899 290
rect -3945 218 -3939 252
rect -3905 218 -3899 252
rect -3945 180 -3899 218
rect -3945 146 -3939 180
rect -3905 146 -3899 180
rect -3945 109 -3899 146
rect -3797 972 -3751 1009
rect -3797 938 -3791 972
rect -3757 938 -3751 972
rect -3797 900 -3751 938
rect -3797 866 -3791 900
rect -3757 866 -3751 900
rect -3797 828 -3751 866
rect -3797 794 -3791 828
rect -3757 794 -3751 828
rect -3797 756 -3751 794
rect -3797 722 -3791 756
rect -3757 722 -3751 756
rect -3797 684 -3751 722
rect -3797 650 -3791 684
rect -3757 650 -3751 684
rect -3797 612 -3751 650
rect -3797 578 -3791 612
rect -3757 578 -3751 612
rect -3797 540 -3751 578
rect -3797 506 -3791 540
rect -3757 506 -3751 540
rect -3797 468 -3751 506
rect -3797 434 -3791 468
rect -3757 434 -3751 468
rect -3797 396 -3751 434
rect -3797 362 -3791 396
rect -3757 362 -3751 396
rect -3797 324 -3751 362
rect -3797 290 -3791 324
rect -3757 290 -3751 324
rect -3797 252 -3751 290
rect -3797 218 -3791 252
rect -3757 218 -3751 252
rect -3797 180 -3751 218
rect -3797 146 -3791 180
rect -3757 146 -3751 180
rect -3797 109 -3751 146
rect -3649 972 -3603 1009
rect -3649 938 -3643 972
rect -3609 938 -3603 972
rect -3649 900 -3603 938
rect -3649 866 -3643 900
rect -3609 866 -3603 900
rect -3649 828 -3603 866
rect -3649 794 -3643 828
rect -3609 794 -3603 828
rect -3649 756 -3603 794
rect -3649 722 -3643 756
rect -3609 722 -3603 756
rect -3649 684 -3603 722
rect -3649 650 -3643 684
rect -3609 650 -3603 684
rect -3649 612 -3603 650
rect -3649 578 -3643 612
rect -3609 578 -3603 612
rect -3649 540 -3603 578
rect -3649 506 -3643 540
rect -3609 506 -3603 540
rect -3649 468 -3603 506
rect -3649 434 -3643 468
rect -3609 434 -3603 468
rect -3649 396 -3603 434
rect -3649 362 -3643 396
rect -3609 362 -3603 396
rect -3649 324 -3603 362
rect -3649 290 -3643 324
rect -3609 290 -3603 324
rect -3649 252 -3603 290
rect -3649 218 -3643 252
rect -3609 218 -3603 252
rect -3649 180 -3603 218
rect -3649 146 -3643 180
rect -3609 146 -3603 180
rect -3649 109 -3603 146
rect -3501 972 -3455 1009
rect -3501 938 -3495 972
rect -3461 938 -3455 972
rect -3501 900 -3455 938
rect -3501 866 -3495 900
rect -3461 866 -3455 900
rect -3501 828 -3455 866
rect -3501 794 -3495 828
rect -3461 794 -3455 828
rect -3501 756 -3455 794
rect -3501 722 -3495 756
rect -3461 722 -3455 756
rect -3501 684 -3455 722
rect -3501 650 -3495 684
rect -3461 650 -3455 684
rect -3501 612 -3455 650
rect -3501 578 -3495 612
rect -3461 578 -3455 612
rect -3501 540 -3455 578
rect -3501 506 -3495 540
rect -3461 506 -3455 540
rect -3501 468 -3455 506
rect -3501 434 -3495 468
rect -3461 434 -3455 468
rect -3501 396 -3455 434
rect -3501 362 -3495 396
rect -3461 362 -3455 396
rect -3501 324 -3455 362
rect -3501 290 -3495 324
rect -3461 290 -3455 324
rect -3501 252 -3455 290
rect -3501 218 -3495 252
rect -3461 218 -3455 252
rect -3501 180 -3455 218
rect -3501 146 -3495 180
rect -3461 146 -3455 180
rect -3501 109 -3455 146
rect -3353 972 -3307 1009
rect -3353 938 -3347 972
rect -3313 938 -3307 972
rect -3353 900 -3307 938
rect -3353 866 -3347 900
rect -3313 866 -3307 900
rect -3353 828 -3307 866
rect -3353 794 -3347 828
rect -3313 794 -3307 828
rect -3353 756 -3307 794
rect -3353 722 -3347 756
rect -3313 722 -3307 756
rect -3353 684 -3307 722
rect -3353 650 -3347 684
rect -3313 650 -3307 684
rect -3353 612 -3307 650
rect -3353 578 -3347 612
rect -3313 578 -3307 612
rect -3353 540 -3307 578
rect -3353 506 -3347 540
rect -3313 506 -3307 540
rect -3353 468 -3307 506
rect -3353 434 -3347 468
rect -3313 434 -3307 468
rect -3353 396 -3307 434
rect -3353 362 -3347 396
rect -3313 362 -3307 396
rect -3353 324 -3307 362
rect -3353 290 -3347 324
rect -3313 290 -3307 324
rect -3353 252 -3307 290
rect -3353 218 -3347 252
rect -3313 218 -3307 252
rect -3353 180 -3307 218
rect -3353 146 -3347 180
rect -3313 146 -3307 180
rect -3353 109 -3307 146
rect -3205 972 -3159 1009
rect -3205 938 -3199 972
rect -3165 938 -3159 972
rect -3205 900 -3159 938
rect -3205 866 -3199 900
rect -3165 866 -3159 900
rect -3205 828 -3159 866
rect -3205 794 -3199 828
rect -3165 794 -3159 828
rect -3205 756 -3159 794
rect -3205 722 -3199 756
rect -3165 722 -3159 756
rect -3205 684 -3159 722
rect -3205 650 -3199 684
rect -3165 650 -3159 684
rect -3205 612 -3159 650
rect -3205 578 -3199 612
rect -3165 578 -3159 612
rect -3205 540 -3159 578
rect -3205 506 -3199 540
rect -3165 506 -3159 540
rect -3205 468 -3159 506
rect -3205 434 -3199 468
rect -3165 434 -3159 468
rect -3205 396 -3159 434
rect -3205 362 -3199 396
rect -3165 362 -3159 396
rect -3205 324 -3159 362
rect -3205 290 -3199 324
rect -3165 290 -3159 324
rect -3205 252 -3159 290
rect -3205 218 -3199 252
rect -3165 218 -3159 252
rect -3205 180 -3159 218
rect -3205 146 -3199 180
rect -3165 146 -3159 180
rect -3205 109 -3159 146
rect -3057 972 -3011 1009
rect -3057 938 -3051 972
rect -3017 938 -3011 972
rect -3057 900 -3011 938
rect -3057 866 -3051 900
rect -3017 866 -3011 900
rect -3057 828 -3011 866
rect -3057 794 -3051 828
rect -3017 794 -3011 828
rect -3057 756 -3011 794
rect -3057 722 -3051 756
rect -3017 722 -3011 756
rect -3057 684 -3011 722
rect -3057 650 -3051 684
rect -3017 650 -3011 684
rect -3057 612 -3011 650
rect -3057 578 -3051 612
rect -3017 578 -3011 612
rect -3057 540 -3011 578
rect -3057 506 -3051 540
rect -3017 506 -3011 540
rect -3057 468 -3011 506
rect -3057 434 -3051 468
rect -3017 434 -3011 468
rect -3057 396 -3011 434
rect -3057 362 -3051 396
rect -3017 362 -3011 396
rect -3057 324 -3011 362
rect -3057 290 -3051 324
rect -3017 290 -3011 324
rect -3057 252 -3011 290
rect -3057 218 -3051 252
rect -3017 218 -3011 252
rect -3057 180 -3011 218
rect -3057 146 -3051 180
rect -3017 146 -3011 180
rect -3057 109 -3011 146
rect -2909 972 -2863 1009
rect -2909 938 -2903 972
rect -2869 938 -2863 972
rect -2909 900 -2863 938
rect -2909 866 -2903 900
rect -2869 866 -2863 900
rect -2909 828 -2863 866
rect -2909 794 -2903 828
rect -2869 794 -2863 828
rect -2909 756 -2863 794
rect -2909 722 -2903 756
rect -2869 722 -2863 756
rect -2909 684 -2863 722
rect -2909 650 -2903 684
rect -2869 650 -2863 684
rect -2909 612 -2863 650
rect -2909 578 -2903 612
rect -2869 578 -2863 612
rect -2909 540 -2863 578
rect -2909 506 -2903 540
rect -2869 506 -2863 540
rect -2909 468 -2863 506
rect -2909 434 -2903 468
rect -2869 434 -2863 468
rect -2909 396 -2863 434
rect -2909 362 -2903 396
rect -2869 362 -2863 396
rect -2909 324 -2863 362
rect -2909 290 -2903 324
rect -2869 290 -2863 324
rect -2909 252 -2863 290
rect -2909 218 -2903 252
rect -2869 218 -2863 252
rect -2909 180 -2863 218
rect -2909 146 -2903 180
rect -2869 146 -2863 180
rect -2909 109 -2863 146
rect -2761 972 -2715 1009
rect -2761 938 -2755 972
rect -2721 938 -2715 972
rect -2761 900 -2715 938
rect -2761 866 -2755 900
rect -2721 866 -2715 900
rect -2761 828 -2715 866
rect -2761 794 -2755 828
rect -2721 794 -2715 828
rect -2761 756 -2715 794
rect -2761 722 -2755 756
rect -2721 722 -2715 756
rect -2761 684 -2715 722
rect -2761 650 -2755 684
rect -2721 650 -2715 684
rect -2761 612 -2715 650
rect -2761 578 -2755 612
rect -2721 578 -2715 612
rect -2761 540 -2715 578
rect -2761 506 -2755 540
rect -2721 506 -2715 540
rect -2761 468 -2715 506
rect -2761 434 -2755 468
rect -2721 434 -2715 468
rect -2761 396 -2715 434
rect -2761 362 -2755 396
rect -2721 362 -2715 396
rect -2761 324 -2715 362
rect -2761 290 -2755 324
rect -2721 290 -2715 324
rect -2761 252 -2715 290
rect -2761 218 -2755 252
rect -2721 218 -2715 252
rect -2761 180 -2715 218
rect -2761 146 -2755 180
rect -2721 146 -2715 180
rect -2761 109 -2715 146
rect -2613 972 -2567 1009
rect -2613 938 -2607 972
rect -2573 938 -2567 972
rect -2613 900 -2567 938
rect -2613 866 -2607 900
rect -2573 866 -2567 900
rect -2613 828 -2567 866
rect -2613 794 -2607 828
rect -2573 794 -2567 828
rect -2613 756 -2567 794
rect -2613 722 -2607 756
rect -2573 722 -2567 756
rect -2613 684 -2567 722
rect -2613 650 -2607 684
rect -2573 650 -2567 684
rect -2613 612 -2567 650
rect -2613 578 -2607 612
rect -2573 578 -2567 612
rect -2613 540 -2567 578
rect -2613 506 -2607 540
rect -2573 506 -2567 540
rect -2613 468 -2567 506
rect -2613 434 -2607 468
rect -2573 434 -2567 468
rect -2613 396 -2567 434
rect -2613 362 -2607 396
rect -2573 362 -2567 396
rect -2613 324 -2567 362
rect -2613 290 -2607 324
rect -2573 290 -2567 324
rect -2613 252 -2567 290
rect -2613 218 -2607 252
rect -2573 218 -2567 252
rect -2613 180 -2567 218
rect -2613 146 -2607 180
rect -2573 146 -2567 180
rect -2613 109 -2567 146
rect -2465 972 -2419 1009
rect -2465 938 -2459 972
rect -2425 938 -2419 972
rect -2465 900 -2419 938
rect -2465 866 -2459 900
rect -2425 866 -2419 900
rect -2465 828 -2419 866
rect -2465 794 -2459 828
rect -2425 794 -2419 828
rect -2465 756 -2419 794
rect -2465 722 -2459 756
rect -2425 722 -2419 756
rect -2465 684 -2419 722
rect -2465 650 -2459 684
rect -2425 650 -2419 684
rect -2465 612 -2419 650
rect -2465 578 -2459 612
rect -2425 578 -2419 612
rect -2465 540 -2419 578
rect -2465 506 -2459 540
rect -2425 506 -2419 540
rect -2465 468 -2419 506
rect -2465 434 -2459 468
rect -2425 434 -2419 468
rect -2465 396 -2419 434
rect -2465 362 -2459 396
rect -2425 362 -2419 396
rect -2465 324 -2419 362
rect -2465 290 -2459 324
rect -2425 290 -2419 324
rect -2465 252 -2419 290
rect -2465 218 -2459 252
rect -2425 218 -2419 252
rect -2465 180 -2419 218
rect -2465 146 -2459 180
rect -2425 146 -2419 180
rect -2465 109 -2419 146
rect -2317 972 -2271 1009
rect -2317 938 -2311 972
rect -2277 938 -2271 972
rect -2317 900 -2271 938
rect -2317 866 -2311 900
rect -2277 866 -2271 900
rect -2317 828 -2271 866
rect -2317 794 -2311 828
rect -2277 794 -2271 828
rect -2317 756 -2271 794
rect -2317 722 -2311 756
rect -2277 722 -2271 756
rect -2317 684 -2271 722
rect -2317 650 -2311 684
rect -2277 650 -2271 684
rect -2317 612 -2271 650
rect -2317 578 -2311 612
rect -2277 578 -2271 612
rect -2317 540 -2271 578
rect -2317 506 -2311 540
rect -2277 506 -2271 540
rect -2317 468 -2271 506
rect -2317 434 -2311 468
rect -2277 434 -2271 468
rect -2317 396 -2271 434
rect -2317 362 -2311 396
rect -2277 362 -2271 396
rect -2317 324 -2271 362
rect -2317 290 -2311 324
rect -2277 290 -2271 324
rect -2317 252 -2271 290
rect -2317 218 -2311 252
rect -2277 218 -2271 252
rect -2317 180 -2271 218
rect -2317 146 -2311 180
rect -2277 146 -2271 180
rect -2317 109 -2271 146
rect -2169 972 -2123 1009
rect -2169 938 -2163 972
rect -2129 938 -2123 972
rect -2169 900 -2123 938
rect -2169 866 -2163 900
rect -2129 866 -2123 900
rect -2169 828 -2123 866
rect -2169 794 -2163 828
rect -2129 794 -2123 828
rect -2169 756 -2123 794
rect -2169 722 -2163 756
rect -2129 722 -2123 756
rect -2169 684 -2123 722
rect -2169 650 -2163 684
rect -2129 650 -2123 684
rect -2169 612 -2123 650
rect -2169 578 -2163 612
rect -2129 578 -2123 612
rect -2169 540 -2123 578
rect -2169 506 -2163 540
rect -2129 506 -2123 540
rect -2169 468 -2123 506
rect -2169 434 -2163 468
rect -2129 434 -2123 468
rect -2169 396 -2123 434
rect -2169 362 -2163 396
rect -2129 362 -2123 396
rect -2169 324 -2123 362
rect -2169 290 -2163 324
rect -2129 290 -2123 324
rect -2169 252 -2123 290
rect -2169 218 -2163 252
rect -2129 218 -2123 252
rect -2169 180 -2123 218
rect -2169 146 -2163 180
rect -2129 146 -2123 180
rect -2169 109 -2123 146
rect -2021 972 -1975 1009
rect -2021 938 -2015 972
rect -1981 938 -1975 972
rect -2021 900 -1975 938
rect -2021 866 -2015 900
rect -1981 866 -1975 900
rect -2021 828 -1975 866
rect -2021 794 -2015 828
rect -1981 794 -1975 828
rect -2021 756 -1975 794
rect -2021 722 -2015 756
rect -1981 722 -1975 756
rect -2021 684 -1975 722
rect -2021 650 -2015 684
rect -1981 650 -1975 684
rect -2021 612 -1975 650
rect -2021 578 -2015 612
rect -1981 578 -1975 612
rect -2021 540 -1975 578
rect -2021 506 -2015 540
rect -1981 506 -1975 540
rect -2021 468 -1975 506
rect -2021 434 -2015 468
rect -1981 434 -1975 468
rect -2021 396 -1975 434
rect -2021 362 -2015 396
rect -1981 362 -1975 396
rect -2021 324 -1975 362
rect -2021 290 -2015 324
rect -1981 290 -1975 324
rect -2021 252 -1975 290
rect -2021 218 -2015 252
rect -1981 218 -1975 252
rect -2021 180 -1975 218
rect -2021 146 -2015 180
rect -1981 146 -1975 180
rect -2021 109 -1975 146
rect -1873 972 -1827 1009
rect -1873 938 -1867 972
rect -1833 938 -1827 972
rect -1873 900 -1827 938
rect -1873 866 -1867 900
rect -1833 866 -1827 900
rect -1873 828 -1827 866
rect -1873 794 -1867 828
rect -1833 794 -1827 828
rect -1873 756 -1827 794
rect -1873 722 -1867 756
rect -1833 722 -1827 756
rect -1873 684 -1827 722
rect -1873 650 -1867 684
rect -1833 650 -1827 684
rect -1873 612 -1827 650
rect -1873 578 -1867 612
rect -1833 578 -1827 612
rect -1873 540 -1827 578
rect -1873 506 -1867 540
rect -1833 506 -1827 540
rect -1873 468 -1827 506
rect -1873 434 -1867 468
rect -1833 434 -1827 468
rect -1873 396 -1827 434
rect -1873 362 -1867 396
rect -1833 362 -1827 396
rect -1873 324 -1827 362
rect -1873 290 -1867 324
rect -1833 290 -1827 324
rect -1873 252 -1827 290
rect -1873 218 -1867 252
rect -1833 218 -1827 252
rect -1873 180 -1827 218
rect -1873 146 -1867 180
rect -1833 146 -1827 180
rect -1873 109 -1827 146
rect -1725 972 -1679 1009
rect -1725 938 -1719 972
rect -1685 938 -1679 972
rect -1725 900 -1679 938
rect -1725 866 -1719 900
rect -1685 866 -1679 900
rect -1725 828 -1679 866
rect -1725 794 -1719 828
rect -1685 794 -1679 828
rect -1725 756 -1679 794
rect -1725 722 -1719 756
rect -1685 722 -1679 756
rect -1725 684 -1679 722
rect -1725 650 -1719 684
rect -1685 650 -1679 684
rect -1725 612 -1679 650
rect -1725 578 -1719 612
rect -1685 578 -1679 612
rect -1725 540 -1679 578
rect -1725 506 -1719 540
rect -1685 506 -1679 540
rect -1725 468 -1679 506
rect -1725 434 -1719 468
rect -1685 434 -1679 468
rect -1725 396 -1679 434
rect -1725 362 -1719 396
rect -1685 362 -1679 396
rect -1725 324 -1679 362
rect -1725 290 -1719 324
rect -1685 290 -1679 324
rect -1725 252 -1679 290
rect -1725 218 -1719 252
rect -1685 218 -1679 252
rect -1725 180 -1679 218
rect -1725 146 -1719 180
rect -1685 146 -1679 180
rect -1725 109 -1679 146
rect -1577 972 -1531 1009
rect -1577 938 -1571 972
rect -1537 938 -1531 972
rect -1577 900 -1531 938
rect -1577 866 -1571 900
rect -1537 866 -1531 900
rect -1577 828 -1531 866
rect -1577 794 -1571 828
rect -1537 794 -1531 828
rect -1577 756 -1531 794
rect -1577 722 -1571 756
rect -1537 722 -1531 756
rect -1577 684 -1531 722
rect -1577 650 -1571 684
rect -1537 650 -1531 684
rect -1577 612 -1531 650
rect -1577 578 -1571 612
rect -1537 578 -1531 612
rect -1577 540 -1531 578
rect -1577 506 -1571 540
rect -1537 506 -1531 540
rect -1577 468 -1531 506
rect -1577 434 -1571 468
rect -1537 434 -1531 468
rect -1577 396 -1531 434
rect -1577 362 -1571 396
rect -1537 362 -1531 396
rect -1577 324 -1531 362
rect -1577 290 -1571 324
rect -1537 290 -1531 324
rect -1577 252 -1531 290
rect -1577 218 -1571 252
rect -1537 218 -1531 252
rect -1577 180 -1531 218
rect -1577 146 -1571 180
rect -1537 146 -1531 180
rect -1577 109 -1531 146
rect -1429 972 -1383 1009
rect -1429 938 -1423 972
rect -1389 938 -1383 972
rect -1429 900 -1383 938
rect -1429 866 -1423 900
rect -1389 866 -1383 900
rect -1429 828 -1383 866
rect -1429 794 -1423 828
rect -1389 794 -1383 828
rect -1429 756 -1383 794
rect -1429 722 -1423 756
rect -1389 722 -1383 756
rect -1429 684 -1383 722
rect -1429 650 -1423 684
rect -1389 650 -1383 684
rect -1429 612 -1383 650
rect -1429 578 -1423 612
rect -1389 578 -1383 612
rect -1429 540 -1383 578
rect -1429 506 -1423 540
rect -1389 506 -1383 540
rect -1429 468 -1383 506
rect -1429 434 -1423 468
rect -1389 434 -1383 468
rect -1429 396 -1383 434
rect -1429 362 -1423 396
rect -1389 362 -1383 396
rect -1429 324 -1383 362
rect -1429 290 -1423 324
rect -1389 290 -1383 324
rect -1429 252 -1383 290
rect -1429 218 -1423 252
rect -1389 218 -1383 252
rect -1429 180 -1383 218
rect -1429 146 -1423 180
rect -1389 146 -1383 180
rect -1429 109 -1383 146
rect -1281 972 -1235 1009
rect -1281 938 -1275 972
rect -1241 938 -1235 972
rect -1281 900 -1235 938
rect -1281 866 -1275 900
rect -1241 866 -1235 900
rect -1281 828 -1235 866
rect -1281 794 -1275 828
rect -1241 794 -1235 828
rect -1281 756 -1235 794
rect -1281 722 -1275 756
rect -1241 722 -1235 756
rect -1281 684 -1235 722
rect -1281 650 -1275 684
rect -1241 650 -1235 684
rect -1281 612 -1235 650
rect -1281 578 -1275 612
rect -1241 578 -1235 612
rect -1281 540 -1235 578
rect -1281 506 -1275 540
rect -1241 506 -1235 540
rect -1281 468 -1235 506
rect -1281 434 -1275 468
rect -1241 434 -1235 468
rect -1281 396 -1235 434
rect -1281 362 -1275 396
rect -1241 362 -1235 396
rect -1281 324 -1235 362
rect -1281 290 -1275 324
rect -1241 290 -1235 324
rect -1281 252 -1235 290
rect -1281 218 -1275 252
rect -1241 218 -1235 252
rect -1281 180 -1235 218
rect -1281 146 -1275 180
rect -1241 146 -1235 180
rect -1281 109 -1235 146
rect -1133 972 -1087 1009
rect -1133 938 -1127 972
rect -1093 938 -1087 972
rect -1133 900 -1087 938
rect -1133 866 -1127 900
rect -1093 866 -1087 900
rect -1133 828 -1087 866
rect -1133 794 -1127 828
rect -1093 794 -1087 828
rect -1133 756 -1087 794
rect -1133 722 -1127 756
rect -1093 722 -1087 756
rect -1133 684 -1087 722
rect -1133 650 -1127 684
rect -1093 650 -1087 684
rect -1133 612 -1087 650
rect -1133 578 -1127 612
rect -1093 578 -1087 612
rect -1133 540 -1087 578
rect -1133 506 -1127 540
rect -1093 506 -1087 540
rect -1133 468 -1087 506
rect -1133 434 -1127 468
rect -1093 434 -1087 468
rect -1133 396 -1087 434
rect -1133 362 -1127 396
rect -1093 362 -1087 396
rect -1133 324 -1087 362
rect -1133 290 -1127 324
rect -1093 290 -1087 324
rect -1133 252 -1087 290
rect -1133 218 -1127 252
rect -1093 218 -1087 252
rect -1133 180 -1087 218
rect -1133 146 -1127 180
rect -1093 146 -1087 180
rect -1133 109 -1087 146
rect -985 972 -939 1009
rect -985 938 -979 972
rect -945 938 -939 972
rect -985 900 -939 938
rect -985 866 -979 900
rect -945 866 -939 900
rect -985 828 -939 866
rect -985 794 -979 828
rect -945 794 -939 828
rect -985 756 -939 794
rect -985 722 -979 756
rect -945 722 -939 756
rect -985 684 -939 722
rect -985 650 -979 684
rect -945 650 -939 684
rect -985 612 -939 650
rect -985 578 -979 612
rect -945 578 -939 612
rect -985 540 -939 578
rect -985 506 -979 540
rect -945 506 -939 540
rect -985 468 -939 506
rect -985 434 -979 468
rect -945 434 -939 468
rect -985 396 -939 434
rect -985 362 -979 396
rect -945 362 -939 396
rect -985 324 -939 362
rect -985 290 -979 324
rect -945 290 -939 324
rect -985 252 -939 290
rect -985 218 -979 252
rect -945 218 -939 252
rect -985 180 -939 218
rect -985 146 -979 180
rect -945 146 -939 180
rect -985 109 -939 146
rect -837 972 -791 1009
rect -837 938 -831 972
rect -797 938 -791 972
rect -837 900 -791 938
rect -837 866 -831 900
rect -797 866 -791 900
rect -837 828 -791 866
rect -837 794 -831 828
rect -797 794 -791 828
rect -837 756 -791 794
rect -837 722 -831 756
rect -797 722 -791 756
rect -837 684 -791 722
rect -837 650 -831 684
rect -797 650 -791 684
rect -837 612 -791 650
rect -837 578 -831 612
rect -797 578 -791 612
rect -837 540 -791 578
rect -837 506 -831 540
rect -797 506 -791 540
rect -837 468 -791 506
rect -837 434 -831 468
rect -797 434 -791 468
rect -837 396 -791 434
rect -837 362 -831 396
rect -797 362 -791 396
rect -837 324 -791 362
rect -837 290 -831 324
rect -797 290 -791 324
rect -837 252 -791 290
rect -837 218 -831 252
rect -797 218 -791 252
rect -837 180 -791 218
rect -837 146 -831 180
rect -797 146 -791 180
rect -837 109 -791 146
rect -689 972 -643 1009
rect -689 938 -683 972
rect -649 938 -643 972
rect -689 900 -643 938
rect -689 866 -683 900
rect -649 866 -643 900
rect -689 828 -643 866
rect -689 794 -683 828
rect -649 794 -643 828
rect -689 756 -643 794
rect -689 722 -683 756
rect -649 722 -643 756
rect -689 684 -643 722
rect -689 650 -683 684
rect -649 650 -643 684
rect -689 612 -643 650
rect -689 578 -683 612
rect -649 578 -643 612
rect -689 540 -643 578
rect -689 506 -683 540
rect -649 506 -643 540
rect -689 468 -643 506
rect -689 434 -683 468
rect -649 434 -643 468
rect -689 396 -643 434
rect -689 362 -683 396
rect -649 362 -643 396
rect -689 324 -643 362
rect -689 290 -683 324
rect -649 290 -643 324
rect -689 252 -643 290
rect -689 218 -683 252
rect -649 218 -643 252
rect -689 180 -643 218
rect -689 146 -683 180
rect -649 146 -643 180
rect -689 109 -643 146
rect -541 972 -495 1009
rect -541 938 -535 972
rect -501 938 -495 972
rect -541 900 -495 938
rect -541 866 -535 900
rect -501 866 -495 900
rect -541 828 -495 866
rect -541 794 -535 828
rect -501 794 -495 828
rect -541 756 -495 794
rect -541 722 -535 756
rect -501 722 -495 756
rect -541 684 -495 722
rect -541 650 -535 684
rect -501 650 -495 684
rect -541 612 -495 650
rect -541 578 -535 612
rect -501 578 -495 612
rect -541 540 -495 578
rect -541 506 -535 540
rect -501 506 -495 540
rect -541 468 -495 506
rect -541 434 -535 468
rect -501 434 -495 468
rect -541 396 -495 434
rect -541 362 -535 396
rect -501 362 -495 396
rect -541 324 -495 362
rect -541 290 -535 324
rect -501 290 -495 324
rect -541 252 -495 290
rect -541 218 -535 252
rect -501 218 -495 252
rect -541 180 -495 218
rect -541 146 -535 180
rect -501 146 -495 180
rect -541 109 -495 146
rect -393 972 -347 1009
rect -393 938 -387 972
rect -353 938 -347 972
rect -393 900 -347 938
rect -393 866 -387 900
rect -353 866 -347 900
rect -393 828 -347 866
rect -393 794 -387 828
rect -353 794 -347 828
rect -393 756 -347 794
rect -393 722 -387 756
rect -353 722 -347 756
rect -393 684 -347 722
rect -393 650 -387 684
rect -353 650 -347 684
rect -393 612 -347 650
rect -393 578 -387 612
rect -353 578 -347 612
rect -393 540 -347 578
rect -393 506 -387 540
rect -353 506 -347 540
rect -393 468 -347 506
rect -393 434 -387 468
rect -353 434 -347 468
rect -393 396 -347 434
rect -393 362 -387 396
rect -353 362 -347 396
rect -393 324 -347 362
rect -393 290 -387 324
rect -353 290 -347 324
rect -393 252 -347 290
rect -393 218 -387 252
rect -353 218 -347 252
rect -393 180 -347 218
rect -393 146 -387 180
rect -353 146 -347 180
rect -393 109 -347 146
rect -245 972 -199 1009
rect -245 938 -239 972
rect -205 938 -199 972
rect -245 900 -199 938
rect -245 866 -239 900
rect -205 866 -199 900
rect -245 828 -199 866
rect -245 794 -239 828
rect -205 794 -199 828
rect -245 756 -199 794
rect -245 722 -239 756
rect -205 722 -199 756
rect -245 684 -199 722
rect -245 650 -239 684
rect -205 650 -199 684
rect -245 612 -199 650
rect -245 578 -239 612
rect -205 578 -199 612
rect -245 540 -199 578
rect -245 506 -239 540
rect -205 506 -199 540
rect -245 468 -199 506
rect -245 434 -239 468
rect -205 434 -199 468
rect -245 396 -199 434
rect -245 362 -239 396
rect -205 362 -199 396
rect -245 324 -199 362
rect -245 290 -239 324
rect -205 290 -199 324
rect -245 252 -199 290
rect -245 218 -239 252
rect -205 218 -199 252
rect -245 180 -199 218
rect -245 146 -239 180
rect -205 146 -199 180
rect -245 109 -199 146
rect -97 972 -51 1009
rect -97 938 -91 972
rect -57 938 -51 972
rect -97 900 -51 938
rect -97 866 -91 900
rect -57 866 -51 900
rect -97 828 -51 866
rect -97 794 -91 828
rect -57 794 -51 828
rect -97 756 -51 794
rect -97 722 -91 756
rect -57 722 -51 756
rect -97 684 -51 722
rect -97 650 -91 684
rect -57 650 -51 684
rect -97 612 -51 650
rect -97 578 -91 612
rect -57 578 -51 612
rect -97 540 -51 578
rect -97 506 -91 540
rect -57 506 -51 540
rect -97 468 -51 506
rect -97 434 -91 468
rect -57 434 -51 468
rect -97 396 -51 434
rect -97 362 -91 396
rect -57 362 -51 396
rect -97 324 -51 362
rect -97 290 -91 324
rect -57 290 -51 324
rect -97 252 -51 290
rect -97 218 -91 252
rect -57 218 -51 252
rect -97 180 -51 218
rect -97 146 -91 180
rect -57 146 -51 180
rect -97 109 -51 146
rect 51 972 97 1009
rect 51 938 57 972
rect 91 938 97 972
rect 51 900 97 938
rect 51 866 57 900
rect 91 866 97 900
rect 51 828 97 866
rect 51 794 57 828
rect 91 794 97 828
rect 51 756 97 794
rect 51 722 57 756
rect 91 722 97 756
rect 51 684 97 722
rect 51 650 57 684
rect 91 650 97 684
rect 51 612 97 650
rect 51 578 57 612
rect 91 578 97 612
rect 51 540 97 578
rect 51 506 57 540
rect 91 506 97 540
rect 51 468 97 506
rect 51 434 57 468
rect 91 434 97 468
rect 51 396 97 434
rect 51 362 57 396
rect 91 362 97 396
rect 51 324 97 362
rect 51 290 57 324
rect 91 290 97 324
rect 51 252 97 290
rect 51 218 57 252
rect 91 218 97 252
rect 51 180 97 218
rect 51 146 57 180
rect 91 146 97 180
rect 51 109 97 146
rect 199 972 245 1009
rect 199 938 205 972
rect 239 938 245 972
rect 199 900 245 938
rect 199 866 205 900
rect 239 866 245 900
rect 199 828 245 866
rect 199 794 205 828
rect 239 794 245 828
rect 199 756 245 794
rect 199 722 205 756
rect 239 722 245 756
rect 199 684 245 722
rect 199 650 205 684
rect 239 650 245 684
rect 199 612 245 650
rect 199 578 205 612
rect 239 578 245 612
rect 199 540 245 578
rect 199 506 205 540
rect 239 506 245 540
rect 199 468 245 506
rect 199 434 205 468
rect 239 434 245 468
rect 199 396 245 434
rect 199 362 205 396
rect 239 362 245 396
rect 199 324 245 362
rect 199 290 205 324
rect 239 290 245 324
rect 199 252 245 290
rect 199 218 205 252
rect 239 218 245 252
rect 199 180 245 218
rect 199 146 205 180
rect 239 146 245 180
rect 199 109 245 146
rect 347 972 393 1009
rect 347 938 353 972
rect 387 938 393 972
rect 347 900 393 938
rect 347 866 353 900
rect 387 866 393 900
rect 347 828 393 866
rect 347 794 353 828
rect 387 794 393 828
rect 347 756 393 794
rect 347 722 353 756
rect 387 722 393 756
rect 347 684 393 722
rect 347 650 353 684
rect 387 650 393 684
rect 347 612 393 650
rect 347 578 353 612
rect 387 578 393 612
rect 347 540 393 578
rect 347 506 353 540
rect 387 506 393 540
rect 347 468 393 506
rect 347 434 353 468
rect 387 434 393 468
rect 347 396 393 434
rect 347 362 353 396
rect 387 362 393 396
rect 347 324 393 362
rect 347 290 353 324
rect 387 290 393 324
rect 347 252 393 290
rect 347 218 353 252
rect 387 218 393 252
rect 347 180 393 218
rect 347 146 353 180
rect 387 146 393 180
rect 347 109 393 146
rect 495 972 541 1009
rect 495 938 501 972
rect 535 938 541 972
rect 495 900 541 938
rect 495 866 501 900
rect 535 866 541 900
rect 495 828 541 866
rect 495 794 501 828
rect 535 794 541 828
rect 495 756 541 794
rect 495 722 501 756
rect 535 722 541 756
rect 495 684 541 722
rect 495 650 501 684
rect 535 650 541 684
rect 495 612 541 650
rect 495 578 501 612
rect 535 578 541 612
rect 495 540 541 578
rect 495 506 501 540
rect 535 506 541 540
rect 495 468 541 506
rect 495 434 501 468
rect 535 434 541 468
rect 495 396 541 434
rect 495 362 501 396
rect 535 362 541 396
rect 495 324 541 362
rect 495 290 501 324
rect 535 290 541 324
rect 495 252 541 290
rect 495 218 501 252
rect 535 218 541 252
rect 495 180 541 218
rect 495 146 501 180
rect 535 146 541 180
rect 495 109 541 146
rect 643 972 689 1009
rect 643 938 649 972
rect 683 938 689 972
rect 643 900 689 938
rect 643 866 649 900
rect 683 866 689 900
rect 643 828 689 866
rect 643 794 649 828
rect 683 794 689 828
rect 643 756 689 794
rect 643 722 649 756
rect 683 722 689 756
rect 643 684 689 722
rect 643 650 649 684
rect 683 650 689 684
rect 643 612 689 650
rect 643 578 649 612
rect 683 578 689 612
rect 643 540 689 578
rect 643 506 649 540
rect 683 506 689 540
rect 643 468 689 506
rect 643 434 649 468
rect 683 434 689 468
rect 643 396 689 434
rect 643 362 649 396
rect 683 362 689 396
rect 643 324 689 362
rect 643 290 649 324
rect 683 290 689 324
rect 643 252 689 290
rect 643 218 649 252
rect 683 218 689 252
rect 643 180 689 218
rect 643 146 649 180
rect 683 146 689 180
rect 643 109 689 146
rect 791 972 837 1009
rect 791 938 797 972
rect 831 938 837 972
rect 791 900 837 938
rect 791 866 797 900
rect 831 866 837 900
rect 791 828 837 866
rect 791 794 797 828
rect 831 794 837 828
rect 791 756 837 794
rect 791 722 797 756
rect 831 722 837 756
rect 791 684 837 722
rect 791 650 797 684
rect 831 650 837 684
rect 791 612 837 650
rect 791 578 797 612
rect 831 578 837 612
rect 791 540 837 578
rect 791 506 797 540
rect 831 506 837 540
rect 791 468 837 506
rect 791 434 797 468
rect 831 434 837 468
rect 791 396 837 434
rect 791 362 797 396
rect 831 362 837 396
rect 791 324 837 362
rect 791 290 797 324
rect 831 290 837 324
rect 791 252 837 290
rect 791 218 797 252
rect 831 218 837 252
rect 791 180 837 218
rect 791 146 797 180
rect 831 146 837 180
rect 791 109 837 146
rect 939 972 985 1009
rect 939 938 945 972
rect 979 938 985 972
rect 939 900 985 938
rect 939 866 945 900
rect 979 866 985 900
rect 939 828 985 866
rect 939 794 945 828
rect 979 794 985 828
rect 939 756 985 794
rect 939 722 945 756
rect 979 722 985 756
rect 939 684 985 722
rect 939 650 945 684
rect 979 650 985 684
rect 939 612 985 650
rect 939 578 945 612
rect 979 578 985 612
rect 939 540 985 578
rect 939 506 945 540
rect 979 506 985 540
rect 939 468 985 506
rect 939 434 945 468
rect 979 434 985 468
rect 939 396 985 434
rect 939 362 945 396
rect 979 362 985 396
rect 939 324 985 362
rect 939 290 945 324
rect 979 290 985 324
rect 939 252 985 290
rect 939 218 945 252
rect 979 218 985 252
rect 939 180 985 218
rect 939 146 945 180
rect 979 146 985 180
rect 939 109 985 146
rect 1087 972 1133 1009
rect 1087 938 1093 972
rect 1127 938 1133 972
rect 1087 900 1133 938
rect 1087 866 1093 900
rect 1127 866 1133 900
rect 1087 828 1133 866
rect 1087 794 1093 828
rect 1127 794 1133 828
rect 1087 756 1133 794
rect 1087 722 1093 756
rect 1127 722 1133 756
rect 1087 684 1133 722
rect 1087 650 1093 684
rect 1127 650 1133 684
rect 1087 612 1133 650
rect 1087 578 1093 612
rect 1127 578 1133 612
rect 1087 540 1133 578
rect 1087 506 1093 540
rect 1127 506 1133 540
rect 1087 468 1133 506
rect 1087 434 1093 468
rect 1127 434 1133 468
rect 1087 396 1133 434
rect 1087 362 1093 396
rect 1127 362 1133 396
rect 1087 324 1133 362
rect 1087 290 1093 324
rect 1127 290 1133 324
rect 1087 252 1133 290
rect 1087 218 1093 252
rect 1127 218 1133 252
rect 1087 180 1133 218
rect 1087 146 1093 180
rect 1127 146 1133 180
rect 1087 109 1133 146
rect 1235 972 1281 1009
rect 1235 938 1241 972
rect 1275 938 1281 972
rect 1235 900 1281 938
rect 1235 866 1241 900
rect 1275 866 1281 900
rect 1235 828 1281 866
rect 1235 794 1241 828
rect 1275 794 1281 828
rect 1235 756 1281 794
rect 1235 722 1241 756
rect 1275 722 1281 756
rect 1235 684 1281 722
rect 1235 650 1241 684
rect 1275 650 1281 684
rect 1235 612 1281 650
rect 1235 578 1241 612
rect 1275 578 1281 612
rect 1235 540 1281 578
rect 1235 506 1241 540
rect 1275 506 1281 540
rect 1235 468 1281 506
rect 1235 434 1241 468
rect 1275 434 1281 468
rect 1235 396 1281 434
rect 1235 362 1241 396
rect 1275 362 1281 396
rect 1235 324 1281 362
rect 1235 290 1241 324
rect 1275 290 1281 324
rect 1235 252 1281 290
rect 1235 218 1241 252
rect 1275 218 1281 252
rect 1235 180 1281 218
rect 1235 146 1241 180
rect 1275 146 1281 180
rect 1235 109 1281 146
rect 1383 972 1429 1009
rect 1383 938 1389 972
rect 1423 938 1429 972
rect 1383 900 1429 938
rect 1383 866 1389 900
rect 1423 866 1429 900
rect 1383 828 1429 866
rect 1383 794 1389 828
rect 1423 794 1429 828
rect 1383 756 1429 794
rect 1383 722 1389 756
rect 1423 722 1429 756
rect 1383 684 1429 722
rect 1383 650 1389 684
rect 1423 650 1429 684
rect 1383 612 1429 650
rect 1383 578 1389 612
rect 1423 578 1429 612
rect 1383 540 1429 578
rect 1383 506 1389 540
rect 1423 506 1429 540
rect 1383 468 1429 506
rect 1383 434 1389 468
rect 1423 434 1429 468
rect 1383 396 1429 434
rect 1383 362 1389 396
rect 1423 362 1429 396
rect 1383 324 1429 362
rect 1383 290 1389 324
rect 1423 290 1429 324
rect 1383 252 1429 290
rect 1383 218 1389 252
rect 1423 218 1429 252
rect 1383 180 1429 218
rect 1383 146 1389 180
rect 1423 146 1429 180
rect 1383 109 1429 146
rect 1531 972 1577 1009
rect 1531 938 1537 972
rect 1571 938 1577 972
rect 1531 900 1577 938
rect 1531 866 1537 900
rect 1571 866 1577 900
rect 1531 828 1577 866
rect 1531 794 1537 828
rect 1571 794 1577 828
rect 1531 756 1577 794
rect 1531 722 1537 756
rect 1571 722 1577 756
rect 1531 684 1577 722
rect 1531 650 1537 684
rect 1571 650 1577 684
rect 1531 612 1577 650
rect 1531 578 1537 612
rect 1571 578 1577 612
rect 1531 540 1577 578
rect 1531 506 1537 540
rect 1571 506 1577 540
rect 1531 468 1577 506
rect 1531 434 1537 468
rect 1571 434 1577 468
rect 1531 396 1577 434
rect 1531 362 1537 396
rect 1571 362 1577 396
rect 1531 324 1577 362
rect 1531 290 1537 324
rect 1571 290 1577 324
rect 1531 252 1577 290
rect 1531 218 1537 252
rect 1571 218 1577 252
rect 1531 180 1577 218
rect 1531 146 1537 180
rect 1571 146 1577 180
rect 1531 109 1577 146
rect 1679 972 1725 1009
rect 1679 938 1685 972
rect 1719 938 1725 972
rect 1679 900 1725 938
rect 1679 866 1685 900
rect 1719 866 1725 900
rect 1679 828 1725 866
rect 1679 794 1685 828
rect 1719 794 1725 828
rect 1679 756 1725 794
rect 1679 722 1685 756
rect 1719 722 1725 756
rect 1679 684 1725 722
rect 1679 650 1685 684
rect 1719 650 1725 684
rect 1679 612 1725 650
rect 1679 578 1685 612
rect 1719 578 1725 612
rect 1679 540 1725 578
rect 1679 506 1685 540
rect 1719 506 1725 540
rect 1679 468 1725 506
rect 1679 434 1685 468
rect 1719 434 1725 468
rect 1679 396 1725 434
rect 1679 362 1685 396
rect 1719 362 1725 396
rect 1679 324 1725 362
rect 1679 290 1685 324
rect 1719 290 1725 324
rect 1679 252 1725 290
rect 1679 218 1685 252
rect 1719 218 1725 252
rect 1679 180 1725 218
rect 1679 146 1685 180
rect 1719 146 1725 180
rect 1679 109 1725 146
rect 1827 972 1873 1009
rect 1827 938 1833 972
rect 1867 938 1873 972
rect 1827 900 1873 938
rect 1827 866 1833 900
rect 1867 866 1873 900
rect 1827 828 1873 866
rect 1827 794 1833 828
rect 1867 794 1873 828
rect 1827 756 1873 794
rect 1827 722 1833 756
rect 1867 722 1873 756
rect 1827 684 1873 722
rect 1827 650 1833 684
rect 1867 650 1873 684
rect 1827 612 1873 650
rect 1827 578 1833 612
rect 1867 578 1873 612
rect 1827 540 1873 578
rect 1827 506 1833 540
rect 1867 506 1873 540
rect 1827 468 1873 506
rect 1827 434 1833 468
rect 1867 434 1873 468
rect 1827 396 1873 434
rect 1827 362 1833 396
rect 1867 362 1873 396
rect 1827 324 1873 362
rect 1827 290 1833 324
rect 1867 290 1873 324
rect 1827 252 1873 290
rect 1827 218 1833 252
rect 1867 218 1873 252
rect 1827 180 1873 218
rect 1827 146 1833 180
rect 1867 146 1873 180
rect 1827 109 1873 146
rect 1975 972 2021 1009
rect 1975 938 1981 972
rect 2015 938 2021 972
rect 1975 900 2021 938
rect 1975 866 1981 900
rect 2015 866 2021 900
rect 1975 828 2021 866
rect 1975 794 1981 828
rect 2015 794 2021 828
rect 1975 756 2021 794
rect 1975 722 1981 756
rect 2015 722 2021 756
rect 1975 684 2021 722
rect 1975 650 1981 684
rect 2015 650 2021 684
rect 1975 612 2021 650
rect 1975 578 1981 612
rect 2015 578 2021 612
rect 1975 540 2021 578
rect 1975 506 1981 540
rect 2015 506 2021 540
rect 1975 468 2021 506
rect 1975 434 1981 468
rect 2015 434 2021 468
rect 1975 396 2021 434
rect 1975 362 1981 396
rect 2015 362 2021 396
rect 1975 324 2021 362
rect 1975 290 1981 324
rect 2015 290 2021 324
rect 1975 252 2021 290
rect 1975 218 1981 252
rect 2015 218 2021 252
rect 1975 180 2021 218
rect 1975 146 1981 180
rect 2015 146 2021 180
rect 1975 109 2021 146
rect 2123 972 2169 1009
rect 2123 938 2129 972
rect 2163 938 2169 972
rect 2123 900 2169 938
rect 2123 866 2129 900
rect 2163 866 2169 900
rect 2123 828 2169 866
rect 2123 794 2129 828
rect 2163 794 2169 828
rect 2123 756 2169 794
rect 2123 722 2129 756
rect 2163 722 2169 756
rect 2123 684 2169 722
rect 2123 650 2129 684
rect 2163 650 2169 684
rect 2123 612 2169 650
rect 2123 578 2129 612
rect 2163 578 2169 612
rect 2123 540 2169 578
rect 2123 506 2129 540
rect 2163 506 2169 540
rect 2123 468 2169 506
rect 2123 434 2129 468
rect 2163 434 2169 468
rect 2123 396 2169 434
rect 2123 362 2129 396
rect 2163 362 2169 396
rect 2123 324 2169 362
rect 2123 290 2129 324
rect 2163 290 2169 324
rect 2123 252 2169 290
rect 2123 218 2129 252
rect 2163 218 2169 252
rect 2123 180 2169 218
rect 2123 146 2129 180
rect 2163 146 2169 180
rect 2123 109 2169 146
rect 2271 972 2317 1009
rect 2271 938 2277 972
rect 2311 938 2317 972
rect 2271 900 2317 938
rect 2271 866 2277 900
rect 2311 866 2317 900
rect 2271 828 2317 866
rect 2271 794 2277 828
rect 2311 794 2317 828
rect 2271 756 2317 794
rect 2271 722 2277 756
rect 2311 722 2317 756
rect 2271 684 2317 722
rect 2271 650 2277 684
rect 2311 650 2317 684
rect 2271 612 2317 650
rect 2271 578 2277 612
rect 2311 578 2317 612
rect 2271 540 2317 578
rect 2271 506 2277 540
rect 2311 506 2317 540
rect 2271 468 2317 506
rect 2271 434 2277 468
rect 2311 434 2317 468
rect 2271 396 2317 434
rect 2271 362 2277 396
rect 2311 362 2317 396
rect 2271 324 2317 362
rect 2271 290 2277 324
rect 2311 290 2317 324
rect 2271 252 2317 290
rect 2271 218 2277 252
rect 2311 218 2317 252
rect 2271 180 2317 218
rect 2271 146 2277 180
rect 2311 146 2317 180
rect 2271 109 2317 146
rect 2419 972 2465 1009
rect 2419 938 2425 972
rect 2459 938 2465 972
rect 2419 900 2465 938
rect 2419 866 2425 900
rect 2459 866 2465 900
rect 2419 828 2465 866
rect 2419 794 2425 828
rect 2459 794 2465 828
rect 2419 756 2465 794
rect 2419 722 2425 756
rect 2459 722 2465 756
rect 2419 684 2465 722
rect 2419 650 2425 684
rect 2459 650 2465 684
rect 2419 612 2465 650
rect 2419 578 2425 612
rect 2459 578 2465 612
rect 2419 540 2465 578
rect 2419 506 2425 540
rect 2459 506 2465 540
rect 2419 468 2465 506
rect 2419 434 2425 468
rect 2459 434 2465 468
rect 2419 396 2465 434
rect 2419 362 2425 396
rect 2459 362 2465 396
rect 2419 324 2465 362
rect 2419 290 2425 324
rect 2459 290 2465 324
rect 2419 252 2465 290
rect 2419 218 2425 252
rect 2459 218 2465 252
rect 2419 180 2465 218
rect 2419 146 2425 180
rect 2459 146 2465 180
rect 2419 109 2465 146
rect 2567 972 2613 1009
rect 2567 938 2573 972
rect 2607 938 2613 972
rect 2567 900 2613 938
rect 2567 866 2573 900
rect 2607 866 2613 900
rect 2567 828 2613 866
rect 2567 794 2573 828
rect 2607 794 2613 828
rect 2567 756 2613 794
rect 2567 722 2573 756
rect 2607 722 2613 756
rect 2567 684 2613 722
rect 2567 650 2573 684
rect 2607 650 2613 684
rect 2567 612 2613 650
rect 2567 578 2573 612
rect 2607 578 2613 612
rect 2567 540 2613 578
rect 2567 506 2573 540
rect 2607 506 2613 540
rect 2567 468 2613 506
rect 2567 434 2573 468
rect 2607 434 2613 468
rect 2567 396 2613 434
rect 2567 362 2573 396
rect 2607 362 2613 396
rect 2567 324 2613 362
rect 2567 290 2573 324
rect 2607 290 2613 324
rect 2567 252 2613 290
rect 2567 218 2573 252
rect 2607 218 2613 252
rect 2567 180 2613 218
rect 2567 146 2573 180
rect 2607 146 2613 180
rect 2567 109 2613 146
rect 2715 972 2761 1009
rect 2715 938 2721 972
rect 2755 938 2761 972
rect 2715 900 2761 938
rect 2715 866 2721 900
rect 2755 866 2761 900
rect 2715 828 2761 866
rect 2715 794 2721 828
rect 2755 794 2761 828
rect 2715 756 2761 794
rect 2715 722 2721 756
rect 2755 722 2761 756
rect 2715 684 2761 722
rect 2715 650 2721 684
rect 2755 650 2761 684
rect 2715 612 2761 650
rect 2715 578 2721 612
rect 2755 578 2761 612
rect 2715 540 2761 578
rect 2715 506 2721 540
rect 2755 506 2761 540
rect 2715 468 2761 506
rect 2715 434 2721 468
rect 2755 434 2761 468
rect 2715 396 2761 434
rect 2715 362 2721 396
rect 2755 362 2761 396
rect 2715 324 2761 362
rect 2715 290 2721 324
rect 2755 290 2761 324
rect 2715 252 2761 290
rect 2715 218 2721 252
rect 2755 218 2761 252
rect 2715 180 2761 218
rect 2715 146 2721 180
rect 2755 146 2761 180
rect 2715 109 2761 146
rect 2863 972 2909 1009
rect 2863 938 2869 972
rect 2903 938 2909 972
rect 2863 900 2909 938
rect 2863 866 2869 900
rect 2903 866 2909 900
rect 2863 828 2909 866
rect 2863 794 2869 828
rect 2903 794 2909 828
rect 2863 756 2909 794
rect 2863 722 2869 756
rect 2903 722 2909 756
rect 2863 684 2909 722
rect 2863 650 2869 684
rect 2903 650 2909 684
rect 2863 612 2909 650
rect 2863 578 2869 612
rect 2903 578 2909 612
rect 2863 540 2909 578
rect 2863 506 2869 540
rect 2903 506 2909 540
rect 2863 468 2909 506
rect 2863 434 2869 468
rect 2903 434 2909 468
rect 2863 396 2909 434
rect 2863 362 2869 396
rect 2903 362 2909 396
rect 2863 324 2909 362
rect 2863 290 2869 324
rect 2903 290 2909 324
rect 2863 252 2909 290
rect 2863 218 2869 252
rect 2903 218 2909 252
rect 2863 180 2909 218
rect 2863 146 2869 180
rect 2903 146 2909 180
rect 2863 109 2909 146
rect 3011 972 3057 1009
rect 3011 938 3017 972
rect 3051 938 3057 972
rect 3011 900 3057 938
rect 3011 866 3017 900
rect 3051 866 3057 900
rect 3011 828 3057 866
rect 3011 794 3017 828
rect 3051 794 3057 828
rect 3011 756 3057 794
rect 3011 722 3017 756
rect 3051 722 3057 756
rect 3011 684 3057 722
rect 3011 650 3017 684
rect 3051 650 3057 684
rect 3011 612 3057 650
rect 3011 578 3017 612
rect 3051 578 3057 612
rect 3011 540 3057 578
rect 3011 506 3017 540
rect 3051 506 3057 540
rect 3011 468 3057 506
rect 3011 434 3017 468
rect 3051 434 3057 468
rect 3011 396 3057 434
rect 3011 362 3017 396
rect 3051 362 3057 396
rect 3011 324 3057 362
rect 3011 290 3017 324
rect 3051 290 3057 324
rect 3011 252 3057 290
rect 3011 218 3017 252
rect 3051 218 3057 252
rect 3011 180 3057 218
rect 3011 146 3017 180
rect 3051 146 3057 180
rect 3011 109 3057 146
rect 3159 972 3205 1009
rect 3159 938 3165 972
rect 3199 938 3205 972
rect 3159 900 3205 938
rect 3159 866 3165 900
rect 3199 866 3205 900
rect 3159 828 3205 866
rect 3159 794 3165 828
rect 3199 794 3205 828
rect 3159 756 3205 794
rect 3159 722 3165 756
rect 3199 722 3205 756
rect 3159 684 3205 722
rect 3159 650 3165 684
rect 3199 650 3205 684
rect 3159 612 3205 650
rect 3159 578 3165 612
rect 3199 578 3205 612
rect 3159 540 3205 578
rect 3159 506 3165 540
rect 3199 506 3205 540
rect 3159 468 3205 506
rect 3159 434 3165 468
rect 3199 434 3205 468
rect 3159 396 3205 434
rect 3159 362 3165 396
rect 3199 362 3205 396
rect 3159 324 3205 362
rect 3159 290 3165 324
rect 3199 290 3205 324
rect 3159 252 3205 290
rect 3159 218 3165 252
rect 3199 218 3205 252
rect 3159 180 3205 218
rect 3159 146 3165 180
rect 3199 146 3205 180
rect 3159 109 3205 146
rect 3307 972 3353 1009
rect 3307 938 3313 972
rect 3347 938 3353 972
rect 3307 900 3353 938
rect 3307 866 3313 900
rect 3347 866 3353 900
rect 3307 828 3353 866
rect 3307 794 3313 828
rect 3347 794 3353 828
rect 3307 756 3353 794
rect 3307 722 3313 756
rect 3347 722 3353 756
rect 3307 684 3353 722
rect 3307 650 3313 684
rect 3347 650 3353 684
rect 3307 612 3353 650
rect 3307 578 3313 612
rect 3347 578 3353 612
rect 3307 540 3353 578
rect 3307 506 3313 540
rect 3347 506 3353 540
rect 3307 468 3353 506
rect 3307 434 3313 468
rect 3347 434 3353 468
rect 3307 396 3353 434
rect 3307 362 3313 396
rect 3347 362 3353 396
rect 3307 324 3353 362
rect 3307 290 3313 324
rect 3347 290 3353 324
rect 3307 252 3353 290
rect 3307 218 3313 252
rect 3347 218 3353 252
rect 3307 180 3353 218
rect 3307 146 3313 180
rect 3347 146 3353 180
rect 3307 109 3353 146
rect 3455 972 3501 1009
rect 3455 938 3461 972
rect 3495 938 3501 972
rect 3455 900 3501 938
rect 3455 866 3461 900
rect 3495 866 3501 900
rect 3455 828 3501 866
rect 3455 794 3461 828
rect 3495 794 3501 828
rect 3455 756 3501 794
rect 3455 722 3461 756
rect 3495 722 3501 756
rect 3455 684 3501 722
rect 3455 650 3461 684
rect 3495 650 3501 684
rect 3455 612 3501 650
rect 3455 578 3461 612
rect 3495 578 3501 612
rect 3455 540 3501 578
rect 3455 506 3461 540
rect 3495 506 3501 540
rect 3455 468 3501 506
rect 3455 434 3461 468
rect 3495 434 3501 468
rect 3455 396 3501 434
rect 3455 362 3461 396
rect 3495 362 3501 396
rect 3455 324 3501 362
rect 3455 290 3461 324
rect 3495 290 3501 324
rect 3455 252 3501 290
rect 3455 218 3461 252
rect 3495 218 3501 252
rect 3455 180 3501 218
rect 3455 146 3461 180
rect 3495 146 3501 180
rect 3455 109 3501 146
rect 3603 972 3649 1009
rect 3603 938 3609 972
rect 3643 938 3649 972
rect 3603 900 3649 938
rect 3603 866 3609 900
rect 3643 866 3649 900
rect 3603 828 3649 866
rect 3603 794 3609 828
rect 3643 794 3649 828
rect 3603 756 3649 794
rect 3603 722 3609 756
rect 3643 722 3649 756
rect 3603 684 3649 722
rect 3603 650 3609 684
rect 3643 650 3649 684
rect 3603 612 3649 650
rect 3603 578 3609 612
rect 3643 578 3649 612
rect 3603 540 3649 578
rect 3603 506 3609 540
rect 3643 506 3649 540
rect 3603 468 3649 506
rect 3603 434 3609 468
rect 3643 434 3649 468
rect 3603 396 3649 434
rect 3603 362 3609 396
rect 3643 362 3649 396
rect 3603 324 3649 362
rect 3603 290 3609 324
rect 3643 290 3649 324
rect 3603 252 3649 290
rect 3603 218 3609 252
rect 3643 218 3649 252
rect 3603 180 3649 218
rect 3603 146 3609 180
rect 3643 146 3649 180
rect 3603 109 3649 146
rect 3751 972 3797 1009
rect 3751 938 3757 972
rect 3791 938 3797 972
rect 3751 900 3797 938
rect 3751 866 3757 900
rect 3791 866 3797 900
rect 3751 828 3797 866
rect 3751 794 3757 828
rect 3791 794 3797 828
rect 3751 756 3797 794
rect 3751 722 3757 756
rect 3791 722 3797 756
rect 3751 684 3797 722
rect 3751 650 3757 684
rect 3791 650 3797 684
rect 3751 612 3797 650
rect 3751 578 3757 612
rect 3791 578 3797 612
rect 3751 540 3797 578
rect 3751 506 3757 540
rect 3791 506 3797 540
rect 3751 468 3797 506
rect 3751 434 3757 468
rect 3791 434 3797 468
rect 3751 396 3797 434
rect 3751 362 3757 396
rect 3791 362 3797 396
rect 3751 324 3797 362
rect 3751 290 3757 324
rect 3791 290 3797 324
rect 3751 252 3797 290
rect 3751 218 3757 252
rect 3791 218 3797 252
rect 3751 180 3797 218
rect 3751 146 3757 180
rect 3791 146 3797 180
rect 3751 109 3797 146
rect 3899 972 3945 1009
rect 3899 938 3905 972
rect 3939 938 3945 972
rect 3899 900 3945 938
rect 3899 866 3905 900
rect 3939 866 3945 900
rect 3899 828 3945 866
rect 3899 794 3905 828
rect 3939 794 3945 828
rect 3899 756 3945 794
rect 3899 722 3905 756
rect 3939 722 3945 756
rect 3899 684 3945 722
rect 3899 650 3905 684
rect 3939 650 3945 684
rect 3899 612 3945 650
rect 3899 578 3905 612
rect 3939 578 3945 612
rect 3899 540 3945 578
rect 3899 506 3905 540
rect 3939 506 3945 540
rect 3899 468 3945 506
rect 3899 434 3905 468
rect 3939 434 3945 468
rect 3899 396 3945 434
rect 3899 362 3905 396
rect 3939 362 3945 396
rect 3899 324 3945 362
rect 3899 290 3905 324
rect 3939 290 3945 324
rect 3899 252 3945 290
rect 3899 218 3905 252
rect 3939 218 3945 252
rect 3899 180 3945 218
rect 3899 146 3905 180
rect 3939 146 3945 180
rect 3899 109 3945 146
rect 4047 972 4093 1009
rect 4047 938 4053 972
rect 4087 938 4093 972
rect 4047 900 4093 938
rect 4047 866 4053 900
rect 4087 866 4093 900
rect 4047 828 4093 866
rect 4047 794 4053 828
rect 4087 794 4093 828
rect 4047 756 4093 794
rect 4047 722 4053 756
rect 4087 722 4093 756
rect 4047 684 4093 722
rect 4047 650 4053 684
rect 4087 650 4093 684
rect 4047 612 4093 650
rect 4047 578 4053 612
rect 4087 578 4093 612
rect 4047 540 4093 578
rect 4047 506 4053 540
rect 4087 506 4093 540
rect 4047 468 4093 506
rect 4047 434 4053 468
rect 4087 434 4093 468
rect 4047 396 4093 434
rect 4047 362 4053 396
rect 4087 362 4093 396
rect 4047 324 4093 362
rect 4047 290 4053 324
rect 4087 290 4093 324
rect 4047 252 4093 290
rect 4047 218 4053 252
rect 4087 218 4093 252
rect 4047 180 4093 218
rect 4047 146 4053 180
rect 4087 146 4093 180
rect 4047 109 4093 146
rect 4195 972 4241 1009
rect 4195 938 4201 972
rect 4235 938 4241 972
rect 4195 900 4241 938
rect 4195 866 4201 900
rect 4235 866 4241 900
rect 4195 828 4241 866
rect 4195 794 4201 828
rect 4235 794 4241 828
rect 4195 756 4241 794
rect 4195 722 4201 756
rect 4235 722 4241 756
rect 4195 684 4241 722
rect 4195 650 4201 684
rect 4235 650 4241 684
rect 4195 612 4241 650
rect 4195 578 4201 612
rect 4235 578 4241 612
rect 4195 540 4241 578
rect 4195 506 4201 540
rect 4235 506 4241 540
rect 4195 468 4241 506
rect 4195 434 4201 468
rect 4235 434 4241 468
rect 4195 396 4241 434
rect 4195 362 4201 396
rect 4235 362 4241 396
rect 4195 324 4241 362
rect 4195 290 4201 324
rect 4235 290 4241 324
rect 4195 252 4241 290
rect 4195 218 4201 252
rect 4235 218 4241 252
rect 4195 180 4241 218
rect 4195 146 4201 180
rect 4235 146 4241 180
rect 4195 109 4241 146
rect 4343 972 4389 1009
rect 4343 938 4349 972
rect 4383 938 4389 972
rect 4343 900 4389 938
rect 4343 866 4349 900
rect 4383 866 4389 900
rect 4343 828 4389 866
rect 4343 794 4349 828
rect 4383 794 4389 828
rect 4343 756 4389 794
rect 4343 722 4349 756
rect 4383 722 4389 756
rect 4343 684 4389 722
rect 4343 650 4349 684
rect 4383 650 4389 684
rect 4343 612 4389 650
rect 4343 578 4349 612
rect 4383 578 4389 612
rect 4343 540 4389 578
rect 4343 506 4349 540
rect 4383 506 4389 540
rect 4343 468 4389 506
rect 4343 434 4349 468
rect 4383 434 4389 468
rect 4343 396 4389 434
rect 4343 362 4349 396
rect 4383 362 4389 396
rect 4343 324 4389 362
rect 4343 290 4349 324
rect 4383 290 4389 324
rect 4343 252 4389 290
rect 4343 218 4349 252
rect 4383 218 4389 252
rect 4343 180 4389 218
rect 4343 146 4349 180
rect 4383 146 4389 180
rect 4343 109 4389 146
rect 4491 972 4537 1009
rect 4491 938 4497 972
rect 4531 938 4537 972
rect 4491 900 4537 938
rect 4491 866 4497 900
rect 4531 866 4537 900
rect 4491 828 4537 866
rect 4491 794 4497 828
rect 4531 794 4537 828
rect 4491 756 4537 794
rect 4491 722 4497 756
rect 4531 722 4537 756
rect 4491 684 4537 722
rect 4491 650 4497 684
rect 4531 650 4537 684
rect 4491 612 4537 650
rect 4491 578 4497 612
rect 4531 578 4537 612
rect 4491 540 4537 578
rect 4491 506 4497 540
rect 4531 506 4537 540
rect 4491 468 4537 506
rect 4491 434 4497 468
rect 4531 434 4537 468
rect 4491 396 4537 434
rect 4491 362 4497 396
rect 4531 362 4537 396
rect 4491 324 4537 362
rect 4491 290 4497 324
rect 4531 290 4537 324
rect 4491 252 4537 290
rect 4491 218 4497 252
rect 4531 218 4537 252
rect 4491 180 4537 218
rect 4491 146 4497 180
rect 4531 146 4537 180
rect 4491 109 4537 146
rect 4639 972 4685 1009
rect 4639 938 4645 972
rect 4679 938 4685 972
rect 4639 900 4685 938
rect 4639 866 4645 900
rect 4679 866 4685 900
rect 4639 828 4685 866
rect 4639 794 4645 828
rect 4679 794 4685 828
rect 4639 756 4685 794
rect 4639 722 4645 756
rect 4679 722 4685 756
rect 4639 684 4685 722
rect 4639 650 4645 684
rect 4679 650 4685 684
rect 4639 612 4685 650
rect 4639 578 4645 612
rect 4679 578 4685 612
rect 4639 540 4685 578
rect 4639 506 4645 540
rect 4679 506 4685 540
rect 4639 468 4685 506
rect 4639 434 4645 468
rect 4679 434 4685 468
rect 4639 396 4685 434
rect 4639 362 4645 396
rect 4679 362 4685 396
rect 4639 324 4685 362
rect 4639 290 4645 324
rect 4679 290 4685 324
rect 4639 252 4685 290
rect 4639 218 4645 252
rect 4679 218 4685 252
rect 4639 180 4685 218
rect 4639 146 4645 180
rect 4679 146 4685 180
rect 4639 109 4685 146
rect 4787 972 4833 1009
rect 4787 938 4793 972
rect 4827 938 4833 972
rect 4787 900 4833 938
rect 4787 866 4793 900
rect 4827 866 4833 900
rect 4787 828 4833 866
rect 4787 794 4793 828
rect 4827 794 4833 828
rect 4787 756 4833 794
rect 4787 722 4793 756
rect 4827 722 4833 756
rect 4787 684 4833 722
rect 4787 650 4793 684
rect 4827 650 4833 684
rect 4787 612 4833 650
rect 4787 578 4793 612
rect 4827 578 4833 612
rect 4787 540 4833 578
rect 4787 506 4793 540
rect 4827 506 4833 540
rect 4787 468 4833 506
rect 4787 434 4793 468
rect 4827 434 4833 468
rect 4787 396 4833 434
rect 4787 362 4793 396
rect 4827 362 4833 396
rect 4787 324 4833 362
rect 4787 290 4793 324
rect 4827 290 4833 324
rect 4787 252 4833 290
rect 4787 218 4793 252
rect 4827 218 4833 252
rect 4787 180 4833 218
rect 4787 146 4793 180
rect 4827 146 4833 180
rect 4787 109 4833 146
rect 4935 972 4981 1009
rect 4935 938 4941 972
rect 4975 938 4981 972
rect 4935 900 4981 938
rect 4935 866 4941 900
rect 4975 866 4981 900
rect 4935 828 4981 866
rect 4935 794 4941 828
rect 4975 794 4981 828
rect 4935 756 4981 794
rect 4935 722 4941 756
rect 4975 722 4981 756
rect 4935 684 4981 722
rect 4935 650 4941 684
rect 4975 650 4981 684
rect 4935 612 4981 650
rect 4935 578 4941 612
rect 4975 578 4981 612
rect 4935 540 4981 578
rect 4935 506 4941 540
rect 4975 506 4981 540
rect 4935 468 4981 506
rect 4935 434 4941 468
rect 4975 434 4981 468
rect 4935 396 4981 434
rect 4935 362 4941 396
rect 4975 362 4981 396
rect 4935 324 4981 362
rect 4935 290 4941 324
rect 4975 290 4981 324
rect 4935 252 4981 290
rect 4935 218 4941 252
rect 4975 218 4981 252
rect 4935 180 4981 218
rect 4935 146 4941 180
rect 4975 146 4981 180
rect 4935 109 4981 146
rect 5083 972 5129 1009
rect 5083 938 5089 972
rect 5123 938 5129 972
rect 5083 900 5129 938
rect 5083 866 5089 900
rect 5123 866 5129 900
rect 5083 828 5129 866
rect 5083 794 5089 828
rect 5123 794 5129 828
rect 5083 756 5129 794
rect 5083 722 5089 756
rect 5123 722 5129 756
rect 5083 684 5129 722
rect 5083 650 5089 684
rect 5123 650 5129 684
rect 5083 612 5129 650
rect 5083 578 5089 612
rect 5123 578 5129 612
rect 5083 540 5129 578
rect 5083 506 5089 540
rect 5123 506 5129 540
rect 5083 468 5129 506
rect 5083 434 5089 468
rect 5123 434 5129 468
rect 5083 396 5129 434
rect 5083 362 5089 396
rect 5123 362 5129 396
rect 5083 324 5129 362
rect 5083 290 5089 324
rect 5123 290 5129 324
rect 5083 252 5129 290
rect 5083 218 5089 252
rect 5123 218 5129 252
rect 5083 180 5129 218
rect 5083 146 5089 180
rect 5123 146 5129 180
rect 5083 109 5129 146
rect 5231 972 5277 1009
rect 5231 938 5237 972
rect 5271 938 5277 972
rect 5231 900 5277 938
rect 5231 866 5237 900
rect 5271 866 5277 900
rect 5231 828 5277 866
rect 5231 794 5237 828
rect 5271 794 5277 828
rect 5231 756 5277 794
rect 5231 722 5237 756
rect 5271 722 5277 756
rect 5231 684 5277 722
rect 5231 650 5237 684
rect 5271 650 5277 684
rect 5231 612 5277 650
rect 5231 578 5237 612
rect 5271 578 5277 612
rect 5231 540 5277 578
rect 5231 506 5237 540
rect 5271 506 5277 540
rect 5231 468 5277 506
rect 5231 434 5237 468
rect 5271 434 5277 468
rect 5231 396 5277 434
rect 5231 362 5237 396
rect 5271 362 5277 396
rect 5231 324 5277 362
rect 5231 290 5237 324
rect 5271 290 5277 324
rect 5231 252 5277 290
rect 5231 218 5237 252
rect 5271 218 5277 252
rect 5231 180 5277 218
rect 5231 146 5237 180
rect 5271 146 5277 180
rect 5231 109 5277 146
rect 5379 972 5425 1009
rect 5379 938 5385 972
rect 5419 938 5425 972
rect 5379 900 5425 938
rect 5379 866 5385 900
rect 5419 866 5425 900
rect 5379 828 5425 866
rect 5379 794 5385 828
rect 5419 794 5425 828
rect 5379 756 5425 794
rect 5379 722 5385 756
rect 5419 722 5425 756
rect 5379 684 5425 722
rect 5379 650 5385 684
rect 5419 650 5425 684
rect 5379 612 5425 650
rect 5379 578 5385 612
rect 5419 578 5425 612
rect 5379 540 5425 578
rect 5379 506 5385 540
rect 5419 506 5425 540
rect 5379 468 5425 506
rect 5379 434 5385 468
rect 5419 434 5425 468
rect 5379 396 5425 434
rect 5379 362 5385 396
rect 5419 362 5425 396
rect 5379 324 5425 362
rect 5379 290 5385 324
rect 5419 290 5425 324
rect 5379 252 5425 290
rect 5379 218 5385 252
rect 5419 218 5425 252
rect 5379 180 5425 218
rect 5379 146 5385 180
rect 5419 146 5425 180
rect 5379 109 5425 146
rect 5527 972 5573 1009
rect 5527 938 5533 972
rect 5567 938 5573 972
rect 5527 900 5573 938
rect 5527 866 5533 900
rect 5567 866 5573 900
rect 5527 828 5573 866
rect 5527 794 5533 828
rect 5567 794 5573 828
rect 5527 756 5573 794
rect 5527 722 5533 756
rect 5567 722 5573 756
rect 5527 684 5573 722
rect 5527 650 5533 684
rect 5567 650 5573 684
rect 5527 612 5573 650
rect 5527 578 5533 612
rect 5567 578 5573 612
rect 5527 540 5573 578
rect 5527 506 5533 540
rect 5567 506 5573 540
rect 5527 468 5573 506
rect 5527 434 5533 468
rect 5567 434 5573 468
rect 5527 396 5573 434
rect 5527 362 5533 396
rect 5567 362 5573 396
rect 5527 324 5573 362
rect 5527 290 5533 324
rect 5567 290 5573 324
rect 5527 252 5573 290
rect 5527 218 5533 252
rect 5567 218 5573 252
rect 5527 180 5573 218
rect 5527 146 5533 180
rect 5567 146 5573 180
rect 5527 109 5573 146
rect -5517 71 -5435 77
rect -5517 37 -5493 71
rect -5459 37 -5435 71
rect -5517 31 -5435 37
rect -5369 71 -5287 77
rect -5369 37 -5345 71
rect -5311 37 -5287 71
rect -5369 31 -5287 37
rect -5221 71 -5139 77
rect -5221 37 -5197 71
rect -5163 37 -5139 71
rect -5221 31 -5139 37
rect -5073 71 -4991 77
rect -5073 37 -5049 71
rect -5015 37 -4991 71
rect -5073 31 -4991 37
rect -4925 71 -4843 77
rect -4925 37 -4901 71
rect -4867 37 -4843 71
rect -4925 31 -4843 37
rect -4777 71 -4695 77
rect -4777 37 -4753 71
rect -4719 37 -4695 71
rect -4777 31 -4695 37
rect -4629 71 -4547 77
rect -4629 37 -4605 71
rect -4571 37 -4547 71
rect -4629 31 -4547 37
rect -4481 71 -4399 77
rect -4481 37 -4457 71
rect -4423 37 -4399 71
rect -4481 31 -4399 37
rect -4333 71 -4251 77
rect -4333 37 -4309 71
rect -4275 37 -4251 71
rect -4333 31 -4251 37
rect -4185 71 -4103 77
rect -4185 37 -4161 71
rect -4127 37 -4103 71
rect -4185 31 -4103 37
rect -4037 71 -3955 77
rect -4037 37 -4013 71
rect -3979 37 -3955 71
rect -4037 31 -3955 37
rect -3889 71 -3807 77
rect -3889 37 -3865 71
rect -3831 37 -3807 71
rect -3889 31 -3807 37
rect -3741 71 -3659 77
rect -3741 37 -3717 71
rect -3683 37 -3659 71
rect -3741 31 -3659 37
rect -3593 71 -3511 77
rect -3593 37 -3569 71
rect -3535 37 -3511 71
rect -3593 31 -3511 37
rect -3445 71 -3363 77
rect -3445 37 -3421 71
rect -3387 37 -3363 71
rect -3445 31 -3363 37
rect -3297 71 -3215 77
rect -3297 37 -3273 71
rect -3239 37 -3215 71
rect -3297 31 -3215 37
rect -3149 71 -3067 77
rect -3149 37 -3125 71
rect -3091 37 -3067 71
rect -3149 31 -3067 37
rect -3001 71 -2919 77
rect -3001 37 -2977 71
rect -2943 37 -2919 71
rect -3001 31 -2919 37
rect -2853 71 -2771 77
rect -2853 37 -2829 71
rect -2795 37 -2771 71
rect -2853 31 -2771 37
rect -2705 71 -2623 77
rect -2705 37 -2681 71
rect -2647 37 -2623 71
rect -2705 31 -2623 37
rect -2557 71 -2475 77
rect -2557 37 -2533 71
rect -2499 37 -2475 71
rect -2557 31 -2475 37
rect -2409 71 -2327 77
rect -2409 37 -2385 71
rect -2351 37 -2327 71
rect -2409 31 -2327 37
rect -2261 71 -2179 77
rect -2261 37 -2237 71
rect -2203 37 -2179 71
rect -2261 31 -2179 37
rect -2113 71 -2031 77
rect -2113 37 -2089 71
rect -2055 37 -2031 71
rect -2113 31 -2031 37
rect -1965 71 -1883 77
rect -1965 37 -1941 71
rect -1907 37 -1883 71
rect -1965 31 -1883 37
rect -1817 71 -1735 77
rect -1817 37 -1793 71
rect -1759 37 -1735 71
rect -1817 31 -1735 37
rect -1669 71 -1587 77
rect -1669 37 -1645 71
rect -1611 37 -1587 71
rect -1669 31 -1587 37
rect -1521 71 -1439 77
rect -1521 37 -1497 71
rect -1463 37 -1439 71
rect -1521 31 -1439 37
rect -1373 71 -1291 77
rect -1373 37 -1349 71
rect -1315 37 -1291 71
rect -1373 31 -1291 37
rect -1225 71 -1143 77
rect -1225 37 -1201 71
rect -1167 37 -1143 71
rect -1225 31 -1143 37
rect -1077 71 -995 77
rect -1077 37 -1053 71
rect -1019 37 -995 71
rect -1077 31 -995 37
rect -929 71 -847 77
rect -929 37 -905 71
rect -871 37 -847 71
rect -929 31 -847 37
rect -781 71 -699 77
rect -781 37 -757 71
rect -723 37 -699 71
rect -781 31 -699 37
rect -633 71 -551 77
rect -633 37 -609 71
rect -575 37 -551 71
rect -633 31 -551 37
rect -485 71 -403 77
rect -485 37 -461 71
rect -427 37 -403 71
rect -485 31 -403 37
rect -337 71 -255 77
rect -337 37 -313 71
rect -279 37 -255 71
rect -337 31 -255 37
rect -189 71 -107 77
rect -189 37 -165 71
rect -131 37 -107 71
rect -189 31 -107 37
rect -41 71 41 77
rect -41 37 -17 71
rect 17 37 41 71
rect -41 31 41 37
rect 107 71 189 77
rect 107 37 131 71
rect 165 37 189 71
rect 107 31 189 37
rect 255 71 337 77
rect 255 37 279 71
rect 313 37 337 71
rect 255 31 337 37
rect 403 71 485 77
rect 403 37 427 71
rect 461 37 485 71
rect 403 31 485 37
rect 551 71 633 77
rect 551 37 575 71
rect 609 37 633 71
rect 551 31 633 37
rect 699 71 781 77
rect 699 37 723 71
rect 757 37 781 71
rect 699 31 781 37
rect 847 71 929 77
rect 847 37 871 71
rect 905 37 929 71
rect 847 31 929 37
rect 995 71 1077 77
rect 995 37 1019 71
rect 1053 37 1077 71
rect 995 31 1077 37
rect 1143 71 1225 77
rect 1143 37 1167 71
rect 1201 37 1225 71
rect 1143 31 1225 37
rect 1291 71 1373 77
rect 1291 37 1315 71
rect 1349 37 1373 71
rect 1291 31 1373 37
rect 1439 71 1521 77
rect 1439 37 1463 71
rect 1497 37 1521 71
rect 1439 31 1521 37
rect 1587 71 1669 77
rect 1587 37 1611 71
rect 1645 37 1669 71
rect 1587 31 1669 37
rect 1735 71 1817 77
rect 1735 37 1759 71
rect 1793 37 1817 71
rect 1735 31 1817 37
rect 1883 71 1965 77
rect 1883 37 1907 71
rect 1941 37 1965 71
rect 1883 31 1965 37
rect 2031 71 2113 77
rect 2031 37 2055 71
rect 2089 37 2113 71
rect 2031 31 2113 37
rect 2179 71 2261 77
rect 2179 37 2203 71
rect 2237 37 2261 71
rect 2179 31 2261 37
rect 2327 71 2409 77
rect 2327 37 2351 71
rect 2385 37 2409 71
rect 2327 31 2409 37
rect 2475 71 2557 77
rect 2475 37 2499 71
rect 2533 37 2557 71
rect 2475 31 2557 37
rect 2623 71 2705 77
rect 2623 37 2647 71
rect 2681 37 2705 71
rect 2623 31 2705 37
rect 2771 71 2853 77
rect 2771 37 2795 71
rect 2829 37 2853 71
rect 2771 31 2853 37
rect 2919 71 3001 77
rect 2919 37 2943 71
rect 2977 37 3001 71
rect 2919 31 3001 37
rect 3067 71 3149 77
rect 3067 37 3091 71
rect 3125 37 3149 71
rect 3067 31 3149 37
rect 3215 71 3297 77
rect 3215 37 3239 71
rect 3273 37 3297 71
rect 3215 31 3297 37
rect 3363 71 3445 77
rect 3363 37 3387 71
rect 3421 37 3445 71
rect 3363 31 3445 37
rect 3511 71 3593 77
rect 3511 37 3535 71
rect 3569 37 3593 71
rect 3511 31 3593 37
rect 3659 71 3741 77
rect 3659 37 3683 71
rect 3717 37 3741 71
rect 3659 31 3741 37
rect 3807 71 3889 77
rect 3807 37 3831 71
rect 3865 37 3889 71
rect 3807 31 3889 37
rect 3955 71 4037 77
rect 3955 37 3979 71
rect 4013 37 4037 71
rect 3955 31 4037 37
rect 4103 71 4185 77
rect 4103 37 4127 71
rect 4161 37 4185 71
rect 4103 31 4185 37
rect 4251 71 4333 77
rect 4251 37 4275 71
rect 4309 37 4333 71
rect 4251 31 4333 37
rect 4399 71 4481 77
rect 4399 37 4423 71
rect 4457 37 4481 71
rect 4399 31 4481 37
rect 4547 71 4629 77
rect 4547 37 4571 71
rect 4605 37 4629 71
rect 4547 31 4629 37
rect 4695 71 4777 77
rect 4695 37 4719 71
rect 4753 37 4777 71
rect 4695 31 4777 37
rect 4843 71 4925 77
rect 4843 37 4867 71
rect 4901 37 4925 71
rect 4843 31 4925 37
rect 4991 71 5073 77
rect 4991 37 5015 71
rect 5049 37 5073 71
rect 4991 31 5073 37
rect 5139 71 5221 77
rect 5139 37 5163 71
rect 5197 37 5221 71
rect 5139 31 5221 37
rect 5287 71 5369 77
rect 5287 37 5311 71
rect 5345 37 5369 71
rect 5287 31 5369 37
rect 5435 71 5517 77
rect 5435 37 5459 71
rect 5493 37 5517 71
rect 5435 31 5517 37
rect -5517 -37 -5435 -31
rect -5517 -71 -5493 -37
rect -5459 -71 -5435 -37
rect -5517 -77 -5435 -71
rect -5369 -37 -5287 -31
rect -5369 -71 -5345 -37
rect -5311 -71 -5287 -37
rect -5369 -77 -5287 -71
rect -5221 -37 -5139 -31
rect -5221 -71 -5197 -37
rect -5163 -71 -5139 -37
rect -5221 -77 -5139 -71
rect -5073 -37 -4991 -31
rect -5073 -71 -5049 -37
rect -5015 -71 -4991 -37
rect -5073 -77 -4991 -71
rect -4925 -37 -4843 -31
rect -4925 -71 -4901 -37
rect -4867 -71 -4843 -37
rect -4925 -77 -4843 -71
rect -4777 -37 -4695 -31
rect -4777 -71 -4753 -37
rect -4719 -71 -4695 -37
rect -4777 -77 -4695 -71
rect -4629 -37 -4547 -31
rect -4629 -71 -4605 -37
rect -4571 -71 -4547 -37
rect -4629 -77 -4547 -71
rect -4481 -37 -4399 -31
rect -4481 -71 -4457 -37
rect -4423 -71 -4399 -37
rect -4481 -77 -4399 -71
rect -4333 -37 -4251 -31
rect -4333 -71 -4309 -37
rect -4275 -71 -4251 -37
rect -4333 -77 -4251 -71
rect -4185 -37 -4103 -31
rect -4185 -71 -4161 -37
rect -4127 -71 -4103 -37
rect -4185 -77 -4103 -71
rect -4037 -37 -3955 -31
rect -4037 -71 -4013 -37
rect -3979 -71 -3955 -37
rect -4037 -77 -3955 -71
rect -3889 -37 -3807 -31
rect -3889 -71 -3865 -37
rect -3831 -71 -3807 -37
rect -3889 -77 -3807 -71
rect -3741 -37 -3659 -31
rect -3741 -71 -3717 -37
rect -3683 -71 -3659 -37
rect -3741 -77 -3659 -71
rect -3593 -37 -3511 -31
rect -3593 -71 -3569 -37
rect -3535 -71 -3511 -37
rect -3593 -77 -3511 -71
rect -3445 -37 -3363 -31
rect -3445 -71 -3421 -37
rect -3387 -71 -3363 -37
rect -3445 -77 -3363 -71
rect -3297 -37 -3215 -31
rect -3297 -71 -3273 -37
rect -3239 -71 -3215 -37
rect -3297 -77 -3215 -71
rect -3149 -37 -3067 -31
rect -3149 -71 -3125 -37
rect -3091 -71 -3067 -37
rect -3149 -77 -3067 -71
rect -3001 -37 -2919 -31
rect -3001 -71 -2977 -37
rect -2943 -71 -2919 -37
rect -3001 -77 -2919 -71
rect -2853 -37 -2771 -31
rect -2853 -71 -2829 -37
rect -2795 -71 -2771 -37
rect -2853 -77 -2771 -71
rect -2705 -37 -2623 -31
rect -2705 -71 -2681 -37
rect -2647 -71 -2623 -37
rect -2705 -77 -2623 -71
rect -2557 -37 -2475 -31
rect -2557 -71 -2533 -37
rect -2499 -71 -2475 -37
rect -2557 -77 -2475 -71
rect -2409 -37 -2327 -31
rect -2409 -71 -2385 -37
rect -2351 -71 -2327 -37
rect -2409 -77 -2327 -71
rect -2261 -37 -2179 -31
rect -2261 -71 -2237 -37
rect -2203 -71 -2179 -37
rect -2261 -77 -2179 -71
rect -2113 -37 -2031 -31
rect -2113 -71 -2089 -37
rect -2055 -71 -2031 -37
rect -2113 -77 -2031 -71
rect -1965 -37 -1883 -31
rect -1965 -71 -1941 -37
rect -1907 -71 -1883 -37
rect -1965 -77 -1883 -71
rect -1817 -37 -1735 -31
rect -1817 -71 -1793 -37
rect -1759 -71 -1735 -37
rect -1817 -77 -1735 -71
rect -1669 -37 -1587 -31
rect -1669 -71 -1645 -37
rect -1611 -71 -1587 -37
rect -1669 -77 -1587 -71
rect -1521 -37 -1439 -31
rect -1521 -71 -1497 -37
rect -1463 -71 -1439 -37
rect -1521 -77 -1439 -71
rect -1373 -37 -1291 -31
rect -1373 -71 -1349 -37
rect -1315 -71 -1291 -37
rect -1373 -77 -1291 -71
rect -1225 -37 -1143 -31
rect -1225 -71 -1201 -37
rect -1167 -71 -1143 -37
rect -1225 -77 -1143 -71
rect -1077 -37 -995 -31
rect -1077 -71 -1053 -37
rect -1019 -71 -995 -37
rect -1077 -77 -995 -71
rect -929 -37 -847 -31
rect -929 -71 -905 -37
rect -871 -71 -847 -37
rect -929 -77 -847 -71
rect -781 -37 -699 -31
rect -781 -71 -757 -37
rect -723 -71 -699 -37
rect -781 -77 -699 -71
rect -633 -37 -551 -31
rect -633 -71 -609 -37
rect -575 -71 -551 -37
rect -633 -77 -551 -71
rect -485 -37 -403 -31
rect -485 -71 -461 -37
rect -427 -71 -403 -37
rect -485 -77 -403 -71
rect -337 -37 -255 -31
rect -337 -71 -313 -37
rect -279 -71 -255 -37
rect -337 -77 -255 -71
rect -189 -37 -107 -31
rect -189 -71 -165 -37
rect -131 -71 -107 -37
rect -189 -77 -107 -71
rect -41 -37 41 -31
rect -41 -71 -17 -37
rect 17 -71 41 -37
rect -41 -77 41 -71
rect 107 -37 189 -31
rect 107 -71 131 -37
rect 165 -71 189 -37
rect 107 -77 189 -71
rect 255 -37 337 -31
rect 255 -71 279 -37
rect 313 -71 337 -37
rect 255 -77 337 -71
rect 403 -37 485 -31
rect 403 -71 427 -37
rect 461 -71 485 -37
rect 403 -77 485 -71
rect 551 -37 633 -31
rect 551 -71 575 -37
rect 609 -71 633 -37
rect 551 -77 633 -71
rect 699 -37 781 -31
rect 699 -71 723 -37
rect 757 -71 781 -37
rect 699 -77 781 -71
rect 847 -37 929 -31
rect 847 -71 871 -37
rect 905 -71 929 -37
rect 847 -77 929 -71
rect 995 -37 1077 -31
rect 995 -71 1019 -37
rect 1053 -71 1077 -37
rect 995 -77 1077 -71
rect 1143 -37 1225 -31
rect 1143 -71 1167 -37
rect 1201 -71 1225 -37
rect 1143 -77 1225 -71
rect 1291 -37 1373 -31
rect 1291 -71 1315 -37
rect 1349 -71 1373 -37
rect 1291 -77 1373 -71
rect 1439 -37 1521 -31
rect 1439 -71 1463 -37
rect 1497 -71 1521 -37
rect 1439 -77 1521 -71
rect 1587 -37 1669 -31
rect 1587 -71 1611 -37
rect 1645 -71 1669 -37
rect 1587 -77 1669 -71
rect 1735 -37 1817 -31
rect 1735 -71 1759 -37
rect 1793 -71 1817 -37
rect 1735 -77 1817 -71
rect 1883 -37 1965 -31
rect 1883 -71 1907 -37
rect 1941 -71 1965 -37
rect 1883 -77 1965 -71
rect 2031 -37 2113 -31
rect 2031 -71 2055 -37
rect 2089 -71 2113 -37
rect 2031 -77 2113 -71
rect 2179 -37 2261 -31
rect 2179 -71 2203 -37
rect 2237 -71 2261 -37
rect 2179 -77 2261 -71
rect 2327 -37 2409 -31
rect 2327 -71 2351 -37
rect 2385 -71 2409 -37
rect 2327 -77 2409 -71
rect 2475 -37 2557 -31
rect 2475 -71 2499 -37
rect 2533 -71 2557 -37
rect 2475 -77 2557 -71
rect 2623 -37 2705 -31
rect 2623 -71 2647 -37
rect 2681 -71 2705 -37
rect 2623 -77 2705 -71
rect 2771 -37 2853 -31
rect 2771 -71 2795 -37
rect 2829 -71 2853 -37
rect 2771 -77 2853 -71
rect 2919 -37 3001 -31
rect 2919 -71 2943 -37
rect 2977 -71 3001 -37
rect 2919 -77 3001 -71
rect 3067 -37 3149 -31
rect 3067 -71 3091 -37
rect 3125 -71 3149 -37
rect 3067 -77 3149 -71
rect 3215 -37 3297 -31
rect 3215 -71 3239 -37
rect 3273 -71 3297 -37
rect 3215 -77 3297 -71
rect 3363 -37 3445 -31
rect 3363 -71 3387 -37
rect 3421 -71 3445 -37
rect 3363 -77 3445 -71
rect 3511 -37 3593 -31
rect 3511 -71 3535 -37
rect 3569 -71 3593 -37
rect 3511 -77 3593 -71
rect 3659 -37 3741 -31
rect 3659 -71 3683 -37
rect 3717 -71 3741 -37
rect 3659 -77 3741 -71
rect 3807 -37 3889 -31
rect 3807 -71 3831 -37
rect 3865 -71 3889 -37
rect 3807 -77 3889 -71
rect 3955 -37 4037 -31
rect 3955 -71 3979 -37
rect 4013 -71 4037 -37
rect 3955 -77 4037 -71
rect 4103 -37 4185 -31
rect 4103 -71 4127 -37
rect 4161 -71 4185 -37
rect 4103 -77 4185 -71
rect 4251 -37 4333 -31
rect 4251 -71 4275 -37
rect 4309 -71 4333 -37
rect 4251 -77 4333 -71
rect 4399 -37 4481 -31
rect 4399 -71 4423 -37
rect 4457 -71 4481 -37
rect 4399 -77 4481 -71
rect 4547 -37 4629 -31
rect 4547 -71 4571 -37
rect 4605 -71 4629 -37
rect 4547 -77 4629 -71
rect 4695 -37 4777 -31
rect 4695 -71 4719 -37
rect 4753 -71 4777 -37
rect 4695 -77 4777 -71
rect 4843 -37 4925 -31
rect 4843 -71 4867 -37
rect 4901 -71 4925 -37
rect 4843 -77 4925 -71
rect 4991 -37 5073 -31
rect 4991 -71 5015 -37
rect 5049 -71 5073 -37
rect 4991 -77 5073 -71
rect 5139 -37 5221 -31
rect 5139 -71 5163 -37
rect 5197 -71 5221 -37
rect 5139 -77 5221 -71
rect 5287 -37 5369 -31
rect 5287 -71 5311 -37
rect 5345 -71 5369 -37
rect 5287 -77 5369 -71
rect 5435 -37 5517 -31
rect 5435 -71 5459 -37
rect 5493 -71 5517 -37
rect 5435 -77 5517 -71
rect -5573 -146 -5527 -109
rect -5573 -180 -5567 -146
rect -5533 -180 -5527 -146
rect -5573 -218 -5527 -180
rect -5573 -252 -5567 -218
rect -5533 -252 -5527 -218
rect -5573 -290 -5527 -252
rect -5573 -324 -5567 -290
rect -5533 -324 -5527 -290
rect -5573 -362 -5527 -324
rect -5573 -396 -5567 -362
rect -5533 -396 -5527 -362
rect -5573 -434 -5527 -396
rect -5573 -468 -5567 -434
rect -5533 -468 -5527 -434
rect -5573 -506 -5527 -468
rect -5573 -540 -5567 -506
rect -5533 -540 -5527 -506
rect -5573 -578 -5527 -540
rect -5573 -612 -5567 -578
rect -5533 -612 -5527 -578
rect -5573 -650 -5527 -612
rect -5573 -684 -5567 -650
rect -5533 -684 -5527 -650
rect -5573 -722 -5527 -684
rect -5573 -756 -5567 -722
rect -5533 -756 -5527 -722
rect -5573 -794 -5527 -756
rect -5573 -828 -5567 -794
rect -5533 -828 -5527 -794
rect -5573 -866 -5527 -828
rect -5573 -900 -5567 -866
rect -5533 -900 -5527 -866
rect -5573 -938 -5527 -900
rect -5573 -972 -5567 -938
rect -5533 -972 -5527 -938
rect -5573 -1009 -5527 -972
rect -5425 -146 -5379 -109
rect -5425 -180 -5419 -146
rect -5385 -180 -5379 -146
rect -5425 -218 -5379 -180
rect -5425 -252 -5419 -218
rect -5385 -252 -5379 -218
rect -5425 -290 -5379 -252
rect -5425 -324 -5419 -290
rect -5385 -324 -5379 -290
rect -5425 -362 -5379 -324
rect -5425 -396 -5419 -362
rect -5385 -396 -5379 -362
rect -5425 -434 -5379 -396
rect -5425 -468 -5419 -434
rect -5385 -468 -5379 -434
rect -5425 -506 -5379 -468
rect -5425 -540 -5419 -506
rect -5385 -540 -5379 -506
rect -5425 -578 -5379 -540
rect -5425 -612 -5419 -578
rect -5385 -612 -5379 -578
rect -5425 -650 -5379 -612
rect -5425 -684 -5419 -650
rect -5385 -684 -5379 -650
rect -5425 -722 -5379 -684
rect -5425 -756 -5419 -722
rect -5385 -756 -5379 -722
rect -5425 -794 -5379 -756
rect -5425 -828 -5419 -794
rect -5385 -828 -5379 -794
rect -5425 -866 -5379 -828
rect -5425 -900 -5419 -866
rect -5385 -900 -5379 -866
rect -5425 -938 -5379 -900
rect -5425 -972 -5419 -938
rect -5385 -972 -5379 -938
rect -5425 -1009 -5379 -972
rect -5277 -146 -5231 -109
rect -5277 -180 -5271 -146
rect -5237 -180 -5231 -146
rect -5277 -218 -5231 -180
rect -5277 -252 -5271 -218
rect -5237 -252 -5231 -218
rect -5277 -290 -5231 -252
rect -5277 -324 -5271 -290
rect -5237 -324 -5231 -290
rect -5277 -362 -5231 -324
rect -5277 -396 -5271 -362
rect -5237 -396 -5231 -362
rect -5277 -434 -5231 -396
rect -5277 -468 -5271 -434
rect -5237 -468 -5231 -434
rect -5277 -506 -5231 -468
rect -5277 -540 -5271 -506
rect -5237 -540 -5231 -506
rect -5277 -578 -5231 -540
rect -5277 -612 -5271 -578
rect -5237 -612 -5231 -578
rect -5277 -650 -5231 -612
rect -5277 -684 -5271 -650
rect -5237 -684 -5231 -650
rect -5277 -722 -5231 -684
rect -5277 -756 -5271 -722
rect -5237 -756 -5231 -722
rect -5277 -794 -5231 -756
rect -5277 -828 -5271 -794
rect -5237 -828 -5231 -794
rect -5277 -866 -5231 -828
rect -5277 -900 -5271 -866
rect -5237 -900 -5231 -866
rect -5277 -938 -5231 -900
rect -5277 -972 -5271 -938
rect -5237 -972 -5231 -938
rect -5277 -1009 -5231 -972
rect -5129 -146 -5083 -109
rect -5129 -180 -5123 -146
rect -5089 -180 -5083 -146
rect -5129 -218 -5083 -180
rect -5129 -252 -5123 -218
rect -5089 -252 -5083 -218
rect -5129 -290 -5083 -252
rect -5129 -324 -5123 -290
rect -5089 -324 -5083 -290
rect -5129 -362 -5083 -324
rect -5129 -396 -5123 -362
rect -5089 -396 -5083 -362
rect -5129 -434 -5083 -396
rect -5129 -468 -5123 -434
rect -5089 -468 -5083 -434
rect -5129 -506 -5083 -468
rect -5129 -540 -5123 -506
rect -5089 -540 -5083 -506
rect -5129 -578 -5083 -540
rect -5129 -612 -5123 -578
rect -5089 -612 -5083 -578
rect -5129 -650 -5083 -612
rect -5129 -684 -5123 -650
rect -5089 -684 -5083 -650
rect -5129 -722 -5083 -684
rect -5129 -756 -5123 -722
rect -5089 -756 -5083 -722
rect -5129 -794 -5083 -756
rect -5129 -828 -5123 -794
rect -5089 -828 -5083 -794
rect -5129 -866 -5083 -828
rect -5129 -900 -5123 -866
rect -5089 -900 -5083 -866
rect -5129 -938 -5083 -900
rect -5129 -972 -5123 -938
rect -5089 -972 -5083 -938
rect -5129 -1009 -5083 -972
rect -4981 -146 -4935 -109
rect -4981 -180 -4975 -146
rect -4941 -180 -4935 -146
rect -4981 -218 -4935 -180
rect -4981 -252 -4975 -218
rect -4941 -252 -4935 -218
rect -4981 -290 -4935 -252
rect -4981 -324 -4975 -290
rect -4941 -324 -4935 -290
rect -4981 -362 -4935 -324
rect -4981 -396 -4975 -362
rect -4941 -396 -4935 -362
rect -4981 -434 -4935 -396
rect -4981 -468 -4975 -434
rect -4941 -468 -4935 -434
rect -4981 -506 -4935 -468
rect -4981 -540 -4975 -506
rect -4941 -540 -4935 -506
rect -4981 -578 -4935 -540
rect -4981 -612 -4975 -578
rect -4941 -612 -4935 -578
rect -4981 -650 -4935 -612
rect -4981 -684 -4975 -650
rect -4941 -684 -4935 -650
rect -4981 -722 -4935 -684
rect -4981 -756 -4975 -722
rect -4941 -756 -4935 -722
rect -4981 -794 -4935 -756
rect -4981 -828 -4975 -794
rect -4941 -828 -4935 -794
rect -4981 -866 -4935 -828
rect -4981 -900 -4975 -866
rect -4941 -900 -4935 -866
rect -4981 -938 -4935 -900
rect -4981 -972 -4975 -938
rect -4941 -972 -4935 -938
rect -4981 -1009 -4935 -972
rect -4833 -146 -4787 -109
rect -4833 -180 -4827 -146
rect -4793 -180 -4787 -146
rect -4833 -218 -4787 -180
rect -4833 -252 -4827 -218
rect -4793 -252 -4787 -218
rect -4833 -290 -4787 -252
rect -4833 -324 -4827 -290
rect -4793 -324 -4787 -290
rect -4833 -362 -4787 -324
rect -4833 -396 -4827 -362
rect -4793 -396 -4787 -362
rect -4833 -434 -4787 -396
rect -4833 -468 -4827 -434
rect -4793 -468 -4787 -434
rect -4833 -506 -4787 -468
rect -4833 -540 -4827 -506
rect -4793 -540 -4787 -506
rect -4833 -578 -4787 -540
rect -4833 -612 -4827 -578
rect -4793 -612 -4787 -578
rect -4833 -650 -4787 -612
rect -4833 -684 -4827 -650
rect -4793 -684 -4787 -650
rect -4833 -722 -4787 -684
rect -4833 -756 -4827 -722
rect -4793 -756 -4787 -722
rect -4833 -794 -4787 -756
rect -4833 -828 -4827 -794
rect -4793 -828 -4787 -794
rect -4833 -866 -4787 -828
rect -4833 -900 -4827 -866
rect -4793 -900 -4787 -866
rect -4833 -938 -4787 -900
rect -4833 -972 -4827 -938
rect -4793 -972 -4787 -938
rect -4833 -1009 -4787 -972
rect -4685 -146 -4639 -109
rect -4685 -180 -4679 -146
rect -4645 -180 -4639 -146
rect -4685 -218 -4639 -180
rect -4685 -252 -4679 -218
rect -4645 -252 -4639 -218
rect -4685 -290 -4639 -252
rect -4685 -324 -4679 -290
rect -4645 -324 -4639 -290
rect -4685 -362 -4639 -324
rect -4685 -396 -4679 -362
rect -4645 -396 -4639 -362
rect -4685 -434 -4639 -396
rect -4685 -468 -4679 -434
rect -4645 -468 -4639 -434
rect -4685 -506 -4639 -468
rect -4685 -540 -4679 -506
rect -4645 -540 -4639 -506
rect -4685 -578 -4639 -540
rect -4685 -612 -4679 -578
rect -4645 -612 -4639 -578
rect -4685 -650 -4639 -612
rect -4685 -684 -4679 -650
rect -4645 -684 -4639 -650
rect -4685 -722 -4639 -684
rect -4685 -756 -4679 -722
rect -4645 -756 -4639 -722
rect -4685 -794 -4639 -756
rect -4685 -828 -4679 -794
rect -4645 -828 -4639 -794
rect -4685 -866 -4639 -828
rect -4685 -900 -4679 -866
rect -4645 -900 -4639 -866
rect -4685 -938 -4639 -900
rect -4685 -972 -4679 -938
rect -4645 -972 -4639 -938
rect -4685 -1009 -4639 -972
rect -4537 -146 -4491 -109
rect -4537 -180 -4531 -146
rect -4497 -180 -4491 -146
rect -4537 -218 -4491 -180
rect -4537 -252 -4531 -218
rect -4497 -252 -4491 -218
rect -4537 -290 -4491 -252
rect -4537 -324 -4531 -290
rect -4497 -324 -4491 -290
rect -4537 -362 -4491 -324
rect -4537 -396 -4531 -362
rect -4497 -396 -4491 -362
rect -4537 -434 -4491 -396
rect -4537 -468 -4531 -434
rect -4497 -468 -4491 -434
rect -4537 -506 -4491 -468
rect -4537 -540 -4531 -506
rect -4497 -540 -4491 -506
rect -4537 -578 -4491 -540
rect -4537 -612 -4531 -578
rect -4497 -612 -4491 -578
rect -4537 -650 -4491 -612
rect -4537 -684 -4531 -650
rect -4497 -684 -4491 -650
rect -4537 -722 -4491 -684
rect -4537 -756 -4531 -722
rect -4497 -756 -4491 -722
rect -4537 -794 -4491 -756
rect -4537 -828 -4531 -794
rect -4497 -828 -4491 -794
rect -4537 -866 -4491 -828
rect -4537 -900 -4531 -866
rect -4497 -900 -4491 -866
rect -4537 -938 -4491 -900
rect -4537 -972 -4531 -938
rect -4497 -972 -4491 -938
rect -4537 -1009 -4491 -972
rect -4389 -146 -4343 -109
rect -4389 -180 -4383 -146
rect -4349 -180 -4343 -146
rect -4389 -218 -4343 -180
rect -4389 -252 -4383 -218
rect -4349 -252 -4343 -218
rect -4389 -290 -4343 -252
rect -4389 -324 -4383 -290
rect -4349 -324 -4343 -290
rect -4389 -362 -4343 -324
rect -4389 -396 -4383 -362
rect -4349 -396 -4343 -362
rect -4389 -434 -4343 -396
rect -4389 -468 -4383 -434
rect -4349 -468 -4343 -434
rect -4389 -506 -4343 -468
rect -4389 -540 -4383 -506
rect -4349 -540 -4343 -506
rect -4389 -578 -4343 -540
rect -4389 -612 -4383 -578
rect -4349 -612 -4343 -578
rect -4389 -650 -4343 -612
rect -4389 -684 -4383 -650
rect -4349 -684 -4343 -650
rect -4389 -722 -4343 -684
rect -4389 -756 -4383 -722
rect -4349 -756 -4343 -722
rect -4389 -794 -4343 -756
rect -4389 -828 -4383 -794
rect -4349 -828 -4343 -794
rect -4389 -866 -4343 -828
rect -4389 -900 -4383 -866
rect -4349 -900 -4343 -866
rect -4389 -938 -4343 -900
rect -4389 -972 -4383 -938
rect -4349 -972 -4343 -938
rect -4389 -1009 -4343 -972
rect -4241 -146 -4195 -109
rect -4241 -180 -4235 -146
rect -4201 -180 -4195 -146
rect -4241 -218 -4195 -180
rect -4241 -252 -4235 -218
rect -4201 -252 -4195 -218
rect -4241 -290 -4195 -252
rect -4241 -324 -4235 -290
rect -4201 -324 -4195 -290
rect -4241 -362 -4195 -324
rect -4241 -396 -4235 -362
rect -4201 -396 -4195 -362
rect -4241 -434 -4195 -396
rect -4241 -468 -4235 -434
rect -4201 -468 -4195 -434
rect -4241 -506 -4195 -468
rect -4241 -540 -4235 -506
rect -4201 -540 -4195 -506
rect -4241 -578 -4195 -540
rect -4241 -612 -4235 -578
rect -4201 -612 -4195 -578
rect -4241 -650 -4195 -612
rect -4241 -684 -4235 -650
rect -4201 -684 -4195 -650
rect -4241 -722 -4195 -684
rect -4241 -756 -4235 -722
rect -4201 -756 -4195 -722
rect -4241 -794 -4195 -756
rect -4241 -828 -4235 -794
rect -4201 -828 -4195 -794
rect -4241 -866 -4195 -828
rect -4241 -900 -4235 -866
rect -4201 -900 -4195 -866
rect -4241 -938 -4195 -900
rect -4241 -972 -4235 -938
rect -4201 -972 -4195 -938
rect -4241 -1009 -4195 -972
rect -4093 -146 -4047 -109
rect -4093 -180 -4087 -146
rect -4053 -180 -4047 -146
rect -4093 -218 -4047 -180
rect -4093 -252 -4087 -218
rect -4053 -252 -4047 -218
rect -4093 -290 -4047 -252
rect -4093 -324 -4087 -290
rect -4053 -324 -4047 -290
rect -4093 -362 -4047 -324
rect -4093 -396 -4087 -362
rect -4053 -396 -4047 -362
rect -4093 -434 -4047 -396
rect -4093 -468 -4087 -434
rect -4053 -468 -4047 -434
rect -4093 -506 -4047 -468
rect -4093 -540 -4087 -506
rect -4053 -540 -4047 -506
rect -4093 -578 -4047 -540
rect -4093 -612 -4087 -578
rect -4053 -612 -4047 -578
rect -4093 -650 -4047 -612
rect -4093 -684 -4087 -650
rect -4053 -684 -4047 -650
rect -4093 -722 -4047 -684
rect -4093 -756 -4087 -722
rect -4053 -756 -4047 -722
rect -4093 -794 -4047 -756
rect -4093 -828 -4087 -794
rect -4053 -828 -4047 -794
rect -4093 -866 -4047 -828
rect -4093 -900 -4087 -866
rect -4053 -900 -4047 -866
rect -4093 -938 -4047 -900
rect -4093 -972 -4087 -938
rect -4053 -972 -4047 -938
rect -4093 -1009 -4047 -972
rect -3945 -146 -3899 -109
rect -3945 -180 -3939 -146
rect -3905 -180 -3899 -146
rect -3945 -218 -3899 -180
rect -3945 -252 -3939 -218
rect -3905 -252 -3899 -218
rect -3945 -290 -3899 -252
rect -3945 -324 -3939 -290
rect -3905 -324 -3899 -290
rect -3945 -362 -3899 -324
rect -3945 -396 -3939 -362
rect -3905 -396 -3899 -362
rect -3945 -434 -3899 -396
rect -3945 -468 -3939 -434
rect -3905 -468 -3899 -434
rect -3945 -506 -3899 -468
rect -3945 -540 -3939 -506
rect -3905 -540 -3899 -506
rect -3945 -578 -3899 -540
rect -3945 -612 -3939 -578
rect -3905 -612 -3899 -578
rect -3945 -650 -3899 -612
rect -3945 -684 -3939 -650
rect -3905 -684 -3899 -650
rect -3945 -722 -3899 -684
rect -3945 -756 -3939 -722
rect -3905 -756 -3899 -722
rect -3945 -794 -3899 -756
rect -3945 -828 -3939 -794
rect -3905 -828 -3899 -794
rect -3945 -866 -3899 -828
rect -3945 -900 -3939 -866
rect -3905 -900 -3899 -866
rect -3945 -938 -3899 -900
rect -3945 -972 -3939 -938
rect -3905 -972 -3899 -938
rect -3945 -1009 -3899 -972
rect -3797 -146 -3751 -109
rect -3797 -180 -3791 -146
rect -3757 -180 -3751 -146
rect -3797 -218 -3751 -180
rect -3797 -252 -3791 -218
rect -3757 -252 -3751 -218
rect -3797 -290 -3751 -252
rect -3797 -324 -3791 -290
rect -3757 -324 -3751 -290
rect -3797 -362 -3751 -324
rect -3797 -396 -3791 -362
rect -3757 -396 -3751 -362
rect -3797 -434 -3751 -396
rect -3797 -468 -3791 -434
rect -3757 -468 -3751 -434
rect -3797 -506 -3751 -468
rect -3797 -540 -3791 -506
rect -3757 -540 -3751 -506
rect -3797 -578 -3751 -540
rect -3797 -612 -3791 -578
rect -3757 -612 -3751 -578
rect -3797 -650 -3751 -612
rect -3797 -684 -3791 -650
rect -3757 -684 -3751 -650
rect -3797 -722 -3751 -684
rect -3797 -756 -3791 -722
rect -3757 -756 -3751 -722
rect -3797 -794 -3751 -756
rect -3797 -828 -3791 -794
rect -3757 -828 -3751 -794
rect -3797 -866 -3751 -828
rect -3797 -900 -3791 -866
rect -3757 -900 -3751 -866
rect -3797 -938 -3751 -900
rect -3797 -972 -3791 -938
rect -3757 -972 -3751 -938
rect -3797 -1009 -3751 -972
rect -3649 -146 -3603 -109
rect -3649 -180 -3643 -146
rect -3609 -180 -3603 -146
rect -3649 -218 -3603 -180
rect -3649 -252 -3643 -218
rect -3609 -252 -3603 -218
rect -3649 -290 -3603 -252
rect -3649 -324 -3643 -290
rect -3609 -324 -3603 -290
rect -3649 -362 -3603 -324
rect -3649 -396 -3643 -362
rect -3609 -396 -3603 -362
rect -3649 -434 -3603 -396
rect -3649 -468 -3643 -434
rect -3609 -468 -3603 -434
rect -3649 -506 -3603 -468
rect -3649 -540 -3643 -506
rect -3609 -540 -3603 -506
rect -3649 -578 -3603 -540
rect -3649 -612 -3643 -578
rect -3609 -612 -3603 -578
rect -3649 -650 -3603 -612
rect -3649 -684 -3643 -650
rect -3609 -684 -3603 -650
rect -3649 -722 -3603 -684
rect -3649 -756 -3643 -722
rect -3609 -756 -3603 -722
rect -3649 -794 -3603 -756
rect -3649 -828 -3643 -794
rect -3609 -828 -3603 -794
rect -3649 -866 -3603 -828
rect -3649 -900 -3643 -866
rect -3609 -900 -3603 -866
rect -3649 -938 -3603 -900
rect -3649 -972 -3643 -938
rect -3609 -972 -3603 -938
rect -3649 -1009 -3603 -972
rect -3501 -146 -3455 -109
rect -3501 -180 -3495 -146
rect -3461 -180 -3455 -146
rect -3501 -218 -3455 -180
rect -3501 -252 -3495 -218
rect -3461 -252 -3455 -218
rect -3501 -290 -3455 -252
rect -3501 -324 -3495 -290
rect -3461 -324 -3455 -290
rect -3501 -362 -3455 -324
rect -3501 -396 -3495 -362
rect -3461 -396 -3455 -362
rect -3501 -434 -3455 -396
rect -3501 -468 -3495 -434
rect -3461 -468 -3455 -434
rect -3501 -506 -3455 -468
rect -3501 -540 -3495 -506
rect -3461 -540 -3455 -506
rect -3501 -578 -3455 -540
rect -3501 -612 -3495 -578
rect -3461 -612 -3455 -578
rect -3501 -650 -3455 -612
rect -3501 -684 -3495 -650
rect -3461 -684 -3455 -650
rect -3501 -722 -3455 -684
rect -3501 -756 -3495 -722
rect -3461 -756 -3455 -722
rect -3501 -794 -3455 -756
rect -3501 -828 -3495 -794
rect -3461 -828 -3455 -794
rect -3501 -866 -3455 -828
rect -3501 -900 -3495 -866
rect -3461 -900 -3455 -866
rect -3501 -938 -3455 -900
rect -3501 -972 -3495 -938
rect -3461 -972 -3455 -938
rect -3501 -1009 -3455 -972
rect -3353 -146 -3307 -109
rect -3353 -180 -3347 -146
rect -3313 -180 -3307 -146
rect -3353 -218 -3307 -180
rect -3353 -252 -3347 -218
rect -3313 -252 -3307 -218
rect -3353 -290 -3307 -252
rect -3353 -324 -3347 -290
rect -3313 -324 -3307 -290
rect -3353 -362 -3307 -324
rect -3353 -396 -3347 -362
rect -3313 -396 -3307 -362
rect -3353 -434 -3307 -396
rect -3353 -468 -3347 -434
rect -3313 -468 -3307 -434
rect -3353 -506 -3307 -468
rect -3353 -540 -3347 -506
rect -3313 -540 -3307 -506
rect -3353 -578 -3307 -540
rect -3353 -612 -3347 -578
rect -3313 -612 -3307 -578
rect -3353 -650 -3307 -612
rect -3353 -684 -3347 -650
rect -3313 -684 -3307 -650
rect -3353 -722 -3307 -684
rect -3353 -756 -3347 -722
rect -3313 -756 -3307 -722
rect -3353 -794 -3307 -756
rect -3353 -828 -3347 -794
rect -3313 -828 -3307 -794
rect -3353 -866 -3307 -828
rect -3353 -900 -3347 -866
rect -3313 -900 -3307 -866
rect -3353 -938 -3307 -900
rect -3353 -972 -3347 -938
rect -3313 -972 -3307 -938
rect -3353 -1009 -3307 -972
rect -3205 -146 -3159 -109
rect -3205 -180 -3199 -146
rect -3165 -180 -3159 -146
rect -3205 -218 -3159 -180
rect -3205 -252 -3199 -218
rect -3165 -252 -3159 -218
rect -3205 -290 -3159 -252
rect -3205 -324 -3199 -290
rect -3165 -324 -3159 -290
rect -3205 -362 -3159 -324
rect -3205 -396 -3199 -362
rect -3165 -396 -3159 -362
rect -3205 -434 -3159 -396
rect -3205 -468 -3199 -434
rect -3165 -468 -3159 -434
rect -3205 -506 -3159 -468
rect -3205 -540 -3199 -506
rect -3165 -540 -3159 -506
rect -3205 -578 -3159 -540
rect -3205 -612 -3199 -578
rect -3165 -612 -3159 -578
rect -3205 -650 -3159 -612
rect -3205 -684 -3199 -650
rect -3165 -684 -3159 -650
rect -3205 -722 -3159 -684
rect -3205 -756 -3199 -722
rect -3165 -756 -3159 -722
rect -3205 -794 -3159 -756
rect -3205 -828 -3199 -794
rect -3165 -828 -3159 -794
rect -3205 -866 -3159 -828
rect -3205 -900 -3199 -866
rect -3165 -900 -3159 -866
rect -3205 -938 -3159 -900
rect -3205 -972 -3199 -938
rect -3165 -972 -3159 -938
rect -3205 -1009 -3159 -972
rect -3057 -146 -3011 -109
rect -3057 -180 -3051 -146
rect -3017 -180 -3011 -146
rect -3057 -218 -3011 -180
rect -3057 -252 -3051 -218
rect -3017 -252 -3011 -218
rect -3057 -290 -3011 -252
rect -3057 -324 -3051 -290
rect -3017 -324 -3011 -290
rect -3057 -362 -3011 -324
rect -3057 -396 -3051 -362
rect -3017 -396 -3011 -362
rect -3057 -434 -3011 -396
rect -3057 -468 -3051 -434
rect -3017 -468 -3011 -434
rect -3057 -506 -3011 -468
rect -3057 -540 -3051 -506
rect -3017 -540 -3011 -506
rect -3057 -578 -3011 -540
rect -3057 -612 -3051 -578
rect -3017 -612 -3011 -578
rect -3057 -650 -3011 -612
rect -3057 -684 -3051 -650
rect -3017 -684 -3011 -650
rect -3057 -722 -3011 -684
rect -3057 -756 -3051 -722
rect -3017 -756 -3011 -722
rect -3057 -794 -3011 -756
rect -3057 -828 -3051 -794
rect -3017 -828 -3011 -794
rect -3057 -866 -3011 -828
rect -3057 -900 -3051 -866
rect -3017 -900 -3011 -866
rect -3057 -938 -3011 -900
rect -3057 -972 -3051 -938
rect -3017 -972 -3011 -938
rect -3057 -1009 -3011 -972
rect -2909 -146 -2863 -109
rect -2909 -180 -2903 -146
rect -2869 -180 -2863 -146
rect -2909 -218 -2863 -180
rect -2909 -252 -2903 -218
rect -2869 -252 -2863 -218
rect -2909 -290 -2863 -252
rect -2909 -324 -2903 -290
rect -2869 -324 -2863 -290
rect -2909 -362 -2863 -324
rect -2909 -396 -2903 -362
rect -2869 -396 -2863 -362
rect -2909 -434 -2863 -396
rect -2909 -468 -2903 -434
rect -2869 -468 -2863 -434
rect -2909 -506 -2863 -468
rect -2909 -540 -2903 -506
rect -2869 -540 -2863 -506
rect -2909 -578 -2863 -540
rect -2909 -612 -2903 -578
rect -2869 -612 -2863 -578
rect -2909 -650 -2863 -612
rect -2909 -684 -2903 -650
rect -2869 -684 -2863 -650
rect -2909 -722 -2863 -684
rect -2909 -756 -2903 -722
rect -2869 -756 -2863 -722
rect -2909 -794 -2863 -756
rect -2909 -828 -2903 -794
rect -2869 -828 -2863 -794
rect -2909 -866 -2863 -828
rect -2909 -900 -2903 -866
rect -2869 -900 -2863 -866
rect -2909 -938 -2863 -900
rect -2909 -972 -2903 -938
rect -2869 -972 -2863 -938
rect -2909 -1009 -2863 -972
rect -2761 -146 -2715 -109
rect -2761 -180 -2755 -146
rect -2721 -180 -2715 -146
rect -2761 -218 -2715 -180
rect -2761 -252 -2755 -218
rect -2721 -252 -2715 -218
rect -2761 -290 -2715 -252
rect -2761 -324 -2755 -290
rect -2721 -324 -2715 -290
rect -2761 -362 -2715 -324
rect -2761 -396 -2755 -362
rect -2721 -396 -2715 -362
rect -2761 -434 -2715 -396
rect -2761 -468 -2755 -434
rect -2721 -468 -2715 -434
rect -2761 -506 -2715 -468
rect -2761 -540 -2755 -506
rect -2721 -540 -2715 -506
rect -2761 -578 -2715 -540
rect -2761 -612 -2755 -578
rect -2721 -612 -2715 -578
rect -2761 -650 -2715 -612
rect -2761 -684 -2755 -650
rect -2721 -684 -2715 -650
rect -2761 -722 -2715 -684
rect -2761 -756 -2755 -722
rect -2721 -756 -2715 -722
rect -2761 -794 -2715 -756
rect -2761 -828 -2755 -794
rect -2721 -828 -2715 -794
rect -2761 -866 -2715 -828
rect -2761 -900 -2755 -866
rect -2721 -900 -2715 -866
rect -2761 -938 -2715 -900
rect -2761 -972 -2755 -938
rect -2721 -972 -2715 -938
rect -2761 -1009 -2715 -972
rect -2613 -146 -2567 -109
rect -2613 -180 -2607 -146
rect -2573 -180 -2567 -146
rect -2613 -218 -2567 -180
rect -2613 -252 -2607 -218
rect -2573 -252 -2567 -218
rect -2613 -290 -2567 -252
rect -2613 -324 -2607 -290
rect -2573 -324 -2567 -290
rect -2613 -362 -2567 -324
rect -2613 -396 -2607 -362
rect -2573 -396 -2567 -362
rect -2613 -434 -2567 -396
rect -2613 -468 -2607 -434
rect -2573 -468 -2567 -434
rect -2613 -506 -2567 -468
rect -2613 -540 -2607 -506
rect -2573 -540 -2567 -506
rect -2613 -578 -2567 -540
rect -2613 -612 -2607 -578
rect -2573 -612 -2567 -578
rect -2613 -650 -2567 -612
rect -2613 -684 -2607 -650
rect -2573 -684 -2567 -650
rect -2613 -722 -2567 -684
rect -2613 -756 -2607 -722
rect -2573 -756 -2567 -722
rect -2613 -794 -2567 -756
rect -2613 -828 -2607 -794
rect -2573 -828 -2567 -794
rect -2613 -866 -2567 -828
rect -2613 -900 -2607 -866
rect -2573 -900 -2567 -866
rect -2613 -938 -2567 -900
rect -2613 -972 -2607 -938
rect -2573 -972 -2567 -938
rect -2613 -1009 -2567 -972
rect -2465 -146 -2419 -109
rect -2465 -180 -2459 -146
rect -2425 -180 -2419 -146
rect -2465 -218 -2419 -180
rect -2465 -252 -2459 -218
rect -2425 -252 -2419 -218
rect -2465 -290 -2419 -252
rect -2465 -324 -2459 -290
rect -2425 -324 -2419 -290
rect -2465 -362 -2419 -324
rect -2465 -396 -2459 -362
rect -2425 -396 -2419 -362
rect -2465 -434 -2419 -396
rect -2465 -468 -2459 -434
rect -2425 -468 -2419 -434
rect -2465 -506 -2419 -468
rect -2465 -540 -2459 -506
rect -2425 -540 -2419 -506
rect -2465 -578 -2419 -540
rect -2465 -612 -2459 -578
rect -2425 -612 -2419 -578
rect -2465 -650 -2419 -612
rect -2465 -684 -2459 -650
rect -2425 -684 -2419 -650
rect -2465 -722 -2419 -684
rect -2465 -756 -2459 -722
rect -2425 -756 -2419 -722
rect -2465 -794 -2419 -756
rect -2465 -828 -2459 -794
rect -2425 -828 -2419 -794
rect -2465 -866 -2419 -828
rect -2465 -900 -2459 -866
rect -2425 -900 -2419 -866
rect -2465 -938 -2419 -900
rect -2465 -972 -2459 -938
rect -2425 -972 -2419 -938
rect -2465 -1009 -2419 -972
rect -2317 -146 -2271 -109
rect -2317 -180 -2311 -146
rect -2277 -180 -2271 -146
rect -2317 -218 -2271 -180
rect -2317 -252 -2311 -218
rect -2277 -252 -2271 -218
rect -2317 -290 -2271 -252
rect -2317 -324 -2311 -290
rect -2277 -324 -2271 -290
rect -2317 -362 -2271 -324
rect -2317 -396 -2311 -362
rect -2277 -396 -2271 -362
rect -2317 -434 -2271 -396
rect -2317 -468 -2311 -434
rect -2277 -468 -2271 -434
rect -2317 -506 -2271 -468
rect -2317 -540 -2311 -506
rect -2277 -540 -2271 -506
rect -2317 -578 -2271 -540
rect -2317 -612 -2311 -578
rect -2277 -612 -2271 -578
rect -2317 -650 -2271 -612
rect -2317 -684 -2311 -650
rect -2277 -684 -2271 -650
rect -2317 -722 -2271 -684
rect -2317 -756 -2311 -722
rect -2277 -756 -2271 -722
rect -2317 -794 -2271 -756
rect -2317 -828 -2311 -794
rect -2277 -828 -2271 -794
rect -2317 -866 -2271 -828
rect -2317 -900 -2311 -866
rect -2277 -900 -2271 -866
rect -2317 -938 -2271 -900
rect -2317 -972 -2311 -938
rect -2277 -972 -2271 -938
rect -2317 -1009 -2271 -972
rect -2169 -146 -2123 -109
rect -2169 -180 -2163 -146
rect -2129 -180 -2123 -146
rect -2169 -218 -2123 -180
rect -2169 -252 -2163 -218
rect -2129 -252 -2123 -218
rect -2169 -290 -2123 -252
rect -2169 -324 -2163 -290
rect -2129 -324 -2123 -290
rect -2169 -362 -2123 -324
rect -2169 -396 -2163 -362
rect -2129 -396 -2123 -362
rect -2169 -434 -2123 -396
rect -2169 -468 -2163 -434
rect -2129 -468 -2123 -434
rect -2169 -506 -2123 -468
rect -2169 -540 -2163 -506
rect -2129 -540 -2123 -506
rect -2169 -578 -2123 -540
rect -2169 -612 -2163 -578
rect -2129 -612 -2123 -578
rect -2169 -650 -2123 -612
rect -2169 -684 -2163 -650
rect -2129 -684 -2123 -650
rect -2169 -722 -2123 -684
rect -2169 -756 -2163 -722
rect -2129 -756 -2123 -722
rect -2169 -794 -2123 -756
rect -2169 -828 -2163 -794
rect -2129 -828 -2123 -794
rect -2169 -866 -2123 -828
rect -2169 -900 -2163 -866
rect -2129 -900 -2123 -866
rect -2169 -938 -2123 -900
rect -2169 -972 -2163 -938
rect -2129 -972 -2123 -938
rect -2169 -1009 -2123 -972
rect -2021 -146 -1975 -109
rect -2021 -180 -2015 -146
rect -1981 -180 -1975 -146
rect -2021 -218 -1975 -180
rect -2021 -252 -2015 -218
rect -1981 -252 -1975 -218
rect -2021 -290 -1975 -252
rect -2021 -324 -2015 -290
rect -1981 -324 -1975 -290
rect -2021 -362 -1975 -324
rect -2021 -396 -2015 -362
rect -1981 -396 -1975 -362
rect -2021 -434 -1975 -396
rect -2021 -468 -2015 -434
rect -1981 -468 -1975 -434
rect -2021 -506 -1975 -468
rect -2021 -540 -2015 -506
rect -1981 -540 -1975 -506
rect -2021 -578 -1975 -540
rect -2021 -612 -2015 -578
rect -1981 -612 -1975 -578
rect -2021 -650 -1975 -612
rect -2021 -684 -2015 -650
rect -1981 -684 -1975 -650
rect -2021 -722 -1975 -684
rect -2021 -756 -2015 -722
rect -1981 -756 -1975 -722
rect -2021 -794 -1975 -756
rect -2021 -828 -2015 -794
rect -1981 -828 -1975 -794
rect -2021 -866 -1975 -828
rect -2021 -900 -2015 -866
rect -1981 -900 -1975 -866
rect -2021 -938 -1975 -900
rect -2021 -972 -2015 -938
rect -1981 -972 -1975 -938
rect -2021 -1009 -1975 -972
rect -1873 -146 -1827 -109
rect -1873 -180 -1867 -146
rect -1833 -180 -1827 -146
rect -1873 -218 -1827 -180
rect -1873 -252 -1867 -218
rect -1833 -252 -1827 -218
rect -1873 -290 -1827 -252
rect -1873 -324 -1867 -290
rect -1833 -324 -1827 -290
rect -1873 -362 -1827 -324
rect -1873 -396 -1867 -362
rect -1833 -396 -1827 -362
rect -1873 -434 -1827 -396
rect -1873 -468 -1867 -434
rect -1833 -468 -1827 -434
rect -1873 -506 -1827 -468
rect -1873 -540 -1867 -506
rect -1833 -540 -1827 -506
rect -1873 -578 -1827 -540
rect -1873 -612 -1867 -578
rect -1833 -612 -1827 -578
rect -1873 -650 -1827 -612
rect -1873 -684 -1867 -650
rect -1833 -684 -1827 -650
rect -1873 -722 -1827 -684
rect -1873 -756 -1867 -722
rect -1833 -756 -1827 -722
rect -1873 -794 -1827 -756
rect -1873 -828 -1867 -794
rect -1833 -828 -1827 -794
rect -1873 -866 -1827 -828
rect -1873 -900 -1867 -866
rect -1833 -900 -1827 -866
rect -1873 -938 -1827 -900
rect -1873 -972 -1867 -938
rect -1833 -972 -1827 -938
rect -1873 -1009 -1827 -972
rect -1725 -146 -1679 -109
rect -1725 -180 -1719 -146
rect -1685 -180 -1679 -146
rect -1725 -218 -1679 -180
rect -1725 -252 -1719 -218
rect -1685 -252 -1679 -218
rect -1725 -290 -1679 -252
rect -1725 -324 -1719 -290
rect -1685 -324 -1679 -290
rect -1725 -362 -1679 -324
rect -1725 -396 -1719 -362
rect -1685 -396 -1679 -362
rect -1725 -434 -1679 -396
rect -1725 -468 -1719 -434
rect -1685 -468 -1679 -434
rect -1725 -506 -1679 -468
rect -1725 -540 -1719 -506
rect -1685 -540 -1679 -506
rect -1725 -578 -1679 -540
rect -1725 -612 -1719 -578
rect -1685 -612 -1679 -578
rect -1725 -650 -1679 -612
rect -1725 -684 -1719 -650
rect -1685 -684 -1679 -650
rect -1725 -722 -1679 -684
rect -1725 -756 -1719 -722
rect -1685 -756 -1679 -722
rect -1725 -794 -1679 -756
rect -1725 -828 -1719 -794
rect -1685 -828 -1679 -794
rect -1725 -866 -1679 -828
rect -1725 -900 -1719 -866
rect -1685 -900 -1679 -866
rect -1725 -938 -1679 -900
rect -1725 -972 -1719 -938
rect -1685 -972 -1679 -938
rect -1725 -1009 -1679 -972
rect -1577 -146 -1531 -109
rect -1577 -180 -1571 -146
rect -1537 -180 -1531 -146
rect -1577 -218 -1531 -180
rect -1577 -252 -1571 -218
rect -1537 -252 -1531 -218
rect -1577 -290 -1531 -252
rect -1577 -324 -1571 -290
rect -1537 -324 -1531 -290
rect -1577 -362 -1531 -324
rect -1577 -396 -1571 -362
rect -1537 -396 -1531 -362
rect -1577 -434 -1531 -396
rect -1577 -468 -1571 -434
rect -1537 -468 -1531 -434
rect -1577 -506 -1531 -468
rect -1577 -540 -1571 -506
rect -1537 -540 -1531 -506
rect -1577 -578 -1531 -540
rect -1577 -612 -1571 -578
rect -1537 -612 -1531 -578
rect -1577 -650 -1531 -612
rect -1577 -684 -1571 -650
rect -1537 -684 -1531 -650
rect -1577 -722 -1531 -684
rect -1577 -756 -1571 -722
rect -1537 -756 -1531 -722
rect -1577 -794 -1531 -756
rect -1577 -828 -1571 -794
rect -1537 -828 -1531 -794
rect -1577 -866 -1531 -828
rect -1577 -900 -1571 -866
rect -1537 -900 -1531 -866
rect -1577 -938 -1531 -900
rect -1577 -972 -1571 -938
rect -1537 -972 -1531 -938
rect -1577 -1009 -1531 -972
rect -1429 -146 -1383 -109
rect -1429 -180 -1423 -146
rect -1389 -180 -1383 -146
rect -1429 -218 -1383 -180
rect -1429 -252 -1423 -218
rect -1389 -252 -1383 -218
rect -1429 -290 -1383 -252
rect -1429 -324 -1423 -290
rect -1389 -324 -1383 -290
rect -1429 -362 -1383 -324
rect -1429 -396 -1423 -362
rect -1389 -396 -1383 -362
rect -1429 -434 -1383 -396
rect -1429 -468 -1423 -434
rect -1389 -468 -1383 -434
rect -1429 -506 -1383 -468
rect -1429 -540 -1423 -506
rect -1389 -540 -1383 -506
rect -1429 -578 -1383 -540
rect -1429 -612 -1423 -578
rect -1389 -612 -1383 -578
rect -1429 -650 -1383 -612
rect -1429 -684 -1423 -650
rect -1389 -684 -1383 -650
rect -1429 -722 -1383 -684
rect -1429 -756 -1423 -722
rect -1389 -756 -1383 -722
rect -1429 -794 -1383 -756
rect -1429 -828 -1423 -794
rect -1389 -828 -1383 -794
rect -1429 -866 -1383 -828
rect -1429 -900 -1423 -866
rect -1389 -900 -1383 -866
rect -1429 -938 -1383 -900
rect -1429 -972 -1423 -938
rect -1389 -972 -1383 -938
rect -1429 -1009 -1383 -972
rect -1281 -146 -1235 -109
rect -1281 -180 -1275 -146
rect -1241 -180 -1235 -146
rect -1281 -218 -1235 -180
rect -1281 -252 -1275 -218
rect -1241 -252 -1235 -218
rect -1281 -290 -1235 -252
rect -1281 -324 -1275 -290
rect -1241 -324 -1235 -290
rect -1281 -362 -1235 -324
rect -1281 -396 -1275 -362
rect -1241 -396 -1235 -362
rect -1281 -434 -1235 -396
rect -1281 -468 -1275 -434
rect -1241 -468 -1235 -434
rect -1281 -506 -1235 -468
rect -1281 -540 -1275 -506
rect -1241 -540 -1235 -506
rect -1281 -578 -1235 -540
rect -1281 -612 -1275 -578
rect -1241 -612 -1235 -578
rect -1281 -650 -1235 -612
rect -1281 -684 -1275 -650
rect -1241 -684 -1235 -650
rect -1281 -722 -1235 -684
rect -1281 -756 -1275 -722
rect -1241 -756 -1235 -722
rect -1281 -794 -1235 -756
rect -1281 -828 -1275 -794
rect -1241 -828 -1235 -794
rect -1281 -866 -1235 -828
rect -1281 -900 -1275 -866
rect -1241 -900 -1235 -866
rect -1281 -938 -1235 -900
rect -1281 -972 -1275 -938
rect -1241 -972 -1235 -938
rect -1281 -1009 -1235 -972
rect -1133 -146 -1087 -109
rect -1133 -180 -1127 -146
rect -1093 -180 -1087 -146
rect -1133 -218 -1087 -180
rect -1133 -252 -1127 -218
rect -1093 -252 -1087 -218
rect -1133 -290 -1087 -252
rect -1133 -324 -1127 -290
rect -1093 -324 -1087 -290
rect -1133 -362 -1087 -324
rect -1133 -396 -1127 -362
rect -1093 -396 -1087 -362
rect -1133 -434 -1087 -396
rect -1133 -468 -1127 -434
rect -1093 -468 -1087 -434
rect -1133 -506 -1087 -468
rect -1133 -540 -1127 -506
rect -1093 -540 -1087 -506
rect -1133 -578 -1087 -540
rect -1133 -612 -1127 -578
rect -1093 -612 -1087 -578
rect -1133 -650 -1087 -612
rect -1133 -684 -1127 -650
rect -1093 -684 -1087 -650
rect -1133 -722 -1087 -684
rect -1133 -756 -1127 -722
rect -1093 -756 -1087 -722
rect -1133 -794 -1087 -756
rect -1133 -828 -1127 -794
rect -1093 -828 -1087 -794
rect -1133 -866 -1087 -828
rect -1133 -900 -1127 -866
rect -1093 -900 -1087 -866
rect -1133 -938 -1087 -900
rect -1133 -972 -1127 -938
rect -1093 -972 -1087 -938
rect -1133 -1009 -1087 -972
rect -985 -146 -939 -109
rect -985 -180 -979 -146
rect -945 -180 -939 -146
rect -985 -218 -939 -180
rect -985 -252 -979 -218
rect -945 -252 -939 -218
rect -985 -290 -939 -252
rect -985 -324 -979 -290
rect -945 -324 -939 -290
rect -985 -362 -939 -324
rect -985 -396 -979 -362
rect -945 -396 -939 -362
rect -985 -434 -939 -396
rect -985 -468 -979 -434
rect -945 -468 -939 -434
rect -985 -506 -939 -468
rect -985 -540 -979 -506
rect -945 -540 -939 -506
rect -985 -578 -939 -540
rect -985 -612 -979 -578
rect -945 -612 -939 -578
rect -985 -650 -939 -612
rect -985 -684 -979 -650
rect -945 -684 -939 -650
rect -985 -722 -939 -684
rect -985 -756 -979 -722
rect -945 -756 -939 -722
rect -985 -794 -939 -756
rect -985 -828 -979 -794
rect -945 -828 -939 -794
rect -985 -866 -939 -828
rect -985 -900 -979 -866
rect -945 -900 -939 -866
rect -985 -938 -939 -900
rect -985 -972 -979 -938
rect -945 -972 -939 -938
rect -985 -1009 -939 -972
rect -837 -146 -791 -109
rect -837 -180 -831 -146
rect -797 -180 -791 -146
rect -837 -218 -791 -180
rect -837 -252 -831 -218
rect -797 -252 -791 -218
rect -837 -290 -791 -252
rect -837 -324 -831 -290
rect -797 -324 -791 -290
rect -837 -362 -791 -324
rect -837 -396 -831 -362
rect -797 -396 -791 -362
rect -837 -434 -791 -396
rect -837 -468 -831 -434
rect -797 -468 -791 -434
rect -837 -506 -791 -468
rect -837 -540 -831 -506
rect -797 -540 -791 -506
rect -837 -578 -791 -540
rect -837 -612 -831 -578
rect -797 -612 -791 -578
rect -837 -650 -791 -612
rect -837 -684 -831 -650
rect -797 -684 -791 -650
rect -837 -722 -791 -684
rect -837 -756 -831 -722
rect -797 -756 -791 -722
rect -837 -794 -791 -756
rect -837 -828 -831 -794
rect -797 -828 -791 -794
rect -837 -866 -791 -828
rect -837 -900 -831 -866
rect -797 -900 -791 -866
rect -837 -938 -791 -900
rect -837 -972 -831 -938
rect -797 -972 -791 -938
rect -837 -1009 -791 -972
rect -689 -146 -643 -109
rect -689 -180 -683 -146
rect -649 -180 -643 -146
rect -689 -218 -643 -180
rect -689 -252 -683 -218
rect -649 -252 -643 -218
rect -689 -290 -643 -252
rect -689 -324 -683 -290
rect -649 -324 -643 -290
rect -689 -362 -643 -324
rect -689 -396 -683 -362
rect -649 -396 -643 -362
rect -689 -434 -643 -396
rect -689 -468 -683 -434
rect -649 -468 -643 -434
rect -689 -506 -643 -468
rect -689 -540 -683 -506
rect -649 -540 -643 -506
rect -689 -578 -643 -540
rect -689 -612 -683 -578
rect -649 -612 -643 -578
rect -689 -650 -643 -612
rect -689 -684 -683 -650
rect -649 -684 -643 -650
rect -689 -722 -643 -684
rect -689 -756 -683 -722
rect -649 -756 -643 -722
rect -689 -794 -643 -756
rect -689 -828 -683 -794
rect -649 -828 -643 -794
rect -689 -866 -643 -828
rect -689 -900 -683 -866
rect -649 -900 -643 -866
rect -689 -938 -643 -900
rect -689 -972 -683 -938
rect -649 -972 -643 -938
rect -689 -1009 -643 -972
rect -541 -146 -495 -109
rect -541 -180 -535 -146
rect -501 -180 -495 -146
rect -541 -218 -495 -180
rect -541 -252 -535 -218
rect -501 -252 -495 -218
rect -541 -290 -495 -252
rect -541 -324 -535 -290
rect -501 -324 -495 -290
rect -541 -362 -495 -324
rect -541 -396 -535 -362
rect -501 -396 -495 -362
rect -541 -434 -495 -396
rect -541 -468 -535 -434
rect -501 -468 -495 -434
rect -541 -506 -495 -468
rect -541 -540 -535 -506
rect -501 -540 -495 -506
rect -541 -578 -495 -540
rect -541 -612 -535 -578
rect -501 -612 -495 -578
rect -541 -650 -495 -612
rect -541 -684 -535 -650
rect -501 -684 -495 -650
rect -541 -722 -495 -684
rect -541 -756 -535 -722
rect -501 -756 -495 -722
rect -541 -794 -495 -756
rect -541 -828 -535 -794
rect -501 -828 -495 -794
rect -541 -866 -495 -828
rect -541 -900 -535 -866
rect -501 -900 -495 -866
rect -541 -938 -495 -900
rect -541 -972 -535 -938
rect -501 -972 -495 -938
rect -541 -1009 -495 -972
rect -393 -146 -347 -109
rect -393 -180 -387 -146
rect -353 -180 -347 -146
rect -393 -218 -347 -180
rect -393 -252 -387 -218
rect -353 -252 -347 -218
rect -393 -290 -347 -252
rect -393 -324 -387 -290
rect -353 -324 -347 -290
rect -393 -362 -347 -324
rect -393 -396 -387 -362
rect -353 -396 -347 -362
rect -393 -434 -347 -396
rect -393 -468 -387 -434
rect -353 -468 -347 -434
rect -393 -506 -347 -468
rect -393 -540 -387 -506
rect -353 -540 -347 -506
rect -393 -578 -347 -540
rect -393 -612 -387 -578
rect -353 -612 -347 -578
rect -393 -650 -347 -612
rect -393 -684 -387 -650
rect -353 -684 -347 -650
rect -393 -722 -347 -684
rect -393 -756 -387 -722
rect -353 -756 -347 -722
rect -393 -794 -347 -756
rect -393 -828 -387 -794
rect -353 -828 -347 -794
rect -393 -866 -347 -828
rect -393 -900 -387 -866
rect -353 -900 -347 -866
rect -393 -938 -347 -900
rect -393 -972 -387 -938
rect -353 -972 -347 -938
rect -393 -1009 -347 -972
rect -245 -146 -199 -109
rect -245 -180 -239 -146
rect -205 -180 -199 -146
rect -245 -218 -199 -180
rect -245 -252 -239 -218
rect -205 -252 -199 -218
rect -245 -290 -199 -252
rect -245 -324 -239 -290
rect -205 -324 -199 -290
rect -245 -362 -199 -324
rect -245 -396 -239 -362
rect -205 -396 -199 -362
rect -245 -434 -199 -396
rect -245 -468 -239 -434
rect -205 -468 -199 -434
rect -245 -506 -199 -468
rect -245 -540 -239 -506
rect -205 -540 -199 -506
rect -245 -578 -199 -540
rect -245 -612 -239 -578
rect -205 -612 -199 -578
rect -245 -650 -199 -612
rect -245 -684 -239 -650
rect -205 -684 -199 -650
rect -245 -722 -199 -684
rect -245 -756 -239 -722
rect -205 -756 -199 -722
rect -245 -794 -199 -756
rect -245 -828 -239 -794
rect -205 -828 -199 -794
rect -245 -866 -199 -828
rect -245 -900 -239 -866
rect -205 -900 -199 -866
rect -245 -938 -199 -900
rect -245 -972 -239 -938
rect -205 -972 -199 -938
rect -245 -1009 -199 -972
rect -97 -146 -51 -109
rect -97 -180 -91 -146
rect -57 -180 -51 -146
rect -97 -218 -51 -180
rect -97 -252 -91 -218
rect -57 -252 -51 -218
rect -97 -290 -51 -252
rect -97 -324 -91 -290
rect -57 -324 -51 -290
rect -97 -362 -51 -324
rect -97 -396 -91 -362
rect -57 -396 -51 -362
rect -97 -434 -51 -396
rect -97 -468 -91 -434
rect -57 -468 -51 -434
rect -97 -506 -51 -468
rect -97 -540 -91 -506
rect -57 -540 -51 -506
rect -97 -578 -51 -540
rect -97 -612 -91 -578
rect -57 -612 -51 -578
rect -97 -650 -51 -612
rect -97 -684 -91 -650
rect -57 -684 -51 -650
rect -97 -722 -51 -684
rect -97 -756 -91 -722
rect -57 -756 -51 -722
rect -97 -794 -51 -756
rect -97 -828 -91 -794
rect -57 -828 -51 -794
rect -97 -866 -51 -828
rect -97 -900 -91 -866
rect -57 -900 -51 -866
rect -97 -938 -51 -900
rect -97 -972 -91 -938
rect -57 -972 -51 -938
rect -97 -1009 -51 -972
rect 51 -146 97 -109
rect 51 -180 57 -146
rect 91 -180 97 -146
rect 51 -218 97 -180
rect 51 -252 57 -218
rect 91 -252 97 -218
rect 51 -290 97 -252
rect 51 -324 57 -290
rect 91 -324 97 -290
rect 51 -362 97 -324
rect 51 -396 57 -362
rect 91 -396 97 -362
rect 51 -434 97 -396
rect 51 -468 57 -434
rect 91 -468 97 -434
rect 51 -506 97 -468
rect 51 -540 57 -506
rect 91 -540 97 -506
rect 51 -578 97 -540
rect 51 -612 57 -578
rect 91 -612 97 -578
rect 51 -650 97 -612
rect 51 -684 57 -650
rect 91 -684 97 -650
rect 51 -722 97 -684
rect 51 -756 57 -722
rect 91 -756 97 -722
rect 51 -794 97 -756
rect 51 -828 57 -794
rect 91 -828 97 -794
rect 51 -866 97 -828
rect 51 -900 57 -866
rect 91 -900 97 -866
rect 51 -938 97 -900
rect 51 -972 57 -938
rect 91 -972 97 -938
rect 51 -1009 97 -972
rect 199 -146 245 -109
rect 199 -180 205 -146
rect 239 -180 245 -146
rect 199 -218 245 -180
rect 199 -252 205 -218
rect 239 -252 245 -218
rect 199 -290 245 -252
rect 199 -324 205 -290
rect 239 -324 245 -290
rect 199 -362 245 -324
rect 199 -396 205 -362
rect 239 -396 245 -362
rect 199 -434 245 -396
rect 199 -468 205 -434
rect 239 -468 245 -434
rect 199 -506 245 -468
rect 199 -540 205 -506
rect 239 -540 245 -506
rect 199 -578 245 -540
rect 199 -612 205 -578
rect 239 -612 245 -578
rect 199 -650 245 -612
rect 199 -684 205 -650
rect 239 -684 245 -650
rect 199 -722 245 -684
rect 199 -756 205 -722
rect 239 -756 245 -722
rect 199 -794 245 -756
rect 199 -828 205 -794
rect 239 -828 245 -794
rect 199 -866 245 -828
rect 199 -900 205 -866
rect 239 -900 245 -866
rect 199 -938 245 -900
rect 199 -972 205 -938
rect 239 -972 245 -938
rect 199 -1009 245 -972
rect 347 -146 393 -109
rect 347 -180 353 -146
rect 387 -180 393 -146
rect 347 -218 393 -180
rect 347 -252 353 -218
rect 387 -252 393 -218
rect 347 -290 393 -252
rect 347 -324 353 -290
rect 387 -324 393 -290
rect 347 -362 393 -324
rect 347 -396 353 -362
rect 387 -396 393 -362
rect 347 -434 393 -396
rect 347 -468 353 -434
rect 387 -468 393 -434
rect 347 -506 393 -468
rect 347 -540 353 -506
rect 387 -540 393 -506
rect 347 -578 393 -540
rect 347 -612 353 -578
rect 387 -612 393 -578
rect 347 -650 393 -612
rect 347 -684 353 -650
rect 387 -684 393 -650
rect 347 -722 393 -684
rect 347 -756 353 -722
rect 387 -756 393 -722
rect 347 -794 393 -756
rect 347 -828 353 -794
rect 387 -828 393 -794
rect 347 -866 393 -828
rect 347 -900 353 -866
rect 387 -900 393 -866
rect 347 -938 393 -900
rect 347 -972 353 -938
rect 387 -972 393 -938
rect 347 -1009 393 -972
rect 495 -146 541 -109
rect 495 -180 501 -146
rect 535 -180 541 -146
rect 495 -218 541 -180
rect 495 -252 501 -218
rect 535 -252 541 -218
rect 495 -290 541 -252
rect 495 -324 501 -290
rect 535 -324 541 -290
rect 495 -362 541 -324
rect 495 -396 501 -362
rect 535 -396 541 -362
rect 495 -434 541 -396
rect 495 -468 501 -434
rect 535 -468 541 -434
rect 495 -506 541 -468
rect 495 -540 501 -506
rect 535 -540 541 -506
rect 495 -578 541 -540
rect 495 -612 501 -578
rect 535 -612 541 -578
rect 495 -650 541 -612
rect 495 -684 501 -650
rect 535 -684 541 -650
rect 495 -722 541 -684
rect 495 -756 501 -722
rect 535 -756 541 -722
rect 495 -794 541 -756
rect 495 -828 501 -794
rect 535 -828 541 -794
rect 495 -866 541 -828
rect 495 -900 501 -866
rect 535 -900 541 -866
rect 495 -938 541 -900
rect 495 -972 501 -938
rect 535 -972 541 -938
rect 495 -1009 541 -972
rect 643 -146 689 -109
rect 643 -180 649 -146
rect 683 -180 689 -146
rect 643 -218 689 -180
rect 643 -252 649 -218
rect 683 -252 689 -218
rect 643 -290 689 -252
rect 643 -324 649 -290
rect 683 -324 689 -290
rect 643 -362 689 -324
rect 643 -396 649 -362
rect 683 -396 689 -362
rect 643 -434 689 -396
rect 643 -468 649 -434
rect 683 -468 689 -434
rect 643 -506 689 -468
rect 643 -540 649 -506
rect 683 -540 689 -506
rect 643 -578 689 -540
rect 643 -612 649 -578
rect 683 -612 689 -578
rect 643 -650 689 -612
rect 643 -684 649 -650
rect 683 -684 689 -650
rect 643 -722 689 -684
rect 643 -756 649 -722
rect 683 -756 689 -722
rect 643 -794 689 -756
rect 643 -828 649 -794
rect 683 -828 689 -794
rect 643 -866 689 -828
rect 643 -900 649 -866
rect 683 -900 689 -866
rect 643 -938 689 -900
rect 643 -972 649 -938
rect 683 -972 689 -938
rect 643 -1009 689 -972
rect 791 -146 837 -109
rect 791 -180 797 -146
rect 831 -180 837 -146
rect 791 -218 837 -180
rect 791 -252 797 -218
rect 831 -252 837 -218
rect 791 -290 837 -252
rect 791 -324 797 -290
rect 831 -324 837 -290
rect 791 -362 837 -324
rect 791 -396 797 -362
rect 831 -396 837 -362
rect 791 -434 837 -396
rect 791 -468 797 -434
rect 831 -468 837 -434
rect 791 -506 837 -468
rect 791 -540 797 -506
rect 831 -540 837 -506
rect 791 -578 837 -540
rect 791 -612 797 -578
rect 831 -612 837 -578
rect 791 -650 837 -612
rect 791 -684 797 -650
rect 831 -684 837 -650
rect 791 -722 837 -684
rect 791 -756 797 -722
rect 831 -756 837 -722
rect 791 -794 837 -756
rect 791 -828 797 -794
rect 831 -828 837 -794
rect 791 -866 837 -828
rect 791 -900 797 -866
rect 831 -900 837 -866
rect 791 -938 837 -900
rect 791 -972 797 -938
rect 831 -972 837 -938
rect 791 -1009 837 -972
rect 939 -146 985 -109
rect 939 -180 945 -146
rect 979 -180 985 -146
rect 939 -218 985 -180
rect 939 -252 945 -218
rect 979 -252 985 -218
rect 939 -290 985 -252
rect 939 -324 945 -290
rect 979 -324 985 -290
rect 939 -362 985 -324
rect 939 -396 945 -362
rect 979 -396 985 -362
rect 939 -434 985 -396
rect 939 -468 945 -434
rect 979 -468 985 -434
rect 939 -506 985 -468
rect 939 -540 945 -506
rect 979 -540 985 -506
rect 939 -578 985 -540
rect 939 -612 945 -578
rect 979 -612 985 -578
rect 939 -650 985 -612
rect 939 -684 945 -650
rect 979 -684 985 -650
rect 939 -722 985 -684
rect 939 -756 945 -722
rect 979 -756 985 -722
rect 939 -794 985 -756
rect 939 -828 945 -794
rect 979 -828 985 -794
rect 939 -866 985 -828
rect 939 -900 945 -866
rect 979 -900 985 -866
rect 939 -938 985 -900
rect 939 -972 945 -938
rect 979 -972 985 -938
rect 939 -1009 985 -972
rect 1087 -146 1133 -109
rect 1087 -180 1093 -146
rect 1127 -180 1133 -146
rect 1087 -218 1133 -180
rect 1087 -252 1093 -218
rect 1127 -252 1133 -218
rect 1087 -290 1133 -252
rect 1087 -324 1093 -290
rect 1127 -324 1133 -290
rect 1087 -362 1133 -324
rect 1087 -396 1093 -362
rect 1127 -396 1133 -362
rect 1087 -434 1133 -396
rect 1087 -468 1093 -434
rect 1127 -468 1133 -434
rect 1087 -506 1133 -468
rect 1087 -540 1093 -506
rect 1127 -540 1133 -506
rect 1087 -578 1133 -540
rect 1087 -612 1093 -578
rect 1127 -612 1133 -578
rect 1087 -650 1133 -612
rect 1087 -684 1093 -650
rect 1127 -684 1133 -650
rect 1087 -722 1133 -684
rect 1087 -756 1093 -722
rect 1127 -756 1133 -722
rect 1087 -794 1133 -756
rect 1087 -828 1093 -794
rect 1127 -828 1133 -794
rect 1087 -866 1133 -828
rect 1087 -900 1093 -866
rect 1127 -900 1133 -866
rect 1087 -938 1133 -900
rect 1087 -972 1093 -938
rect 1127 -972 1133 -938
rect 1087 -1009 1133 -972
rect 1235 -146 1281 -109
rect 1235 -180 1241 -146
rect 1275 -180 1281 -146
rect 1235 -218 1281 -180
rect 1235 -252 1241 -218
rect 1275 -252 1281 -218
rect 1235 -290 1281 -252
rect 1235 -324 1241 -290
rect 1275 -324 1281 -290
rect 1235 -362 1281 -324
rect 1235 -396 1241 -362
rect 1275 -396 1281 -362
rect 1235 -434 1281 -396
rect 1235 -468 1241 -434
rect 1275 -468 1281 -434
rect 1235 -506 1281 -468
rect 1235 -540 1241 -506
rect 1275 -540 1281 -506
rect 1235 -578 1281 -540
rect 1235 -612 1241 -578
rect 1275 -612 1281 -578
rect 1235 -650 1281 -612
rect 1235 -684 1241 -650
rect 1275 -684 1281 -650
rect 1235 -722 1281 -684
rect 1235 -756 1241 -722
rect 1275 -756 1281 -722
rect 1235 -794 1281 -756
rect 1235 -828 1241 -794
rect 1275 -828 1281 -794
rect 1235 -866 1281 -828
rect 1235 -900 1241 -866
rect 1275 -900 1281 -866
rect 1235 -938 1281 -900
rect 1235 -972 1241 -938
rect 1275 -972 1281 -938
rect 1235 -1009 1281 -972
rect 1383 -146 1429 -109
rect 1383 -180 1389 -146
rect 1423 -180 1429 -146
rect 1383 -218 1429 -180
rect 1383 -252 1389 -218
rect 1423 -252 1429 -218
rect 1383 -290 1429 -252
rect 1383 -324 1389 -290
rect 1423 -324 1429 -290
rect 1383 -362 1429 -324
rect 1383 -396 1389 -362
rect 1423 -396 1429 -362
rect 1383 -434 1429 -396
rect 1383 -468 1389 -434
rect 1423 -468 1429 -434
rect 1383 -506 1429 -468
rect 1383 -540 1389 -506
rect 1423 -540 1429 -506
rect 1383 -578 1429 -540
rect 1383 -612 1389 -578
rect 1423 -612 1429 -578
rect 1383 -650 1429 -612
rect 1383 -684 1389 -650
rect 1423 -684 1429 -650
rect 1383 -722 1429 -684
rect 1383 -756 1389 -722
rect 1423 -756 1429 -722
rect 1383 -794 1429 -756
rect 1383 -828 1389 -794
rect 1423 -828 1429 -794
rect 1383 -866 1429 -828
rect 1383 -900 1389 -866
rect 1423 -900 1429 -866
rect 1383 -938 1429 -900
rect 1383 -972 1389 -938
rect 1423 -972 1429 -938
rect 1383 -1009 1429 -972
rect 1531 -146 1577 -109
rect 1531 -180 1537 -146
rect 1571 -180 1577 -146
rect 1531 -218 1577 -180
rect 1531 -252 1537 -218
rect 1571 -252 1577 -218
rect 1531 -290 1577 -252
rect 1531 -324 1537 -290
rect 1571 -324 1577 -290
rect 1531 -362 1577 -324
rect 1531 -396 1537 -362
rect 1571 -396 1577 -362
rect 1531 -434 1577 -396
rect 1531 -468 1537 -434
rect 1571 -468 1577 -434
rect 1531 -506 1577 -468
rect 1531 -540 1537 -506
rect 1571 -540 1577 -506
rect 1531 -578 1577 -540
rect 1531 -612 1537 -578
rect 1571 -612 1577 -578
rect 1531 -650 1577 -612
rect 1531 -684 1537 -650
rect 1571 -684 1577 -650
rect 1531 -722 1577 -684
rect 1531 -756 1537 -722
rect 1571 -756 1577 -722
rect 1531 -794 1577 -756
rect 1531 -828 1537 -794
rect 1571 -828 1577 -794
rect 1531 -866 1577 -828
rect 1531 -900 1537 -866
rect 1571 -900 1577 -866
rect 1531 -938 1577 -900
rect 1531 -972 1537 -938
rect 1571 -972 1577 -938
rect 1531 -1009 1577 -972
rect 1679 -146 1725 -109
rect 1679 -180 1685 -146
rect 1719 -180 1725 -146
rect 1679 -218 1725 -180
rect 1679 -252 1685 -218
rect 1719 -252 1725 -218
rect 1679 -290 1725 -252
rect 1679 -324 1685 -290
rect 1719 -324 1725 -290
rect 1679 -362 1725 -324
rect 1679 -396 1685 -362
rect 1719 -396 1725 -362
rect 1679 -434 1725 -396
rect 1679 -468 1685 -434
rect 1719 -468 1725 -434
rect 1679 -506 1725 -468
rect 1679 -540 1685 -506
rect 1719 -540 1725 -506
rect 1679 -578 1725 -540
rect 1679 -612 1685 -578
rect 1719 -612 1725 -578
rect 1679 -650 1725 -612
rect 1679 -684 1685 -650
rect 1719 -684 1725 -650
rect 1679 -722 1725 -684
rect 1679 -756 1685 -722
rect 1719 -756 1725 -722
rect 1679 -794 1725 -756
rect 1679 -828 1685 -794
rect 1719 -828 1725 -794
rect 1679 -866 1725 -828
rect 1679 -900 1685 -866
rect 1719 -900 1725 -866
rect 1679 -938 1725 -900
rect 1679 -972 1685 -938
rect 1719 -972 1725 -938
rect 1679 -1009 1725 -972
rect 1827 -146 1873 -109
rect 1827 -180 1833 -146
rect 1867 -180 1873 -146
rect 1827 -218 1873 -180
rect 1827 -252 1833 -218
rect 1867 -252 1873 -218
rect 1827 -290 1873 -252
rect 1827 -324 1833 -290
rect 1867 -324 1873 -290
rect 1827 -362 1873 -324
rect 1827 -396 1833 -362
rect 1867 -396 1873 -362
rect 1827 -434 1873 -396
rect 1827 -468 1833 -434
rect 1867 -468 1873 -434
rect 1827 -506 1873 -468
rect 1827 -540 1833 -506
rect 1867 -540 1873 -506
rect 1827 -578 1873 -540
rect 1827 -612 1833 -578
rect 1867 -612 1873 -578
rect 1827 -650 1873 -612
rect 1827 -684 1833 -650
rect 1867 -684 1873 -650
rect 1827 -722 1873 -684
rect 1827 -756 1833 -722
rect 1867 -756 1873 -722
rect 1827 -794 1873 -756
rect 1827 -828 1833 -794
rect 1867 -828 1873 -794
rect 1827 -866 1873 -828
rect 1827 -900 1833 -866
rect 1867 -900 1873 -866
rect 1827 -938 1873 -900
rect 1827 -972 1833 -938
rect 1867 -972 1873 -938
rect 1827 -1009 1873 -972
rect 1975 -146 2021 -109
rect 1975 -180 1981 -146
rect 2015 -180 2021 -146
rect 1975 -218 2021 -180
rect 1975 -252 1981 -218
rect 2015 -252 2021 -218
rect 1975 -290 2021 -252
rect 1975 -324 1981 -290
rect 2015 -324 2021 -290
rect 1975 -362 2021 -324
rect 1975 -396 1981 -362
rect 2015 -396 2021 -362
rect 1975 -434 2021 -396
rect 1975 -468 1981 -434
rect 2015 -468 2021 -434
rect 1975 -506 2021 -468
rect 1975 -540 1981 -506
rect 2015 -540 2021 -506
rect 1975 -578 2021 -540
rect 1975 -612 1981 -578
rect 2015 -612 2021 -578
rect 1975 -650 2021 -612
rect 1975 -684 1981 -650
rect 2015 -684 2021 -650
rect 1975 -722 2021 -684
rect 1975 -756 1981 -722
rect 2015 -756 2021 -722
rect 1975 -794 2021 -756
rect 1975 -828 1981 -794
rect 2015 -828 2021 -794
rect 1975 -866 2021 -828
rect 1975 -900 1981 -866
rect 2015 -900 2021 -866
rect 1975 -938 2021 -900
rect 1975 -972 1981 -938
rect 2015 -972 2021 -938
rect 1975 -1009 2021 -972
rect 2123 -146 2169 -109
rect 2123 -180 2129 -146
rect 2163 -180 2169 -146
rect 2123 -218 2169 -180
rect 2123 -252 2129 -218
rect 2163 -252 2169 -218
rect 2123 -290 2169 -252
rect 2123 -324 2129 -290
rect 2163 -324 2169 -290
rect 2123 -362 2169 -324
rect 2123 -396 2129 -362
rect 2163 -396 2169 -362
rect 2123 -434 2169 -396
rect 2123 -468 2129 -434
rect 2163 -468 2169 -434
rect 2123 -506 2169 -468
rect 2123 -540 2129 -506
rect 2163 -540 2169 -506
rect 2123 -578 2169 -540
rect 2123 -612 2129 -578
rect 2163 -612 2169 -578
rect 2123 -650 2169 -612
rect 2123 -684 2129 -650
rect 2163 -684 2169 -650
rect 2123 -722 2169 -684
rect 2123 -756 2129 -722
rect 2163 -756 2169 -722
rect 2123 -794 2169 -756
rect 2123 -828 2129 -794
rect 2163 -828 2169 -794
rect 2123 -866 2169 -828
rect 2123 -900 2129 -866
rect 2163 -900 2169 -866
rect 2123 -938 2169 -900
rect 2123 -972 2129 -938
rect 2163 -972 2169 -938
rect 2123 -1009 2169 -972
rect 2271 -146 2317 -109
rect 2271 -180 2277 -146
rect 2311 -180 2317 -146
rect 2271 -218 2317 -180
rect 2271 -252 2277 -218
rect 2311 -252 2317 -218
rect 2271 -290 2317 -252
rect 2271 -324 2277 -290
rect 2311 -324 2317 -290
rect 2271 -362 2317 -324
rect 2271 -396 2277 -362
rect 2311 -396 2317 -362
rect 2271 -434 2317 -396
rect 2271 -468 2277 -434
rect 2311 -468 2317 -434
rect 2271 -506 2317 -468
rect 2271 -540 2277 -506
rect 2311 -540 2317 -506
rect 2271 -578 2317 -540
rect 2271 -612 2277 -578
rect 2311 -612 2317 -578
rect 2271 -650 2317 -612
rect 2271 -684 2277 -650
rect 2311 -684 2317 -650
rect 2271 -722 2317 -684
rect 2271 -756 2277 -722
rect 2311 -756 2317 -722
rect 2271 -794 2317 -756
rect 2271 -828 2277 -794
rect 2311 -828 2317 -794
rect 2271 -866 2317 -828
rect 2271 -900 2277 -866
rect 2311 -900 2317 -866
rect 2271 -938 2317 -900
rect 2271 -972 2277 -938
rect 2311 -972 2317 -938
rect 2271 -1009 2317 -972
rect 2419 -146 2465 -109
rect 2419 -180 2425 -146
rect 2459 -180 2465 -146
rect 2419 -218 2465 -180
rect 2419 -252 2425 -218
rect 2459 -252 2465 -218
rect 2419 -290 2465 -252
rect 2419 -324 2425 -290
rect 2459 -324 2465 -290
rect 2419 -362 2465 -324
rect 2419 -396 2425 -362
rect 2459 -396 2465 -362
rect 2419 -434 2465 -396
rect 2419 -468 2425 -434
rect 2459 -468 2465 -434
rect 2419 -506 2465 -468
rect 2419 -540 2425 -506
rect 2459 -540 2465 -506
rect 2419 -578 2465 -540
rect 2419 -612 2425 -578
rect 2459 -612 2465 -578
rect 2419 -650 2465 -612
rect 2419 -684 2425 -650
rect 2459 -684 2465 -650
rect 2419 -722 2465 -684
rect 2419 -756 2425 -722
rect 2459 -756 2465 -722
rect 2419 -794 2465 -756
rect 2419 -828 2425 -794
rect 2459 -828 2465 -794
rect 2419 -866 2465 -828
rect 2419 -900 2425 -866
rect 2459 -900 2465 -866
rect 2419 -938 2465 -900
rect 2419 -972 2425 -938
rect 2459 -972 2465 -938
rect 2419 -1009 2465 -972
rect 2567 -146 2613 -109
rect 2567 -180 2573 -146
rect 2607 -180 2613 -146
rect 2567 -218 2613 -180
rect 2567 -252 2573 -218
rect 2607 -252 2613 -218
rect 2567 -290 2613 -252
rect 2567 -324 2573 -290
rect 2607 -324 2613 -290
rect 2567 -362 2613 -324
rect 2567 -396 2573 -362
rect 2607 -396 2613 -362
rect 2567 -434 2613 -396
rect 2567 -468 2573 -434
rect 2607 -468 2613 -434
rect 2567 -506 2613 -468
rect 2567 -540 2573 -506
rect 2607 -540 2613 -506
rect 2567 -578 2613 -540
rect 2567 -612 2573 -578
rect 2607 -612 2613 -578
rect 2567 -650 2613 -612
rect 2567 -684 2573 -650
rect 2607 -684 2613 -650
rect 2567 -722 2613 -684
rect 2567 -756 2573 -722
rect 2607 -756 2613 -722
rect 2567 -794 2613 -756
rect 2567 -828 2573 -794
rect 2607 -828 2613 -794
rect 2567 -866 2613 -828
rect 2567 -900 2573 -866
rect 2607 -900 2613 -866
rect 2567 -938 2613 -900
rect 2567 -972 2573 -938
rect 2607 -972 2613 -938
rect 2567 -1009 2613 -972
rect 2715 -146 2761 -109
rect 2715 -180 2721 -146
rect 2755 -180 2761 -146
rect 2715 -218 2761 -180
rect 2715 -252 2721 -218
rect 2755 -252 2761 -218
rect 2715 -290 2761 -252
rect 2715 -324 2721 -290
rect 2755 -324 2761 -290
rect 2715 -362 2761 -324
rect 2715 -396 2721 -362
rect 2755 -396 2761 -362
rect 2715 -434 2761 -396
rect 2715 -468 2721 -434
rect 2755 -468 2761 -434
rect 2715 -506 2761 -468
rect 2715 -540 2721 -506
rect 2755 -540 2761 -506
rect 2715 -578 2761 -540
rect 2715 -612 2721 -578
rect 2755 -612 2761 -578
rect 2715 -650 2761 -612
rect 2715 -684 2721 -650
rect 2755 -684 2761 -650
rect 2715 -722 2761 -684
rect 2715 -756 2721 -722
rect 2755 -756 2761 -722
rect 2715 -794 2761 -756
rect 2715 -828 2721 -794
rect 2755 -828 2761 -794
rect 2715 -866 2761 -828
rect 2715 -900 2721 -866
rect 2755 -900 2761 -866
rect 2715 -938 2761 -900
rect 2715 -972 2721 -938
rect 2755 -972 2761 -938
rect 2715 -1009 2761 -972
rect 2863 -146 2909 -109
rect 2863 -180 2869 -146
rect 2903 -180 2909 -146
rect 2863 -218 2909 -180
rect 2863 -252 2869 -218
rect 2903 -252 2909 -218
rect 2863 -290 2909 -252
rect 2863 -324 2869 -290
rect 2903 -324 2909 -290
rect 2863 -362 2909 -324
rect 2863 -396 2869 -362
rect 2903 -396 2909 -362
rect 2863 -434 2909 -396
rect 2863 -468 2869 -434
rect 2903 -468 2909 -434
rect 2863 -506 2909 -468
rect 2863 -540 2869 -506
rect 2903 -540 2909 -506
rect 2863 -578 2909 -540
rect 2863 -612 2869 -578
rect 2903 -612 2909 -578
rect 2863 -650 2909 -612
rect 2863 -684 2869 -650
rect 2903 -684 2909 -650
rect 2863 -722 2909 -684
rect 2863 -756 2869 -722
rect 2903 -756 2909 -722
rect 2863 -794 2909 -756
rect 2863 -828 2869 -794
rect 2903 -828 2909 -794
rect 2863 -866 2909 -828
rect 2863 -900 2869 -866
rect 2903 -900 2909 -866
rect 2863 -938 2909 -900
rect 2863 -972 2869 -938
rect 2903 -972 2909 -938
rect 2863 -1009 2909 -972
rect 3011 -146 3057 -109
rect 3011 -180 3017 -146
rect 3051 -180 3057 -146
rect 3011 -218 3057 -180
rect 3011 -252 3017 -218
rect 3051 -252 3057 -218
rect 3011 -290 3057 -252
rect 3011 -324 3017 -290
rect 3051 -324 3057 -290
rect 3011 -362 3057 -324
rect 3011 -396 3017 -362
rect 3051 -396 3057 -362
rect 3011 -434 3057 -396
rect 3011 -468 3017 -434
rect 3051 -468 3057 -434
rect 3011 -506 3057 -468
rect 3011 -540 3017 -506
rect 3051 -540 3057 -506
rect 3011 -578 3057 -540
rect 3011 -612 3017 -578
rect 3051 -612 3057 -578
rect 3011 -650 3057 -612
rect 3011 -684 3017 -650
rect 3051 -684 3057 -650
rect 3011 -722 3057 -684
rect 3011 -756 3017 -722
rect 3051 -756 3057 -722
rect 3011 -794 3057 -756
rect 3011 -828 3017 -794
rect 3051 -828 3057 -794
rect 3011 -866 3057 -828
rect 3011 -900 3017 -866
rect 3051 -900 3057 -866
rect 3011 -938 3057 -900
rect 3011 -972 3017 -938
rect 3051 -972 3057 -938
rect 3011 -1009 3057 -972
rect 3159 -146 3205 -109
rect 3159 -180 3165 -146
rect 3199 -180 3205 -146
rect 3159 -218 3205 -180
rect 3159 -252 3165 -218
rect 3199 -252 3205 -218
rect 3159 -290 3205 -252
rect 3159 -324 3165 -290
rect 3199 -324 3205 -290
rect 3159 -362 3205 -324
rect 3159 -396 3165 -362
rect 3199 -396 3205 -362
rect 3159 -434 3205 -396
rect 3159 -468 3165 -434
rect 3199 -468 3205 -434
rect 3159 -506 3205 -468
rect 3159 -540 3165 -506
rect 3199 -540 3205 -506
rect 3159 -578 3205 -540
rect 3159 -612 3165 -578
rect 3199 -612 3205 -578
rect 3159 -650 3205 -612
rect 3159 -684 3165 -650
rect 3199 -684 3205 -650
rect 3159 -722 3205 -684
rect 3159 -756 3165 -722
rect 3199 -756 3205 -722
rect 3159 -794 3205 -756
rect 3159 -828 3165 -794
rect 3199 -828 3205 -794
rect 3159 -866 3205 -828
rect 3159 -900 3165 -866
rect 3199 -900 3205 -866
rect 3159 -938 3205 -900
rect 3159 -972 3165 -938
rect 3199 -972 3205 -938
rect 3159 -1009 3205 -972
rect 3307 -146 3353 -109
rect 3307 -180 3313 -146
rect 3347 -180 3353 -146
rect 3307 -218 3353 -180
rect 3307 -252 3313 -218
rect 3347 -252 3353 -218
rect 3307 -290 3353 -252
rect 3307 -324 3313 -290
rect 3347 -324 3353 -290
rect 3307 -362 3353 -324
rect 3307 -396 3313 -362
rect 3347 -396 3353 -362
rect 3307 -434 3353 -396
rect 3307 -468 3313 -434
rect 3347 -468 3353 -434
rect 3307 -506 3353 -468
rect 3307 -540 3313 -506
rect 3347 -540 3353 -506
rect 3307 -578 3353 -540
rect 3307 -612 3313 -578
rect 3347 -612 3353 -578
rect 3307 -650 3353 -612
rect 3307 -684 3313 -650
rect 3347 -684 3353 -650
rect 3307 -722 3353 -684
rect 3307 -756 3313 -722
rect 3347 -756 3353 -722
rect 3307 -794 3353 -756
rect 3307 -828 3313 -794
rect 3347 -828 3353 -794
rect 3307 -866 3353 -828
rect 3307 -900 3313 -866
rect 3347 -900 3353 -866
rect 3307 -938 3353 -900
rect 3307 -972 3313 -938
rect 3347 -972 3353 -938
rect 3307 -1009 3353 -972
rect 3455 -146 3501 -109
rect 3455 -180 3461 -146
rect 3495 -180 3501 -146
rect 3455 -218 3501 -180
rect 3455 -252 3461 -218
rect 3495 -252 3501 -218
rect 3455 -290 3501 -252
rect 3455 -324 3461 -290
rect 3495 -324 3501 -290
rect 3455 -362 3501 -324
rect 3455 -396 3461 -362
rect 3495 -396 3501 -362
rect 3455 -434 3501 -396
rect 3455 -468 3461 -434
rect 3495 -468 3501 -434
rect 3455 -506 3501 -468
rect 3455 -540 3461 -506
rect 3495 -540 3501 -506
rect 3455 -578 3501 -540
rect 3455 -612 3461 -578
rect 3495 -612 3501 -578
rect 3455 -650 3501 -612
rect 3455 -684 3461 -650
rect 3495 -684 3501 -650
rect 3455 -722 3501 -684
rect 3455 -756 3461 -722
rect 3495 -756 3501 -722
rect 3455 -794 3501 -756
rect 3455 -828 3461 -794
rect 3495 -828 3501 -794
rect 3455 -866 3501 -828
rect 3455 -900 3461 -866
rect 3495 -900 3501 -866
rect 3455 -938 3501 -900
rect 3455 -972 3461 -938
rect 3495 -972 3501 -938
rect 3455 -1009 3501 -972
rect 3603 -146 3649 -109
rect 3603 -180 3609 -146
rect 3643 -180 3649 -146
rect 3603 -218 3649 -180
rect 3603 -252 3609 -218
rect 3643 -252 3649 -218
rect 3603 -290 3649 -252
rect 3603 -324 3609 -290
rect 3643 -324 3649 -290
rect 3603 -362 3649 -324
rect 3603 -396 3609 -362
rect 3643 -396 3649 -362
rect 3603 -434 3649 -396
rect 3603 -468 3609 -434
rect 3643 -468 3649 -434
rect 3603 -506 3649 -468
rect 3603 -540 3609 -506
rect 3643 -540 3649 -506
rect 3603 -578 3649 -540
rect 3603 -612 3609 -578
rect 3643 -612 3649 -578
rect 3603 -650 3649 -612
rect 3603 -684 3609 -650
rect 3643 -684 3649 -650
rect 3603 -722 3649 -684
rect 3603 -756 3609 -722
rect 3643 -756 3649 -722
rect 3603 -794 3649 -756
rect 3603 -828 3609 -794
rect 3643 -828 3649 -794
rect 3603 -866 3649 -828
rect 3603 -900 3609 -866
rect 3643 -900 3649 -866
rect 3603 -938 3649 -900
rect 3603 -972 3609 -938
rect 3643 -972 3649 -938
rect 3603 -1009 3649 -972
rect 3751 -146 3797 -109
rect 3751 -180 3757 -146
rect 3791 -180 3797 -146
rect 3751 -218 3797 -180
rect 3751 -252 3757 -218
rect 3791 -252 3797 -218
rect 3751 -290 3797 -252
rect 3751 -324 3757 -290
rect 3791 -324 3797 -290
rect 3751 -362 3797 -324
rect 3751 -396 3757 -362
rect 3791 -396 3797 -362
rect 3751 -434 3797 -396
rect 3751 -468 3757 -434
rect 3791 -468 3797 -434
rect 3751 -506 3797 -468
rect 3751 -540 3757 -506
rect 3791 -540 3797 -506
rect 3751 -578 3797 -540
rect 3751 -612 3757 -578
rect 3791 -612 3797 -578
rect 3751 -650 3797 -612
rect 3751 -684 3757 -650
rect 3791 -684 3797 -650
rect 3751 -722 3797 -684
rect 3751 -756 3757 -722
rect 3791 -756 3797 -722
rect 3751 -794 3797 -756
rect 3751 -828 3757 -794
rect 3791 -828 3797 -794
rect 3751 -866 3797 -828
rect 3751 -900 3757 -866
rect 3791 -900 3797 -866
rect 3751 -938 3797 -900
rect 3751 -972 3757 -938
rect 3791 -972 3797 -938
rect 3751 -1009 3797 -972
rect 3899 -146 3945 -109
rect 3899 -180 3905 -146
rect 3939 -180 3945 -146
rect 3899 -218 3945 -180
rect 3899 -252 3905 -218
rect 3939 -252 3945 -218
rect 3899 -290 3945 -252
rect 3899 -324 3905 -290
rect 3939 -324 3945 -290
rect 3899 -362 3945 -324
rect 3899 -396 3905 -362
rect 3939 -396 3945 -362
rect 3899 -434 3945 -396
rect 3899 -468 3905 -434
rect 3939 -468 3945 -434
rect 3899 -506 3945 -468
rect 3899 -540 3905 -506
rect 3939 -540 3945 -506
rect 3899 -578 3945 -540
rect 3899 -612 3905 -578
rect 3939 -612 3945 -578
rect 3899 -650 3945 -612
rect 3899 -684 3905 -650
rect 3939 -684 3945 -650
rect 3899 -722 3945 -684
rect 3899 -756 3905 -722
rect 3939 -756 3945 -722
rect 3899 -794 3945 -756
rect 3899 -828 3905 -794
rect 3939 -828 3945 -794
rect 3899 -866 3945 -828
rect 3899 -900 3905 -866
rect 3939 -900 3945 -866
rect 3899 -938 3945 -900
rect 3899 -972 3905 -938
rect 3939 -972 3945 -938
rect 3899 -1009 3945 -972
rect 4047 -146 4093 -109
rect 4047 -180 4053 -146
rect 4087 -180 4093 -146
rect 4047 -218 4093 -180
rect 4047 -252 4053 -218
rect 4087 -252 4093 -218
rect 4047 -290 4093 -252
rect 4047 -324 4053 -290
rect 4087 -324 4093 -290
rect 4047 -362 4093 -324
rect 4047 -396 4053 -362
rect 4087 -396 4093 -362
rect 4047 -434 4093 -396
rect 4047 -468 4053 -434
rect 4087 -468 4093 -434
rect 4047 -506 4093 -468
rect 4047 -540 4053 -506
rect 4087 -540 4093 -506
rect 4047 -578 4093 -540
rect 4047 -612 4053 -578
rect 4087 -612 4093 -578
rect 4047 -650 4093 -612
rect 4047 -684 4053 -650
rect 4087 -684 4093 -650
rect 4047 -722 4093 -684
rect 4047 -756 4053 -722
rect 4087 -756 4093 -722
rect 4047 -794 4093 -756
rect 4047 -828 4053 -794
rect 4087 -828 4093 -794
rect 4047 -866 4093 -828
rect 4047 -900 4053 -866
rect 4087 -900 4093 -866
rect 4047 -938 4093 -900
rect 4047 -972 4053 -938
rect 4087 -972 4093 -938
rect 4047 -1009 4093 -972
rect 4195 -146 4241 -109
rect 4195 -180 4201 -146
rect 4235 -180 4241 -146
rect 4195 -218 4241 -180
rect 4195 -252 4201 -218
rect 4235 -252 4241 -218
rect 4195 -290 4241 -252
rect 4195 -324 4201 -290
rect 4235 -324 4241 -290
rect 4195 -362 4241 -324
rect 4195 -396 4201 -362
rect 4235 -396 4241 -362
rect 4195 -434 4241 -396
rect 4195 -468 4201 -434
rect 4235 -468 4241 -434
rect 4195 -506 4241 -468
rect 4195 -540 4201 -506
rect 4235 -540 4241 -506
rect 4195 -578 4241 -540
rect 4195 -612 4201 -578
rect 4235 -612 4241 -578
rect 4195 -650 4241 -612
rect 4195 -684 4201 -650
rect 4235 -684 4241 -650
rect 4195 -722 4241 -684
rect 4195 -756 4201 -722
rect 4235 -756 4241 -722
rect 4195 -794 4241 -756
rect 4195 -828 4201 -794
rect 4235 -828 4241 -794
rect 4195 -866 4241 -828
rect 4195 -900 4201 -866
rect 4235 -900 4241 -866
rect 4195 -938 4241 -900
rect 4195 -972 4201 -938
rect 4235 -972 4241 -938
rect 4195 -1009 4241 -972
rect 4343 -146 4389 -109
rect 4343 -180 4349 -146
rect 4383 -180 4389 -146
rect 4343 -218 4389 -180
rect 4343 -252 4349 -218
rect 4383 -252 4389 -218
rect 4343 -290 4389 -252
rect 4343 -324 4349 -290
rect 4383 -324 4389 -290
rect 4343 -362 4389 -324
rect 4343 -396 4349 -362
rect 4383 -396 4389 -362
rect 4343 -434 4389 -396
rect 4343 -468 4349 -434
rect 4383 -468 4389 -434
rect 4343 -506 4389 -468
rect 4343 -540 4349 -506
rect 4383 -540 4389 -506
rect 4343 -578 4389 -540
rect 4343 -612 4349 -578
rect 4383 -612 4389 -578
rect 4343 -650 4389 -612
rect 4343 -684 4349 -650
rect 4383 -684 4389 -650
rect 4343 -722 4389 -684
rect 4343 -756 4349 -722
rect 4383 -756 4389 -722
rect 4343 -794 4389 -756
rect 4343 -828 4349 -794
rect 4383 -828 4389 -794
rect 4343 -866 4389 -828
rect 4343 -900 4349 -866
rect 4383 -900 4389 -866
rect 4343 -938 4389 -900
rect 4343 -972 4349 -938
rect 4383 -972 4389 -938
rect 4343 -1009 4389 -972
rect 4491 -146 4537 -109
rect 4491 -180 4497 -146
rect 4531 -180 4537 -146
rect 4491 -218 4537 -180
rect 4491 -252 4497 -218
rect 4531 -252 4537 -218
rect 4491 -290 4537 -252
rect 4491 -324 4497 -290
rect 4531 -324 4537 -290
rect 4491 -362 4537 -324
rect 4491 -396 4497 -362
rect 4531 -396 4537 -362
rect 4491 -434 4537 -396
rect 4491 -468 4497 -434
rect 4531 -468 4537 -434
rect 4491 -506 4537 -468
rect 4491 -540 4497 -506
rect 4531 -540 4537 -506
rect 4491 -578 4537 -540
rect 4491 -612 4497 -578
rect 4531 -612 4537 -578
rect 4491 -650 4537 -612
rect 4491 -684 4497 -650
rect 4531 -684 4537 -650
rect 4491 -722 4537 -684
rect 4491 -756 4497 -722
rect 4531 -756 4537 -722
rect 4491 -794 4537 -756
rect 4491 -828 4497 -794
rect 4531 -828 4537 -794
rect 4491 -866 4537 -828
rect 4491 -900 4497 -866
rect 4531 -900 4537 -866
rect 4491 -938 4537 -900
rect 4491 -972 4497 -938
rect 4531 -972 4537 -938
rect 4491 -1009 4537 -972
rect 4639 -146 4685 -109
rect 4639 -180 4645 -146
rect 4679 -180 4685 -146
rect 4639 -218 4685 -180
rect 4639 -252 4645 -218
rect 4679 -252 4685 -218
rect 4639 -290 4685 -252
rect 4639 -324 4645 -290
rect 4679 -324 4685 -290
rect 4639 -362 4685 -324
rect 4639 -396 4645 -362
rect 4679 -396 4685 -362
rect 4639 -434 4685 -396
rect 4639 -468 4645 -434
rect 4679 -468 4685 -434
rect 4639 -506 4685 -468
rect 4639 -540 4645 -506
rect 4679 -540 4685 -506
rect 4639 -578 4685 -540
rect 4639 -612 4645 -578
rect 4679 -612 4685 -578
rect 4639 -650 4685 -612
rect 4639 -684 4645 -650
rect 4679 -684 4685 -650
rect 4639 -722 4685 -684
rect 4639 -756 4645 -722
rect 4679 -756 4685 -722
rect 4639 -794 4685 -756
rect 4639 -828 4645 -794
rect 4679 -828 4685 -794
rect 4639 -866 4685 -828
rect 4639 -900 4645 -866
rect 4679 -900 4685 -866
rect 4639 -938 4685 -900
rect 4639 -972 4645 -938
rect 4679 -972 4685 -938
rect 4639 -1009 4685 -972
rect 4787 -146 4833 -109
rect 4787 -180 4793 -146
rect 4827 -180 4833 -146
rect 4787 -218 4833 -180
rect 4787 -252 4793 -218
rect 4827 -252 4833 -218
rect 4787 -290 4833 -252
rect 4787 -324 4793 -290
rect 4827 -324 4833 -290
rect 4787 -362 4833 -324
rect 4787 -396 4793 -362
rect 4827 -396 4833 -362
rect 4787 -434 4833 -396
rect 4787 -468 4793 -434
rect 4827 -468 4833 -434
rect 4787 -506 4833 -468
rect 4787 -540 4793 -506
rect 4827 -540 4833 -506
rect 4787 -578 4833 -540
rect 4787 -612 4793 -578
rect 4827 -612 4833 -578
rect 4787 -650 4833 -612
rect 4787 -684 4793 -650
rect 4827 -684 4833 -650
rect 4787 -722 4833 -684
rect 4787 -756 4793 -722
rect 4827 -756 4833 -722
rect 4787 -794 4833 -756
rect 4787 -828 4793 -794
rect 4827 -828 4833 -794
rect 4787 -866 4833 -828
rect 4787 -900 4793 -866
rect 4827 -900 4833 -866
rect 4787 -938 4833 -900
rect 4787 -972 4793 -938
rect 4827 -972 4833 -938
rect 4787 -1009 4833 -972
rect 4935 -146 4981 -109
rect 4935 -180 4941 -146
rect 4975 -180 4981 -146
rect 4935 -218 4981 -180
rect 4935 -252 4941 -218
rect 4975 -252 4981 -218
rect 4935 -290 4981 -252
rect 4935 -324 4941 -290
rect 4975 -324 4981 -290
rect 4935 -362 4981 -324
rect 4935 -396 4941 -362
rect 4975 -396 4981 -362
rect 4935 -434 4981 -396
rect 4935 -468 4941 -434
rect 4975 -468 4981 -434
rect 4935 -506 4981 -468
rect 4935 -540 4941 -506
rect 4975 -540 4981 -506
rect 4935 -578 4981 -540
rect 4935 -612 4941 -578
rect 4975 -612 4981 -578
rect 4935 -650 4981 -612
rect 4935 -684 4941 -650
rect 4975 -684 4981 -650
rect 4935 -722 4981 -684
rect 4935 -756 4941 -722
rect 4975 -756 4981 -722
rect 4935 -794 4981 -756
rect 4935 -828 4941 -794
rect 4975 -828 4981 -794
rect 4935 -866 4981 -828
rect 4935 -900 4941 -866
rect 4975 -900 4981 -866
rect 4935 -938 4981 -900
rect 4935 -972 4941 -938
rect 4975 -972 4981 -938
rect 4935 -1009 4981 -972
rect 5083 -146 5129 -109
rect 5083 -180 5089 -146
rect 5123 -180 5129 -146
rect 5083 -218 5129 -180
rect 5083 -252 5089 -218
rect 5123 -252 5129 -218
rect 5083 -290 5129 -252
rect 5083 -324 5089 -290
rect 5123 -324 5129 -290
rect 5083 -362 5129 -324
rect 5083 -396 5089 -362
rect 5123 -396 5129 -362
rect 5083 -434 5129 -396
rect 5083 -468 5089 -434
rect 5123 -468 5129 -434
rect 5083 -506 5129 -468
rect 5083 -540 5089 -506
rect 5123 -540 5129 -506
rect 5083 -578 5129 -540
rect 5083 -612 5089 -578
rect 5123 -612 5129 -578
rect 5083 -650 5129 -612
rect 5083 -684 5089 -650
rect 5123 -684 5129 -650
rect 5083 -722 5129 -684
rect 5083 -756 5089 -722
rect 5123 -756 5129 -722
rect 5083 -794 5129 -756
rect 5083 -828 5089 -794
rect 5123 -828 5129 -794
rect 5083 -866 5129 -828
rect 5083 -900 5089 -866
rect 5123 -900 5129 -866
rect 5083 -938 5129 -900
rect 5083 -972 5089 -938
rect 5123 -972 5129 -938
rect 5083 -1009 5129 -972
rect 5231 -146 5277 -109
rect 5231 -180 5237 -146
rect 5271 -180 5277 -146
rect 5231 -218 5277 -180
rect 5231 -252 5237 -218
rect 5271 -252 5277 -218
rect 5231 -290 5277 -252
rect 5231 -324 5237 -290
rect 5271 -324 5277 -290
rect 5231 -362 5277 -324
rect 5231 -396 5237 -362
rect 5271 -396 5277 -362
rect 5231 -434 5277 -396
rect 5231 -468 5237 -434
rect 5271 -468 5277 -434
rect 5231 -506 5277 -468
rect 5231 -540 5237 -506
rect 5271 -540 5277 -506
rect 5231 -578 5277 -540
rect 5231 -612 5237 -578
rect 5271 -612 5277 -578
rect 5231 -650 5277 -612
rect 5231 -684 5237 -650
rect 5271 -684 5277 -650
rect 5231 -722 5277 -684
rect 5231 -756 5237 -722
rect 5271 -756 5277 -722
rect 5231 -794 5277 -756
rect 5231 -828 5237 -794
rect 5271 -828 5277 -794
rect 5231 -866 5277 -828
rect 5231 -900 5237 -866
rect 5271 -900 5277 -866
rect 5231 -938 5277 -900
rect 5231 -972 5237 -938
rect 5271 -972 5277 -938
rect 5231 -1009 5277 -972
rect 5379 -146 5425 -109
rect 5379 -180 5385 -146
rect 5419 -180 5425 -146
rect 5379 -218 5425 -180
rect 5379 -252 5385 -218
rect 5419 -252 5425 -218
rect 5379 -290 5425 -252
rect 5379 -324 5385 -290
rect 5419 -324 5425 -290
rect 5379 -362 5425 -324
rect 5379 -396 5385 -362
rect 5419 -396 5425 -362
rect 5379 -434 5425 -396
rect 5379 -468 5385 -434
rect 5419 -468 5425 -434
rect 5379 -506 5425 -468
rect 5379 -540 5385 -506
rect 5419 -540 5425 -506
rect 5379 -578 5425 -540
rect 5379 -612 5385 -578
rect 5419 -612 5425 -578
rect 5379 -650 5425 -612
rect 5379 -684 5385 -650
rect 5419 -684 5425 -650
rect 5379 -722 5425 -684
rect 5379 -756 5385 -722
rect 5419 -756 5425 -722
rect 5379 -794 5425 -756
rect 5379 -828 5385 -794
rect 5419 -828 5425 -794
rect 5379 -866 5425 -828
rect 5379 -900 5385 -866
rect 5419 -900 5425 -866
rect 5379 -938 5425 -900
rect 5379 -972 5385 -938
rect 5419 -972 5425 -938
rect 5379 -1009 5425 -972
rect 5527 -146 5573 -109
rect 5527 -180 5533 -146
rect 5567 -180 5573 -146
rect 5527 -218 5573 -180
rect 5527 -252 5533 -218
rect 5567 -252 5573 -218
rect 5527 -290 5573 -252
rect 5527 -324 5533 -290
rect 5567 -324 5573 -290
rect 5527 -362 5573 -324
rect 5527 -396 5533 -362
rect 5567 -396 5573 -362
rect 5527 -434 5573 -396
rect 5527 -468 5533 -434
rect 5567 -468 5573 -434
rect 5527 -506 5573 -468
rect 5527 -540 5533 -506
rect 5567 -540 5573 -506
rect 5527 -578 5573 -540
rect 5527 -612 5533 -578
rect 5567 -612 5573 -578
rect 5527 -650 5573 -612
rect 5527 -684 5533 -650
rect 5567 -684 5573 -650
rect 5527 -722 5573 -684
rect 5527 -756 5533 -722
rect 5567 -756 5573 -722
rect 5527 -794 5573 -756
rect 5527 -828 5533 -794
rect 5567 -828 5573 -794
rect 5527 -866 5573 -828
rect 5527 -900 5533 -866
rect 5567 -900 5573 -866
rect 5527 -938 5573 -900
rect 5527 -972 5533 -938
rect 5567 -972 5573 -938
rect 5527 -1009 5573 -972
rect -5517 -1047 -5435 -1041
rect -5517 -1081 -5493 -1047
rect -5459 -1081 -5435 -1047
rect -5517 -1087 -5435 -1081
rect -5369 -1047 -5287 -1041
rect -5369 -1081 -5345 -1047
rect -5311 -1081 -5287 -1047
rect -5369 -1087 -5287 -1081
rect -5221 -1047 -5139 -1041
rect -5221 -1081 -5197 -1047
rect -5163 -1081 -5139 -1047
rect -5221 -1087 -5139 -1081
rect -5073 -1047 -4991 -1041
rect -5073 -1081 -5049 -1047
rect -5015 -1081 -4991 -1047
rect -5073 -1087 -4991 -1081
rect -4925 -1047 -4843 -1041
rect -4925 -1081 -4901 -1047
rect -4867 -1081 -4843 -1047
rect -4925 -1087 -4843 -1081
rect -4777 -1047 -4695 -1041
rect -4777 -1081 -4753 -1047
rect -4719 -1081 -4695 -1047
rect -4777 -1087 -4695 -1081
rect -4629 -1047 -4547 -1041
rect -4629 -1081 -4605 -1047
rect -4571 -1081 -4547 -1047
rect -4629 -1087 -4547 -1081
rect -4481 -1047 -4399 -1041
rect -4481 -1081 -4457 -1047
rect -4423 -1081 -4399 -1047
rect -4481 -1087 -4399 -1081
rect -4333 -1047 -4251 -1041
rect -4333 -1081 -4309 -1047
rect -4275 -1081 -4251 -1047
rect -4333 -1087 -4251 -1081
rect -4185 -1047 -4103 -1041
rect -4185 -1081 -4161 -1047
rect -4127 -1081 -4103 -1047
rect -4185 -1087 -4103 -1081
rect -4037 -1047 -3955 -1041
rect -4037 -1081 -4013 -1047
rect -3979 -1081 -3955 -1047
rect -4037 -1087 -3955 -1081
rect -3889 -1047 -3807 -1041
rect -3889 -1081 -3865 -1047
rect -3831 -1081 -3807 -1047
rect -3889 -1087 -3807 -1081
rect -3741 -1047 -3659 -1041
rect -3741 -1081 -3717 -1047
rect -3683 -1081 -3659 -1047
rect -3741 -1087 -3659 -1081
rect -3593 -1047 -3511 -1041
rect -3593 -1081 -3569 -1047
rect -3535 -1081 -3511 -1047
rect -3593 -1087 -3511 -1081
rect -3445 -1047 -3363 -1041
rect -3445 -1081 -3421 -1047
rect -3387 -1081 -3363 -1047
rect -3445 -1087 -3363 -1081
rect -3297 -1047 -3215 -1041
rect -3297 -1081 -3273 -1047
rect -3239 -1081 -3215 -1047
rect -3297 -1087 -3215 -1081
rect -3149 -1047 -3067 -1041
rect -3149 -1081 -3125 -1047
rect -3091 -1081 -3067 -1047
rect -3149 -1087 -3067 -1081
rect -3001 -1047 -2919 -1041
rect -3001 -1081 -2977 -1047
rect -2943 -1081 -2919 -1047
rect -3001 -1087 -2919 -1081
rect -2853 -1047 -2771 -1041
rect -2853 -1081 -2829 -1047
rect -2795 -1081 -2771 -1047
rect -2853 -1087 -2771 -1081
rect -2705 -1047 -2623 -1041
rect -2705 -1081 -2681 -1047
rect -2647 -1081 -2623 -1047
rect -2705 -1087 -2623 -1081
rect -2557 -1047 -2475 -1041
rect -2557 -1081 -2533 -1047
rect -2499 -1081 -2475 -1047
rect -2557 -1087 -2475 -1081
rect -2409 -1047 -2327 -1041
rect -2409 -1081 -2385 -1047
rect -2351 -1081 -2327 -1047
rect -2409 -1087 -2327 -1081
rect -2261 -1047 -2179 -1041
rect -2261 -1081 -2237 -1047
rect -2203 -1081 -2179 -1047
rect -2261 -1087 -2179 -1081
rect -2113 -1047 -2031 -1041
rect -2113 -1081 -2089 -1047
rect -2055 -1081 -2031 -1047
rect -2113 -1087 -2031 -1081
rect -1965 -1047 -1883 -1041
rect -1965 -1081 -1941 -1047
rect -1907 -1081 -1883 -1047
rect -1965 -1087 -1883 -1081
rect -1817 -1047 -1735 -1041
rect -1817 -1081 -1793 -1047
rect -1759 -1081 -1735 -1047
rect -1817 -1087 -1735 -1081
rect -1669 -1047 -1587 -1041
rect -1669 -1081 -1645 -1047
rect -1611 -1081 -1587 -1047
rect -1669 -1087 -1587 -1081
rect -1521 -1047 -1439 -1041
rect -1521 -1081 -1497 -1047
rect -1463 -1081 -1439 -1047
rect -1521 -1087 -1439 -1081
rect -1373 -1047 -1291 -1041
rect -1373 -1081 -1349 -1047
rect -1315 -1081 -1291 -1047
rect -1373 -1087 -1291 -1081
rect -1225 -1047 -1143 -1041
rect -1225 -1081 -1201 -1047
rect -1167 -1081 -1143 -1047
rect -1225 -1087 -1143 -1081
rect -1077 -1047 -995 -1041
rect -1077 -1081 -1053 -1047
rect -1019 -1081 -995 -1047
rect -1077 -1087 -995 -1081
rect -929 -1047 -847 -1041
rect -929 -1081 -905 -1047
rect -871 -1081 -847 -1047
rect -929 -1087 -847 -1081
rect -781 -1047 -699 -1041
rect -781 -1081 -757 -1047
rect -723 -1081 -699 -1047
rect -781 -1087 -699 -1081
rect -633 -1047 -551 -1041
rect -633 -1081 -609 -1047
rect -575 -1081 -551 -1047
rect -633 -1087 -551 -1081
rect -485 -1047 -403 -1041
rect -485 -1081 -461 -1047
rect -427 -1081 -403 -1047
rect -485 -1087 -403 -1081
rect -337 -1047 -255 -1041
rect -337 -1081 -313 -1047
rect -279 -1081 -255 -1047
rect -337 -1087 -255 -1081
rect -189 -1047 -107 -1041
rect -189 -1081 -165 -1047
rect -131 -1081 -107 -1047
rect -189 -1087 -107 -1081
rect -41 -1047 41 -1041
rect -41 -1081 -17 -1047
rect 17 -1081 41 -1047
rect -41 -1087 41 -1081
rect 107 -1047 189 -1041
rect 107 -1081 131 -1047
rect 165 -1081 189 -1047
rect 107 -1087 189 -1081
rect 255 -1047 337 -1041
rect 255 -1081 279 -1047
rect 313 -1081 337 -1047
rect 255 -1087 337 -1081
rect 403 -1047 485 -1041
rect 403 -1081 427 -1047
rect 461 -1081 485 -1047
rect 403 -1087 485 -1081
rect 551 -1047 633 -1041
rect 551 -1081 575 -1047
rect 609 -1081 633 -1047
rect 551 -1087 633 -1081
rect 699 -1047 781 -1041
rect 699 -1081 723 -1047
rect 757 -1081 781 -1047
rect 699 -1087 781 -1081
rect 847 -1047 929 -1041
rect 847 -1081 871 -1047
rect 905 -1081 929 -1047
rect 847 -1087 929 -1081
rect 995 -1047 1077 -1041
rect 995 -1081 1019 -1047
rect 1053 -1081 1077 -1047
rect 995 -1087 1077 -1081
rect 1143 -1047 1225 -1041
rect 1143 -1081 1167 -1047
rect 1201 -1081 1225 -1047
rect 1143 -1087 1225 -1081
rect 1291 -1047 1373 -1041
rect 1291 -1081 1315 -1047
rect 1349 -1081 1373 -1047
rect 1291 -1087 1373 -1081
rect 1439 -1047 1521 -1041
rect 1439 -1081 1463 -1047
rect 1497 -1081 1521 -1047
rect 1439 -1087 1521 -1081
rect 1587 -1047 1669 -1041
rect 1587 -1081 1611 -1047
rect 1645 -1081 1669 -1047
rect 1587 -1087 1669 -1081
rect 1735 -1047 1817 -1041
rect 1735 -1081 1759 -1047
rect 1793 -1081 1817 -1047
rect 1735 -1087 1817 -1081
rect 1883 -1047 1965 -1041
rect 1883 -1081 1907 -1047
rect 1941 -1081 1965 -1047
rect 1883 -1087 1965 -1081
rect 2031 -1047 2113 -1041
rect 2031 -1081 2055 -1047
rect 2089 -1081 2113 -1047
rect 2031 -1087 2113 -1081
rect 2179 -1047 2261 -1041
rect 2179 -1081 2203 -1047
rect 2237 -1081 2261 -1047
rect 2179 -1087 2261 -1081
rect 2327 -1047 2409 -1041
rect 2327 -1081 2351 -1047
rect 2385 -1081 2409 -1047
rect 2327 -1087 2409 -1081
rect 2475 -1047 2557 -1041
rect 2475 -1081 2499 -1047
rect 2533 -1081 2557 -1047
rect 2475 -1087 2557 -1081
rect 2623 -1047 2705 -1041
rect 2623 -1081 2647 -1047
rect 2681 -1081 2705 -1047
rect 2623 -1087 2705 -1081
rect 2771 -1047 2853 -1041
rect 2771 -1081 2795 -1047
rect 2829 -1081 2853 -1047
rect 2771 -1087 2853 -1081
rect 2919 -1047 3001 -1041
rect 2919 -1081 2943 -1047
rect 2977 -1081 3001 -1047
rect 2919 -1087 3001 -1081
rect 3067 -1047 3149 -1041
rect 3067 -1081 3091 -1047
rect 3125 -1081 3149 -1047
rect 3067 -1087 3149 -1081
rect 3215 -1047 3297 -1041
rect 3215 -1081 3239 -1047
rect 3273 -1081 3297 -1047
rect 3215 -1087 3297 -1081
rect 3363 -1047 3445 -1041
rect 3363 -1081 3387 -1047
rect 3421 -1081 3445 -1047
rect 3363 -1087 3445 -1081
rect 3511 -1047 3593 -1041
rect 3511 -1081 3535 -1047
rect 3569 -1081 3593 -1047
rect 3511 -1087 3593 -1081
rect 3659 -1047 3741 -1041
rect 3659 -1081 3683 -1047
rect 3717 -1081 3741 -1047
rect 3659 -1087 3741 -1081
rect 3807 -1047 3889 -1041
rect 3807 -1081 3831 -1047
rect 3865 -1081 3889 -1047
rect 3807 -1087 3889 -1081
rect 3955 -1047 4037 -1041
rect 3955 -1081 3979 -1047
rect 4013 -1081 4037 -1047
rect 3955 -1087 4037 -1081
rect 4103 -1047 4185 -1041
rect 4103 -1081 4127 -1047
rect 4161 -1081 4185 -1047
rect 4103 -1087 4185 -1081
rect 4251 -1047 4333 -1041
rect 4251 -1081 4275 -1047
rect 4309 -1081 4333 -1047
rect 4251 -1087 4333 -1081
rect 4399 -1047 4481 -1041
rect 4399 -1081 4423 -1047
rect 4457 -1081 4481 -1047
rect 4399 -1087 4481 -1081
rect 4547 -1047 4629 -1041
rect 4547 -1081 4571 -1047
rect 4605 -1081 4629 -1047
rect 4547 -1087 4629 -1081
rect 4695 -1047 4777 -1041
rect 4695 -1081 4719 -1047
rect 4753 -1081 4777 -1047
rect 4695 -1087 4777 -1081
rect 4843 -1047 4925 -1041
rect 4843 -1081 4867 -1047
rect 4901 -1081 4925 -1047
rect 4843 -1087 4925 -1081
rect 4991 -1047 5073 -1041
rect 4991 -1081 5015 -1047
rect 5049 -1081 5073 -1047
rect 4991 -1087 5073 -1081
rect 5139 -1047 5221 -1041
rect 5139 -1081 5163 -1047
rect 5197 -1081 5221 -1047
rect 5139 -1087 5221 -1081
rect 5287 -1047 5369 -1041
rect 5287 -1081 5311 -1047
rect 5345 -1081 5369 -1047
rect 5287 -1087 5369 -1081
rect 5435 -1047 5517 -1041
rect 5435 -1081 5459 -1047
rect 5493 -1081 5517 -1047
rect 5435 -1087 5517 -1081
<< properties >>
string FIXED_BBOX -5664 -1166 5664 1166
<< end >>
