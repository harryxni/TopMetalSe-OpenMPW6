magic
tech sky130A
magscale 1 2
timestamp 1654643737
<< pwell >>
rect 514 -6906 2166 -6274
rect 3514 -6906 5166 -6274
rect 6514 -6906 8166 -6274
<< nmoslvt >>
rect 540 -6800 2140 -6400
rect 3540 -6800 5140 -6400
rect 6540 -6800 8140 -6400
<< ndiff >>
rect 540 -6333 2140 -6300
rect 540 -6367 575 -6333
rect 609 -6367 643 -6333
rect 677 -6367 711 -6333
rect 745 -6367 779 -6333
rect 813 -6367 847 -6333
rect 881 -6367 915 -6333
rect 949 -6367 983 -6333
rect 1017 -6367 1051 -6333
rect 1085 -6367 1119 -6333
rect 1153 -6367 1187 -6333
rect 1221 -6367 1255 -6333
rect 1289 -6367 1323 -6333
rect 1357 -6367 1391 -6333
rect 1425 -6367 1459 -6333
rect 1493 -6367 1527 -6333
rect 1561 -6367 1595 -6333
rect 1629 -6367 1663 -6333
rect 1697 -6367 1731 -6333
rect 1765 -6367 1799 -6333
rect 1833 -6367 1867 -6333
rect 1901 -6367 1935 -6333
rect 1969 -6367 2003 -6333
rect 2037 -6367 2071 -6333
rect 2105 -6367 2140 -6333
rect 540 -6400 2140 -6367
rect 3540 -6333 5140 -6300
rect 3540 -6367 3575 -6333
rect 3609 -6367 3643 -6333
rect 3677 -6367 3711 -6333
rect 3745 -6367 3779 -6333
rect 3813 -6367 3847 -6333
rect 3881 -6367 3915 -6333
rect 3949 -6367 3983 -6333
rect 4017 -6367 4051 -6333
rect 4085 -6367 4119 -6333
rect 4153 -6367 4187 -6333
rect 4221 -6367 4255 -6333
rect 4289 -6367 4323 -6333
rect 4357 -6367 4391 -6333
rect 4425 -6367 4459 -6333
rect 4493 -6367 4527 -6333
rect 4561 -6367 4595 -6333
rect 4629 -6367 4663 -6333
rect 4697 -6367 4731 -6333
rect 4765 -6367 4799 -6333
rect 4833 -6367 4867 -6333
rect 4901 -6367 4935 -6333
rect 4969 -6367 5003 -6333
rect 5037 -6367 5071 -6333
rect 5105 -6367 5140 -6333
rect 3540 -6400 5140 -6367
rect 6540 -6333 8140 -6300
rect 6540 -6367 6575 -6333
rect 6609 -6367 6643 -6333
rect 6677 -6367 6711 -6333
rect 6745 -6367 6779 -6333
rect 6813 -6367 6847 -6333
rect 6881 -6367 6915 -6333
rect 6949 -6367 6983 -6333
rect 7017 -6367 7051 -6333
rect 7085 -6367 7119 -6333
rect 7153 -6367 7187 -6333
rect 7221 -6367 7255 -6333
rect 7289 -6367 7323 -6333
rect 7357 -6367 7391 -6333
rect 7425 -6367 7459 -6333
rect 7493 -6367 7527 -6333
rect 7561 -6367 7595 -6333
rect 7629 -6367 7663 -6333
rect 7697 -6367 7731 -6333
rect 7765 -6367 7799 -6333
rect 7833 -6367 7867 -6333
rect 7901 -6367 7935 -6333
rect 7969 -6367 8003 -6333
rect 8037 -6367 8071 -6333
rect 8105 -6367 8140 -6333
rect 6540 -6400 8140 -6367
rect 540 -6833 2140 -6800
rect 540 -6867 575 -6833
rect 609 -6867 643 -6833
rect 677 -6867 711 -6833
rect 745 -6867 779 -6833
rect 813 -6867 847 -6833
rect 881 -6867 915 -6833
rect 949 -6867 983 -6833
rect 1017 -6867 1051 -6833
rect 1085 -6867 1119 -6833
rect 1153 -6867 1187 -6833
rect 1221 -6867 1255 -6833
rect 1289 -6867 1323 -6833
rect 1357 -6867 1391 -6833
rect 1425 -6867 1459 -6833
rect 1493 -6867 1527 -6833
rect 1561 -6867 1595 -6833
rect 1629 -6867 1663 -6833
rect 1697 -6867 1731 -6833
rect 1765 -6867 1799 -6833
rect 1833 -6867 1867 -6833
rect 1901 -6867 1935 -6833
rect 1969 -6867 2003 -6833
rect 2037 -6867 2071 -6833
rect 2105 -6867 2140 -6833
rect 540 -6880 2140 -6867
rect 3540 -6833 5140 -6800
rect 3540 -6867 3575 -6833
rect 3609 -6867 3643 -6833
rect 3677 -6867 3711 -6833
rect 3745 -6867 3779 -6833
rect 3813 -6867 3847 -6833
rect 3881 -6867 3915 -6833
rect 3949 -6867 3983 -6833
rect 4017 -6867 4051 -6833
rect 4085 -6867 4119 -6833
rect 4153 -6867 4187 -6833
rect 4221 -6867 4255 -6833
rect 4289 -6867 4323 -6833
rect 4357 -6867 4391 -6833
rect 4425 -6867 4459 -6833
rect 4493 -6867 4527 -6833
rect 4561 -6867 4595 -6833
rect 4629 -6867 4663 -6833
rect 4697 -6867 4731 -6833
rect 4765 -6867 4799 -6833
rect 4833 -6867 4867 -6833
rect 4901 -6867 4935 -6833
rect 4969 -6867 5003 -6833
rect 5037 -6867 5071 -6833
rect 5105 -6867 5140 -6833
rect 3540 -6880 5140 -6867
rect 6540 -6833 8140 -6800
rect 6540 -6867 6575 -6833
rect 6609 -6867 6643 -6833
rect 6677 -6867 6711 -6833
rect 6745 -6867 6779 -6833
rect 6813 -6867 6847 -6833
rect 6881 -6867 6915 -6833
rect 6949 -6867 6983 -6833
rect 7017 -6867 7051 -6833
rect 7085 -6867 7119 -6833
rect 7153 -6867 7187 -6833
rect 7221 -6867 7255 -6833
rect 7289 -6867 7323 -6833
rect 7357 -6867 7391 -6833
rect 7425 -6867 7459 -6833
rect 7493 -6867 7527 -6833
rect 7561 -6867 7595 -6833
rect 7629 -6867 7663 -6833
rect 7697 -6867 7731 -6833
rect 7765 -6867 7799 -6833
rect 7833 -6867 7867 -6833
rect 7901 -6867 7935 -6833
rect 7969 -6867 8003 -6833
rect 8037 -6867 8071 -6833
rect 8105 -6867 8140 -6833
rect 6540 -6880 8140 -6867
<< ndiffc >>
rect 575 -6367 609 -6333
rect 643 -6367 677 -6333
rect 711 -6367 745 -6333
rect 779 -6367 813 -6333
rect 847 -6367 881 -6333
rect 915 -6367 949 -6333
rect 983 -6367 1017 -6333
rect 1051 -6367 1085 -6333
rect 1119 -6367 1153 -6333
rect 1187 -6367 1221 -6333
rect 1255 -6367 1289 -6333
rect 1323 -6367 1357 -6333
rect 1391 -6367 1425 -6333
rect 1459 -6367 1493 -6333
rect 1527 -6367 1561 -6333
rect 1595 -6367 1629 -6333
rect 1663 -6367 1697 -6333
rect 1731 -6367 1765 -6333
rect 1799 -6367 1833 -6333
rect 1867 -6367 1901 -6333
rect 1935 -6367 1969 -6333
rect 2003 -6367 2037 -6333
rect 2071 -6367 2105 -6333
rect 3575 -6367 3609 -6333
rect 3643 -6367 3677 -6333
rect 3711 -6367 3745 -6333
rect 3779 -6367 3813 -6333
rect 3847 -6367 3881 -6333
rect 3915 -6367 3949 -6333
rect 3983 -6367 4017 -6333
rect 4051 -6367 4085 -6333
rect 4119 -6367 4153 -6333
rect 4187 -6367 4221 -6333
rect 4255 -6367 4289 -6333
rect 4323 -6367 4357 -6333
rect 4391 -6367 4425 -6333
rect 4459 -6367 4493 -6333
rect 4527 -6367 4561 -6333
rect 4595 -6367 4629 -6333
rect 4663 -6367 4697 -6333
rect 4731 -6367 4765 -6333
rect 4799 -6367 4833 -6333
rect 4867 -6367 4901 -6333
rect 4935 -6367 4969 -6333
rect 5003 -6367 5037 -6333
rect 5071 -6367 5105 -6333
rect 6575 -6367 6609 -6333
rect 6643 -6367 6677 -6333
rect 6711 -6367 6745 -6333
rect 6779 -6367 6813 -6333
rect 6847 -6367 6881 -6333
rect 6915 -6367 6949 -6333
rect 6983 -6367 7017 -6333
rect 7051 -6367 7085 -6333
rect 7119 -6367 7153 -6333
rect 7187 -6367 7221 -6333
rect 7255 -6367 7289 -6333
rect 7323 -6367 7357 -6333
rect 7391 -6367 7425 -6333
rect 7459 -6367 7493 -6333
rect 7527 -6367 7561 -6333
rect 7595 -6367 7629 -6333
rect 7663 -6367 7697 -6333
rect 7731 -6367 7765 -6333
rect 7799 -6367 7833 -6333
rect 7867 -6367 7901 -6333
rect 7935 -6367 7969 -6333
rect 8003 -6367 8037 -6333
rect 8071 -6367 8105 -6333
rect 575 -6867 609 -6833
rect 643 -6867 677 -6833
rect 711 -6867 745 -6833
rect 779 -6867 813 -6833
rect 847 -6867 881 -6833
rect 915 -6867 949 -6833
rect 983 -6867 1017 -6833
rect 1051 -6867 1085 -6833
rect 1119 -6867 1153 -6833
rect 1187 -6867 1221 -6833
rect 1255 -6867 1289 -6833
rect 1323 -6867 1357 -6833
rect 1391 -6867 1425 -6833
rect 1459 -6867 1493 -6833
rect 1527 -6867 1561 -6833
rect 1595 -6867 1629 -6833
rect 1663 -6867 1697 -6833
rect 1731 -6867 1765 -6833
rect 1799 -6867 1833 -6833
rect 1867 -6867 1901 -6833
rect 1935 -6867 1969 -6833
rect 2003 -6867 2037 -6833
rect 2071 -6867 2105 -6833
rect 3575 -6867 3609 -6833
rect 3643 -6867 3677 -6833
rect 3711 -6867 3745 -6833
rect 3779 -6867 3813 -6833
rect 3847 -6867 3881 -6833
rect 3915 -6867 3949 -6833
rect 3983 -6867 4017 -6833
rect 4051 -6867 4085 -6833
rect 4119 -6867 4153 -6833
rect 4187 -6867 4221 -6833
rect 4255 -6867 4289 -6833
rect 4323 -6867 4357 -6833
rect 4391 -6867 4425 -6833
rect 4459 -6867 4493 -6833
rect 4527 -6867 4561 -6833
rect 4595 -6867 4629 -6833
rect 4663 -6867 4697 -6833
rect 4731 -6867 4765 -6833
rect 4799 -6867 4833 -6833
rect 4867 -6867 4901 -6833
rect 4935 -6867 4969 -6833
rect 5003 -6867 5037 -6833
rect 5071 -6867 5105 -6833
rect 6575 -6867 6609 -6833
rect 6643 -6867 6677 -6833
rect 6711 -6867 6745 -6833
rect 6779 -6867 6813 -6833
rect 6847 -6867 6881 -6833
rect 6915 -6867 6949 -6833
rect 6983 -6867 7017 -6833
rect 7051 -6867 7085 -6833
rect 7119 -6867 7153 -6833
rect 7187 -6867 7221 -6833
rect 7255 -6867 7289 -6833
rect 7323 -6867 7357 -6833
rect 7391 -6867 7425 -6833
rect 7459 -6867 7493 -6833
rect 7527 -6867 7561 -6833
rect 7595 -6867 7629 -6833
rect 7663 -6867 7697 -6833
rect 7731 -6867 7765 -6833
rect 7799 -6867 7833 -6833
rect 7867 -6867 7901 -6833
rect 7935 -6867 7969 -6833
rect 8003 -6867 8037 -6833
rect 8071 -6867 8105 -6833
<< poly >>
rect 510 -6490 540 -6400
rect 220 -6515 540 -6490
rect 220 -6685 245 -6515
rect 415 -6685 540 -6515
rect 220 -6710 540 -6685
rect 510 -6800 540 -6710
rect 2140 -6800 2170 -6400
rect 3510 -6490 3540 -6400
rect 3220 -6515 3540 -6490
rect 3220 -6685 3245 -6515
rect 3415 -6685 3540 -6515
rect 3220 -6710 3540 -6685
rect 3510 -6800 3540 -6710
rect 5140 -6800 5170 -6400
rect 6510 -6490 6540 -6400
rect 6220 -6515 6540 -6490
rect 6220 -6685 6245 -6515
rect 6415 -6685 6540 -6515
rect 6220 -6710 6540 -6685
rect 6510 -6800 6540 -6710
rect 8140 -6800 8170 -6400
<< polycont >>
rect 245 -6685 415 -6515
rect 3245 -6685 3415 -6515
rect 6245 -6685 6415 -6515
<< locali >>
rect 540 -6243 2140 -6230
rect 540 -6277 567 -6243
rect 601 -6277 639 -6243
rect 673 -6277 711 -6243
rect 745 -6277 783 -6243
rect 817 -6277 855 -6243
rect 889 -6277 927 -6243
rect 961 -6277 999 -6243
rect 1033 -6277 1071 -6243
rect 1105 -6277 1143 -6243
rect 1177 -6277 1215 -6243
rect 1249 -6277 1287 -6243
rect 1321 -6277 1359 -6243
rect 1393 -6277 1431 -6243
rect 1465 -6277 1503 -6243
rect 1537 -6277 1575 -6243
rect 1609 -6277 1647 -6243
rect 1681 -6277 1719 -6243
rect 1753 -6277 1791 -6243
rect 1825 -6277 1863 -6243
rect 1897 -6277 1935 -6243
rect 1969 -6277 2007 -6243
rect 2041 -6277 2079 -6243
rect 2113 -6277 2140 -6243
rect 540 -6333 2140 -6277
rect 540 -6367 575 -6333
rect 609 -6367 643 -6333
rect 677 -6367 711 -6333
rect 745 -6367 779 -6333
rect 813 -6367 847 -6333
rect 881 -6367 915 -6333
rect 949 -6367 983 -6333
rect 1017 -6367 1051 -6333
rect 1085 -6367 1119 -6333
rect 1153 -6367 1187 -6333
rect 1221 -6367 1255 -6333
rect 1289 -6367 1323 -6333
rect 1357 -6367 1391 -6333
rect 1425 -6367 1459 -6333
rect 1493 -6367 1527 -6333
rect 1561 -6367 1595 -6333
rect 1629 -6367 1663 -6333
rect 1697 -6367 1731 -6333
rect 1765 -6367 1799 -6333
rect 1833 -6367 1867 -6333
rect 1901 -6367 1935 -6333
rect 1969 -6367 2003 -6333
rect 2037 -6367 2071 -6333
rect 2105 -6367 2140 -6333
rect 540 -6380 2140 -6367
rect 3540 -6243 5140 -6230
rect 3540 -6277 3567 -6243
rect 3601 -6277 3639 -6243
rect 3673 -6277 3711 -6243
rect 3745 -6277 3783 -6243
rect 3817 -6277 3855 -6243
rect 3889 -6277 3927 -6243
rect 3961 -6277 3999 -6243
rect 4033 -6277 4071 -6243
rect 4105 -6277 4143 -6243
rect 4177 -6277 4215 -6243
rect 4249 -6277 4287 -6243
rect 4321 -6277 4359 -6243
rect 4393 -6277 4431 -6243
rect 4465 -6277 4503 -6243
rect 4537 -6277 4575 -6243
rect 4609 -6277 4647 -6243
rect 4681 -6277 4719 -6243
rect 4753 -6277 4791 -6243
rect 4825 -6277 4863 -6243
rect 4897 -6277 4935 -6243
rect 4969 -6277 5007 -6243
rect 5041 -6277 5079 -6243
rect 5113 -6277 5140 -6243
rect 3540 -6333 5140 -6277
rect 3540 -6367 3575 -6333
rect 3609 -6367 3643 -6333
rect 3677 -6367 3711 -6333
rect 3745 -6367 3779 -6333
rect 3813 -6367 3847 -6333
rect 3881 -6367 3915 -6333
rect 3949 -6367 3983 -6333
rect 4017 -6367 4051 -6333
rect 4085 -6367 4119 -6333
rect 4153 -6367 4187 -6333
rect 4221 -6367 4255 -6333
rect 4289 -6367 4323 -6333
rect 4357 -6367 4391 -6333
rect 4425 -6367 4459 -6333
rect 4493 -6367 4527 -6333
rect 4561 -6367 4595 -6333
rect 4629 -6367 4663 -6333
rect 4697 -6367 4731 -6333
rect 4765 -6367 4799 -6333
rect 4833 -6367 4867 -6333
rect 4901 -6367 4935 -6333
rect 4969 -6367 5003 -6333
rect 5037 -6367 5071 -6333
rect 5105 -6367 5140 -6333
rect 3540 -6380 5140 -6367
rect 6540 -6243 8140 -6230
rect 6540 -6277 6567 -6243
rect 6601 -6277 6639 -6243
rect 6673 -6277 6711 -6243
rect 6745 -6277 6783 -6243
rect 6817 -6277 6855 -6243
rect 6889 -6277 6927 -6243
rect 6961 -6277 6999 -6243
rect 7033 -6277 7071 -6243
rect 7105 -6277 7143 -6243
rect 7177 -6277 7215 -6243
rect 7249 -6277 7287 -6243
rect 7321 -6277 7359 -6243
rect 7393 -6277 7431 -6243
rect 7465 -6277 7503 -6243
rect 7537 -6277 7575 -6243
rect 7609 -6277 7647 -6243
rect 7681 -6277 7719 -6243
rect 7753 -6277 7791 -6243
rect 7825 -6277 7863 -6243
rect 7897 -6277 7935 -6243
rect 7969 -6277 8007 -6243
rect 8041 -6277 8079 -6243
rect 8113 -6277 8140 -6243
rect 6540 -6333 8140 -6277
rect 6540 -6367 6575 -6333
rect 6609 -6367 6643 -6333
rect 6677 -6367 6711 -6333
rect 6745 -6367 6779 -6333
rect 6813 -6367 6847 -6333
rect 6881 -6367 6915 -6333
rect 6949 -6367 6983 -6333
rect 7017 -6367 7051 -6333
rect 7085 -6367 7119 -6333
rect 7153 -6367 7187 -6333
rect 7221 -6367 7255 -6333
rect 7289 -6367 7323 -6333
rect 7357 -6367 7391 -6333
rect 7425 -6367 7459 -6333
rect 7493 -6367 7527 -6333
rect 7561 -6367 7595 -6333
rect 7629 -6367 7663 -6333
rect 7697 -6367 7731 -6333
rect 7765 -6367 7799 -6333
rect 7833 -6367 7867 -6333
rect 7901 -6367 7935 -6333
rect 7969 -6367 8003 -6333
rect 8037 -6367 8071 -6333
rect 8105 -6367 8140 -6333
rect 6540 -6380 8140 -6367
rect 220 -6511 440 -6490
rect 220 -6689 241 -6511
rect 419 -6689 440 -6511
rect 220 -6710 440 -6689
rect 3220 -6511 3440 -6490
rect 3220 -6689 3241 -6511
rect 3419 -6689 3440 -6511
rect 3220 -6710 3440 -6689
rect 6220 -6511 6440 -6490
rect 6220 -6689 6241 -6511
rect 6419 -6689 6440 -6511
rect 6220 -6710 6440 -6689
rect 540 -6833 2140 -6800
rect 540 -6867 575 -6833
rect 609 -6867 643 -6833
rect 677 -6867 711 -6833
rect 745 -6867 779 -6833
rect 813 -6867 847 -6833
rect 881 -6867 915 -6833
rect 949 -6867 983 -6833
rect 1017 -6867 1051 -6833
rect 1085 -6867 1119 -6833
rect 1153 -6867 1187 -6833
rect 1221 -6867 1255 -6833
rect 1289 -6867 1323 -6833
rect 1357 -6867 1391 -6833
rect 1425 -6867 1459 -6833
rect 1493 -6867 1527 -6833
rect 1561 -6867 1595 -6833
rect 1629 -6867 1663 -6833
rect 1697 -6867 1731 -6833
rect 1765 -6867 1799 -6833
rect 1833 -6867 1867 -6833
rect 1901 -6867 1935 -6833
rect 1969 -6867 2003 -6833
rect 2037 -6867 2071 -6833
rect 2105 -6867 2140 -6833
rect 540 -6933 2140 -6867
rect 540 -6967 567 -6933
rect 601 -6967 639 -6933
rect 673 -6967 711 -6933
rect 745 -6967 783 -6933
rect 817 -6967 855 -6933
rect 889 -6967 927 -6933
rect 961 -6967 999 -6933
rect 1033 -6967 1071 -6933
rect 1105 -6967 1143 -6933
rect 1177 -6967 1215 -6933
rect 1249 -6967 1287 -6933
rect 1321 -6967 1359 -6933
rect 1393 -6967 1431 -6933
rect 1465 -6967 1503 -6933
rect 1537 -6967 1575 -6933
rect 1609 -6967 1647 -6933
rect 1681 -6967 1719 -6933
rect 1753 -6967 1791 -6933
rect 1825 -6967 1863 -6933
rect 1897 -6967 1935 -6933
rect 1969 -6967 2007 -6933
rect 2041 -6967 2079 -6933
rect 2113 -6967 2140 -6933
rect 540 -7000 2140 -6967
rect 3540 -6833 5140 -6800
rect 3540 -6867 3575 -6833
rect 3609 -6867 3643 -6833
rect 3677 -6867 3711 -6833
rect 3745 -6867 3779 -6833
rect 3813 -6867 3847 -6833
rect 3881 -6867 3915 -6833
rect 3949 -6867 3983 -6833
rect 4017 -6867 4051 -6833
rect 4085 -6867 4119 -6833
rect 4153 -6867 4187 -6833
rect 4221 -6867 4255 -6833
rect 4289 -6867 4323 -6833
rect 4357 -6867 4391 -6833
rect 4425 -6867 4459 -6833
rect 4493 -6867 4527 -6833
rect 4561 -6867 4595 -6833
rect 4629 -6867 4663 -6833
rect 4697 -6867 4731 -6833
rect 4765 -6867 4799 -6833
rect 4833 -6867 4867 -6833
rect 4901 -6867 4935 -6833
rect 4969 -6867 5003 -6833
rect 5037 -6867 5071 -6833
rect 5105 -6867 5140 -6833
rect 3540 -6933 5140 -6867
rect 3540 -6967 3567 -6933
rect 3601 -6967 3639 -6933
rect 3673 -6967 3711 -6933
rect 3745 -6967 3783 -6933
rect 3817 -6967 3855 -6933
rect 3889 -6967 3927 -6933
rect 3961 -6967 3999 -6933
rect 4033 -6967 4071 -6933
rect 4105 -6967 4143 -6933
rect 4177 -6967 4215 -6933
rect 4249 -6967 4287 -6933
rect 4321 -6967 4359 -6933
rect 4393 -6967 4431 -6933
rect 4465 -6967 4503 -6933
rect 4537 -6967 4575 -6933
rect 4609 -6967 4647 -6933
rect 4681 -6967 4719 -6933
rect 4753 -6967 4791 -6933
rect 4825 -6967 4863 -6933
rect 4897 -6967 4935 -6933
rect 4969 -6967 5007 -6933
rect 5041 -6967 5079 -6933
rect 5113 -6967 5140 -6933
rect 3540 -7000 5140 -6967
rect 6540 -6833 8140 -6800
rect 6540 -6867 6575 -6833
rect 6609 -6867 6643 -6833
rect 6677 -6867 6711 -6833
rect 6745 -6867 6779 -6833
rect 6813 -6867 6847 -6833
rect 6881 -6867 6915 -6833
rect 6949 -6867 6983 -6833
rect 7017 -6867 7051 -6833
rect 7085 -6867 7119 -6833
rect 7153 -6867 7187 -6833
rect 7221 -6867 7255 -6833
rect 7289 -6867 7323 -6833
rect 7357 -6867 7391 -6833
rect 7425 -6867 7459 -6833
rect 7493 -6867 7527 -6833
rect 7561 -6867 7595 -6833
rect 7629 -6867 7663 -6833
rect 7697 -6867 7731 -6833
rect 7765 -6867 7799 -6833
rect 7833 -6867 7867 -6833
rect 7901 -6867 7935 -6833
rect 7969 -6867 8003 -6833
rect 8037 -6867 8071 -6833
rect 8105 -6867 8140 -6833
rect 6540 -6933 8140 -6867
rect 6540 -6967 6567 -6933
rect 6601 -6967 6639 -6933
rect 6673 -6967 6711 -6933
rect 6745 -6967 6783 -6933
rect 6817 -6967 6855 -6933
rect 6889 -6967 6927 -6933
rect 6961 -6967 6999 -6933
rect 7033 -6967 7071 -6933
rect 7105 -6967 7143 -6933
rect 7177 -6967 7215 -6933
rect 7249 -6967 7287 -6933
rect 7321 -6967 7359 -6933
rect 7393 -6967 7431 -6933
rect 7465 -6967 7503 -6933
rect 7537 -6967 7575 -6933
rect 7609 -6967 7647 -6933
rect 7681 -6967 7719 -6933
rect 7753 -6967 7791 -6933
rect 7825 -6967 7863 -6933
rect 7897 -6967 7935 -6933
rect 7969 -6967 8007 -6933
rect 8041 -6967 8079 -6933
rect 8113 -6967 8140 -6933
rect 6540 -7000 8140 -6967
<< viali >>
rect 567 -6277 601 -6243
rect 639 -6277 673 -6243
rect 711 -6277 745 -6243
rect 783 -6277 817 -6243
rect 855 -6277 889 -6243
rect 927 -6277 961 -6243
rect 999 -6277 1033 -6243
rect 1071 -6277 1105 -6243
rect 1143 -6277 1177 -6243
rect 1215 -6277 1249 -6243
rect 1287 -6277 1321 -6243
rect 1359 -6277 1393 -6243
rect 1431 -6277 1465 -6243
rect 1503 -6277 1537 -6243
rect 1575 -6277 1609 -6243
rect 1647 -6277 1681 -6243
rect 1719 -6277 1753 -6243
rect 1791 -6277 1825 -6243
rect 1863 -6277 1897 -6243
rect 1935 -6277 1969 -6243
rect 2007 -6277 2041 -6243
rect 2079 -6277 2113 -6243
rect 3567 -6277 3601 -6243
rect 3639 -6277 3673 -6243
rect 3711 -6277 3745 -6243
rect 3783 -6277 3817 -6243
rect 3855 -6277 3889 -6243
rect 3927 -6277 3961 -6243
rect 3999 -6277 4033 -6243
rect 4071 -6277 4105 -6243
rect 4143 -6277 4177 -6243
rect 4215 -6277 4249 -6243
rect 4287 -6277 4321 -6243
rect 4359 -6277 4393 -6243
rect 4431 -6277 4465 -6243
rect 4503 -6277 4537 -6243
rect 4575 -6277 4609 -6243
rect 4647 -6277 4681 -6243
rect 4719 -6277 4753 -6243
rect 4791 -6277 4825 -6243
rect 4863 -6277 4897 -6243
rect 4935 -6277 4969 -6243
rect 5007 -6277 5041 -6243
rect 5079 -6277 5113 -6243
rect 6567 -6277 6601 -6243
rect 6639 -6277 6673 -6243
rect 6711 -6277 6745 -6243
rect 6783 -6277 6817 -6243
rect 6855 -6277 6889 -6243
rect 6927 -6277 6961 -6243
rect 6999 -6277 7033 -6243
rect 7071 -6277 7105 -6243
rect 7143 -6277 7177 -6243
rect 7215 -6277 7249 -6243
rect 7287 -6277 7321 -6243
rect 7359 -6277 7393 -6243
rect 7431 -6277 7465 -6243
rect 7503 -6277 7537 -6243
rect 7575 -6277 7609 -6243
rect 7647 -6277 7681 -6243
rect 7719 -6277 7753 -6243
rect 7791 -6277 7825 -6243
rect 7863 -6277 7897 -6243
rect 7935 -6277 7969 -6243
rect 8007 -6277 8041 -6243
rect 8079 -6277 8113 -6243
rect 241 -6515 419 -6511
rect 241 -6685 245 -6515
rect 245 -6685 415 -6515
rect 415 -6685 419 -6515
rect 241 -6689 419 -6685
rect 3241 -6515 3419 -6511
rect 3241 -6685 3245 -6515
rect 3245 -6685 3415 -6515
rect 3415 -6685 3419 -6515
rect 3241 -6689 3419 -6685
rect 6241 -6515 6419 -6511
rect 6241 -6685 6245 -6515
rect 6245 -6685 6415 -6515
rect 6415 -6685 6419 -6515
rect 6241 -6689 6419 -6685
rect 567 -6967 601 -6933
rect 639 -6967 673 -6933
rect 711 -6967 745 -6933
rect 783 -6967 817 -6933
rect 855 -6967 889 -6933
rect 927 -6967 961 -6933
rect 999 -6967 1033 -6933
rect 1071 -6967 1105 -6933
rect 1143 -6967 1177 -6933
rect 1215 -6967 1249 -6933
rect 1287 -6967 1321 -6933
rect 1359 -6967 1393 -6933
rect 1431 -6967 1465 -6933
rect 1503 -6967 1537 -6933
rect 1575 -6967 1609 -6933
rect 1647 -6967 1681 -6933
rect 1719 -6967 1753 -6933
rect 1791 -6967 1825 -6933
rect 1863 -6967 1897 -6933
rect 1935 -6967 1969 -6933
rect 2007 -6967 2041 -6933
rect 2079 -6967 2113 -6933
rect 3567 -6967 3601 -6933
rect 3639 -6967 3673 -6933
rect 3711 -6967 3745 -6933
rect 3783 -6967 3817 -6933
rect 3855 -6967 3889 -6933
rect 3927 -6967 3961 -6933
rect 3999 -6967 4033 -6933
rect 4071 -6967 4105 -6933
rect 4143 -6967 4177 -6933
rect 4215 -6967 4249 -6933
rect 4287 -6967 4321 -6933
rect 4359 -6967 4393 -6933
rect 4431 -6967 4465 -6933
rect 4503 -6967 4537 -6933
rect 4575 -6967 4609 -6933
rect 4647 -6967 4681 -6933
rect 4719 -6967 4753 -6933
rect 4791 -6967 4825 -6933
rect 4863 -6967 4897 -6933
rect 4935 -6967 4969 -6933
rect 5007 -6967 5041 -6933
rect 5079 -6967 5113 -6933
rect 6567 -6967 6601 -6933
rect 6639 -6967 6673 -6933
rect 6711 -6967 6745 -6933
rect 6783 -6967 6817 -6933
rect 6855 -6967 6889 -6933
rect 6927 -6967 6961 -6933
rect 6999 -6967 7033 -6933
rect 7071 -6967 7105 -6933
rect 7143 -6967 7177 -6933
rect 7215 -6967 7249 -6933
rect 7287 -6967 7321 -6933
rect 7359 -6967 7393 -6933
rect 7431 -6967 7465 -6933
rect 7503 -6967 7537 -6933
rect 7575 -6967 7609 -6933
rect 7647 -6967 7681 -6933
rect 7719 -6967 7753 -6933
rect 7791 -6967 7825 -6933
rect 7863 -6967 7897 -6933
rect 7935 -6967 7969 -6933
rect 8007 -6967 8041 -6933
rect 8079 -6967 8113 -6933
<< metal1 >>
rect -1770 3431 8000 3460
rect -1770 3379 -1745 3431
rect -1693 3379 -1681 3431
rect -1629 3379 -1617 3431
rect -1565 3379 -1553 3431
rect -1501 3379 -1489 3431
rect -1437 3379 -1425 3431
rect -1373 3379 -1361 3431
rect -1309 3379 -1297 3431
rect -1245 3379 -1233 3431
rect -1181 3379 -1169 3431
rect -1117 3379 -1105 3431
rect -1053 3379 -1041 3431
rect -989 3379 -977 3431
rect -925 3379 69 3431
rect 121 3379 3069 3431
rect 3121 3379 6069 3431
rect 6121 3379 8000 3431
rect -1770 3350 8000 3379
rect -2000 2970 -1800 2990
rect -2000 2880 40 2970
rect -2000 2820 0 2880
rect -2000 -30 -1800 2820
rect -1600 1551 0 1570
rect -1600 1499 -1566 1551
rect -1514 1499 -1502 1551
rect -1450 1499 -1438 1551
rect -1386 1499 -1374 1551
rect -1322 1499 -1310 1551
rect -1258 1499 -1246 1551
rect -1194 1499 -522 1551
rect -470 1499 -458 1551
rect -406 1499 -394 1551
rect -342 1499 -330 1551
rect -278 1499 0 1551
rect -1600 1480 0 1499
rect 9400 180 9600 3030
rect 9000 30 9600 180
rect -2000 -120 40 -30
rect -2000 -180 0 -120
rect -2000 -3030 -1800 -180
rect -1600 -1449 0 -1430
rect -1600 -1501 -1566 -1449
rect -1514 -1501 -1502 -1449
rect -1450 -1501 -1438 -1449
rect -1386 -1501 -1374 -1449
rect -1322 -1501 -1310 -1449
rect -1258 -1501 -1246 -1449
rect -1194 -1501 -522 -1449
rect -470 -1501 -458 -1449
rect -406 -1501 -394 -1449
rect -342 -1501 -330 -1449
rect -278 -1501 0 -1449
rect -1600 -1520 0 -1501
rect 9400 -2820 9600 30
rect 9000 -2970 9600 -2820
rect -2000 -3120 40 -3030
rect -2000 -3180 0 -3120
rect -2000 -6000 -1800 -3180
rect -1600 -4449 0 -4430
rect -1600 -4501 -1566 -4449
rect -1514 -4501 -1502 -4449
rect -1450 -4501 -1438 -4449
rect -1386 -4501 -1374 -4449
rect -1322 -4501 -1310 -4449
rect -1258 -4501 -1246 -4449
rect -1194 -4501 -522 -4449
rect -470 -4501 -458 -4449
rect -406 -4501 -394 -4449
rect -342 -4501 -330 -4449
rect -278 -4501 0 -4449
rect -1600 -4520 0 -4501
rect 9400 -5820 9600 -2970
rect 2860 -5910 3000 -5830
rect 9000 -5970 9600 -5820
rect 540 -6139 2140 -6130
rect 540 -6191 578 -6139
rect 630 -6191 642 -6139
rect 694 -6191 706 -6139
rect 758 -6191 770 -6139
rect 822 -6191 834 -6139
rect 886 -6191 898 -6139
rect 950 -6191 962 -6139
rect 1014 -6191 1026 -6139
rect 1078 -6191 1090 -6139
rect 1142 -6191 1154 -6139
rect 1206 -6191 1218 -6139
rect 1270 -6191 1282 -6139
rect 1334 -6191 1346 -6139
rect 1398 -6191 1410 -6139
rect 1462 -6191 1474 -6139
rect 1526 -6191 1538 -6139
rect 1590 -6191 1602 -6139
rect 1654 -6191 1666 -6139
rect 1718 -6191 1730 -6139
rect 1782 -6191 1794 -6139
rect 1846 -6191 1858 -6139
rect 1910 -6191 1922 -6139
rect 1974 -6191 1986 -6139
rect 2038 -6191 2050 -6139
rect 2102 -6191 2140 -6139
rect 540 -6243 2140 -6191
rect 540 -6277 567 -6243
rect 601 -6277 639 -6243
rect 673 -6277 711 -6243
rect 745 -6277 783 -6243
rect 817 -6277 855 -6243
rect 889 -6277 927 -6243
rect 961 -6277 999 -6243
rect 1033 -6277 1071 -6243
rect 1105 -6277 1143 -6243
rect 1177 -6277 1215 -6243
rect 1249 -6277 1287 -6243
rect 1321 -6277 1359 -6243
rect 1393 -6277 1431 -6243
rect 1465 -6277 1503 -6243
rect 1537 -6277 1575 -6243
rect 1609 -6277 1647 -6243
rect 1681 -6277 1719 -6243
rect 1753 -6277 1791 -6243
rect 1825 -6277 1863 -6243
rect 1897 -6277 1935 -6243
rect 1969 -6277 2007 -6243
rect 2041 -6277 2079 -6243
rect 2113 -6277 2140 -6243
rect 540 -6300 2140 -6277
rect 3540 -6139 5140 -6130
rect 3540 -6191 3578 -6139
rect 3630 -6191 3642 -6139
rect 3694 -6191 3706 -6139
rect 3758 -6191 3770 -6139
rect 3822 -6191 3834 -6139
rect 3886 -6191 3898 -6139
rect 3950 -6191 3962 -6139
rect 4014 -6191 4026 -6139
rect 4078 -6191 4090 -6139
rect 4142 -6191 4154 -6139
rect 4206 -6191 4218 -6139
rect 4270 -6191 4282 -6139
rect 4334 -6191 4346 -6139
rect 4398 -6191 4410 -6139
rect 4462 -6191 4474 -6139
rect 4526 -6191 4538 -6139
rect 4590 -6191 4602 -6139
rect 4654 -6191 4666 -6139
rect 4718 -6191 4730 -6139
rect 4782 -6191 4794 -6139
rect 4846 -6191 4858 -6139
rect 4910 -6191 4922 -6139
rect 4974 -6191 4986 -6139
rect 5038 -6191 5050 -6139
rect 5102 -6191 5140 -6139
rect 3540 -6243 5140 -6191
rect 3540 -6277 3567 -6243
rect 3601 -6277 3639 -6243
rect 3673 -6277 3711 -6243
rect 3745 -6277 3783 -6243
rect 3817 -6277 3855 -6243
rect 3889 -6277 3927 -6243
rect 3961 -6277 3999 -6243
rect 4033 -6277 4071 -6243
rect 4105 -6277 4143 -6243
rect 4177 -6277 4215 -6243
rect 4249 -6277 4287 -6243
rect 4321 -6277 4359 -6243
rect 4393 -6277 4431 -6243
rect 4465 -6277 4503 -6243
rect 4537 -6277 4575 -6243
rect 4609 -6277 4647 -6243
rect 4681 -6277 4719 -6243
rect 4753 -6277 4791 -6243
rect 4825 -6277 4863 -6243
rect 4897 -6277 4935 -6243
rect 4969 -6277 5007 -6243
rect 5041 -6277 5079 -6243
rect 5113 -6277 5140 -6243
rect 3540 -6300 5140 -6277
rect 6540 -6139 8140 -6130
rect 6540 -6191 6578 -6139
rect 6630 -6191 6642 -6139
rect 6694 -6191 6706 -6139
rect 6758 -6191 6770 -6139
rect 6822 -6191 6834 -6139
rect 6886 -6191 6898 -6139
rect 6950 -6191 6962 -6139
rect 7014 -6191 7026 -6139
rect 7078 -6191 7090 -6139
rect 7142 -6191 7154 -6139
rect 7206 -6191 7218 -6139
rect 7270 -6191 7282 -6139
rect 7334 -6191 7346 -6139
rect 7398 -6191 7410 -6139
rect 7462 -6191 7474 -6139
rect 7526 -6191 7538 -6139
rect 7590 -6191 7602 -6139
rect 7654 -6191 7666 -6139
rect 7718 -6191 7730 -6139
rect 7782 -6191 7794 -6139
rect 7846 -6191 7858 -6139
rect 7910 -6191 7922 -6139
rect 7974 -6191 7986 -6139
rect 8038 -6191 8050 -6139
rect 8102 -6191 8140 -6139
rect 6540 -6243 8140 -6191
rect 6540 -6277 6567 -6243
rect 6601 -6277 6639 -6243
rect 6673 -6277 6711 -6243
rect 6745 -6277 6783 -6243
rect 6817 -6277 6855 -6243
rect 6889 -6277 6927 -6243
rect 6961 -6277 6999 -6243
rect 7033 -6277 7071 -6243
rect 7105 -6277 7143 -6243
rect 7177 -6277 7215 -6243
rect 7249 -6277 7287 -6243
rect 7321 -6277 7359 -6243
rect 7393 -6277 7431 -6243
rect 7465 -6277 7503 -6243
rect 7537 -6277 7575 -6243
rect 7609 -6277 7647 -6243
rect 7681 -6277 7719 -6243
rect 7753 -6277 7791 -6243
rect 7825 -6277 7863 -6243
rect 7897 -6277 7935 -6243
rect 7969 -6277 8007 -6243
rect 8041 -6277 8079 -6243
rect 8113 -6277 8140 -6243
rect 6540 -6300 8140 -6277
rect 220 -6510 440 -6490
rect 220 -6690 240 -6510
rect 420 -6690 440 -6510
rect 220 -6710 440 -6690
rect 3220 -6510 3440 -6490
rect 3220 -6690 3240 -6510
rect 3420 -6690 3440 -6510
rect 3220 -6710 3440 -6690
rect 6220 -6510 6440 -6490
rect 6220 -6690 6240 -6510
rect 6420 -6690 6440 -6510
rect 6220 -6710 6440 -6690
rect 540 -6933 9740 -6900
rect 540 -6967 567 -6933
rect 601 -6942 639 -6933
rect 673 -6942 711 -6933
rect 745 -6942 783 -6933
rect 817 -6942 855 -6933
rect 889 -6942 927 -6933
rect 961 -6942 999 -6933
rect 1033 -6942 1071 -6933
rect 1105 -6942 1143 -6933
rect 1177 -6942 1215 -6933
rect 1249 -6942 1287 -6933
rect 1321 -6942 1359 -6933
rect 1393 -6942 1431 -6933
rect 1465 -6942 1503 -6933
rect 1537 -6942 1575 -6933
rect 1609 -6942 1647 -6933
rect 1681 -6942 1719 -6933
rect 1753 -6942 1791 -6933
rect 1825 -6942 1863 -6933
rect 1897 -6942 1935 -6933
rect 1969 -6942 2007 -6933
rect 2041 -6942 2079 -6933
rect 2113 -6942 3567 -6933
rect 3601 -6942 3639 -6933
rect 3673 -6942 3711 -6933
rect 3745 -6942 3783 -6933
rect 3817 -6942 3855 -6933
rect 3889 -6942 3927 -6933
rect 3961 -6942 3999 -6933
rect 4033 -6942 4071 -6933
rect 4105 -6942 4143 -6933
rect 4177 -6942 4215 -6933
rect 4249 -6942 4287 -6933
rect 4321 -6942 4359 -6933
rect 4393 -6942 4431 -6933
rect 4465 -6942 4503 -6933
rect 4537 -6942 4575 -6933
rect 4609 -6942 4647 -6933
rect 4681 -6942 4719 -6933
rect 4753 -6942 4791 -6933
rect 4825 -6942 4863 -6933
rect 4897 -6942 4935 -6933
rect 4969 -6942 5007 -6933
rect 5041 -6942 5079 -6933
rect 5113 -6942 6567 -6933
rect 6601 -6942 6639 -6933
rect 6673 -6942 6711 -6933
rect 6745 -6942 6783 -6933
rect 6817 -6942 6855 -6933
rect 6889 -6942 6927 -6933
rect 6961 -6942 6999 -6933
rect 7033 -6942 7071 -6933
rect 7105 -6942 7143 -6933
rect 7177 -6942 7215 -6933
rect 7249 -6942 7287 -6933
rect 7321 -6942 7359 -6933
rect 7393 -6942 7431 -6933
rect 7465 -6942 7503 -6933
rect 7537 -6942 7575 -6933
rect 7609 -6942 7647 -6933
rect 7681 -6942 7719 -6933
rect 7753 -6942 7791 -6933
rect 7825 -6942 7863 -6933
rect 7897 -6942 7935 -6933
rect 7969 -6942 8007 -6933
rect 8041 -6942 8079 -6933
rect 8113 -6942 9740 -6933
rect 540 -7058 580 -6967
rect 9720 -7058 9740 -6942
rect 540 -7100 9740 -7058
<< via1 >>
rect -1745 3379 -1693 3431
rect -1681 3379 -1629 3431
rect -1617 3379 -1565 3431
rect -1553 3379 -1501 3431
rect -1489 3379 -1437 3431
rect -1425 3379 -1373 3431
rect -1361 3379 -1309 3431
rect -1297 3379 -1245 3431
rect -1233 3379 -1181 3431
rect -1169 3379 -1117 3431
rect -1105 3379 -1053 3431
rect -1041 3379 -989 3431
rect -977 3379 -925 3431
rect 69 3379 121 3431
rect 3069 3379 3121 3431
rect 6069 3379 6121 3431
rect -1566 1499 -1514 1551
rect -1502 1499 -1450 1551
rect -1438 1499 -1386 1551
rect -1374 1499 -1322 1551
rect -1310 1499 -1258 1551
rect -1246 1499 -1194 1551
rect -522 1499 -470 1551
rect -458 1499 -406 1551
rect -394 1499 -342 1551
rect -330 1499 -278 1551
rect -1566 -1501 -1514 -1449
rect -1502 -1501 -1450 -1449
rect -1438 -1501 -1386 -1449
rect -1374 -1501 -1322 -1449
rect -1310 -1501 -1258 -1449
rect -1246 -1501 -1194 -1449
rect -522 -1501 -470 -1449
rect -458 -1501 -406 -1449
rect -394 -1501 -342 -1449
rect -330 -1501 -278 -1449
rect -1566 -4501 -1514 -4449
rect -1502 -4501 -1450 -4449
rect -1438 -4501 -1386 -4449
rect -1374 -4501 -1322 -4449
rect -1310 -4501 -1258 -4449
rect -1246 -4501 -1194 -4449
rect -522 -4501 -470 -4449
rect -458 -4501 -406 -4449
rect -394 -4501 -342 -4449
rect -330 -4501 -278 -4449
rect 578 -6191 630 -6139
rect 642 -6191 694 -6139
rect 706 -6191 758 -6139
rect 770 -6191 822 -6139
rect 834 -6191 886 -6139
rect 898 -6191 950 -6139
rect 962 -6191 1014 -6139
rect 1026 -6191 1078 -6139
rect 1090 -6191 1142 -6139
rect 1154 -6191 1206 -6139
rect 1218 -6191 1270 -6139
rect 1282 -6191 1334 -6139
rect 1346 -6191 1398 -6139
rect 1410 -6191 1462 -6139
rect 1474 -6191 1526 -6139
rect 1538 -6191 1590 -6139
rect 1602 -6191 1654 -6139
rect 1666 -6191 1718 -6139
rect 1730 -6191 1782 -6139
rect 1794 -6191 1846 -6139
rect 1858 -6191 1910 -6139
rect 1922 -6191 1974 -6139
rect 1986 -6191 2038 -6139
rect 2050 -6191 2102 -6139
rect 3578 -6191 3630 -6139
rect 3642 -6191 3694 -6139
rect 3706 -6191 3758 -6139
rect 3770 -6191 3822 -6139
rect 3834 -6191 3886 -6139
rect 3898 -6191 3950 -6139
rect 3962 -6191 4014 -6139
rect 4026 -6191 4078 -6139
rect 4090 -6191 4142 -6139
rect 4154 -6191 4206 -6139
rect 4218 -6191 4270 -6139
rect 4282 -6191 4334 -6139
rect 4346 -6191 4398 -6139
rect 4410 -6191 4462 -6139
rect 4474 -6191 4526 -6139
rect 4538 -6191 4590 -6139
rect 4602 -6191 4654 -6139
rect 4666 -6191 4718 -6139
rect 4730 -6191 4782 -6139
rect 4794 -6191 4846 -6139
rect 4858 -6191 4910 -6139
rect 4922 -6191 4974 -6139
rect 4986 -6191 5038 -6139
rect 5050 -6191 5102 -6139
rect 6578 -6191 6630 -6139
rect 6642 -6191 6694 -6139
rect 6706 -6191 6758 -6139
rect 6770 -6191 6822 -6139
rect 6834 -6191 6886 -6139
rect 6898 -6191 6950 -6139
rect 6962 -6191 7014 -6139
rect 7026 -6191 7078 -6139
rect 7090 -6191 7142 -6139
rect 7154 -6191 7206 -6139
rect 7218 -6191 7270 -6139
rect 7282 -6191 7334 -6139
rect 7346 -6191 7398 -6139
rect 7410 -6191 7462 -6139
rect 7474 -6191 7526 -6139
rect 7538 -6191 7590 -6139
rect 7602 -6191 7654 -6139
rect 7666 -6191 7718 -6139
rect 7730 -6191 7782 -6139
rect 7794 -6191 7846 -6139
rect 7858 -6191 7910 -6139
rect 7922 -6191 7974 -6139
rect 7986 -6191 8038 -6139
rect 8050 -6191 8102 -6139
rect 240 -6511 420 -6510
rect 240 -6689 241 -6511
rect 241 -6689 419 -6511
rect 419 -6689 420 -6511
rect 240 -6690 420 -6689
rect 3240 -6511 3420 -6510
rect 3240 -6689 3241 -6511
rect 3241 -6689 3419 -6511
rect 3419 -6689 3420 -6511
rect 3240 -6690 3420 -6689
rect 6240 -6511 6420 -6510
rect 6240 -6689 6241 -6511
rect 6241 -6689 6419 -6511
rect 6419 -6689 6420 -6511
rect 6240 -6690 6420 -6689
rect 580 -6967 601 -6942
rect 601 -6967 639 -6942
rect 639 -6967 673 -6942
rect 673 -6967 711 -6942
rect 711 -6967 745 -6942
rect 745 -6967 783 -6942
rect 783 -6967 817 -6942
rect 817 -6967 855 -6942
rect 855 -6967 889 -6942
rect 889 -6967 927 -6942
rect 927 -6967 961 -6942
rect 961 -6967 999 -6942
rect 999 -6967 1033 -6942
rect 1033 -6967 1071 -6942
rect 1071 -6967 1105 -6942
rect 1105 -6967 1143 -6942
rect 1143 -6967 1177 -6942
rect 1177 -6967 1215 -6942
rect 1215 -6967 1249 -6942
rect 1249 -6967 1287 -6942
rect 1287 -6967 1321 -6942
rect 1321 -6967 1359 -6942
rect 1359 -6967 1393 -6942
rect 1393 -6967 1431 -6942
rect 1431 -6967 1465 -6942
rect 1465 -6967 1503 -6942
rect 1503 -6967 1537 -6942
rect 1537 -6967 1575 -6942
rect 1575 -6967 1609 -6942
rect 1609 -6967 1647 -6942
rect 1647 -6967 1681 -6942
rect 1681 -6967 1719 -6942
rect 1719 -6967 1753 -6942
rect 1753 -6967 1791 -6942
rect 1791 -6967 1825 -6942
rect 1825 -6967 1863 -6942
rect 1863 -6967 1897 -6942
rect 1897 -6967 1935 -6942
rect 1935 -6967 1969 -6942
rect 1969 -6967 2007 -6942
rect 2007 -6967 2041 -6942
rect 2041 -6967 2079 -6942
rect 2079 -6967 2113 -6942
rect 2113 -6967 3567 -6942
rect 3567 -6967 3601 -6942
rect 3601 -6967 3639 -6942
rect 3639 -6967 3673 -6942
rect 3673 -6967 3711 -6942
rect 3711 -6967 3745 -6942
rect 3745 -6967 3783 -6942
rect 3783 -6967 3817 -6942
rect 3817 -6967 3855 -6942
rect 3855 -6967 3889 -6942
rect 3889 -6967 3927 -6942
rect 3927 -6967 3961 -6942
rect 3961 -6967 3999 -6942
rect 3999 -6967 4033 -6942
rect 4033 -6967 4071 -6942
rect 4071 -6967 4105 -6942
rect 4105 -6967 4143 -6942
rect 4143 -6967 4177 -6942
rect 4177 -6967 4215 -6942
rect 4215 -6967 4249 -6942
rect 4249 -6967 4287 -6942
rect 4287 -6967 4321 -6942
rect 4321 -6967 4359 -6942
rect 4359 -6967 4393 -6942
rect 4393 -6967 4431 -6942
rect 4431 -6967 4465 -6942
rect 4465 -6967 4503 -6942
rect 4503 -6967 4537 -6942
rect 4537 -6967 4575 -6942
rect 4575 -6967 4609 -6942
rect 4609 -6967 4647 -6942
rect 4647 -6967 4681 -6942
rect 4681 -6967 4719 -6942
rect 4719 -6967 4753 -6942
rect 4753 -6967 4791 -6942
rect 4791 -6967 4825 -6942
rect 4825 -6967 4863 -6942
rect 4863 -6967 4897 -6942
rect 4897 -6967 4935 -6942
rect 4935 -6967 4969 -6942
rect 4969 -6967 5007 -6942
rect 5007 -6967 5041 -6942
rect 5041 -6967 5079 -6942
rect 5079 -6967 5113 -6942
rect 5113 -6967 6567 -6942
rect 6567 -6967 6601 -6942
rect 6601 -6967 6639 -6942
rect 6639 -6967 6673 -6942
rect 6673 -6967 6711 -6942
rect 6711 -6967 6745 -6942
rect 6745 -6967 6783 -6942
rect 6783 -6967 6817 -6942
rect 6817 -6967 6855 -6942
rect 6855 -6967 6889 -6942
rect 6889 -6967 6927 -6942
rect 6927 -6967 6961 -6942
rect 6961 -6967 6999 -6942
rect 6999 -6967 7033 -6942
rect 7033 -6967 7071 -6942
rect 7071 -6967 7105 -6942
rect 7105 -6967 7143 -6942
rect 7143 -6967 7177 -6942
rect 7177 -6967 7215 -6942
rect 7215 -6967 7249 -6942
rect 7249 -6967 7287 -6942
rect 7287 -6967 7321 -6942
rect 7321 -6967 7359 -6942
rect 7359 -6967 7393 -6942
rect 7393 -6967 7431 -6942
rect 7431 -6967 7465 -6942
rect 7465 -6967 7503 -6942
rect 7503 -6967 7537 -6942
rect 7537 -6967 7575 -6942
rect 7575 -6967 7609 -6942
rect 7609 -6967 7647 -6942
rect 7647 -6967 7681 -6942
rect 7681 -6967 7719 -6942
rect 7719 -6967 7753 -6942
rect 7753 -6967 7791 -6942
rect 7791 -6967 7825 -6942
rect 7825 -6967 7863 -6942
rect 7863 -6967 7897 -6942
rect 7897 -6967 7935 -6942
rect 7935 -6967 7969 -6942
rect 7969 -6967 8007 -6942
rect 8007 -6967 8041 -6942
rect 8041 -6967 8079 -6942
rect 8079 -6967 8113 -6942
rect 8113 -6967 9720 -6942
rect 580 -7058 9720 -6967
<< metal2 >>
rect 0 4040 9000 4150
rect -3000 3431 -890 3460
rect -3000 3379 -1745 3431
rect -1693 3379 -1681 3431
rect -1629 3379 -1617 3431
rect -1565 3379 -1553 3431
rect -1501 3379 -1489 3431
rect -1437 3379 -1425 3431
rect -1373 3379 -1361 3431
rect -1309 3379 -1297 3431
rect -1245 3379 -1233 3431
rect -1181 3379 -1169 3431
rect -1117 3379 -1105 3431
rect -1053 3379 -1041 3431
rect -989 3379 -977 3431
rect -925 3379 -890 3431
rect -3000 3350 -890 3379
rect -3000 1551 -1000 1570
rect -3000 1499 -1566 1551
rect -1514 1499 -1502 1551
rect -1450 1499 -1438 1551
rect -1386 1499 -1374 1551
rect -1322 1499 -1310 1551
rect -1258 1499 -1246 1551
rect -1194 1499 -1000 1551
rect -3000 1480 -1000 1499
rect -750 223 -640 4000
rect 480 3633 590 3660
rect 60 3460 130 3600
rect 480 3577 507 3633
rect 563 3577 590 3633
rect 480 3550 590 3577
rect 40 3431 150 3460
rect 40 3379 69 3431
rect 121 3379 150 3431
rect 40 3350 150 3379
rect 60 3000 130 3350
rect 500 3000 570 3550
rect 1020 3000 1090 4040
rect 3480 3633 3590 3660
rect 3060 3460 3130 3600
rect 3480 3577 3507 3633
rect 3563 3577 3590 3633
rect 3480 3550 3590 3577
rect 3040 3431 3150 3460
rect 3040 3379 3069 3431
rect 3121 3379 3150 3431
rect 3040 3350 3150 3379
rect 3060 3000 3130 3350
rect 3500 3000 3570 3550
rect 4020 3000 4090 4040
rect 6480 3633 6590 3660
rect 6060 3460 6130 3600
rect 6480 3577 6507 3633
rect 6563 3577 6590 3633
rect 6480 3550 6590 3577
rect 6040 3431 6150 3460
rect 6040 3379 6069 3431
rect 6121 3379 6150 3431
rect 6040 3350 6150 3379
rect 6060 3000 6130 3350
rect 6500 3000 6570 3550
rect 7020 3000 7090 4040
rect -560 1553 -260 1570
rect -560 1551 -508 1553
rect -452 1551 -428 1553
rect -372 1551 -348 1553
rect -292 1551 -260 1553
rect -560 1499 -522 1551
rect -278 1499 -260 1551
rect -560 1497 -508 1499
rect -452 1497 -428 1499
rect -372 1497 -348 1499
rect -292 1497 -260 1499
rect -560 1480 -260 1497
rect -750 167 -723 223
rect -667 167 -640 223
rect -3000 -1449 -1000 -1430
rect -3000 -1501 -1566 -1449
rect -1514 -1501 -1502 -1449
rect -1450 -1501 -1438 -1449
rect -1386 -1501 -1374 -1449
rect -1322 -1501 -1310 -1449
rect -1258 -1501 -1246 -1449
rect -1194 -1501 -1000 -1449
rect -3000 -1520 -1000 -1501
rect -750 -2777 -640 167
rect -560 -1447 -260 -1430
rect -560 -1449 -508 -1447
rect -452 -1449 -428 -1447
rect -372 -1449 -348 -1447
rect -292 -1449 -260 -1447
rect -560 -1501 -522 -1449
rect -278 -1501 -260 -1449
rect -560 -1503 -508 -1501
rect -452 -1503 -428 -1501
rect -372 -1503 -348 -1501
rect -292 -1503 -260 -1501
rect -560 -1520 -260 -1503
rect -750 -2833 -723 -2777
rect -667 -2833 -640 -2777
rect -3000 -4449 -1000 -4430
rect -3000 -4501 -1566 -4449
rect -1514 -4501 -1502 -4449
rect -1450 -4501 -1438 -4449
rect -1386 -4501 -1374 -4449
rect -1322 -4501 -1310 -4449
rect -1258 -4501 -1246 -4449
rect -1194 -4501 -1000 -4449
rect -3000 -4520 -1000 -4501
rect -750 -5777 -640 -2833
rect -560 -4447 -260 -4430
rect -560 -4449 -508 -4447
rect -452 -4449 -428 -4447
rect -372 -4449 -348 -4447
rect -292 -4449 -260 -4447
rect -560 -4501 -522 -4449
rect -278 -4501 -260 -4449
rect -560 -4503 -508 -4501
rect -452 -4503 -428 -4501
rect -372 -4503 -348 -4501
rect -292 -4503 -260 -4501
rect -560 -4520 -260 -4503
rect -750 -5833 -723 -5777
rect -667 -5833 -640 -5777
rect -750 -6000 -640 -5833
rect 540 -6102 2780 -6060
rect 540 -6139 592 -6102
rect 648 -6139 672 -6102
rect 728 -6139 752 -6102
rect 808 -6139 832 -6102
rect 888 -6139 912 -6102
rect 968 -6139 992 -6102
rect 1048 -6139 1072 -6102
rect 1128 -6139 1152 -6102
rect 1208 -6139 1232 -6102
rect 1288 -6139 1312 -6102
rect 1368 -6139 1392 -6102
rect 1448 -6139 1472 -6102
rect 1528 -6139 1552 -6102
rect 1608 -6139 1632 -6102
rect 1688 -6139 1712 -6102
rect 1768 -6139 1792 -6102
rect 1848 -6139 1872 -6102
rect 1928 -6139 1952 -6102
rect 2008 -6139 2032 -6102
rect 2088 -6139 2112 -6102
rect 540 -6191 578 -6139
rect 822 -6158 832 -6139
rect 888 -6158 898 -6139
rect 1142 -6158 1152 -6139
rect 1208 -6158 1218 -6139
rect 1462 -6158 1472 -6139
rect 1528 -6158 1538 -6139
rect 1782 -6158 1792 -6139
rect 1848 -6158 1858 -6139
rect 2102 -6158 2112 -6139
rect 2168 -6158 2192 -6102
rect 2248 -6158 2272 -6102
rect 2328 -6158 2352 -6102
rect 2408 -6158 2432 -6102
rect 2488 -6158 2512 -6102
rect 2568 -6158 2592 -6102
rect 2648 -6158 2672 -6102
rect 2728 -6158 2780 -6102
rect 630 -6191 642 -6158
rect 694 -6191 706 -6158
rect 758 -6191 770 -6158
rect 822 -6191 834 -6158
rect 886 -6191 898 -6158
rect 950 -6191 962 -6158
rect 1014 -6191 1026 -6158
rect 1078 -6191 1090 -6158
rect 1142 -6191 1154 -6158
rect 1206 -6191 1218 -6158
rect 1270 -6191 1282 -6158
rect 1334 -6191 1346 -6158
rect 1398 -6191 1410 -6158
rect 1462 -6191 1474 -6158
rect 1526 -6191 1538 -6158
rect 1590 -6191 1602 -6158
rect 1654 -6191 1666 -6158
rect 1718 -6191 1730 -6158
rect 1782 -6191 1794 -6158
rect 1846 -6191 1858 -6158
rect 1910 -6191 1922 -6158
rect 1974 -6191 1986 -6158
rect 2038 -6191 2050 -6158
rect 2102 -6191 2780 -6158
rect 540 -6200 2780 -6191
rect 3540 -6102 5780 -6060
rect 3540 -6139 3592 -6102
rect 3648 -6139 3672 -6102
rect 3728 -6139 3752 -6102
rect 3808 -6139 3832 -6102
rect 3888 -6139 3912 -6102
rect 3968 -6139 3992 -6102
rect 4048 -6139 4072 -6102
rect 4128 -6139 4152 -6102
rect 4208 -6139 4232 -6102
rect 4288 -6139 4312 -6102
rect 4368 -6139 4392 -6102
rect 4448 -6139 4472 -6102
rect 4528 -6139 4552 -6102
rect 4608 -6139 4632 -6102
rect 4688 -6139 4712 -6102
rect 4768 -6139 4792 -6102
rect 4848 -6139 4872 -6102
rect 4928 -6139 4952 -6102
rect 5008 -6139 5032 -6102
rect 5088 -6139 5112 -6102
rect 3540 -6191 3578 -6139
rect 3822 -6158 3832 -6139
rect 3888 -6158 3898 -6139
rect 4142 -6158 4152 -6139
rect 4208 -6158 4218 -6139
rect 4462 -6158 4472 -6139
rect 4528 -6158 4538 -6139
rect 4782 -6158 4792 -6139
rect 4848 -6158 4858 -6139
rect 5102 -6158 5112 -6139
rect 5168 -6158 5192 -6102
rect 5248 -6158 5272 -6102
rect 5328 -6158 5352 -6102
rect 5408 -6158 5432 -6102
rect 5488 -6158 5512 -6102
rect 5568 -6158 5592 -6102
rect 5648 -6158 5672 -6102
rect 5728 -6158 5780 -6102
rect 3630 -6191 3642 -6158
rect 3694 -6191 3706 -6158
rect 3758 -6191 3770 -6158
rect 3822 -6191 3834 -6158
rect 3886 -6191 3898 -6158
rect 3950 -6191 3962 -6158
rect 4014 -6191 4026 -6158
rect 4078 -6191 4090 -6158
rect 4142 -6191 4154 -6158
rect 4206 -6191 4218 -6158
rect 4270 -6191 4282 -6158
rect 4334 -6191 4346 -6158
rect 4398 -6191 4410 -6158
rect 4462 -6191 4474 -6158
rect 4526 -6191 4538 -6158
rect 4590 -6191 4602 -6158
rect 4654 -6191 4666 -6158
rect 4718 -6191 4730 -6158
rect 4782 -6191 4794 -6158
rect 4846 -6191 4858 -6158
rect 4910 -6191 4922 -6158
rect 4974 -6191 4986 -6158
rect 5038 -6191 5050 -6158
rect 5102 -6191 5780 -6158
rect 3540 -6200 5780 -6191
rect 6540 -6102 8780 -6060
rect 6540 -6139 6592 -6102
rect 6648 -6139 6672 -6102
rect 6728 -6139 6752 -6102
rect 6808 -6139 6832 -6102
rect 6888 -6139 6912 -6102
rect 6968 -6139 6992 -6102
rect 7048 -6139 7072 -6102
rect 7128 -6139 7152 -6102
rect 7208 -6139 7232 -6102
rect 7288 -6139 7312 -6102
rect 7368 -6139 7392 -6102
rect 7448 -6139 7472 -6102
rect 7528 -6139 7552 -6102
rect 7608 -6139 7632 -6102
rect 7688 -6139 7712 -6102
rect 7768 -6139 7792 -6102
rect 7848 -6139 7872 -6102
rect 7928 -6139 7952 -6102
rect 8008 -6139 8032 -6102
rect 8088 -6139 8112 -6102
rect 6540 -6191 6578 -6139
rect 6822 -6158 6832 -6139
rect 6888 -6158 6898 -6139
rect 7142 -6158 7152 -6139
rect 7208 -6158 7218 -6139
rect 7462 -6158 7472 -6139
rect 7528 -6158 7538 -6139
rect 7782 -6158 7792 -6139
rect 7848 -6158 7858 -6139
rect 8102 -6158 8112 -6139
rect 8168 -6158 8192 -6102
rect 8248 -6158 8272 -6102
rect 8328 -6158 8352 -6102
rect 8408 -6158 8432 -6102
rect 8488 -6158 8512 -6102
rect 8568 -6158 8592 -6102
rect 8648 -6158 8672 -6102
rect 8728 -6158 8780 -6102
rect 6630 -6191 6642 -6158
rect 6694 -6191 6706 -6158
rect 6758 -6191 6770 -6158
rect 6822 -6191 6834 -6158
rect 6886 -6191 6898 -6158
rect 6950 -6191 6962 -6158
rect 7014 -6191 7026 -6158
rect 7078 -6191 7090 -6158
rect 7142 -6191 7154 -6158
rect 7206 -6191 7218 -6158
rect 7270 -6191 7282 -6158
rect 7334 -6191 7346 -6158
rect 7398 -6191 7410 -6158
rect 7462 -6191 7474 -6158
rect 7526 -6191 7538 -6158
rect 7590 -6191 7602 -6158
rect 7654 -6191 7666 -6158
rect 7718 -6191 7730 -6158
rect 7782 -6191 7794 -6158
rect 7846 -6191 7858 -6158
rect 7910 -6191 7922 -6158
rect 7974 -6191 7986 -6158
rect 8038 -6191 8050 -6158
rect 8102 -6191 8780 -6158
rect 6540 -6200 8780 -6191
rect 220 -6510 440 -6490
rect 220 -6690 240 -6510
rect 420 -6690 440 -6510
rect 220 -6710 440 -6690
rect 3220 -6510 3440 -6490
rect 3220 -6690 3240 -6510
rect 3420 -6690 3440 -6510
rect 3220 -6710 3440 -6690
rect 6220 -6510 6440 -6490
rect 6220 -6690 6240 -6510
rect 6420 -6690 6440 -6510
rect 6220 -6710 6440 -6690
rect 540 -6942 9740 -6900
rect 540 -7058 580 -6942
rect 9720 -7058 9740 -6942
rect 540 -7100 9740 -7058
<< via2 >>
rect 507 3577 563 3633
rect 3507 3577 3563 3633
rect 6507 3577 6563 3633
rect -508 1551 -452 1553
rect -428 1551 -372 1553
rect -348 1551 -292 1553
rect -508 1499 -470 1551
rect -470 1499 -458 1551
rect -458 1499 -452 1551
rect -428 1499 -406 1551
rect -406 1499 -394 1551
rect -394 1499 -372 1551
rect -348 1499 -342 1551
rect -342 1499 -330 1551
rect -330 1499 -292 1551
rect -508 1497 -452 1499
rect -428 1497 -372 1499
rect -348 1497 -292 1499
rect -723 167 -667 223
rect -508 -1449 -452 -1447
rect -428 -1449 -372 -1447
rect -348 -1449 -292 -1447
rect -508 -1501 -470 -1449
rect -470 -1501 -458 -1449
rect -458 -1501 -452 -1449
rect -428 -1501 -406 -1449
rect -406 -1501 -394 -1449
rect -394 -1501 -372 -1449
rect -348 -1501 -342 -1449
rect -342 -1501 -330 -1449
rect -330 -1501 -292 -1449
rect -508 -1503 -452 -1501
rect -428 -1503 -372 -1501
rect -348 -1503 -292 -1501
rect -723 -2833 -667 -2777
rect -508 -4449 -452 -4447
rect -428 -4449 -372 -4447
rect -348 -4449 -292 -4447
rect -508 -4501 -470 -4449
rect -470 -4501 -458 -4449
rect -458 -4501 -452 -4449
rect -428 -4501 -406 -4449
rect -406 -4501 -394 -4449
rect -394 -4501 -372 -4449
rect -348 -4501 -342 -4449
rect -342 -4501 -330 -4449
rect -330 -4501 -292 -4449
rect -508 -4503 -452 -4501
rect -428 -4503 -372 -4501
rect -348 -4503 -292 -4501
rect -723 -5833 -667 -5777
rect 592 -6139 648 -6102
rect 672 -6139 728 -6102
rect 752 -6139 808 -6102
rect 832 -6139 888 -6102
rect 912 -6139 968 -6102
rect 992 -6139 1048 -6102
rect 1072 -6139 1128 -6102
rect 1152 -6139 1208 -6102
rect 1232 -6139 1288 -6102
rect 1312 -6139 1368 -6102
rect 1392 -6139 1448 -6102
rect 1472 -6139 1528 -6102
rect 1552 -6139 1608 -6102
rect 1632 -6139 1688 -6102
rect 1712 -6139 1768 -6102
rect 1792 -6139 1848 -6102
rect 1872 -6139 1928 -6102
rect 1952 -6139 2008 -6102
rect 2032 -6139 2088 -6102
rect 592 -6158 630 -6139
rect 630 -6158 642 -6139
rect 642 -6158 648 -6139
rect 672 -6158 694 -6139
rect 694 -6158 706 -6139
rect 706 -6158 728 -6139
rect 752 -6158 758 -6139
rect 758 -6158 770 -6139
rect 770 -6158 808 -6139
rect 832 -6158 834 -6139
rect 834 -6158 886 -6139
rect 886 -6158 888 -6139
rect 912 -6158 950 -6139
rect 950 -6158 962 -6139
rect 962 -6158 968 -6139
rect 992 -6158 1014 -6139
rect 1014 -6158 1026 -6139
rect 1026 -6158 1048 -6139
rect 1072 -6158 1078 -6139
rect 1078 -6158 1090 -6139
rect 1090 -6158 1128 -6139
rect 1152 -6158 1154 -6139
rect 1154 -6158 1206 -6139
rect 1206 -6158 1208 -6139
rect 1232 -6158 1270 -6139
rect 1270 -6158 1282 -6139
rect 1282 -6158 1288 -6139
rect 1312 -6158 1334 -6139
rect 1334 -6158 1346 -6139
rect 1346 -6158 1368 -6139
rect 1392 -6158 1398 -6139
rect 1398 -6158 1410 -6139
rect 1410 -6158 1448 -6139
rect 1472 -6158 1474 -6139
rect 1474 -6158 1526 -6139
rect 1526 -6158 1528 -6139
rect 1552 -6158 1590 -6139
rect 1590 -6158 1602 -6139
rect 1602 -6158 1608 -6139
rect 1632 -6158 1654 -6139
rect 1654 -6158 1666 -6139
rect 1666 -6158 1688 -6139
rect 1712 -6158 1718 -6139
rect 1718 -6158 1730 -6139
rect 1730 -6158 1768 -6139
rect 1792 -6158 1794 -6139
rect 1794 -6158 1846 -6139
rect 1846 -6158 1848 -6139
rect 1872 -6158 1910 -6139
rect 1910 -6158 1922 -6139
rect 1922 -6158 1928 -6139
rect 1952 -6158 1974 -6139
rect 1974 -6158 1986 -6139
rect 1986 -6158 2008 -6139
rect 2032 -6158 2038 -6139
rect 2038 -6158 2050 -6139
rect 2050 -6158 2088 -6139
rect 2112 -6158 2168 -6102
rect 2192 -6158 2248 -6102
rect 2272 -6158 2328 -6102
rect 2352 -6158 2408 -6102
rect 2432 -6158 2488 -6102
rect 2512 -6158 2568 -6102
rect 2592 -6158 2648 -6102
rect 2672 -6158 2728 -6102
rect 3592 -6139 3648 -6102
rect 3672 -6139 3728 -6102
rect 3752 -6139 3808 -6102
rect 3832 -6139 3888 -6102
rect 3912 -6139 3968 -6102
rect 3992 -6139 4048 -6102
rect 4072 -6139 4128 -6102
rect 4152 -6139 4208 -6102
rect 4232 -6139 4288 -6102
rect 4312 -6139 4368 -6102
rect 4392 -6139 4448 -6102
rect 4472 -6139 4528 -6102
rect 4552 -6139 4608 -6102
rect 4632 -6139 4688 -6102
rect 4712 -6139 4768 -6102
rect 4792 -6139 4848 -6102
rect 4872 -6139 4928 -6102
rect 4952 -6139 5008 -6102
rect 5032 -6139 5088 -6102
rect 3592 -6158 3630 -6139
rect 3630 -6158 3642 -6139
rect 3642 -6158 3648 -6139
rect 3672 -6158 3694 -6139
rect 3694 -6158 3706 -6139
rect 3706 -6158 3728 -6139
rect 3752 -6158 3758 -6139
rect 3758 -6158 3770 -6139
rect 3770 -6158 3808 -6139
rect 3832 -6158 3834 -6139
rect 3834 -6158 3886 -6139
rect 3886 -6158 3888 -6139
rect 3912 -6158 3950 -6139
rect 3950 -6158 3962 -6139
rect 3962 -6158 3968 -6139
rect 3992 -6158 4014 -6139
rect 4014 -6158 4026 -6139
rect 4026 -6158 4048 -6139
rect 4072 -6158 4078 -6139
rect 4078 -6158 4090 -6139
rect 4090 -6158 4128 -6139
rect 4152 -6158 4154 -6139
rect 4154 -6158 4206 -6139
rect 4206 -6158 4208 -6139
rect 4232 -6158 4270 -6139
rect 4270 -6158 4282 -6139
rect 4282 -6158 4288 -6139
rect 4312 -6158 4334 -6139
rect 4334 -6158 4346 -6139
rect 4346 -6158 4368 -6139
rect 4392 -6158 4398 -6139
rect 4398 -6158 4410 -6139
rect 4410 -6158 4448 -6139
rect 4472 -6158 4474 -6139
rect 4474 -6158 4526 -6139
rect 4526 -6158 4528 -6139
rect 4552 -6158 4590 -6139
rect 4590 -6158 4602 -6139
rect 4602 -6158 4608 -6139
rect 4632 -6158 4654 -6139
rect 4654 -6158 4666 -6139
rect 4666 -6158 4688 -6139
rect 4712 -6158 4718 -6139
rect 4718 -6158 4730 -6139
rect 4730 -6158 4768 -6139
rect 4792 -6158 4794 -6139
rect 4794 -6158 4846 -6139
rect 4846 -6158 4848 -6139
rect 4872 -6158 4910 -6139
rect 4910 -6158 4922 -6139
rect 4922 -6158 4928 -6139
rect 4952 -6158 4974 -6139
rect 4974 -6158 4986 -6139
rect 4986 -6158 5008 -6139
rect 5032 -6158 5038 -6139
rect 5038 -6158 5050 -6139
rect 5050 -6158 5088 -6139
rect 5112 -6158 5168 -6102
rect 5192 -6158 5248 -6102
rect 5272 -6158 5328 -6102
rect 5352 -6158 5408 -6102
rect 5432 -6158 5488 -6102
rect 5512 -6158 5568 -6102
rect 5592 -6158 5648 -6102
rect 5672 -6158 5728 -6102
rect 6592 -6139 6648 -6102
rect 6672 -6139 6728 -6102
rect 6752 -6139 6808 -6102
rect 6832 -6139 6888 -6102
rect 6912 -6139 6968 -6102
rect 6992 -6139 7048 -6102
rect 7072 -6139 7128 -6102
rect 7152 -6139 7208 -6102
rect 7232 -6139 7288 -6102
rect 7312 -6139 7368 -6102
rect 7392 -6139 7448 -6102
rect 7472 -6139 7528 -6102
rect 7552 -6139 7608 -6102
rect 7632 -6139 7688 -6102
rect 7712 -6139 7768 -6102
rect 7792 -6139 7848 -6102
rect 7872 -6139 7928 -6102
rect 7952 -6139 8008 -6102
rect 8032 -6139 8088 -6102
rect 6592 -6158 6630 -6139
rect 6630 -6158 6642 -6139
rect 6642 -6158 6648 -6139
rect 6672 -6158 6694 -6139
rect 6694 -6158 6706 -6139
rect 6706 -6158 6728 -6139
rect 6752 -6158 6758 -6139
rect 6758 -6158 6770 -6139
rect 6770 -6158 6808 -6139
rect 6832 -6158 6834 -6139
rect 6834 -6158 6886 -6139
rect 6886 -6158 6888 -6139
rect 6912 -6158 6950 -6139
rect 6950 -6158 6962 -6139
rect 6962 -6158 6968 -6139
rect 6992 -6158 7014 -6139
rect 7014 -6158 7026 -6139
rect 7026 -6158 7048 -6139
rect 7072 -6158 7078 -6139
rect 7078 -6158 7090 -6139
rect 7090 -6158 7128 -6139
rect 7152 -6158 7154 -6139
rect 7154 -6158 7206 -6139
rect 7206 -6158 7208 -6139
rect 7232 -6158 7270 -6139
rect 7270 -6158 7282 -6139
rect 7282 -6158 7288 -6139
rect 7312 -6158 7334 -6139
rect 7334 -6158 7346 -6139
rect 7346 -6158 7368 -6139
rect 7392 -6158 7398 -6139
rect 7398 -6158 7410 -6139
rect 7410 -6158 7448 -6139
rect 7472 -6158 7474 -6139
rect 7474 -6158 7526 -6139
rect 7526 -6158 7528 -6139
rect 7552 -6158 7590 -6139
rect 7590 -6158 7602 -6139
rect 7602 -6158 7608 -6139
rect 7632 -6158 7654 -6139
rect 7654 -6158 7666 -6139
rect 7666 -6158 7688 -6139
rect 7712 -6158 7718 -6139
rect 7718 -6158 7730 -6139
rect 7730 -6158 7768 -6139
rect 7792 -6158 7794 -6139
rect 7794 -6158 7846 -6139
rect 7846 -6158 7848 -6139
rect 7872 -6158 7910 -6139
rect 7910 -6158 7922 -6139
rect 7922 -6158 7928 -6139
rect 7952 -6158 7974 -6139
rect 7974 -6158 7986 -6139
rect 7986 -6158 8008 -6139
rect 8032 -6158 8038 -6139
rect 8038 -6158 8050 -6139
rect 8050 -6158 8088 -6139
rect 8112 -6158 8168 -6102
rect 8192 -6158 8248 -6102
rect 8272 -6158 8328 -6102
rect 8352 -6158 8408 -6102
rect 8432 -6158 8488 -6102
rect 8512 -6158 8568 -6102
rect 8592 -6158 8648 -6102
rect 8672 -6158 8728 -6102
rect 262 -6668 398 -6532
rect 3262 -6668 3398 -6532
rect 6262 -6668 6398 -6532
<< metal3 >>
rect -1200 2840 -1110 5000
rect 480 3637 590 3660
rect 480 3573 503 3637
rect 567 3573 590 3637
rect 480 3550 590 3573
rect 3480 3637 3590 3660
rect 3480 3573 3503 3637
rect 3567 3573 3590 3637
rect 3480 3550 3590 3573
rect 6480 3637 6590 3660
rect 6480 3573 6503 3637
rect 6567 3573 6590 3637
rect 6480 3550 6590 3573
rect -1200 2750 200 2840
rect -1200 -160 -1110 2750
rect -480 2550 -370 2560
rect -560 2537 520 2550
rect -560 2473 -457 2537
rect -393 2473 520 2537
rect -560 2460 520 2473
rect -480 2450 -370 2460
rect -560 1553 440 1570
rect -560 1497 -508 1553
rect -452 1497 -428 1553
rect -372 1497 -348 1553
rect -292 1497 440 1553
rect -560 1480 440 1497
rect -760 223 40 250
rect -760 167 -723 223
rect -667 167 40 223
rect -760 160 40 167
rect -750 140 -640 160
rect -1200 -250 200 -160
rect -1200 -3160 -1110 -250
rect -480 -450 -370 -440
rect -560 -463 520 -450
rect -560 -527 -457 -463
rect -393 -527 520 -463
rect -560 -540 520 -527
rect -480 -550 -370 -540
rect -560 -1447 440 -1430
rect -560 -1503 -508 -1447
rect -452 -1503 -428 -1447
rect -372 -1503 -348 -1447
rect -292 -1503 440 -1447
rect -560 -1520 440 -1503
rect -760 -2777 40 -2750
rect -760 -2833 -723 -2777
rect -667 -2833 40 -2777
rect -760 -2840 40 -2833
rect -750 -2860 -640 -2840
rect -1200 -3250 200 -3160
rect -1200 -4000 -1110 -3250
rect -480 -3450 -370 -3440
rect -560 -3463 520 -3450
rect -560 -3527 -457 -3463
rect -393 -3527 520 -3463
rect -560 -3540 520 -3527
rect -480 -3550 -370 -3540
rect -560 -4447 440 -4430
rect -560 -4503 -508 -4447
rect -452 -4503 -428 -4447
rect -372 -4503 -348 -4447
rect -292 -4503 440 -4447
rect -560 -4520 440 -4503
rect -760 -5777 40 -5750
rect -760 -5833 -723 -5777
rect -667 -5833 40 -5777
rect -760 -5840 40 -5833
rect -750 -5860 -640 -5840
rect 540 -6098 2780 -6060
rect 540 -6162 588 -6098
rect 652 -6162 668 -6098
rect 732 -6162 748 -6098
rect 812 -6162 828 -6098
rect 892 -6162 908 -6098
rect 972 -6162 988 -6098
rect 1052 -6162 1068 -6098
rect 1132 -6162 1148 -6098
rect 1212 -6162 1228 -6098
rect 1292 -6162 1308 -6098
rect 1372 -6162 1388 -6098
rect 1452 -6162 1468 -6098
rect 1532 -6162 1548 -6098
rect 1612 -6162 1628 -6098
rect 1692 -6162 1708 -6098
rect 1772 -6162 1788 -6098
rect 1852 -6162 1868 -6098
rect 1932 -6162 1948 -6098
rect 2012 -6162 2028 -6098
rect 2092 -6162 2108 -6098
rect 2172 -6162 2188 -6098
rect 2252 -6162 2268 -6098
rect 2332 -6162 2348 -6098
rect 2412 -6162 2428 -6098
rect 2492 -6162 2508 -6098
rect 2572 -6162 2588 -6098
rect 2652 -6162 2668 -6098
rect 2732 -6162 2780 -6098
rect 540 -6200 2780 -6162
rect 3540 -6098 5780 -6060
rect 3540 -6162 3588 -6098
rect 3652 -6162 3668 -6098
rect 3732 -6162 3748 -6098
rect 3812 -6162 3828 -6098
rect 3892 -6162 3908 -6098
rect 3972 -6162 3988 -6098
rect 4052 -6162 4068 -6098
rect 4132 -6162 4148 -6098
rect 4212 -6162 4228 -6098
rect 4292 -6162 4308 -6098
rect 4372 -6162 4388 -6098
rect 4452 -6162 4468 -6098
rect 4532 -6162 4548 -6098
rect 4612 -6162 4628 -6098
rect 4692 -6162 4708 -6098
rect 4772 -6162 4788 -6098
rect 4852 -6162 4868 -6098
rect 4932 -6162 4948 -6098
rect 5012 -6162 5028 -6098
rect 5092 -6162 5108 -6098
rect 5172 -6162 5188 -6098
rect 5252 -6162 5268 -6098
rect 5332 -6162 5348 -6098
rect 5412 -6162 5428 -6098
rect 5492 -6162 5508 -6098
rect 5572 -6162 5588 -6098
rect 5652 -6162 5668 -6098
rect 5732 -6162 5780 -6098
rect 3540 -6200 5780 -6162
rect 6540 -6098 8780 -6060
rect 6540 -6162 6588 -6098
rect 6652 -6162 6668 -6098
rect 6732 -6162 6748 -6098
rect 6812 -6162 6828 -6098
rect 6892 -6162 6908 -6098
rect 6972 -6162 6988 -6098
rect 7052 -6162 7068 -6098
rect 7132 -6162 7148 -6098
rect 7212 -6162 7228 -6098
rect 7292 -6162 7308 -6098
rect 7372 -6162 7388 -6098
rect 7452 -6162 7468 -6098
rect 7532 -6162 7548 -6098
rect 7612 -6162 7628 -6098
rect 7692 -6162 7708 -6098
rect 7772 -6162 7788 -6098
rect 7852 -6162 7868 -6098
rect 7932 -6162 7948 -6098
rect 8012 -6162 8028 -6098
rect 8092 -6162 8108 -6098
rect 8172 -6162 8188 -6098
rect 8252 -6162 8268 -6098
rect 8332 -6162 8348 -6098
rect 8412 -6162 8428 -6098
rect 8492 -6162 8508 -6098
rect 8572 -6162 8588 -6098
rect 8652 -6162 8668 -6098
rect 8732 -6162 8780 -6098
rect 6540 -6200 8780 -6162
rect 220 -6528 440 -6490
rect 220 -6672 258 -6528
rect 402 -6672 440 -6528
rect 220 -6710 440 -6672
rect 3220 -6528 3440 -6490
rect 3220 -6672 3258 -6528
rect 3402 -6672 3440 -6528
rect 3220 -6710 3440 -6672
rect 6220 -6528 6440 -6490
rect 6220 -6672 6258 -6528
rect 6402 -6672 6440 -6528
rect 6220 -6710 6440 -6672
<< via3 >>
rect 503 3633 567 3637
rect 503 3577 507 3633
rect 507 3577 563 3633
rect 563 3577 567 3633
rect 503 3573 567 3577
rect 3503 3633 3567 3637
rect 3503 3577 3507 3633
rect 3507 3577 3563 3633
rect 3563 3577 3567 3633
rect 3503 3573 3567 3577
rect 6503 3633 6567 3637
rect 6503 3577 6507 3633
rect 6507 3577 6563 3633
rect 6563 3577 6567 3633
rect 6503 3573 6567 3577
rect -457 2473 -393 2537
rect -457 -527 -393 -463
rect -457 -3527 -393 -3463
rect 588 -6102 652 -6098
rect 588 -6158 592 -6102
rect 592 -6158 648 -6102
rect 648 -6158 652 -6102
rect 588 -6162 652 -6158
rect 668 -6102 732 -6098
rect 668 -6158 672 -6102
rect 672 -6158 728 -6102
rect 728 -6158 732 -6102
rect 668 -6162 732 -6158
rect 748 -6102 812 -6098
rect 748 -6158 752 -6102
rect 752 -6158 808 -6102
rect 808 -6158 812 -6102
rect 748 -6162 812 -6158
rect 828 -6102 892 -6098
rect 828 -6158 832 -6102
rect 832 -6158 888 -6102
rect 888 -6158 892 -6102
rect 828 -6162 892 -6158
rect 908 -6102 972 -6098
rect 908 -6158 912 -6102
rect 912 -6158 968 -6102
rect 968 -6158 972 -6102
rect 908 -6162 972 -6158
rect 988 -6102 1052 -6098
rect 988 -6158 992 -6102
rect 992 -6158 1048 -6102
rect 1048 -6158 1052 -6102
rect 988 -6162 1052 -6158
rect 1068 -6102 1132 -6098
rect 1068 -6158 1072 -6102
rect 1072 -6158 1128 -6102
rect 1128 -6158 1132 -6102
rect 1068 -6162 1132 -6158
rect 1148 -6102 1212 -6098
rect 1148 -6158 1152 -6102
rect 1152 -6158 1208 -6102
rect 1208 -6158 1212 -6102
rect 1148 -6162 1212 -6158
rect 1228 -6102 1292 -6098
rect 1228 -6158 1232 -6102
rect 1232 -6158 1288 -6102
rect 1288 -6158 1292 -6102
rect 1228 -6162 1292 -6158
rect 1308 -6102 1372 -6098
rect 1308 -6158 1312 -6102
rect 1312 -6158 1368 -6102
rect 1368 -6158 1372 -6102
rect 1308 -6162 1372 -6158
rect 1388 -6102 1452 -6098
rect 1388 -6158 1392 -6102
rect 1392 -6158 1448 -6102
rect 1448 -6158 1452 -6102
rect 1388 -6162 1452 -6158
rect 1468 -6102 1532 -6098
rect 1468 -6158 1472 -6102
rect 1472 -6158 1528 -6102
rect 1528 -6158 1532 -6102
rect 1468 -6162 1532 -6158
rect 1548 -6102 1612 -6098
rect 1548 -6158 1552 -6102
rect 1552 -6158 1608 -6102
rect 1608 -6158 1612 -6102
rect 1548 -6162 1612 -6158
rect 1628 -6102 1692 -6098
rect 1628 -6158 1632 -6102
rect 1632 -6158 1688 -6102
rect 1688 -6158 1692 -6102
rect 1628 -6162 1692 -6158
rect 1708 -6102 1772 -6098
rect 1708 -6158 1712 -6102
rect 1712 -6158 1768 -6102
rect 1768 -6158 1772 -6102
rect 1708 -6162 1772 -6158
rect 1788 -6102 1852 -6098
rect 1788 -6158 1792 -6102
rect 1792 -6158 1848 -6102
rect 1848 -6158 1852 -6102
rect 1788 -6162 1852 -6158
rect 1868 -6102 1932 -6098
rect 1868 -6158 1872 -6102
rect 1872 -6158 1928 -6102
rect 1928 -6158 1932 -6102
rect 1868 -6162 1932 -6158
rect 1948 -6102 2012 -6098
rect 1948 -6158 1952 -6102
rect 1952 -6158 2008 -6102
rect 2008 -6158 2012 -6102
rect 1948 -6162 2012 -6158
rect 2028 -6102 2092 -6098
rect 2028 -6158 2032 -6102
rect 2032 -6158 2088 -6102
rect 2088 -6158 2092 -6102
rect 2028 -6162 2092 -6158
rect 2108 -6102 2172 -6098
rect 2108 -6158 2112 -6102
rect 2112 -6158 2168 -6102
rect 2168 -6158 2172 -6102
rect 2108 -6162 2172 -6158
rect 2188 -6102 2252 -6098
rect 2188 -6158 2192 -6102
rect 2192 -6158 2248 -6102
rect 2248 -6158 2252 -6102
rect 2188 -6162 2252 -6158
rect 2268 -6102 2332 -6098
rect 2268 -6158 2272 -6102
rect 2272 -6158 2328 -6102
rect 2328 -6158 2332 -6102
rect 2268 -6162 2332 -6158
rect 2348 -6102 2412 -6098
rect 2348 -6158 2352 -6102
rect 2352 -6158 2408 -6102
rect 2408 -6158 2412 -6102
rect 2348 -6162 2412 -6158
rect 2428 -6102 2492 -6098
rect 2428 -6158 2432 -6102
rect 2432 -6158 2488 -6102
rect 2488 -6158 2492 -6102
rect 2428 -6162 2492 -6158
rect 2508 -6102 2572 -6098
rect 2508 -6158 2512 -6102
rect 2512 -6158 2568 -6102
rect 2568 -6158 2572 -6102
rect 2508 -6162 2572 -6158
rect 2588 -6102 2652 -6098
rect 2588 -6158 2592 -6102
rect 2592 -6158 2648 -6102
rect 2648 -6158 2652 -6102
rect 2588 -6162 2652 -6158
rect 2668 -6102 2732 -6098
rect 2668 -6158 2672 -6102
rect 2672 -6158 2728 -6102
rect 2728 -6158 2732 -6102
rect 2668 -6162 2732 -6158
rect 3588 -6102 3652 -6098
rect 3588 -6158 3592 -6102
rect 3592 -6158 3648 -6102
rect 3648 -6158 3652 -6102
rect 3588 -6162 3652 -6158
rect 3668 -6102 3732 -6098
rect 3668 -6158 3672 -6102
rect 3672 -6158 3728 -6102
rect 3728 -6158 3732 -6102
rect 3668 -6162 3732 -6158
rect 3748 -6102 3812 -6098
rect 3748 -6158 3752 -6102
rect 3752 -6158 3808 -6102
rect 3808 -6158 3812 -6102
rect 3748 -6162 3812 -6158
rect 3828 -6102 3892 -6098
rect 3828 -6158 3832 -6102
rect 3832 -6158 3888 -6102
rect 3888 -6158 3892 -6102
rect 3828 -6162 3892 -6158
rect 3908 -6102 3972 -6098
rect 3908 -6158 3912 -6102
rect 3912 -6158 3968 -6102
rect 3968 -6158 3972 -6102
rect 3908 -6162 3972 -6158
rect 3988 -6102 4052 -6098
rect 3988 -6158 3992 -6102
rect 3992 -6158 4048 -6102
rect 4048 -6158 4052 -6102
rect 3988 -6162 4052 -6158
rect 4068 -6102 4132 -6098
rect 4068 -6158 4072 -6102
rect 4072 -6158 4128 -6102
rect 4128 -6158 4132 -6102
rect 4068 -6162 4132 -6158
rect 4148 -6102 4212 -6098
rect 4148 -6158 4152 -6102
rect 4152 -6158 4208 -6102
rect 4208 -6158 4212 -6102
rect 4148 -6162 4212 -6158
rect 4228 -6102 4292 -6098
rect 4228 -6158 4232 -6102
rect 4232 -6158 4288 -6102
rect 4288 -6158 4292 -6102
rect 4228 -6162 4292 -6158
rect 4308 -6102 4372 -6098
rect 4308 -6158 4312 -6102
rect 4312 -6158 4368 -6102
rect 4368 -6158 4372 -6102
rect 4308 -6162 4372 -6158
rect 4388 -6102 4452 -6098
rect 4388 -6158 4392 -6102
rect 4392 -6158 4448 -6102
rect 4448 -6158 4452 -6102
rect 4388 -6162 4452 -6158
rect 4468 -6102 4532 -6098
rect 4468 -6158 4472 -6102
rect 4472 -6158 4528 -6102
rect 4528 -6158 4532 -6102
rect 4468 -6162 4532 -6158
rect 4548 -6102 4612 -6098
rect 4548 -6158 4552 -6102
rect 4552 -6158 4608 -6102
rect 4608 -6158 4612 -6102
rect 4548 -6162 4612 -6158
rect 4628 -6102 4692 -6098
rect 4628 -6158 4632 -6102
rect 4632 -6158 4688 -6102
rect 4688 -6158 4692 -6102
rect 4628 -6162 4692 -6158
rect 4708 -6102 4772 -6098
rect 4708 -6158 4712 -6102
rect 4712 -6158 4768 -6102
rect 4768 -6158 4772 -6102
rect 4708 -6162 4772 -6158
rect 4788 -6102 4852 -6098
rect 4788 -6158 4792 -6102
rect 4792 -6158 4848 -6102
rect 4848 -6158 4852 -6102
rect 4788 -6162 4852 -6158
rect 4868 -6102 4932 -6098
rect 4868 -6158 4872 -6102
rect 4872 -6158 4928 -6102
rect 4928 -6158 4932 -6102
rect 4868 -6162 4932 -6158
rect 4948 -6102 5012 -6098
rect 4948 -6158 4952 -6102
rect 4952 -6158 5008 -6102
rect 5008 -6158 5012 -6102
rect 4948 -6162 5012 -6158
rect 5028 -6102 5092 -6098
rect 5028 -6158 5032 -6102
rect 5032 -6158 5088 -6102
rect 5088 -6158 5092 -6102
rect 5028 -6162 5092 -6158
rect 5108 -6102 5172 -6098
rect 5108 -6158 5112 -6102
rect 5112 -6158 5168 -6102
rect 5168 -6158 5172 -6102
rect 5108 -6162 5172 -6158
rect 5188 -6102 5252 -6098
rect 5188 -6158 5192 -6102
rect 5192 -6158 5248 -6102
rect 5248 -6158 5252 -6102
rect 5188 -6162 5252 -6158
rect 5268 -6102 5332 -6098
rect 5268 -6158 5272 -6102
rect 5272 -6158 5328 -6102
rect 5328 -6158 5332 -6102
rect 5268 -6162 5332 -6158
rect 5348 -6102 5412 -6098
rect 5348 -6158 5352 -6102
rect 5352 -6158 5408 -6102
rect 5408 -6158 5412 -6102
rect 5348 -6162 5412 -6158
rect 5428 -6102 5492 -6098
rect 5428 -6158 5432 -6102
rect 5432 -6158 5488 -6102
rect 5488 -6158 5492 -6102
rect 5428 -6162 5492 -6158
rect 5508 -6102 5572 -6098
rect 5508 -6158 5512 -6102
rect 5512 -6158 5568 -6102
rect 5568 -6158 5572 -6102
rect 5508 -6162 5572 -6158
rect 5588 -6102 5652 -6098
rect 5588 -6158 5592 -6102
rect 5592 -6158 5648 -6102
rect 5648 -6158 5652 -6102
rect 5588 -6162 5652 -6158
rect 5668 -6102 5732 -6098
rect 5668 -6158 5672 -6102
rect 5672 -6158 5728 -6102
rect 5728 -6158 5732 -6102
rect 5668 -6162 5732 -6158
rect 6588 -6102 6652 -6098
rect 6588 -6158 6592 -6102
rect 6592 -6158 6648 -6102
rect 6648 -6158 6652 -6102
rect 6588 -6162 6652 -6158
rect 6668 -6102 6732 -6098
rect 6668 -6158 6672 -6102
rect 6672 -6158 6728 -6102
rect 6728 -6158 6732 -6102
rect 6668 -6162 6732 -6158
rect 6748 -6102 6812 -6098
rect 6748 -6158 6752 -6102
rect 6752 -6158 6808 -6102
rect 6808 -6158 6812 -6102
rect 6748 -6162 6812 -6158
rect 6828 -6102 6892 -6098
rect 6828 -6158 6832 -6102
rect 6832 -6158 6888 -6102
rect 6888 -6158 6892 -6102
rect 6828 -6162 6892 -6158
rect 6908 -6102 6972 -6098
rect 6908 -6158 6912 -6102
rect 6912 -6158 6968 -6102
rect 6968 -6158 6972 -6102
rect 6908 -6162 6972 -6158
rect 6988 -6102 7052 -6098
rect 6988 -6158 6992 -6102
rect 6992 -6158 7048 -6102
rect 7048 -6158 7052 -6102
rect 6988 -6162 7052 -6158
rect 7068 -6102 7132 -6098
rect 7068 -6158 7072 -6102
rect 7072 -6158 7128 -6102
rect 7128 -6158 7132 -6102
rect 7068 -6162 7132 -6158
rect 7148 -6102 7212 -6098
rect 7148 -6158 7152 -6102
rect 7152 -6158 7208 -6102
rect 7208 -6158 7212 -6102
rect 7148 -6162 7212 -6158
rect 7228 -6102 7292 -6098
rect 7228 -6158 7232 -6102
rect 7232 -6158 7288 -6102
rect 7288 -6158 7292 -6102
rect 7228 -6162 7292 -6158
rect 7308 -6102 7372 -6098
rect 7308 -6158 7312 -6102
rect 7312 -6158 7368 -6102
rect 7368 -6158 7372 -6102
rect 7308 -6162 7372 -6158
rect 7388 -6102 7452 -6098
rect 7388 -6158 7392 -6102
rect 7392 -6158 7448 -6102
rect 7448 -6158 7452 -6102
rect 7388 -6162 7452 -6158
rect 7468 -6102 7532 -6098
rect 7468 -6158 7472 -6102
rect 7472 -6158 7528 -6102
rect 7528 -6158 7532 -6102
rect 7468 -6162 7532 -6158
rect 7548 -6102 7612 -6098
rect 7548 -6158 7552 -6102
rect 7552 -6158 7608 -6102
rect 7608 -6158 7612 -6102
rect 7548 -6162 7612 -6158
rect 7628 -6102 7692 -6098
rect 7628 -6158 7632 -6102
rect 7632 -6158 7688 -6102
rect 7688 -6158 7692 -6102
rect 7628 -6162 7692 -6158
rect 7708 -6102 7772 -6098
rect 7708 -6158 7712 -6102
rect 7712 -6158 7768 -6102
rect 7768 -6158 7772 -6102
rect 7708 -6162 7772 -6158
rect 7788 -6102 7852 -6098
rect 7788 -6158 7792 -6102
rect 7792 -6158 7848 -6102
rect 7848 -6158 7852 -6102
rect 7788 -6162 7852 -6158
rect 7868 -6102 7932 -6098
rect 7868 -6158 7872 -6102
rect 7872 -6158 7928 -6102
rect 7928 -6158 7932 -6102
rect 7868 -6162 7932 -6158
rect 7948 -6102 8012 -6098
rect 7948 -6158 7952 -6102
rect 7952 -6158 8008 -6102
rect 8008 -6158 8012 -6102
rect 7948 -6162 8012 -6158
rect 8028 -6102 8092 -6098
rect 8028 -6158 8032 -6102
rect 8032 -6158 8088 -6102
rect 8088 -6158 8092 -6102
rect 8028 -6162 8092 -6158
rect 8108 -6102 8172 -6098
rect 8108 -6158 8112 -6102
rect 8112 -6158 8168 -6102
rect 8168 -6158 8172 -6102
rect 8108 -6162 8172 -6158
rect 8188 -6102 8252 -6098
rect 8188 -6158 8192 -6102
rect 8192 -6158 8248 -6102
rect 8248 -6158 8252 -6102
rect 8188 -6162 8252 -6158
rect 8268 -6102 8332 -6098
rect 8268 -6158 8272 -6102
rect 8272 -6158 8328 -6102
rect 8328 -6158 8332 -6102
rect 8268 -6162 8332 -6158
rect 8348 -6102 8412 -6098
rect 8348 -6158 8352 -6102
rect 8352 -6158 8408 -6102
rect 8408 -6158 8412 -6102
rect 8348 -6162 8412 -6158
rect 8428 -6102 8492 -6098
rect 8428 -6158 8432 -6102
rect 8432 -6158 8488 -6102
rect 8488 -6158 8492 -6102
rect 8428 -6162 8492 -6158
rect 8508 -6102 8572 -6098
rect 8508 -6158 8512 -6102
rect 8512 -6158 8568 -6102
rect 8568 -6158 8572 -6102
rect 8508 -6162 8572 -6158
rect 8588 -6102 8652 -6098
rect 8588 -6158 8592 -6102
rect 8592 -6158 8648 -6102
rect 8648 -6158 8652 -6102
rect 8588 -6162 8652 -6158
rect 8668 -6102 8732 -6098
rect 8668 -6158 8672 -6102
rect 8672 -6158 8728 -6102
rect 8728 -6158 8732 -6102
rect 8668 -6162 8732 -6158
rect 258 -6532 402 -6528
rect 258 -6668 262 -6532
rect 262 -6668 398 -6532
rect 398 -6668 402 -6532
rect 258 -6672 402 -6668
rect 3258 -6532 3402 -6528
rect 3258 -6668 3262 -6532
rect 3262 -6668 3398 -6532
rect 3398 -6668 3402 -6532
rect 3258 -6672 3402 -6668
rect 6258 -6532 6402 -6528
rect 6258 -6668 6262 -6532
rect 6262 -6668 6398 -6532
rect 6398 -6668 6402 -6532
rect 6258 -6672 6402 -6668
<< metal4 >>
rect -3000 3637 8200 3660
rect -3000 3573 503 3637
rect 567 3573 3503 3637
rect 3567 3573 6503 3637
rect 6567 3573 8200 3637
rect -3000 3550 8200 3573
rect -480 2537 -370 2600
rect -480 2473 -457 2537
rect -393 2473 -370 2537
rect -480 -463 -370 2473
rect -480 -527 -457 -463
rect -393 -527 -370 -463
rect -480 -3463 -370 -527
rect -480 -3527 -457 -3463
rect -393 -3527 -370 -3463
rect -480 -7600 -370 -3527
rect 2630 -6060 2780 -6000
rect 5630 -6060 5780 -6000
rect 8630 -6060 8780 -6000
rect 540 -6098 2780 -6060
rect 540 -6162 588 -6098
rect 652 -6162 668 -6098
rect 732 -6162 748 -6098
rect 812 -6162 828 -6098
rect 892 -6162 908 -6098
rect 972 -6162 988 -6098
rect 1052 -6162 1068 -6098
rect 1132 -6162 1148 -6098
rect 1212 -6162 1228 -6098
rect 1292 -6162 1308 -6098
rect 1372 -6162 1388 -6098
rect 1452 -6162 1468 -6098
rect 1532 -6162 1548 -6098
rect 1612 -6162 1628 -6098
rect 1692 -6162 1708 -6098
rect 1772 -6162 1788 -6098
rect 1852 -6162 1868 -6098
rect 1932 -6162 1948 -6098
rect 2012 -6162 2028 -6098
rect 2092 -6162 2108 -6098
rect 2172 -6162 2188 -6098
rect 2252 -6162 2268 -6098
rect 2332 -6162 2348 -6098
rect 2412 -6162 2428 -6098
rect 2492 -6162 2508 -6098
rect 2572 -6162 2588 -6098
rect 2652 -6162 2668 -6098
rect 2732 -6162 2780 -6098
rect 540 -6200 2780 -6162
rect 3540 -6098 5780 -6060
rect 3540 -6162 3588 -6098
rect 3652 -6162 3668 -6098
rect 3732 -6162 3748 -6098
rect 3812 -6162 3828 -6098
rect 3892 -6162 3908 -6098
rect 3972 -6162 3988 -6098
rect 4052 -6162 4068 -6098
rect 4132 -6162 4148 -6098
rect 4212 -6162 4228 -6098
rect 4292 -6162 4308 -6098
rect 4372 -6162 4388 -6098
rect 4452 -6162 4468 -6098
rect 4532 -6162 4548 -6098
rect 4612 -6162 4628 -6098
rect 4692 -6162 4708 -6098
rect 4772 -6162 4788 -6098
rect 4852 -6162 4868 -6098
rect 4932 -6162 4948 -6098
rect 5012 -6162 5028 -6098
rect 5092 -6162 5108 -6098
rect 5172 -6162 5188 -6098
rect 5252 -6162 5268 -6098
rect 5332 -6162 5348 -6098
rect 5412 -6162 5428 -6098
rect 5492 -6162 5508 -6098
rect 5572 -6162 5588 -6098
rect 5652 -6162 5668 -6098
rect 5732 -6162 5780 -6098
rect 3540 -6200 5780 -6162
rect 6540 -6098 8780 -6060
rect 6540 -6162 6588 -6098
rect 6652 -6162 6668 -6098
rect 6732 -6162 6748 -6098
rect 6812 -6162 6828 -6098
rect 6892 -6162 6908 -6098
rect 6972 -6162 6988 -6098
rect 7052 -6162 7068 -6098
rect 7132 -6162 7148 -6098
rect 7212 -6162 7228 -6098
rect 7292 -6162 7308 -6098
rect 7372 -6162 7388 -6098
rect 7452 -6162 7468 -6098
rect 7532 -6162 7548 -6098
rect 7612 -6162 7628 -6098
rect 7692 -6162 7708 -6098
rect 7772 -6162 7788 -6098
rect 7852 -6162 7868 -6098
rect 7932 -6162 7948 -6098
rect 8012 -6162 8028 -6098
rect 8092 -6162 8108 -6098
rect 8172 -6162 8188 -6098
rect 8252 -6162 8268 -6098
rect 8332 -6162 8348 -6098
rect 8412 -6162 8428 -6098
rect 8492 -6162 8508 -6098
rect 8572 -6162 8588 -6098
rect 8652 -6162 8668 -6098
rect 8732 -6162 8780 -6098
rect 6540 -6200 8780 -6162
rect 220 -6528 440 -6490
rect 220 -6672 258 -6528
rect 402 -6672 440 -6528
rect 220 -7100 440 -6672
rect 3220 -6528 3440 -6490
rect 3220 -6672 3258 -6528
rect 3402 -6672 3440 -6528
rect 3220 -7100 3440 -6672
rect 6220 -6528 6440 -6490
rect 6220 -6672 6258 -6528
rect 6402 -6672 6440 -6528
rect 6220 -7100 6440 -6672
<< metal5 >>
rect -2000 2840 0 3160
rect 1040 1040 1240 1240
rect 4040 1040 4240 1240
rect 7040 1040 7240 1240
rect 1040 -1960 1240 -1760
rect 4040 -1960 4240 -1760
rect 7040 -1960 7240 -1760
rect 1040 -4960 1240 -4760
rect 4040 -4960 4240 -4760
rect 7040 -4960 7240 -4760
use pixel  pixel_0
timestamp 1654643737
transform 1 0 -800 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_1
timestamp 1654643737
transform 1 0 -3800 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_2
timestamp 1654643737
transform 1 0 -800 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_3
timestamp 1654643737
transform 1 0 -3800 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_4
timestamp 1654643737
transform 1 0 2200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_5
timestamp 1654643737
transform 1 0 2200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_6
timestamp 1654643737
transform 1 0 -800 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_7
timestamp 1654643737
transform 1 0 -3800 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_8
timestamp 1654643737
transform 1 0 2200 0 1 2700
box 3640 -2860 6960 460
<< labels >>
rlabel metal2 s 3500 3000 3570 3600 4 VBIAS
port 1 nsew
rlabel metal2 s 3060 3000 3130 3600 4 VREF
port 2 nsew
rlabel metal2 s 4020 3000 4090 3600 4 NB2
port 3 nsew
rlabel metal2 s 6500 3000 6570 3600 4 VBIAS
port 1 nsew
rlabel metal2 s 6060 3000 6130 3600 4 VREF
port 2 nsew
rlabel metal2 s 7020 3000 7090 3600 4 NB2
port 3 nsew
rlabel metal1 s -560 -120 40 -30 4 VDD
port 4 nsew
rlabel metal3 s -560 -250 40 -160 4 SF_IB
port 5 nsew
rlabel metal3 s -560 -540 40 -450 4 CSA_VREF
port 6 nsew
rlabel metal3 s -560 -2840 40 -2750 4 NB1
port 7 nsew
rlabel metal1 s 9000 -2970 9600 -2880 4 GND
port 8 nsew
rlabel metal1 s -560 -3120 40 -3030 4 VDD
port 4 nsew
rlabel metal3 s -560 -3250 40 -3160 4 SF_IB
port 5 nsew
rlabel metal3 s -560 -3540 40 -3450 4 CSA_VREF
port 6 nsew
rlabel metal3 s -560 -5840 40 -5750 4 NB1
port 7 nsew
rlabel metal1 s 9000 -5970 9600 -5880 4 GND
port 8 nsew
rlabel metal2 s 500 3000 570 3600 4 VBIAS
port 1 nsew
rlabel metal4 s -1000 3550 -1000 3550 4 VBIAS
port 1 nsew
rlabel metal4 s -3000 3605 -3000 3605 4 VBIAS
port 1 nsew
rlabel metal2 s 60 3000 130 3600 4 VREF
port 2 nsew
rlabel metal1 s -1000 3350 -1000 3350 4 VREF
port 2 nsew
rlabel metal2 s -3000 3400 -3000 3400 4 VREF
port 2 nsew
rlabel metal2 s 1020 3000 1090 3600 4 NB2
port 3 nsew
rlabel metal2 s 0 4040 0 4040 4 NB2
port 3 nsew
rlabel metal1 s -560 2880 40 2970 4 VDD
port 4 nsew
rlabel metal1 s -2000 0 -2000 0 4 VDD
port 4 nsew
rlabel metal3 s -560 2750 40 2840 4 SF_IB
port 5 nsew
rlabel metal3 s -560 2460 40 2550 4 CSA_VREF
port 6 nsew
rlabel metal4 s -480 -7600 -480 -7600 4 CSA_VREF
port 6 nsew
rlabel metal3 s -560 160 40 250 4 NB1
port 7 nsew
rlabel metal2 s -740 3560 -740 3560 4 NB1
port 7 nsew
rlabel metal3 s -560 1480 40 1570 4 ROW_SEL0
port 9 nsew
rlabel metal2 s -3000 1480 -3000 1480 4 ROW_SEL0
port 9 nsew
rlabel metal2 s -3000 1525 -3000 1525 4 ROW_SEL0
port 9 nsew
rlabel metal1 s 9000 30 9600 120 4 GND
port 8 nsew
rlabel metal1 s 9400 30 9400 30 4 GND
port 8 nsew
rlabel metal3 s -560 -1520 40 -1430 4 ROW_SEL1
port 10 nsew
rlabel metal2 s -3000 -1520 -3000 -1520 4 ROW_SEL1
port 10 nsew
rlabel metal2 s -3000 -1475 -3000 -1475 4 ROW_SEL1
port 10 nsew
rlabel metal3 s -560 -4520 40 -4430 4 ROW_SEL2
port 11 nsew
rlabel metal2 s -3000 -4520 -3000 -4520 4 ROW_SEL2
port 11 nsew
rlabel metal2 s -3000 -4475 -3000 -4475 4 ROW_SEL2
port 11 nsew
rlabel metal5 s 1040 1040 1240 1240 4 PIX0_IN
port 12 nsew
rlabel metal5 s -2000 2840 -2000 2840 4 GRING
port 13 nsew
rlabel metal5 s 4040 1040 4240 1240 4 PIX1_IN
port 14 nsew
rlabel metal5 s 7040 1040 7240 1240 4 PIX2_IN
port 15 nsew
rlabel metal5 s 1040 -1960 1240 -1760 4 PIX3_IN
port 16 nsew
rlabel metal5 s 4040 -1960 4240 -1760 4 PIX4_IN
port 17 nsew
rlabel metal5 s 7040 -1960 7240 -1760 4 PIX5_IN
port 18 nsew
rlabel metal5 s 1040 -4960 1240 -4760 4 PIX6_IN
port 19 nsew
rlabel metal4 s 2630 -6200 2780 -6000 4 PIX_OUT0
port 20 nsew
rlabel metal4 s 220 -7100 440 -6700 4 COL_SEL0
port 21 nsew
rlabel metal5 s 4040 -4960 4240 -4760 4 PIX7_IN
port 22 nsew
rlabel metal4 s 5630 -6200 5780 -6000 4 PIX_OUT1
port 23 nsew
rlabel metal4 s 3220 -7100 3440 -6700 4 COL_SEL1
port 24 nsew
rlabel metal5 s 7040 -4960 7240 -4760 4 PIX8_IN
port 25 nsew
rlabel metal4 s 8630 -6200 8780 -6000 4 PIX_OUT2
port 26 nsew
rlabel metal2 s 8940 -7100 8940 -7100 4 ARRAY_OUT
port 27 nsew
rlabel metal4 s 6220 -7100 6440 -6700 4 COL_SEL2
port 28 nsew
<< end >>
