magic
tech sky130A
magscale 1 2
timestamp 1654639008
<< nwell >>
rect 1010 -1030 1930 -510
<< pmoslvt >>
rect 1280 -960 1480 -760
<< nmoslvt >>
rect 2360 -1410 2560 -1170
rect 2870 -1410 3070 -1170
rect 3230 -1330 4830 -930
rect 5230 -1330 6830 -930
<< ndiff >>
rect 3230 -810 4830 -790
rect 3230 -910 3250 -810
rect 4810 -910 4830 -810
rect 3230 -930 4830 -910
rect 5230 -810 6830 -790
rect 5230 -910 5250 -810
rect 6810 -910 6830 -810
rect 5230 -930 6830 -910
rect 2360 -1110 2560 -1100
rect 2360 -1150 2380 -1110
rect 2540 -1150 2560 -1110
rect 2360 -1170 2560 -1150
rect 2870 -1110 3070 -1100
rect 2870 -1150 2890 -1110
rect 3050 -1150 3070 -1110
rect 2870 -1170 3070 -1150
rect 3230 -1350 4830 -1330
rect 2360 -1430 2560 -1410
rect 2360 -1470 2380 -1430
rect 2540 -1470 2560 -1430
rect 2360 -1480 2560 -1470
rect 2870 -1430 3070 -1410
rect 2870 -1470 2890 -1430
rect 3050 -1470 3070 -1430
rect 3230 -1450 3250 -1350
rect 4810 -1450 4830 -1350
rect 3230 -1460 4830 -1450
rect 5230 -1350 6830 -1330
rect 5230 -1450 5250 -1350
rect 6810 -1450 6830 -1350
rect 5230 -1460 6830 -1450
rect 2870 -1480 3070 -1470
<< pdiff >>
rect 1190 -780 1280 -760
rect 1190 -940 1200 -780
rect 1260 -940 1280 -780
rect 1190 -960 1280 -940
rect 1480 -780 1590 -760
rect 1480 -940 1500 -780
rect 1560 -940 1590 -780
rect 1480 -960 1590 -940
<< ndiffc >>
rect 3250 -910 4810 -810
rect 5250 -910 6810 -810
rect 2380 -1150 2540 -1110
rect 2890 -1150 3050 -1110
rect 2380 -1470 2540 -1430
rect 2890 -1470 3050 -1430
rect 3250 -1450 4810 -1350
rect 5250 -1450 6810 -1350
<< pdiffc >>
rect 1200 -940 1260 -780
rect 1500 -940 1560 -780
<< psubdiff >>
rect 5230 -1490 6830 -1460
rect 5230 -1580 5260 -1490
rect 6800 -1580 6830 -1490
rect 5230 -1600 6830 -1580
<< nsubdiff >>
rect 1090 -790 1190 -760
rect 1090 -930 1110 -790
rect 1160 -930 1190 -790
rect 1090 -960 1190 -930
<< psubdiffcont >>
rect 5260 -1580 6800 -1490
<< nsubdiffcont >>
rect 1110 -930 1160 -790
<< poly >>
rect 1280 -760 1480 -730
rect 1280 -990 1480 -960
rect 1280 -1050 1360 -990
rect 1280 -1110 1290 -1050
rect 1350 -1110 1360 -1050
rect 1280 -1130 1360 -1110
rect 2330 -1330 2360 -1170
rect 2230 -1340 2360 -1330
rect 2230 -1400 2250 -1340
rect 2310 -1400 2360 -1340
rect 2230 -1410 2360 -1400
rect 2560 -1410 2590 -1170
rect 2840 -1330 2870 -1170
rect 2740 -1340 2870 -1330
rect 2740 -1400 2760 -1340
rect 2820 -1400 2870 -1340
rect 2740 -1410 2870 -1400
rect 3070 -1410 3100 -1170
rect 3200 -1330 3230 -930
rect 4830 -1180 4860 -930
rect 4830 -1200 5020 -1180
rect 4830 -1310 4890 -1200
rect 5000 -1310 5020 -1200
rect 4830 -1330 5020 -1310
rect 5200 -1330 5230 -930
rect 6830 -1180 6860 -930
rect 6830 -1200 7020 -1180
rect 6830 -1310 6890 -1200
rect 7000 -1310 7020 -1200
rect 6830 -1330 7020 -1310
<< polycont >>
rect 1290 -1110 1350 -1050
rect 2250 -1400 2310 -1340
rect 2760 -1400 2820 -1340
rect 4890 -1310 5000 -1200
rect 6890 -1310 7000 -1200
<< locali >>
rect 1090 -610 1190 -600
rect 1090 -770 1190 -740
rect 1090 -780 1280 -770
rect 1090 -790 1200 -780
rect 1090 -930 1110 -790
rect 1160 -930 1200 -790
rect 1090 -940 1200 -930
rect 1260 -940 1280 -780
rect 1090 -950 1280 -940
rect 1480 -780 1580 -770
rect 1480 -940 1500 -780
rect 1560 -940 1580 -780
rect 3230 -810 5150 -790
rect 3230 -910 3250 -810
rect 4810 -910 5150 -810
rect 5230 -810 7150 -790
rect 5230 -910 5250 -810
rect 6810 -910 7150 -810
rect 1480 -950 1580 -940
rect 1500 -1040 1580 -950
rect 1090 -1050 1580 -1040
rect 1090 -1120 1110 -1050
rect 1200 -1110 1290 -1050
rect 1350 -1110 1470 -1050
rect 1200 -1120 1470 -1110
rect 1090 -1130 1580 -1120
rect 2250 -1150 2380 -1090
rect 2540 -1150 2560 -1090
rect 2760 -1150 2890 -1090
rect 3050 -1150 3070 -1090
rect 2250 -1330 2310 -1150
rect 2760 -1330 2820 -1150
rect 5040 -1200 5150 -910
rect 7040 -1200 7150 -910
rect 4860 -1310 4890 -1200
rect 5000 -1210 5150 -1200
rect 5120 -1300 5150 -1210
rect 5000 -1310 5150 -1300
rect 6860 -1310 6890 -1200
rect 7000 -1210 7150 -1200
rect 7120 -1300 7150 -1210
rect 7000 -1310 7150 -1300
rect 2180 -1340 2310 -1330
rect 2220 -1400 2250 -1340
rect 2180 -1410 2310 -1400
rect 2600 -1340 2820 -1330
rect 2600 -1400 2620 -1340
rect 2730 -1400 2760 -1340
rect 2600 -1410 2820 -1400
rect 3230 -1350 4820 -1330
rect 2250 -1420 2310 -1410
rect 2360 -1430 2560 -1410
rect 2760 -1420 2820 -1410
rect 2360 -1470 2380 -1430
rect 2540 -1470 2560 -1430
rect 2360 -1550 2560 -1470
rect 2360 -1680 2370 -1550
rect 2550 -1680 2560 -1550
rect 2360 -1690 2560 -1680
rect 2870 -1430 3070 -1410
rect 2870 -1470 2890 -1430
rect 3050 -1470 3070 -1430
rect 2870 -1550 3070 -1470
rect 2870 -1680 2880 -1550
rect 3060 -1680 3070 -1550
rect 2870 -1690 3070 -1680
rect 3230 -1450 3250 -1350
rect 4810 -1450 4820 -1350
rect 3230 -1460 4820 -1450
rect 5230 -1350 6820 -1330
rect 5230 -1450 5250 -1350
rect 6810 -1450 6820 -1350
rect 3230 -1550 4830 -1460
rect 3230 -1920 3250 -1550
rect 4810 -1920 4830 -1550
rect 3230 -1940 4830 -1920
rect 5230 -1476 6820 -1450
rect 5230 -1490 6830 -1476
rect 5230 -1540 5260 -1490
rect 6800 -1540 6830 -1490
rect 5230 -1930 5250 -1540
rect 6810 -1930 6830 -1540
rect 5230 -1950 6830 -1930
<< viali >>
rect 1090 -740 1190 -610
rect 3250 -900 4810 -810
rect 5250 -900 6810 -810
rect 1110 -1120 1200 -1050
rect 1470 -1120 1580 -1050
rect 2380 -1110 2540 -1090
rect 2380 -1130 2540 -1110
rect 2890 -1110 3050 -1090
rect 2890 -1140 3050 -1110
rect 4890 -1300 5000 -1210
rect 5000 -1300 5120 -1210
rect 6890 -1300 7000 -1210
rect 7000 -1300 7120 -1210
rect 2110 -1400 2220 -1340
rect 2620 -1400 2730 -1340
rect 2370 -1680 2550 -1550
rect 2880 -1680 3060 -1550
rect 3250 -1920 4810 -1550
rect 5250 -1580 5260 -1540
rect 5260 -1580 6800 -1540
rect 6800 -1580 6810 -1540
rect 5250 -1930 6810 -1580
<< metal1 >>
rect 860 -610 1930 -220
rect 860 -740 1090 -610
rect 1190 -740 1930 -610
rect 860 -750 1930 -740
rect 2360 -680 2560 -674
rect 820 -1050 1220 -1040
rect 820 -1120 840 -1050
rect 1200 -1120 1220 -1050
rect 820 -1130 1220 -1120
rect 1450 -1050 1930 -1040
rect 1450 -1120 1460 -1050
rect 1910 -1120 1930 -1050
rect 1450 -1130 1930 -1120
rect 2360 -1090 2560 -880
rect 2360 -1130 2380 -1090
rect 2540 -1130 2560 -1090
rect 2360 -1150 2560 -1130
rect 2870 -680 3070 -674
rect 2870 -1090 3070 -880
rect 3230 -800 4830 -790
rect 3230 -900 3250 -800
rect 4810 -900 4830 -800
rect 3230 -910 4830 -900
rect 5230 -800 6830 -790
rect 5230 -900 5250 -800
rect 6810 -900 6830 -800
rect 5230 -910 6830 -900
rect 2870 -1140 2890 -1090
rect 3050 -1140 3070 -1090
rect 2870 -1150 3070 -1140
rect 4860 -1210 5150 -1200
rect 4860 -1300 4890 -1210
rect 5130 -1300 5150 -1210
rect 4860 -1310 5150 -1300
rect 6860 -1210 7150 -1200
rect 6860 -1300 6890 -1210
rect 7130 -1300 7150 -1210
rect 6860 -1310 7150 -1300
rect 2090 -1340 2310 -1330
rect 2090 -1400 2100 -1340
rect 2280 -1400 2310 -1340
rect 2090 -1410 2310 -1400
rect 2600 -1340 2820 -1330
rect 2600 -1400 2610 -1340
rect 2790 -1400 2820 -1340
rect 2600 -1410 2820 -1400
rect 1530 -1540 7180 -1530
rect 1530 -1550 5250 -1540
rect 1530 -1680 2370 -1550
rect 2550 -1680 2880 -1550
rect 3060 -1680 3250 -1550
rect 1530 -1920 3250 -1680
rect 4810 -1920 5250 -1550
rect 1530 -1930 5250 -1920
rect 6810 -1930 7180 -1540
rect 1530 -2170 7180 -1930
<< via1 >>
rect 2360 -880 2560 -680
rect 840 -1120 1110 -1050
rect 1110 -1120 1200 -1050
rect 1460 -1120 1470 -1050
rect 1470 -1120 1580 -1050
rect 1580 -1120 1910 -1050
rect 2870 -880 3070 -680
rect 3250 -810 4810 -800
rect 3250 -900 4810 -810
rect 5250 -810 6810 -800
rect 5250 -900 6810 -810
rect 4890 -1300 5120 -1210
rect 5120 -1300 5130 -1210
rect 6890 -1300 7120 -1210
rect 7120 -1300 7130 -1210
rect 2100 -1400 2110 -1340
rect 2110 -1400 2220 -1340
rect 2220 -1400 2280 -1340
rect 2610 -1400 2620 -1340
rect 2620 -1400 2730 -1340
rect 2730 -1400 2790 -1340
<< metal2 >>
rect 2350 -680 2570 -670
rect 2350 -880 2360 -680
rect 2560 -880 2570 -680
rect 2350 -890 2570 -880
rect 2860 -680 3080 -670
rect 2860 -880 2870 -680
rect 3070 -880 3080 -680
rect 2860 -890 3080 -880
rect 3230 -800 4830 -790
rect 3230 -900 3250 -800
rect 4810 -900 4830 -800
rect 3230 -910 4830 -900
rect 5230 -800 6830 -790
rect 5230 -900 5250 -800
rect 6810 -900 6830 -800
rect 5230 -910 6830 -900
rect 790 -1050 1220 -1040
rect 790 -1120 840 -1050
rect 1200 -1120 1220 -1050
rect 790 -1130 1220 -1120
rect 1450 -1050 1930 -1040
rect 1450 -1120 1460 -1050
rect 1910 -1120 1930 -1050
rect 1450 -1130 1930 -1120
rect 4860 -1210 5150 -1200
rect 4860 -1300 4890 -1210
rect 5130 -1300 5150 -1210
rect 4860 -1310 5150 -1300
rect 6860 -1210 7150 -1200
rect 6860 -1300 6890 -1210
rect 7130 -1300 7150 -1210
rect 6860 -1310 7150 -1300
rect 2090 -1340 2310 -1330
rect 2090 -1400 2100 -1340
rect 2280 -1400 2310 -1340
rect 2090 -1410 2310 -1400
rect 2600 -1340 2820 -1330
rect 2600 -1400 2610 -1340
rect 2790 -1400 2820 -1340
rect 2600 -1410 2820 -1400
rect 2090 -2235 2180 -1410
rect 2600 -2225 2690 -1410
rect 5040 -2205 5150 -1310
rect 7040 -2205 7150 -1310
<< via2 >>
rect 2360 -880 2560 -680
rect 2870 -880 3070 -680
rect 3250 -900 4810 -800
rect 5250 -900 6810 -800
rect 1470 -1120 1910 -1050
<< metal3 >>
rect 2360 -670 2560 -370
rect 2870 -670 3070 -370
rect 2350 -680 2570 -670
rect 2350 -880 2360 -680
rect 2560 -880 2570 -680
rect 2350 -890 2570 -880
rect 2860 -680 3080 -670
rect 2860 -880 2870 -680
rect 3070 -880 3080 -680
rect 2860 -890 3080 -880
rect 3230 -800 4830 -680
rect 3230 -900 3250 -800
rect 4810 -900 4830 -800
rect 3230 -910 4830 -900
rect 5230 -800 6830 -680
rect 5230 -900 5250 -800
rect 6810 -900 6830 -800
rect 5230 -910 6830 -900
rect 1450 -1050 1930 -1040
rect 1450 -1120 1470 -1050
rect 1910 -1120 1930 -1050
rect 1450 -1130 1930 -1120
rect 1840 -2236 1930 -1130
<< labels >>
rlabel metal1 870 -670 870 -670 1 VDD
port 1 n
rlabel metal2 2130 -1630 2130 -1630 1 NB1
port 4 n
rlabel metal2 2640 -1630 2640 -1630 1 NB2
port 5 n
rlabel metal2 5090 -1630 5090 -1630 1 OUT_IB
port 6 n
rlabel metal2 7100 -1630 7100 -1630 1 AMP_IB
port 7 n
rlabel metal1 1650 -1540 1650 -1540 1 GND
port 12 n
rlabel metal3 1840 -2236 1930 -2200 1 SF_IB
port 13 n
<< end >>
