* NGSPICE file created from opampjulia.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_VXTF3X VSUBS a_n385_n600# a_1039_n600# a_1097_n697#
+ a_n1631_n600# a_n919_n600# a_n1751_n697# a_683_n600# a_741_n697# a_1217_n600# a_n683_n697#
+ a_n563_n600# a_n1039_n697# a_29_n697# a_1275_n697# a_861_n600# a_n741_n600# a_n861_n697#
+ a_1453_n697# a_1395_n600# a_n1217_n697# a_207_n697# a_n1097_n600# a_149_n600# a_n29_n600#
+ a_n149_n697# a_1631_n697# a_1573_n600# w_n1947_n819# a_n1275_n600# a_327_n600# a_n1395_n697#
+ a_385_n697# a_n327_n697# a_n1809_n600# a_n207_n600# a_919_n697# a_1751_n600# a_n1573_n697#
+ a_n1453_n600# a_505_n600# a_563_n697# a_n505_n697#
X0 a_505_n600# a_385_n697# a_327_n600# w_n1947_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X1 a_149_n600# a_29_n697# a_n29_n600# w_n1947_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X2 a_1751_n600# a_1631_n697# a_1573_n600# w_n1947_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X3 a_1573_n600# a_1453_n697# a_1395_n600# w_n1947_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X4 a_1395_n600# a_1275_n697# a_1217_n600# w_n1947_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X5 a_1217_n600# a_1097_n697# a_1039_n600# w_n1947_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X6 a_n1097_n600# a_n1217_n697# a_n1275_n600# w_n1947_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X7 a_1039_n600# a_919_n697# a_861_n600# w_n1947_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X8 a_n919_n600# a_n1039_n697# a_n1097_n600# w_n1947_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X9 a_n385_n600# a_n505_n697# a_n563_n600# w_n1947_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X10 a_n1631_n600# a_n1751_n697# a_n1809_n600# w_n1947_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X11 a_n207_n600# a_n327_n697# a_n385_n600# w_n1947_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X12 a_n1453_n600# a_n1573_n697# a_n1631_n600# w_n1947_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X13 a_n1275_n600# a_n1395_n697# a_n1453_n600# w_n1947_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X14 a_n29_n600# a_n149_n697# a_n207_n600# w_n1947_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X15 a_n741_n600# a_n861_n697# a_n919_n600# w_n1947_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X16 a_n563_n600# a_n683_n697# a_n741_n600# w_n1947_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X17 a_327_n600# a_207_n697# a_149_n600# w_n1947_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X18 a_861_n600# a_741_n697# a_683_n600# w_n1947_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X19 a_683_n600# a_563_n697# a_505_n600# w_n1947_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
.ends

.subckt sky130_fd_pr__nfet_01v8_PGN2UQ VSUBS a_n29_527# a_207_439# a_149_527# a_n505_n815#
+ a_n385_n727# a_327_527# a_505_527# a_n207_527# a_29_n397# a_149_n309# a_n29_n309#
+ a_n149_439# a_n563_n727# a_207_21# a_n327_439# a_n385_109# a_29_n815# a_n505_439#
+ a_385_21# a_n563_109# a_327_n309# a_207_n397# a_n207_n309# a_385_439# a_n149_n397#
+ a_149_n727# a_207_n815# a_n29_n727# a_505_n309# a_n149_21# a_29_21# a_n29_109# a_n149_n815#
+ a_n385_527# a_n563_527# a_149_109# a_385_n397# a_327_109# a_n327_n397# a_n385_n309#
+ a_327_n727# a_n327_21# a_505_109# a_n207_n727# a_n207_109# a_385_n815# a_n327_n815#
+ w_n701_n937# a_29_439# a_n563_n309# a_n505_21# a_n505_n397# a_505_n727#
X0 a_n207_109# a_n327_21# a_n385_109# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=600000u
X1 a_505_109# a_385_21# a_327_109# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=600000u
X2 a_327_n727# a_207_n815# a_149_n727# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=600000u
X3 a_327_109# a_207_21# a_149_109# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=600000u
X4 a_505_n727# a_385_n815# a_327_n727# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=600000u
X5 a_149_n727# a_29_n815# a_n29_n727# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=600000u
X6 a_n207_527# a_n327_439# a_n385_527# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=600000u
X7 a_505_527# a_385_439# a_327_527# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=600000u
X8 a_327_527# a_207_439# a_149_527# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=600000u
X9 a_n385_109# a_n505_21# a_n563_109# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=600000u
X10 a_n385_n309# a_n505_n397# a_n563_n309# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=600000u
X11 a_149_109# a_29_21# a_n29_109# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=600000u
X12 a_n207_n309# a_n327_n397# a_n385_n309# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=600000u
X13 a_n29_109# a_n149_21# a_n207_109# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=600000u
X14 a_n29_n309# a_n149_n397# a_n207_n309# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=600000u
X15 a_327_n309# a_207_n397# a_149_n309# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=600000u
X16 a_n385_527# a_n505_439# a_n563_527# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=600000u
X17 a_n385_n727# a_n505_n815# a_n563_n727# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=600000u
X18 a_n29_527# a_n149_439# a_n207_527# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=600000u
X19 a_149_527# a_29_439# a_n29_527# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=600000u
X20 a_n207_n727# a_n327_n815# a_n385_n727# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=600000u
X21 a_n29_n727# a_n149_n815# a_n207_n727# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=600000u
X22 a_505_n309# a_385_n397# a_327_n309# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=600000u
X23 a_149_n309# a_29_n397# a_n29_n309# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=600000u
.ends

.subckt sky130_fd_pr__pfet_01v8_VXT95W a_n7091_21# a_n1573_n1415# VSUBS a_n5311_21#
+ a_n2107_21# a_n6557_n1415# a_149_n1318# a_n3233_n1318# a_3233_n1415# a_n3945_n1318#
+ a_7327_21# a_2285_118# a_6557_118# a_3945_n1415# a_2641_n1318# a_7625_n1318# a_n385_n1318#
+ a_n6557_21# a_n6259_118# a_1275_21# a_n6081_118# a_n3175_n1415# a_2463_118# a_6735_118#
+ a_n3887_n1415# a_n1987_118# a_5547_n1415# a_n5547_n1318# a_3945_21# a_n6437_118#
+ a_n2165_118# a_385_n1415# a_4243_n1318# a_n683_21# a_3055_21# a_4955_n1318# a_2819_118#
+ a_n2285_21# a_2641_118# a_6913_118# a_n6201_n1415# a_505_n1318# a_n7861_n1318# a_n6913_n1415#
+ a_7861_n1415# a_5725_21# a_n6615_118# a_n2343_118# a_n5489_n1415# a_n2165_n1318#
+ a_n4955_21# a_919_21# a_n1929_n1415# a_n1217_n1415# a_2165_n1415# a_2877_n1415#
+ a_n741_n1318# a_n2877_n1318# a_1573_n1318# a_n7149_n1318# a_7149_n1415# a_n4065_21#
+ a_n29_118# a_6557_n1318# a_n7091_n1415# a_7505_21# a_n2521_118# a_n3531_n1415# a_n6735_21#
+ a_n5903_n1318# a_n683_n1415# a_741_n1415# a_5903_n1415# a_149_118# a_1453_21# a_3887_118#
+ a_4479_n1415# a_n4479_n1318# a_4065_118# a_7981_118# a_3887_n1318# a_3175_n1318#
+ a_n3589_118# a_n6081_n1318# a_2699_21# a_n8039_118# a_n7683_118# a_n5845_n1415#
+ a_n5133_n1415# a_6081_n1415# a_6793_n1415# a_n6793_n1318# a_327_118# a_2521_n1415#
+ a_n2521_n1318# a_n861_21# a_3233_21# a_n29_n1318# a_n7505_n1318# a_7505_n1415# a_n2463_21#
+ a_4243_118# a_1097_n1415# a_6201_n1318# a_n1097_n1318# a_6913_n1318# a_7683_21#
+ a_n3767_118# a_4479_21# a_5903_21# a_n7861_118# a_5489_n1318# a_5013_21# a_505_118#
+ a_1929_n1318# a_1217_n1318# a_n1929_21# a_n2463_n1415# a_n4243_21# a_207_21# a_4421_118#
+ a_n7447_n1415# a_n4123_n1318# a_n1039_21# a_4123_n1415# a_4835_n1415# a_7091_n1318#
+ a_n4835_n1318# a_6259_21# a_n3945_118# a_3531_n1318# a_n4123_118# a_n207_118# a_n327_n1415#
+ a_n5489_21# a_n6913_21# a_n3709_21# a_n6023_21# a_1631_21# a_n4065_n1415# a_n4301_118#
+ a_5489_118# a_n4777_n1415# a_1453_n1415# a_n1453_n1318# a_n7269_21# a_6437_n1415#
+ a_n6437_n1318# a_2877_21# a_5133_n1318# a_5191_21# a_5845_n1318# a_683_n1318# a_3411_21#
+ a_1395_118# a_5667_118# a_385_21# a_n2641_21# a_n7803_n1415# a_n5369_118# a_n1097_118#
+ a_n1395_n1415# a_4657_21# a_7861_21# a_n5191_118# a_n6379_n1415# a_n2107_n1415#
+ a_3055_n1415# a_n3055_n1318# a_n2819_n1415# a_3767_n1415# a_n3767_n1318# a_n8039_n1318#
+ a_n3887_21# a_1573_118# a_5845_118# a_2463_n1318# a_6023_118# a_7447_n1318# a_n4421_21#
+ a_n1217_21# a_n5547_118# a_n1275_118# a_n4421_n1415# a_6437_21# a_1929_118# a_n5667_21#
+ a_1751_118# a_2107_118# a_29_n1415# a_n6201_21# a_6201_118# a_5369_n1415# a_n5369_n1318#
+ a_n5725_118# a_n1453_118# a_1809_n1415# a_4777_n1318# a_4065_n1318# a_n1809_n1318#
+ a_n1751_n1415# a_n7447_21# a_n6735_n1415# a_n6023_n1415# a_327_n1318# a_n7683_n1318#
+ a_7683_n1415# a_3411_n1415# a_n3411_n1318# a_2165_21# a_n1809_118# a_n1631_118#
+ a_n5903_118# a_7091_118# a_7269_118# a_n1039_n1415# a_n563_n1318# a_n1395_21# a_563_21#
+ a_2699_n1415# a_7803_n1318# a_n2699_n1318# a_1395_n1318# a_6379_n1318# a_4835_21#
+ a_2997_118# a_2819_n1318# a_2107_n1318# a_3175_118# a_7447_118# a_n3353_n1415# a_n5013_n1318#
+ a_n3175_21# a_n2699_118# a_5013_n1415# a_5725_n1415# a_n5725_n1318# a_n7149_118#
+ a_n6793_118# a_563_n1415# a_4421_n1318# a_6615_21# a_29_21# a_n5845_21# a_n149_21#
+ a_3353_118# a_7625_118# a_n2877_118# a_n7327_118# a_n6971_118# a_n3055_118# a_n5667_n1415#
+ a_n2343_n1318# a_2343_n1415# a_3709_118# a_1751_n1318# a_n7327_n1318# a_7327_n1415#
+ a_n7625_21# a_3531_118# a_7803_118# a_6735_n1318# a_6023_n1318# a_n7981_n1415# a_n207_n1318#
+ a_2343_21# a_n7505_118# a_n3233_118# a_1039_n1318# a_n919_n1318# a_741_21# a_n1573_21#
+ a_n2997_n1415# a_n2285_n1415# a_n861_n1415# a_6793_21# a_n7269_n1415# a_1809_21#
+ a_3589_21# a_n3709_n1415# a_4657_n1415# a_n4657_n1318# a_4123_21# a_n3411_118# a_4599_118#
+ a_3353_n1318# a_n149_n1415# a_n3353_21# a_207_n1415# a_n5311_n1415# a_919_n1415#
+ a_n6971_n1318# a_683_118# a_6971_n1415# a_5369_21# a_4777_118# a_n4599_21# a_n4599_n1415#
+ a_n1275_n1318# a_n2819_21# a_n327_21# a_1275_n1415# a_1987_n1415# a_n1987_n1318#
+ a_n5133_21# a_n4479_118# a_6259_n1415# a_n6259_n1318# a_n385_118# a_5667_n1318#
+ a_7149_21# a_861_118# a_1039_118# a_4955_118# a_n2641_n1415# a_n7803_21# a_n6379_21#
+ a_5133_118# a_n7625_n1415# w_n8177_n1537# a_1987_21# a_4301_n1415# a_n4301_n1318#
+ a_n4657_118# a_7981_n1318# a_1097_21# a_2521_21# a_n563_118# a_n505_n1415# a_3589_n1415#
+ a_n3589_n1318# a_n1751_21# a_1217_118# a_2997_n1318# a_2285_n1318# a_5311_118# a_7269_n1318#
+ a_3767_21# a_6971_21# a_3709_n1318# a_n5191_n1318# a_6081_21# a_n5013_118# a_n4835_118#
+ a_n919_118# a_n4955_n1415# a_n4243_n1415# a_5191_n1415# a_n2997_21# a_4301_21# a_n741_118#
+ a_1631_n1415# a_n1631_n1318# a_6615_n1415# a_n6615_n1318# a_n3531_21# a_5311_n1318#
+ a_861_n1318# a_5547_21# a_n7981_21# a_6379_118# a_4599_n1318# a_n4777_21# a_n505_21#
X0 a_4243_118# a_4123_21# a_4065_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X1 a_4777_n1318# a_4657_n1415# a_4599_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X2 a_n1097_n1318# a_n1217_n1415# a_n1275_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X3 a_3353_118# a_3233_21# a_3175_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X4 a_n4301_n1318# a_n4421_n1415# a_n4479_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X5 a_2463_118# a_2343_21# a_2285_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X6 a_7981_n1318# a_7861_n1415# a_7803_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X7 a_1573_118# a_1453_21# a_1395_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X8 a_4599_n1318# a_4479_n1415# a_4421_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X9 a_149_n1318# a_29_n1415# a_n29_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X10 a_n919_n1318# a_n1039_n1415# a_n1097_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X11 a_n7861_118# a_n7981_21# a_n8039_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X12 a_n2877_n1318# a_n2997_n1415# a_n3055_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X13 a_n919_118# a_n1039_21# a_n1097_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X14 a_7803_n1318# a_7683_n1415# a_7625_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X15 a_4065_n1318# a_3945_n1415# a_3887_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X16 a_n4123_n1318# a_n4243_n1415# a_n4301_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X17 a_n741_n1318# a_n861_n1415# a_n919_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X18 a_n7683_118# a_n7803_21# a_n7861_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X19 a_n6793_118# a_n6913_21# a_n6971_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X20 a_1217_118# a_1097_21# a_1039_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X21 a_3887_n1318# a_3767_n1415# a_3709_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X22 a_n3945_n1318# a_n4065_n1415# a_n4123_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X23 a_7981_118# a_7861_21# a_7803_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X24 a_5133_n1318# a_5013_n1415# a_4955_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X25 a_n563_n1318# a_n683_n1415# a_n741_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X26 a_n3411_n1318# a_n3531_n1415# a_n3589_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X27 a_7091_118# a_6971_21# a_6913_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X28 a_7091_n1318# a_6971_n1415# a_6913_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X29 a_n563_118# a_n683_21# a_n741_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X30 a_n7327_118# a_n7447_21# a_n7505_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X31 a_6023_118# a_5903_21# a_5845_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X32 a_n7683_n1318# a_n7803_n1415# a_n7861_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X33 a_n6437_118# a_n6557_21# a_n6615_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X34 a_n385_118# a_n505_21# a_n563_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X35 a_3709_n1318# a_3589_n1415# a_3531_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X36 a_n5547_118# a_n5667_21# a_n5725_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X37 a_n3233_n1318# a_n3353_n1415# a_n3411_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X38 a_n4657_118# a_n4777_21# a_n4835_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X39 a_6913_n1318# a_6793_n1415# a_6735_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X40 a_n6971_n1318# a_n7091_n1415# a_n7149_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X41 a_4421_n1318# a_4301_n1415# a_4243_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X42 a_n3767_118# a_n3887_21# a_n3945_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X43 a_n2877_118# a_n2997_21# a_n3055_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X44 a_683_118# a_563_21# a_505_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X45 a_n7505_n1318# a_n7625_n1415# a_n7683_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X46 a_7447_118# a_7327_21# a_7269_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X47 a_n3589_118# a_n3709_21# a_n3767_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X48 a_n2699_118# a_n2819_21# a_n2877_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X49 a_149_118# a_29_21# a_n29_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X50 a_6557_118# a_6437_21# a_6379_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X51 a_2997_n1318# a_2877_n1415# a_2819_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X52 a_n3055_n1318# a_n3175_n1415# a_n3233_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X53 a_n1809_118# a_n1929_21# a_n1987_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X54 a_n29_118# a_n149_21# a_n207_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X55 a_5667_118# a_5547_21# a_5489_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X56 a_4243_n1318# a_4123_n1415# a_4065_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X57 a_4777_118# a_4657_21# a_4599_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X58 a_n2521_n1318# a_n2641_n1415# a_n2699_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X59 a_327_n1318# a_207_n1415# a_149_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X60 a_3887_118# a_3767_21# a_3709_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X61 a_n3589_n1318# a_n3709_n1415# a_n3767_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X62 a_n7327_n1318# a_n7447_n1415# a_n7505_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X63 a_n6081_118# a_n6201_21# a_n6259_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X64 a_2997_118# a_2877_21# a_2819_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X65 a_n5191_118# a_n5311_21# a_n5369_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X66 a_2107_118# a_1987_21# a_1929_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X67 a_n6793_n1318# a_n6913_n1415# a_n6971_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X68 a_2819_n1318# a_2699_n1415# a_2641_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X69 a_n4301_118# a_n4421_21# a_n4479_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X70 a_n2343_n1318# a_n2463_n1415# a_n2521_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X71 a_n3411_118# a_n3531_21# a_n3589_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X72 a_1929_118# a_1809_21# a_1751_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X73 a_n2521_118# a_n2641_21# a_n2699_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X74 a_3531_n1318# a_3411_n1415# a_3353_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X75 a_n7149_n1318# a_n7269_n1415# a_n7327_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X76 a_n1631_118# a_n1751_21# a_n1809_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X77 a_n6615_n1318# a_n6735_n1415# a_n6793_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X78 a_4421_118# a_4301_21# a_4243_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X79 a_2107_n1318# a_1987_n1415# a_1929_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X80 a_n2165_n1318# a_n2285_n1415# a_n2343_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X81 a_3353_n1318# a_3233_n1415# a_3175_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X82 a_3531_118# a_3411_21# a_3353_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X83 a_n1631_n1318# a_n1751_n1415# a_n1809_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X84 a_n3945_118# a_n4065_21# a_n4123_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X85 a_2641_118# a_2521_21# a_2463_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X86 a_n3055_118# a_n3175_21# a_n3233_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X87 a_n2699_n1318# a_n2819_n1415# a_n2877_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X88 a_1751_118# a_1631_21# a_1573_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X89 a_n6437_n1318# a_n6557_n1415# a_n6615_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X90 a_n2165_118# a_n2285_21# a_n2343_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X91 a_7625_n1318# a_7505_n1415# a_7447_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X92 a_n1275_118# a_n1395_21# a_n1453_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X93 a_3175_n1318# a_3055_n1415# a_2997_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X94 a_n1987_118# a_n2107_21# a_n2165_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X95 a_n1453_n1318# a_n1573_n1415# a_n1631_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X96 a_n1097_118# a_n1217_21# a_n1275_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X97 a_2641_n1318# a_2521_n1415# a_2463_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X98 a_n6259_n1318# a_n6379_n1415# a_n6437_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X99 a_3175_118# a_3055_21# a_2997_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X100 a_7447_n1318# a_7327_n1415# a_7269_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X101 a_n385_n1318# a_n505_n1415# a_n563_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X102 a_n5725_n1318# a_n5845_n1415# a_n5903_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X103 a_2285_118# a_2165_21# a_2107_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X104 a_1395_118# a_1275_21# a_1217_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X105 a_n1275_n1318# a_n1395_n1415# a_n1453_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X106 a_6201_n1318# a_6081_n1415# a_6023_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X107 a_2463_n1318# a_2343_n1415# a_2285_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X108 a_1039_118# a_919_21# a_861_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X109 a_7269_n1318# a_7149_n1415# a_7091_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X110 a_n1809_n1318# a_n1929_n1415# a_n1987_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X111 a_n741_118# a_n861_21# a_n919_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X112 a_n207_n1318# a_n327_n1415# a_n385_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X113 a_n5547_n1318# a_n5667_n1415# a_n5725_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X114 a_6735_n1318# a_6615_n1415# a_6557_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X115 a_n7505_118# a_n7625_21# a_n7683_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X116 a_n6615_118# a_n6735_21# a_n6793_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X117 a_2285_n1318# a_2165_n1415# a_2107_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X118 a_n5725_118# a_n5845_21# a_n5903_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X119 a_1751_n1318# a_1631_n1415# a_1573_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X120 a_n4835_118# a_n4955_21# a_n5013_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X121 a_n29_n1318# a_n149_n1415# a_n207_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X122 a_n5369_n1318# a_n5489_n1415# a_n5547_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X123 a_7803_118# a_7683_21# a_7625_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X124 a_6557_n1318# a_6437_n1415# a_6379_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X125 a_861_118# a_741_21# a_683_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X126 a_6913_118# a_6793_21# a_6735_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X127 a_n4835_n1318# a_n4955_n1415# a_n5013_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X128 a_6023_n1318# a_5903_n1415# a_5845_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X129 a_n6081_n1318# a_n6201_n1415# a_n6259_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X130 a_7625_118# a_7505_21# a_7447_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X131 a_6735_118# a_6615_21# a_6557_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X132 a_n7149_118# a_n7269_21# a_n7327_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X133 a_5845_118# a_5725_21# a_5667_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X134 a_5311_n1318# a_5191_n1415# a_5133_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X135 a_1573_n1318# a_1453_n1415# a_1395_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X136 a_n6259_118# a_n6379_21# a_n6437_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X137 a_n207_118# a_n327_21# a_n385_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X138 a_4955_118# a_4835_21# a_4777_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X139 a_n5369_118# a_n5489_21# a_n5547_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X140 a_6379_n1318# a_6259_n1415# a_6201_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X141 a_n4657_n1318# a_n4777_n1415# a_n4835_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X142 a_4065_118# a_3945_21# a_3887_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X143 a_861_n1318# a_741_n1415# a_683_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X144 a_n4479_118# a_n4599_21# a_n4657_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X145 a_5845_n1318# a_5725_n1415# a_5667_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X146 a_n5903_n1318# a_n6023_n1415# a_n6081_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X147 a_n7861_n1318# a_n7981_n1415# a_n8039_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X148 a_505_118# a_385_21# a_327_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X149 a_1395_n1318# a_1275_n1415# a_1217_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X150 a_7269_118# a_7149_21# a_7091_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X151 a_327_118# a_207_21# a_149_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X152 a_6379_118# a_6259_21# a_6201_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X153 a_683_n1318# a_563_n1415# a_505_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X154 a_n4479_n1318# a_n4599_n1415# a_n4657_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X155 a_n6971_118# a_n7091_21# a_n7149_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X156 a_5489_118# a_5369_21# a_5311_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X157 a_5667_n1318# a_5547_n1415# a_5489_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X158 a_1929_n1318# a_1809_n1415# a_1751_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X159 a_n1987_n1318# a_n2107_n1415# a_n2165_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X160 a_4599_118# a_4479_21# a_4421_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X161 a_n5191_n1318# a_n5311_n1415# a_n5369_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X162 a_3709_118# a_3589_21# a_3531_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X163 a_1217_n1318# a_1097_n1415# a_1039_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X164 a_n5903_118# a_n6023_21# a_n6081_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X165 a_2819_118# a_2699_21# a_2641_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X166 a_n5013_118# a_n5133_21# a_n5191_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X167 a_n4123_118# a_n4243_21# a_n4301_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X168 a_505_n1318# a_385_n1415# a_327_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X169 a_5489_n1318# a_5369_n1415# a_5311_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X170 a_n3767_n1318# a_n3887_n1415# a_n3945_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X171 a_n3233_118# a_n3353_21# a_n3411_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X172 a_6201_118# a_6081_21# a_6023_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X173 a_4955_n1318# a_4835_n1415# a_4777_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X174 a_n5013_n1318# a_n5133_n1415# a_n5191_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X175 a_n2343_118# a_n2463_21# a_n2521_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X176 a_1039_n1318# a_919_n1415# a_861_n1318# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X177 a_n1453_118# a_n1573_21# a_n1631_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X178 a_5311_118# a_5191_21# a_5133_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X179 a_5133_118# a_5013_21# a_4955_118# w_n8177_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
.ends

.subckt sky130_fd_pr__nfet_01v8_XGTW7K VSUBS a_n1275_109# a_n861_n1397# a_1275_21#
+ a_n1453_109# a_1751_109# a_n149_n1397# a_207_n1397# a_919_n1397# a_n1809_n1309#
+ a_1275_n1397# a_327_n1309# a_n683_21# a_n1809_109# a_n1631_109# a_n563_n1309# a_1395_n1309#
+ a_919_21# a_n505_n1397# a_1631_n1397# a_1453_21# a_1751_n1309# a_n861_21# a_n1573_n1397#
+ a_n919_n1309# a_n207_n1309# a_1039_n1309# a_n1039_21# a_207_21# a_683_109# a_n385_109#
+ a_385_n1397# a_n1275_n1309# a_1631_21# a_861_109# a_1039_109# a_n1217_n1397# a_385_21#
+ a_n563_109# a_1217_109# a_n919_109# a_n741_109# a_n683_n1397# a_741_n1397# a_n1631_n1309#
+ a_n1217_21# a_861_n1309# a_149_n1309# a_1097_n1397# a_n385_n1309# a_n1395_21# a_563_21#
+ a_n327_n1397# a_1453_n1397# a_505_n1309# a_n149_21# a_29_21# a_n29_109# a_n741_n1309#
+ a_1573_n1309# a_n1395_n1397# a_149_109# a_n1573_21# a_741_21# a_327_109# a_29_n1397#
+ a_n1751_n1397# a_n1097_n1309# a_n29_n1309# a_n327_21# a_505_109# a_n1039_n1397#
+ a_1217_n1309# a_n207_109# a_1097_21# a_563_n1397# a_n1751_21# a_n1453_n1309# a_683_n1309#
+ a_n1097_109# a_1395_109# w_n1947_n1519# a_n505_21# a_1573_109#
X0 a_n207_109# a_n327_21# a_n385_109# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X1 a_1573_n1309# a_1453_n1397# a_1395_n1309# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X2 a_861_n1309# a_741_n1397# a_683_n1309# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X3 a_505_109# a_385_21# a_327_109# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X4 a_1395_n1309# a_1275_n1397# a_1217_n1309# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X5 a_327_109# a_207_21# a_149_109# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X6 a_683_n1309# a_563_n1397# a_505_n1309# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X7 a_1217_n1309# a_1097_n1397# a_1039_n1309# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X8 a_505_n1309# a_385_n1397# a_327_n1309# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X9 a_1039_n1309# a_919_n1397# a_861_n1309# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X10 a_n1453_109# a_n1573_21# a_n1631_109# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X11 a_n1097_n1309# a_n1217_n1397# a_n1275_n1309# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X12 a_1573_109# a_1453_21# a_1395_109# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X13 a_n919_n1309# a_n1039_n1397# a_n1097_n1309# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X14 a_149_n1309# a_29_n1397# a_n29_n1309# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X15 a_n919_109# a_n1039_21# a_n1097_109# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X16 a_n741_n1309# a_n861_n1397# a_n919_n1309# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X17 a_1217_109# a_1097_21# a_1039_109# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X18 a_n563_n1309# a_n683_n1397# a_n741_n1309# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X19 a_n563_109# a_n683_21# a_n741_109# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X20 a_n385_109# a_n505_21# a_n563_109# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X21 a_683_109# a_563_21# a_505_109# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X22 a_149_109# a_29_21# a_n29_109# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X23 a_n29_109# a_n149_21# a_n207_109# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X24 a_327_n1309# a_207_n1397# a_149_n1309# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X25 a_n1631_109# a_n1751_21# a_n1809_109# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X26 a_1751_109# a_1631_21# a_1573_109# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X27 a_n1631_n1309# a_n1751_n1397# a_n1809_n1309# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X28 a_n1275_109# a_n1395_21# a_n1453_109# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X29 a_n1097_109# a_n1217_21# a_n1275_109# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X30 a_n1453_n1309# a_n1573_n1397# a_n1631_n1309# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X31 a_n385_n1309# a_n505_n1397# a_n563_n1309# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X32 a_1039_109# a_919_21# a_861_109# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X33 a_1395_109# a_1275_21# a_1217_109# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X34 a_n1275_n1309# a_n1395_n1397# a_n1453_n1309# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X35 a_n741_109# a_n861_21# a_n919_109# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X36 a_n207_n1309# a_n327_n1397# a_n385_n1309# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X37 a_n29_n1309# a_n149_n1397# a_n207_n1309# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X38 a_1751_n1309# a_1631_n1397# a_1573_n1309# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X39 a_861_109# a_741_21# a_683_109# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
.ends

.subckt sky130_fd_pr__nfet_01v8_X8JY7K VSUBS a_n1217_n688# a_n385_n600# a_1039_n600#
+ a_207_n688# a_n149_n688# a_n1631_n600# a_n919_n600# a_683_n600# a_1631_n688# a_1217_n600#
+ a_n1395_n688# a_n563_n600# a_385_n688# a_n327_n688# a_919_n688# a_861_n600# a_n741_n600#
+ a_n1573_n688# a_1395_n600# a_563_n688# a_n505_n688# a_n1097_n600# a_149_n600# a_n29_n600#
+ a_1097_n688# a_n1751_n688# a_741_n688# a_1573_n600# a_n1275_n600# a_327_n600# a_n683_n688#
+ a_29_n688# a_1275_n688# a_n1039_n688# a_n1809_n600# a_n207_n600# a_1751_n600# a_n1453_n600#
+ a_505_n600# w_n1947_n810# a_n861_n688# a_1453_n688#
X0 a_n385_n600# a_n505_n688# a_n563_n600# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X1 a_n1631_n600# a_n1751_n688# a_n1809_n600# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X2 a_n207_n600# a_n327_n688# a_n385_n600# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X3 a_n1453_n600# a_n1573_n688# a_n1631_n600# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X4 a_n29_n600# a_n149_n688# a_n207_n600# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X5 a_n1275_n600# a_n1395_n688# a_n1453_n600# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X6 a_n741_n600# a_n861_n688# a_n919_n600# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X7 a_n563_n600# a_n683_n688# a_n741_n600# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X8 a_327_n600# a_207_n688# a_149_n600# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X9 a_683_n600# a_563_n688# a_505_n600# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X10 a_861_n600# a_741_n688# a_683_n600# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X11 a_505_n600# a_385_n688# a_327_n600# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X12 a_149_n600# a_29_n688# a_n29_n600# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X13 a_1751_n600# a_1631_n688# a_1573_n600# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X14 a_1573_n600# a_1453_n688# a_1395_n600# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X15 a_1217_n600# a_1097_n688# a_1039_n600# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X16 a_1395_n600# a_1275_n688# a_1217_n600# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X17 a_n1097_n600# a_n1217_n688# a_n1275_n600# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X18 a_1039_n600# a_919_n688# a_861_n600# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
X19 a_n919_n600# a_n1039_n688# a_n1097_n600# VSUBS sky130_fd_pr__nfet_01v8 w=6e+06u l=600000u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_BLS9H9 VSUBS c1_n1841_n1500# m3_n1941_n1600#
X0 c1_n1841_n1500# m3_n1941_n1600# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.755e+07u
.ends

.subckt sky130_fd_pr__pfet_01v8_VXTQ3X VSUBS a_n1631_n600# a_n919_n600# a_1217_n600#
+ a_n563_n600# a_861_n600# w_n1769_n819# a_149_n600# a_1573_n600# a_n1275_n600# a_n207_n600#
+ a_505_n600#
X0 a_505_n600# a_385_n697# a_327_n600# w_n1769_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X1 a_149_n600# a_29_n697# a_n29_n600# w_n1769_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X2 a_1573_n600# a_1453_n697# a_1395_n600# w_n1769_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X3 a_1395_n600# a_1275_n697# a_1217_n600# w_n1769_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X4 a_1217_n600# a_1097_n697# a_1039_n600# w_n1769_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X5 a_n1097_n600# a_n1217_n697# a_n1275_n600# w_n1769_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X6 a_1039_n600# a_919_n697# a_861_n600# w_n1769_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X7 a_n919_n600# a_n1039_n697# a_n1097_n600# w_n1769_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X8 a_n385_n600# a_n505_n697# a_n563_n600# w_n1769_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X9 a_n207_n600# a_n327_n697# a_n385_n600# w_n1769_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X10 a_n1453_n600# a_n1573_n697# a_n1631_n600# w_n1769_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X11 a_n1275_n600# a_n1395_n697# a_n1453_n600# w_n1769_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X12 a_n29_n600# a_n149_n697# a_n207_n600# w_n1769_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X13 a_n741_n600# a_n861_n697# a_n919_n600# w_n1769_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X14 a_n563_n600# a_n683_n697# a_n741_n600# w_n1769_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X15 a_327_n600# a_207_n697# a_149_n600# w_n1769_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X16 a_861_n600# a_741_n697# a_683_n600# w_n1769_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X17 a_683_n600# a_563_n697# a_505_n600# w_n1769_n819# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
.ends

.subckt sky130_fd_pr__pfet_01v8_JXF9S2 a_2076_21# a_3500_21# a_3264_n1318# VSUBS a_474_21#
+ a_3976_n1318# a_n2730_21# a_n1364_118# a_118_n1415# a_n2610_n1318# a_1840_118# a_2610_n1415#
+ a_n3976_21# a_n1542_118# a_n1186_n1318# a_n1898_n1318# a_1186_n1415# a_n3086_21#
+ a_n1306_21# a_1898_n1415# a_n60_n1415# a_1306_n1318# a_n2552_n1415# a_n1720_118#
+ a_3086_118# a_3620_n1318# a_n416_n1415# a_2196_n1318# a_3264_118# a_2254_21# a_n2788_118#
+ a_n1542_n1318# a_1542_n1415# a_n1484_21# a_652_21# a_772_n1318# a_3442_118# a_n2966_118#
+ a_n3264_21# a_n3144_118# a_n1484_n1415# a_n3144_n1318# a_3144_n1415# a_2552_n1318#
+ a_n3856_n1318# a_3856_n1415# a_n2908_n1415# a_3620_118# a_n238_21# a_n3322_118#
+ a_n296_n1318# a_594_118# a_n3086_n1415# a_n3798_n1415# a_1898_21# a_n3500_118# a_296_n1415#
+ a_2432_21# a_830_21# a_n296_118# a_n1662_21# a_772_118# a_n1840_n1415# a_416_n1318#
+ a_n3500_n1318# a_3678_21# a_3500_n1415# a_1008_21# a_n652_n1318# a_n2076_n1318#
+ a_n2788_n1318# a_2076_n1415# a_n1128_n1415# a_n474_118# a_1484_n1318# a_2788_n1415#
+ a_n3442_21# a_950_118# a_1128_118# a_2908_n1318# a_n3442_n1415# a_n2908_21# a_n416_21#
+ a_n652_118# a_n594_n1415# a_n2018_21# a_652_n1415# a_1306_118# a_3086_n1318# a_3798_n1318#
+ a_n1008_118# a_60_n1318# a_n830_118# a_1186_21# a_2610_21# a_n2432_n1318# a_2432_n1415#
+ a_n60_21# a_n1840_21# a_1840_n1318# a_2196_118# a_3856_21# a_n594_21# a_1128_n1318#
+ a_n2374_n1415# a_n3620_21# a_n2196_21# a_n950_n1415# a_2374_118# a_n4034_n1318#
+ a_3442_n1318# a_n1898_118# a_n2076_118# a_n238_n1415# a_2552_118# a_n1364_n1318#
+ a_1364_n1415# a_n2254_118# a_60_118# a_2908_118# a_1364_21# a_2730_118# a_594_n1318#
+ a_n2730_n1415# a_n2432_118# a_n772_21# a_3144_21# a_n3678_n1318# a_n2018_n1415#
+ a_2374_n1318# a_3678_n1415# a_n2374_21# a_n2610_118# a_3798_118# a_n1720_n1318#
+ a_1720_n1415# a_238_118# a_118_21# a_3976_118# a_950_n1318# a_n1008_n1318# a_1008_n1415#
+ a_n3678_118# a_n1662_n1415# a_416_118# a_238_n1318# a_n3322_n1318# a_3322_n1415#
+ a_1542_21# a_2730_n1318# a_n3856_118# a_n474_n1318# a_n4034_118# a_n118_118# a_2788_21#
+ a_2018_n1318# a_n950_21# a_3322_21# a_n3264_n1415# a_296_21# a_n3976_n1415# a_n2552_21#
+ a_474_n1415# a_n3798_21# a_n1128_21# a_n830_n1318# a_n2254_n1318# a_2254_n1415#
+ a_n1306_n1415# a_n2966_n1318# a_2966_n1415# a_1662_n1318# a_1484_118# a_1720_21#
+ a_n118_n1318# w_n4172_n1537# a_n3620_n1415# a_n1186_118# a_n772_n1415# a_n2196_n1415#
+ a_830_n1415# a_2966_21# a_1662_118# a_2018_118#
X0 a_n2788_118# a_n2908_21# a_n2966_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X1 a_n118_118# a_n238_21# a_n296_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X2 a_n1008_n1318# a_n1128_n1415# a_n1186_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X3 a_3086_118# a_2966_21# a_2908_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X4 a_3976_118# a_3856_21# a_3798_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X5 a_238_118# a_118_21# a_60_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X6 a_416_118# a_296_21# a_238_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X7 a_n652_n1318# a_n772_n1415# a_n830_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X8 a_3976_n1318# a_3856_n1415# a_3798_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X9 a_n3144_118# a_n3264_21# a_n3322_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X10 a_2730_118# a_2610_21# a_2552_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X11 a_3620_118# a_3500_21# a_3442_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X12 a_n3322_n1318# a_n3442_n1415# a_n3500_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X13 a_n474_n1318# a_n594_n1415# a_n652_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X14 a_3798_n1318# a_3678_n1415# a_3620_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X15 a_n2254_118# a_n2374_21# a_n2432_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X16 a_n1364_118# a_n1484_21# a_n1542_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X17 a_1840_118# a_1720_21# a_1662_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X18 a_n1186_118# a_n1306_21# a_n1364_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X19 a_n3144_n1318# a_n3264_n1415# a_n3322_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X20 a_1128_n1318# a_1008_n1415# a_950_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X21 a_3086_n1318# a_2966_n1415# a_2908_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X22 a_2374_118# a_2254_21# a_2196_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X23 a_3264_118# a_3144_21# a_3086_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X24 a_n830_n1318# a_n950_n1415# a_n1008_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X25 a_1484_118# a_1364_21# a_1306_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X26 a_n2966_n1318# a_n3086_n1415# a_n3144_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X27 a_2908_n1318# a_2788_n1415# a_2730_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X28 a_n2432_n1318# a_n2552_n1415# a_n2610_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X29 a_238_n1318# a_118_n1415# a_60_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X30 a_3620_n1318# a_3500_n1415# a_3442_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X31 a_n3500_n1318# a_n3620_n1415# a_n3678_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X32 a_n2254_n1318# a_n2374_n1415# a_n2432_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X33 a_3442_n1318# a_3322_n1415# a_3264_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X34 a_n474_118# a_n594_21# a_n652_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X35 a_950_118# a_830_21# a_772_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X36 a_n2788_n1318# a_n2908_n1415# a_n2966_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X37 a_n296_118# a_n416_21# a_n474_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X38 a_n2076_n1318# a_n2196_n1415# a_n2254_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X39 a_2018_n1318# a_1898_n1415# a_1840_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X40 a_3264_n1318# a_3144_n1415# a_3086_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X41 a_n2610_n1318# a_n2730_n1415# a_n2788_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X42 a_n1542_n1318# a_n1662_n1415# a_n1720_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X43 a_2730_n1318# a_2610_n1415# a_2552_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X44 a_n3678_118# a_n3798_21# a_n3856_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X45 a_594_118# a_474_21# a_416_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X46 a_n3500_118# a_n3620_21# a_n3678_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X47 a_n2610_118# a_n2730_21# a_n2788_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X48 a_n1720_118# a_n1840_21# a_n1898_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X49 a_n1364_n1318# a_n1484_n1415# a_n1542_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X50 a_2552_n1318# a_2432_n1415# a_2374_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X51 a_3798_118# a_3678_21# a_3620_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X52 a_n296_n1318# a_n416_n1415# a_n474_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X53 a_2018_118# a_1898_21# a_1840_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X54 a_2908_118# a_2788_21# a_2730_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X55 a_2374_n1318# a_2254_n1415# a_2196_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X56 a_n3322_118# a_n3442_21# a_n3500_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X57 a_n2432_118# a_n2552_21# a_n2610_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X58 a_n1720_n1318# a_n1840_n1415# a_n1898_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X59 a_n118_n1318# a_n238_n1415# a_n296_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X60 a_1840_n1318# a_1720_n1415# a_1662_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X61 a_n1542_118# a_n1662_21# a_n1720_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X62 a_2196_n1318# a_2076_n1415# a_2018_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X63 a_3442_118# a_3322_21# a_3264_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X64 a_1662_n1318# a_1542_n1415# a_1484_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X65 a_n2966_118# a_n3086_21# a_n3144_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X66 a_n2076_118# a_n2196_21# a_n2254_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X67 a_1662_118# a_1542_21# a_1484_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X68 a_2552_118# a_2432_21# a_2374_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X69 a_950_n1318# a_830_n1415# a_772_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X70 a_n1898_118# a_n2018_21# a_n2076_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X71 a_60_118# a_n60_21# a_n118_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X72 a_1484_n1318# a_1364_n1415# a_1306_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X73 a_n1008_118# a_n1128_21# a_n1186_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X74 a_n830_118# a_n950_21# a_n1008_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X75 a_772_n1318# a_652_n1415# a_594_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X76 a_1306_118# a_1186_21# a_1128_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X77 a_2196_118# a_2076_21# a_2018_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X78 a_60_n1318# a_n60_n1415# a_n118_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X79 a_1306_n1318# a_1186_n1415# a_1128_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X80 a_1128_118# a_1008_21# a_950_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X81 a_n3856_n1318# a_n3976_n1415# a_n4034_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X82 a_n1898_n1318# a_n2018_n1415# a_n2076_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X83 a_594_n1318# a_474_n1415# a_416_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X84 a_n652_118# a_n772_21# a_n830_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X85 a_n3678_n1318# a_n3798_n1415# a_n3856_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X86 a_416_n1318# a_296_n1415# a_238_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X87 a_n3856_118# a_n3976_21# a_n4034_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X88 a_772_118# a_652_21# a_594_118# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
X89 a_n1186_n1318# a_n1306_n1415# a_n1364_n1318# w_n4172_n1537# sky130_fd_pr__pfet_01v8 w=6e+06u l=600000u
.ends


* Top level circuit opampjulia

Xsky130_fd_pr__pfet_01v8_VXTF3X_1 VSUBS m1_52340_n69842# m1_52340_n69842# m1_60836_n71396#
+ vp vp m1_60836_n71396# m1_52340_n69842# m1_60836_n71396# vp m1_60836_n71396# vp
+ m1_60836_n71396# m1_60836_n71396# m1_60836_n71396# vp m1_52340_n69842# m1_60836_n71396#
+ m1_60836_n71396# m1_52340_n69842# m1_60836_n71396# m1_60836_n71396# m1_52340_n69842#
+ vp m1_52340_n69842# m1_60836_n71396# m1_60836_n71396# vp w_56149_n71520# vp m1_52340_n69842#
+ m1_60836_n71396# m1_60836_n71396# m1_60836_n71396# m1_52340_n69842# vp m1_60836_n71396#
+ m1_52340_n69842# m1_60836_n71396# m1_52340_n69842# vp m1_60836_n71396# m1_60836_n71396#
+ sky130_fd_pr__pfet_01v8_VXTF3X
Xsky130_fd_pr__nfet_01v8_PGN2UQ_0 VSUBS m3_67376_n80074# m1_68118_n71254# m1_68118_n71254#
+ m1_68118_n71254# m3_67376_n80074# m3_67376_n80074# m1_68118_n71254# m1_68118_n71254#
+ m1_68118_n71254# m1_68118_n71254# m3_67376_n80074# m1_68118_n71254# m1_68118_n71254#
+ m1_68118_n71254# m1_68118_n71254# m3_67376_n80074# m1_68118_n71254# m1_68118_n71254#
+ m1_68118_n71254# m1_68118_n71254# m3_67376_n80074# m1_68118_n71254# m1_68118_n71254#
+ m1_68118_n71254# m1_68118_n71254# m1_68118_n71254# m1_68118_n71254# m3_67376_n80074#
+ m1_68118_n71254# m1_68118_n71254# m1_68118_n71254# m3_67376_n80074# m1_68118_n71254#
+ m3_67376_n80074# m1_68118_n71254# m1_68118_n71254# m1_68118_n71254# m3_67376_n80074#
+ m1_68118_n71254# m3_67376_n80074# m3_67376_n80074# m1_68118_n71254# m1_68118_n71254#
+ m1_68118_n71254# m1_68118_n71254# m1_68118_n71254# m1_68118_n71254# VSUBS m1_68118_n71254#
+ m1_68118_n71254# m1_68118_n71254# m1_68118_n71254# m1_68118_n71254# sky130_fd_pr__nfet_01v8_PGN2UQ
Xsky130_fd_pr__pfet_01v8_VXT95W_1 m1_60836_n71396# m1_60836_n71396# VSUBS m1_60836_n71396#
+ m1_60836_n71396# m1_60836_n71396# m1_68118_n71254# vout m1_60836_n71396# vout m1_60836_n71396#
+ m1_68118_n71254# m1_68118_n71254# m1_60836_n71396# m1_68118_n71254# m1_68118_n71254#
+ vout m1_60836_n71396# m1_68118_n71254# m1_60836_n71396# vout m1_60836_n71396# vout
+ vout m1_60836_n71396# m1_68118_n71254# m1_60836_n71396# m1_68118_n71254# m1_60836_n71396#
+ vout vout m1_60836_n71396# vout m1_60836_n71396# m1_60836_n71396# vout vout m1_60836_n71396#
+ m1_68118_n71254# m1_68118_n71254# m1_60836_n71396# m1_68118_n71254# vout m1_60836_n71396#
+ m1_60836_n71396# m1_60836_n71396# m1_68118_n71254# m1_68118_n71254# m1_60836_n71396#
+ vout m1_60836_n71396# m1_60836_n71396# m1_60836_n71396# m1_60836_n71396# m1_60836_n71396#
+ m1_60836_n71396# vout vout m1_68118_n71254# vout m1_60836_n71396# m1_60836_n71396#
+ vout m1_68118_n71254# m1_60836_n71396# m1_60836_n71396# vout m1_60836_n71396# m1_60836_n71396#
+ m1_68118_n71254# m1_60836_n71396# m1_60836_n71396# m1_60836_n71396# m1_68118_n71254#
+ m1_60836_n71396# vout m1_60836_n71396# m1_68118_n71254# m1_68118_n71254# m1_68118_n71254#
+ vout vout vout vout m1_60836_n71396# m1_68118_n71254# m1_68118_n71254# m1_60836_n71396#
+ m1_60836_n71396# m1_60836_n71396# m1_60836_n71396# vout vout m1_60836_n71396# vout
+ m1_60836_n71396# m1_60836_n71396# vout vout m1_60836_n71396# m1_60836_n71396# vout
+ m1_60836_n71396# m1_68118_n71254# vout m1_68118_n71254# m1_60836_n71396# m1_68118_n71254#
+ m1_60836_n71396# m1_60836_n71396# vout m1_68118_n71254# m1_60836_n71396# m1_68118_n71254#
+ m1_68118_n71254# m1_68118_n71254# m1_60836_n71396# m1_60836_n71396# m1_60836_n71396#
+ m1_60836_n71396# m1_68118_n71254# m1_60836_n71396# m1_68118_n71254# m1_60836_n71396#
+ m1_60836_n71396# m1_60836_n71396# vout m1_68118_n71254# m1_60836_n71396# vout vout
+ m1_68118_n71254# m1_68118_n71254# m1_60836_n71396# m1_60836_n71396# m1_60836_n71396#
+ m1_60836_n71396# m1_60836_n71396# m1_60836_n71396# m1_60836_n71396# vout m1_68118_n71254#
+ m1_60836_n71396# m1_60836_n71396# vout m1_60836_n71396# m1_60836_n71396# vout m1_60836_n71396#
+ m1_68118_n71254# m1_60836_n71396# m1_68118_n71254# vout m1_60836_n71396# vout vout
+ m1_60836_n71396# m1_60836_n71396# m1_60836_n71396# vout vout m1_60836_n71396# m1_60836_n71396#
+ m1_60836_n71396# m1_68118_n71254# m1_60836_n71396# m1_60836_n71396# m1_60836_n71396#
+ m1_68118_n71254# m1_60836_n71396# m1_60836_n71396# m1_68118_n71254# m1_68118_n71254#
+ m1_60836_n71396# m1_68118_n71254# m1_68118_n71254# vout vout vout m1_60836_n71396#
+ m1_60836_n71396# m1_68118_n71254# m1_68118_n71254# m1_60836_n71396# m1_60836_n71396#
+ m1_68118_n71254# m1_60836_n71396# vout vout m1_60836_n71396# m1_60836_n71396# m1_68118_n71254#
+ m1_60836_n71396# vout vout vout m1_60836_n71396# m1_68118_n71254# m1_68118_n71254#
+ vout m1_60836_n71396# m1_60836_n71396# m1_60836_n71396# m1_60836_n71396# vout m1_68118_n71254#
+ m1_60836_n71396# m1_60836_n71396# m1_68118_n71254# m1_60836_n71396# vout m1_68118_n71254#
+ m1_68118_n71254# vout m1_68118_n71254# m1_60836_n71396# m1_68118_n71254# m1_60836_n71396#
+ m1_60836_n71396# m1_60836_n71396# vout m1_68118_n71254# vout vout m1_60836_n71396#
+ m1_68118_n71254# vout vout vout vout m1_60836_n71396# vout m1_60836_n71396# m1_68118_n71254#
+ m1_60836_n71396# m1_60836_n71396# vout vout vout m1_60836_n71396# m1_68118_n71254#
+ m1_60836_n71396# m1_60836_n71396# m1_60836_n71396# m1_60836_n71396# m1_68118_n71254#
+ m1_68118_n71254# vout m1_68118_n71254# m1_68118_n71254# m1_68118_n71254# m1_60836_n71396#
+ m1_68118_n71254# m1_60836_n71396# m1_68118_n71254# vout m1_68118_n71254# m1_60836_n71396#
+ m1_60836_n71396# vout vout vout vout m1_60836_n71396# m1_68118_n71254# m1_60836_n71396#
+ vout vout vout m1_68118_n71254# m1_60836_n71396# m1_60836_n71396# m1_60836_n71396#
+ m1_60836_n71396# m1_60836_n71396# m1_60836_n71396# m1_60836_n71396# m1_60836_n71396#
+ m1_60836_n71396# m1_60836_n71396# m1_60836_n71396# vout m1_60836_n71396# m1_68118_n71254#
+ vout m1_68118_n71254# m1_60836_n71396# m1_60836_n71396# m1_60836_n71396# m1_60836_n71396#
+ m1_60836_n71396# m1_68118_n71254# vout m1_60836_n71396# m1_60836_n71396# m1_68118_n71254#
+ m1_60836_n71396# m1_60836_n71396# m1_68118_n71254# m1_60836_n71396# m1_60836_n71396#
+ m1_60836_n71396# m1_60836_n71396# m1_68118_n71254# m1_60836_n71396# m1_68118_n71254#
+ m1_60836_n71396# m1_68118_n71254# vout vout m1_60836_n71396# m1_68118_n71254# vout
+ vout m1_60836_n71396# m1_60836_n71396# m1_60836_n71396# m1_68118_n71254# m1_60836_n71396#
+ w_56149_n71520# m1_60836_n71396# m1_60836_n71396# vout vout m1_68118_n71254# m1_60836_n71396#
+ m1_60836_n71396# m1_68118_n71254# m1_60836_n71396# m1_60836_n71396# vout m1_60836_n71396#
+ m1_68118_n71254# m1_68118_n71254# m1_68118_n71254# vout m1_68118_n71254# m1_60836_n71396#
+ m1_60836_n71396# m1_68118_n71254# m1_68118_n71254# m1_60836_n71396# vout m1_68118_n71254#
+ m1_68118_n71254# m1_60836_n71396# m1_60836_n71396# m1_60836_n71396# m1_60836_n71396#
+ m1_60836_n71396# vout m1_60836_n71396# m1_68118_n71254# m1_60836_n71396# m1_68118_n71254#
+ m1_60836_n71396# vout m1_68118_n71254# m1_60836_n71396# m1_60836_n71396# vout vout
+ m1_60836_n71396# m1_60836_n71396# sky130_fd_pr__pfet_01v8_VXT95W
Xsky130_fd_pr__nfet_01v8_XGTW7K_0 VSUBS vout m1_68118_n71254# m1_68118_n71254# m2_54836_n91946#
+ m2_54836_n91946# m1_68118_n71254# m1_68118_n71254# m1_68118_n71254# m2_54836_n91946#
+ m1_68118_n71254# m2_54836_n91946# m1_68118_n71254# m2_54836_n91946# vout vout m2_54836_n91946#
+ m1_68118_n71254# m1_68118_n71254# m1_68118_n71254# m1_68118_n71254# m2_54836_n91946#
+ m1_68118_n71254# m1_68118_n71254# vout vout m2_54836_n91946# m1_68118_n71254# m1_68118_n71254#
+ m2_54836_n91946# m2_54836_n91946# m1_68118_n71254# vout m1_68118_n71254# vout m2_54836_n91946#
+ m1_68118_n71254# m1_68118_n71254# vout vout vout m2_54836_n91946# m1_68118_n71254#
+ m1_68118_n71254# vout m1_68118_n71254# vout vout m1_68118_n71254# m2_54836_n91946#
+ m1_68118_n71254# m1_68118_n71254# m1_68118_n71254# m1_68118_n71254# vout m1_68118_n71254#
+ m1_68118_n71254# m2_54836_n91946# m2_54836_n91946# vout m1_68118_n71254# vout m1_68118_n71254#
+ m1_68118_n71254# m2_54836_n91946# m1_68118_n71254# m1_68118_n71254# m2_54836_n91946#
+ m2_54836_n91946# m1_68118_n71254# vout m1_68118_n71254# vout vout m1_68118_n71254#
+ m1_68118_n71254# m1_68118_n71254# m2_54836_n91946# m2_54836_n91946# m2_54836_n91946#
+ m2_54836_n91946# VSUBS m1_68118_n71254# vout sky130_fd_pr__nfet_01v8_XGTW7K
Xsky130_fd_pr__nfet_01v8_X8JY7K_0 VSUBS m1_56974_n89276# m2_54836_n91946# m2_54836_n91946#
+ m1_58392_n89276# m1_58036_n89280# m1_56454_n79854# m1_56454_n79854# m2_54836_n91946#
+ m1_59820_n89280# m1_56454_n79854# m1_56796_n89276# m1_56454_n79854# m1_58590_n89280#
+ m1_57880_n89280# m1_59108_n89284# m1_56454_n79854# m2_54836_n91946# m1_56608_n89276#
+ m2_54836_n91946# m1_58750_n89282# m1_57676_n89276# m2_54836_n91946# m1_56454_n79854#
+ m2_54836_n91946# m1_59294_n89282# m1_56438_n89278# m1_58942_n89282# m1_56454_n79854#
+ m1_56454_n79854# m2_54836_n91946# m1_57522_n89276# m1_58232_n89280# m1_59464_n89280#
+ m1_57156_n89284# m2_54836_n91946# m1_56454_n79854# m2_54836_n91946# m2_54836_n91946#
+ m1_56454_n79854# VSUBS m1_57334_n89282# m1_59654_n89288# sky130_fd_pr__nfet_01v8_X8JY7K
Xsky130_fd_pr__nfet_01v8_XGTW7K_1 VSUBS vout m1_68118_n71254# m1_68118_n71254# m2_54836_n91946#
+ m2_54836_n91946# m1_68118_n71254# m1_68118_n71254# m1_68118_n71254# m2_54836_n91946#
+ m1_68118_n71254# m2_54836_n91946# m1_68118_n71254# m2_54836_n91946# vout vout m2_54836_n91946#
+ m1_68118_n71254# m1_68118_n71254# m1_68118_n71254# m1_68118_n71254# m2_54836_n91946#
+ m1_68118_n71254# m1_68118_n71254# vout vout m2_54836_n91946# m1_68118_n71254# m1_68118_n71254#
+ m2_54836_n91946# m2_54836_n91946# m1_68118_n71254# vout m1_68118_n71254# vout m2_54836_n91946#
+ m1_68118_n71254# m1_68118_n71254# vout vout vout m2_54836_n91946# m1_68118_n71254#
+ m1_68118_n71254# vout m1_68118_n71254# vout vout m1_68118_n71254# m2_54836_n91946#
+ m1_68118_n71254# m1_68118_n71254# m1_68118_n71254# m1_68118_n71254# vout m1_68118_n71254#
+ m1_68118_n71254# m2_54836_n91946# m2_54836_n91946# vout m1_68118_n71254# vout m1_68118_n71254#
+ m1_68118_n71254# m2_54836_n91946# m1_68118_n71254# m1_68118_n71254# m2_54836_n91946#
+ m2_54836_n91946# m1_68118_n71254# vout m1_68118_n71254# vout vout m1_68118_n71254#
+ m1_68118_n71254# m1_68118_n71254# m2_54836_n91946# m2_54836_n91946# m2_54836_n91946#
+ m2_54836_n91946# VSUBS m1_68118_n71254# vout sky130_fd_pr__nfet_01v8_XGTW7K
Xsky130_fd_pr__nfet_01v8_XGTW7K_2 VSUBS vout m1_68118_n71254# m1_68118_n71254# m2_54836_n91946#
+ m2_54836_n91946# m1_68118_n71254# m1_68118_n71254# m1_68118_n71254# m2_54836_n91946#
+ m1_68118_n71254# m2_54836_n91946# m1_68118_n71254# m2_54836_n91946# vout vout m2_54836_n91946#
+ m1_68118_n71254# m1_68118_n71254# m1_68118_n71254# m1_68118_n71254# m2_54836_n91946#
+ m1_68118_n71254# m1_68118_n71254# vout vout m2_54836_n91946# m1_68118_n71254# m1_68118_n71254#
+ m2_54836_n91946# m2_54836_n91946# m1_68118_n71254# vout m1_68118_n71254# vout m2_54836_n91946#
+ m1_68118_n71254# m1_68118_n71254# vout vout vout m2_54836_n91946# m1_68118_n71254#
+ m1_68118_n71254# vout m1_68118_n71254# vout vout m1_68118_n71254# m2_54836_n91946#
+ m1_68118_n71254# m1_68118_n71254# m1_68118_n71254# m1_68118_n71254# vout m1_68118_n71254#
+ m1_68118_n71254# m2_54836_n91946# m2_54836_n91946# vout m1_68118_n71254# vout m1_68118_n71254#
+ m1_68118_n71254# m2_54836_n91946# m1_68118_n71254# m1_68118_n71254# m2_54836_n91946#
+ m2_54836_n91946# m1_68118_n71254# vout m1_68118_n71254# vout vout m1_68118_n71254#
+ m1_68118_n71254# m1_68118_n71254# m2_54836_n91946# m2_54836_n91946# m2_54836_n91946#
+ m2_54836_n91946# VSUBS m1_68118_n71254# vout sky130_fd_pr__nfet_01v8_XGTW7K
Xsky130_fd_pr__nfet_01v8_X8JY7K_1 VSUBS m1_61404_n89284# m2_54836_n91946# m2_54836_n91946#
+ m1_62820_n89278# m1_62468_n89280# m1_68118_n71254# m1_68118_n71254# m2_54836_n91946#
+ m1_64252_n89282# m1_68118_n71254# m1_61242_n89282# m1_68118_n71254# m1_63018_n89282#
+ m1_62298_n89276# m1_63538_n89284# m1_68118_n71254# m2_54836_n91946# m1_61044_n89278#
+ m2_54836_n91946# m1_63192_n89290# m1_62110_n89282# m2_54836_n91946# m1_68118_n71254#
+ m2_54836_n91946# m1_63728_n89284# m1_60882_n89280# m1_63368_n89282# m1_68118_n71254#
+ m1_68118_n71254# m2_54836_n91946# m1_61944_n89280# m1_62662_n89276# m1_63898_n89276#
+ m1_61590_n89288# m2_54836_n91946# m1_68118_n71254# m2_54836_n91946# m2_54836_n91946#
+ m1_68118_n71254# VSUBS m1_61766_n89286# m1_64086_n89280# sky130_fd_pr__nfet_01v8_X8JY7K
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_0 VSUBS vout m3_67376_n80074# sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_1 VSUBS vout m3_67376_n80074# sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_2 VSUBS vout m3_67376_n80074# sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_3 VSUBS vout m3_67376_n80074# sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_4 VSUBS vout m3_67376_n80074# sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__pfet_01v8_VXTQ3X_1 VSUBS m1_52340_n69842# m1_52340_n69842# m1_52340_n69842#
+ m1_52340_n69842# m1_52340_n69842# w_56149_n71520# m1_52340_n69842# m1_52340_n69842#
+ m1_52340_n69842# m1_52340_n69842# m1_52340_n69842# sky130_fd_pr__pfet_01v8_VXTQ3X
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_5 VSUBS vout m3_67376_n80074# sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__pfet_01v8_JXF9S2_0 vin_n vin_n m1_63586_n76008# VSUBS vin_n m1_64296_n76008#
+ vin_n m1_56454_n79854# vin_n vp m1_62178_n74550# vin_n vin_n vp vp vp vin_n vin_n
+ vin_n vin_n vin_n vp vin_n m1_56454_n79854# vp m1_63942_n76006# vin_n m1_62520_n76010#
+ m1_63602_n74546# vin_n m1_56454_n79854# vp vin_n vin_n vin_n m1_61096_n76012# vp
+ vp vin_n m1_56454_n79854# vin_n m1_56454_n79854# vin_n m1_62872_n76012# m1_56454_n79854#
+ vin_n vin_n m1_63958_n74544# vin_n vp m1_60028_n76012# vp vin_n vin_n vin_n m1_56454_n79854#
+ vin_n vin_n vin_n m1_60044_n74550# vin_n m1_61112_n74550# vin_n m1_60742_n76008#
+ m1_56454_n79854# vin_n vin_n vin_n m1_56454_n79854# m1_56454_n79854# m1_56454_n79854#
+ vin_n vin_n vp m1_61802_n76012# vin_n vin_n vp m1_61468_n74548# m1_63230_n76006#
+ vin_n vin_n vin_n m1_56454_n79854# vin_n vin_n vin_n vp vp vp m1_56454_n79854# m1_60380_n76016#
+ vp vin_n vin_n m1_56454_n79854# vin_n vin_n vin_n m1_62162_n76012# m1_62536_n74548#
+ vin_n vin_n m1_61452_n76010# vin_n vin_n vin_n vin_n vp vp vp vp m1_56454_n79854#
+ vin_n m1_62888_n74550# m1_56454_n79854# vin_n vp m1_60396_n74554# m1_63246_n74544#
+ vin_n vp vp vin_n m1_56454_n79854# vin_n vin_n vp vin_n vp vin_n vin_n vp vp m1_56454_n79854#
+ vin_n vp vin_n m1_64312_n74546# vp m1_56454_n79854# vin_n vp vin_n m1_60758_n74546#
+ vp vp vin_n vin_n vp m1_56454_n79854# vp vp vp vin_n vp vin_n vin_n vin_n vin_n
+ vin_n vin_n vin_n vin_n vin_n vp vp vin_n vin_n vp vin_n vp m1_61818_n74550# vin_n
+ vp w_56149_n71520# vin_n vp vin_n vin_n vin_n vin_n vp vp sky130_fd_pr__pfet_01v8_JXF9S2
Xsky130_fd_pr__pfet_01v8_JXF9S2_1 vin_n vin_n m1_63576_n79858# VSUBS vin_n m1_64286_n79858#
+ vin_n m1_56454_n79854# vin_n vp m1_62168_n78400# vin_n vin_n vp vp vp vin_n vin_n
+ vin_n vin_n vin_n vp vin_n m1_56454_n79854# vp m1_63932_n79856# vin_n m1_62510_n79860#
+ m1_63592_n78396# vin_n m1_56454_n79854# vp vin_n vin_n vin_n m1_61086_n79862# vp
+ vp vin_n m1_56454_n79854# vin_n m1_56454_n79854# vin_n m1_62862_n79862# m1_56454_n79854#
+ vin_n vin_n m1_63948_n78394# vin_n vp m1_60018_n79862# vp vin_n vin_n vin_n m1_56454_n79854#
+ vin_n vin_n vin_n m1_60034_n78400# vin_n m1_61102_n78400# vin_n m1_60732_n79858#
+ m1_56454_n79854# vin_n vin_n vin_n m1_56454_n79854# m1_56454_n79854# m1_56454_n79854#
+ vin_n vin_n vp m1_61792_n79862# vin_n vin_n vp m1_61458_n78398# m1_63220_n79856#
+ vin_n vin_n vin_n m1_56454_n79854# vin_n vin_n vin_n vp vp vp m1_56454_n79854# m1_60370_n79866#
+ vp vin_n vin_n m1_56454_n79854# vin_n vin_n vin_n m1_62152_n79862# m1_62526_n78398#
+ vin_n vin_n m1_61442_n79860# vin_n vin_n vin_n vin_n vp vp vp vp m1_56454_n79854#
+ vin_n m1_62878_n78400# m1_56454_n79854# vin_n vp m1_60386_n78404# m1_63236_n78394#
+ vin_n vp vp vin_n m1_56454_n79854# vin_n vin_n vp vin_n vp vin_n vin_n vp vp m1_56454_n79854#
+ vin_n vp vin_n m1_64302_n78396# vp m1_56454_n79854# vin_n vp vin_n m1_60748_n78396#
+ vp vp vin_n vin_n vp m1_56454_n79854# vp vp vp vin_n vp vin_n vin_n vin_n vin_n
+ vin_n vin_n vin_n vin_n vin_n vp vp vin_n vin_n vp vin_n vp m1_61808_n78400# vin_n
+ vp w_56149_n71520# vin_n vp vin_n vin_n vin_n vin_n vp vp sky130_fd_pr__pfet_01v8_JXF9S2
Xsky130_fd_pr__pfet_01v8_JXF9S2_2 vin_p vin_p m1_68118_n71254# VSUBS vin_p m1_68118_n71254#
+ vin_p m1_58976_n82362# vin_p vp m1_68118_n71254# vin_p vin_p vp vp vp vin_p vin_p
+ vin_p vin_p vin_p vp vin_p m1_58620_n82364# vp m1_68118_n71254# vin_p m1_68118_n71254#
+ m1_68118_n71254# vin_p m1_57548_n82362# vp vin_p vin_p vin_p m1_68118_n71254# vp
+ vp vin_p m1_57192_n82370# vin_p m1_57176_n83832# vin_p m1_68118_n71254# m1_56464_n83820#
+ vin_p vin_p m1_68118_n71254# vin_p vp m1_60028_n83828# vp vin_p vin_p vin_p m1_56842_n82358#
+ vin_p vin_p vin_p m1_60044_n82366# vin_p m1_68118_n71254# vin_p m1_60742_n83824#
+ m1_56826_n83820# vin_p vin_p vin_p m1_59672_n83824# m1_58250_n83832# m1_57532_n83824#
+ vin_p vin_p vp m1_68118_n71254# vin_p vin_p vp m1_68118_n71254# m1_68118_n71254#
+ vin_p vin_p vin_p m1_59688_n82362# vin_p vin_p vin_p vp vp vp m1_59334_n82362# m1_60380_n83832#
+ vp vin_p vin_p m1_57890_n83828# vin_p vin_p vin_p m1_68118_n71254# m1_68118_n71254#
+ vin_p vin_p m1_68118_n71254# vin_p vin_p vin_p vin_p vp vp vp vp m1_58266_n82370#
+ vin_p m1_68118_n71254# m1_58960_n83824# vin_p vp m1_60396_n82370# m1_68118_n71254#
+ vin_p vp vp vin_p m1_57906_n82366# vin_p vin_p vp vin_p vp vin_p vin_p vp vp m1_58604_n83826#
+ vin_p vp vin_p m1_68118_n71254# vp m1_59318_n83824# vin_p vp vin_p m1_60758_n82362#
+ vp vp vin_p vin_p vp m1_56480_n82358# vp vp vp vin_p vp vin_p vin_p vin_p vin_p
+ vin_p vin_p vin_p vin_p vin_p vp vp vin_p vin_p vp vin_p vp m1_68118_n71254# vin_p
+ vp w_56149_n71520# vin_p vp vin_p vin_p vin_p vin_p vp vp sky130_fd_pr__pfet_01v8_JXF9S2
Xsky130_fd_pr__pfet_01v8_JXF9S2_3 vin_p vin_p m1_68118_n71254# VSUBS vin_p m1_68118_n71254#
+ vin_p m1_58948_n86182# vin_p vp m1_68118_n71254# vin_p vin_p vp vp vp vin_p vin_p
+ vin_p vin_p vin_p vp vin_p m1_58592_n86184# vp m1_68118_n71254# vin_p m1_68118_n71254#
+ m1_68118_n71254# vin_p m1_57520_n86182# vp vin_p vin_p vin_p m1_68118_n71254# vp
+ vp vin_p m1_57164_n86190# vin_p m1_57148_n87652# vin_p m1_68118_n71254# m1_56436_n87640#
+ vin_p vin_p m1_68118_n71254# vin_p vp m1_60000_n87648# vp vin_p vin_p vin_p m1_56814_n86178#
+ vin_p vin_p vin_p m1_60016_n86186# vin_p m1_68118_n71254# vin_p m1_60714_n87644#
+ m1_56798_n87640# vin_p vin_p vin_p m1_59644_n87644# m1_58222_n87652# m1_57504_n87644#
+ vin_p vin_p vp m1_68118_n71254# vin_p vin_p vp m1_68118_n71254# m1_68118_n71254#
+ vin_p vin_p vin_p m1_59660_n86182# vin_p vin_p vin_p vp vp vp m1_59306_n86182# m1_60352_n87652#
+ vp vin_p vin_p m1_57862_n87648# vin_p vin_p vin_p m1_68118_n71254# m1_68118_n71254#
+ vin_p vin_p m1_68118_n71254# vin_p vin_p vin_p vin_p vp vp vp vp m1_58238_n86190#
+ vin_p m1_68118_n71254# m1_58932_n87644# vin_p vp m1_60368_n86190# m1_68118_n71254#
+ vin_p vp vp vin_p m1_57878_n86186# vin_p vin_p vp vin_p vp vin_p vin_p vp vp m1_58576_n87646#
+ vin_p vp vin_p m1_68118_n71254# vp m1_59290_n87644# vin_p vp vin_p m1_60730_n86182#
+ vp vp vin_p vin_p vp m1_56452_n86178# vp vp vp vin_p vp vin_p vin_p vin_p vin_p
+ vin_p vin_p vin_p vin_p vin_p vp vp vin_p vin_p vp vin_p vp m1_68118_n71254# vin_p
+ vp w_56149_n71520# vin_p vp vin_p vin_p vin_p vin_p vp vp sky130_fd_pr__pfet_01v8_JXF9S2
.end

