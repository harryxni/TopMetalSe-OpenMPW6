magic
tech sky130A
magscale 1 2
timestamp 1608321738
<< nwell >>
rect 748 688 1804 1280
rect 96 470 1804 688
<< pwell >>
rect 564 848 650 886
rect 564 754 650 792
<< nmos >>
rect 96 924 126 1092
rect 238 816 454 846
rect 276 288 306 372
rect 476 288 506 372
rect 676 288 706 372
rect 876 288 906 372
rect 1076 288 1106 372
rect 1276 288 1306 372
rect 1476 132 1506 372
rect 1680 266 1710 374
<< pmos >>
rect 1140 922 1170 1090
rect 1376 1054 1406 1138
rect 786 806 1002 836
rect 276 506 306 590
rect 476 506 506 590
rect 676 506 706 590
rect 876 506 906 590
rect 1076 506 1106 590
rect 1276 506 1306 590
rect 1476 506 1506 986
rect 1680 506 1710 722
<< ndiff >>
rect 38 1047 96 1092
rect 38 1013 50 1047
rect 84 1013 96 1047
rect 38 975 96 1013
rect 38 941 50 975
rect 84 941 96 975
rect 38 924 96 941
rect 126 1046 184 1092
rect 126 1012 138 1046
rect 172 1012 184 1046
rect 126 975 184 1012
rect 126 941 138 975
rect 172 941 184 975
rect 126 924 184 941
rect 238 892 454 904
rect 238 858 254 892
rect 288 858 322 892
rect 356 858 390 892
rect 424 858 454 892
rect 238 846 454 858
rect 238 804 454 816
rect 238 770 246 804
rect 280 770 314 804
rect 348 770 382 804
rect 416 770 454 804
rect 238 758 454 770
rect 218 346 276 372
rect 218 312 230 346
rect 264 312 276 346
rect 218 288 276 312
rect 306 346 364 372
rect 306 312 318 346
rect 352 312 364 346
rect 306 288 364 312
rect 418 346 476 372
rect 418 312 430 346
rect 464 312 476 346
rect 418 288 476 312
rect 506 346 564 372
rect 506 312 518 346
rect 552 312 564 346
rect 506 288 564 312
rect 618 346 676 372
rect 618 312 630 346
rect 664 312 676 346
rect 618 288 676 312
rect 706 346 764 372
rect 706 312 718 346
rect 752 312 764 346
rect 706 288 764 312
rect 818 346 876 372
rect 818 312 830 346
rect 864 312 876 346
rect 818 288 876 312
rect 906 346 964 372
rect 906 312 918 346
rect 952 312 964 346
rect 906 288 964 312
rect 1018 346 1076 372
rect 1018 312 1030 346
rect 1064 312 1076 346
rect 1018 288 1076 312
rect 1106 346 1164 372
rect 1106 312 1118 346
rect 1152 312 1164 346
rect 1106 288 1164 312
rect 1218 346 1276 372
rect 1218 312 1230 346
rect 1264 312 1276 346
rect 1218 288 1276 312
rect 1306 346 1364 372
rect 1306 312 1318 346
rect 1352 312 1364 346
rect 1306 288 1364 312
rect 1418 346 1476 372
rect 1418 312 1430 346
rect 1464 312 1476 346
rect 1418 278 1476 312
rect 1418 244 1430 278
rect 1464 244 1476 278
rect 1418 210 1476 244
rect 1418 176 1430 210
rect 1464 176 1476 210
rect 1418 132 1476 176
rect 1506 346 1564 372
rect 1506 312 1518 346
rect 1552 312 1564 346
rect 1506 278 1564 312
rect 1506 244 1518 278
rect 1552 244 1564 278
rect 1622 334 1680 374
rect 1622 300 1634 334
rect 1668 300 1680 334
rect 1622 266 1680 300
rect 1710 334 1768 374
rect 1710 300 1722 334
rect 1756 300 1768 334
rect 1710 266 1768 300
rect 1506 210 1564 244
rect 1506 176 1518 210
rect 1552 176 1564 210
rect 1506 132 1564 176
<< pdiff >>
rect 1310 1112 1376 1138
rect 1082 1074 1140 1090
rect 1082 1040 1094 1074
rect 1128 1040 1140 1074
rect 1082 1006 1140 1040
rect 1082 972 1094 1006
rect 1128 972 1140 1006
rect 1082 922 1140 972
rect 1170 1082 1228 1090
rect 1170 1048 1182 1082
rect 1216 1048 1228 1082
rect 1310 1078 1326 1112
rect 1360 1078 1376 1112
rect 1310 1054 1376 1078
rect 1406 1112 1472 1138
rect 1406 1078 1422 1112
rect 1456 1078 1472 1112
rect 1406 1054 1472 1078
rect 1170 1014 1228 1048
rect 1170 980 1182 1014
rect 1216 980 1228 1014
rect 1170 922 1228 980
rect 786 882 1002 894
rect 786 848 802 882
rect 836 848 870 882
rect 904 848 938 882
rect 972 848 1002 882
rect 786 836 1002 848
rect 1418 902 1476 986
rect 1418 868 1430 902
rect 1464 868 1476 902
rect 1418 818 1476 868
rect 786 794 1002 806
rect 786 760 802 794
rect 836 760 870 794
rect 904 760 938 794
rect 972 760 1002 794
rect 786 748 1002 760
rect 1418 784 1430 818
rect 1464 784 1476 818
rect 1418 734 1476 784
rect 1418 700 1430 734
rect 1464 700 1476 734
rect 1418 650 1476 700
rect 1418 616 1430 650
rect 1464 616 1476 650
rect 218 566 276 590
rect 218 532 230 566
rect 264 532 276 566
rect 218 506 276 532
rect 306 566 364 590
rect 306 532 318 566
rect 352 532 364 566
rect 306 506 364 532
rect 418 566 476 590
rect 418 532 430 566
rect 464 532 476 566
rect 418 506 476 532
rect 506 566 564 590
rect 506 532 518 566
rect 552 532 564 566
rect 506 506 564 532
rect 618 566 676 590
rect 618 532 630 566
rect 664 532 676 566
rect 618 506 676 532
rect 706 566 764 590
rect 706 532 718 566
rect 752 532 764 566
rect 706 506 764 532
rect 818 566 876 590
rect 818 532 830 566
rect 864 532 876 566
rect 818 506 876 532
rect 906 566 964 590
rect 906 532 918 566
rect 952 532 964 566
rect 906 506 964 532
rect 1018 566 1076 590
rect 1018 532 1030 566
rect 1064 532 1076 566
rect 1018 506 1076 532
rect 1106 566 1164 590
rect 1106 532 1118 566
rect 1152 532 1164 566
rect 1106 506 1164 532
rect 1218 566 1276 590
rect 1218 532 1230 566
rect 1264 532 1276 566
rect 1218 506 1276 532
rect 1306 566 1364 590
rect 1306 532 1318 566
rect 1352 532 1364 566
rect 1306 506 1364 532
rect 1418 566 1476 616
rect 1418 532 1430 566
rect 1464 532 1476 566
rect 1418 506 1476 532
rect 1506 902 1566 986
rect 1506 868 1518 902
rect 1552 868 1566 902
rect 1506 818 1566 868
rect 1506 784 1518 818
rect 1552 784 1566 818
rect 1506 734 1566 784
rect 1506 700 1518 734
rect 1552 700 1566 734
rect 1506 650 1566 700
rect 1506 616 1518 650
rect 1552 616 1566 650
rect 1506 566 1566 616
rect 1506 532 1518 566
rect 1552 532 1566 566
rect 1506 506 1566 532
rect 1622 709 1680 722
rect 1622 675 1634 709
rect 1668 675 1680 709
rect 1622 637 1680 675
rect 1622 603 1634 637
rect 1668 603 1680 637
rect 1622 566 1680 603
rect 1622 532 1634 566
rect 1668 532 1680 566
rect 1622 506 1680 532
rect 1710 696 1768 722
rect 1710 662 1722 696
rect 1756 662 1768 696
rect 1710 625 1768 662
rect 1710 591 1722 625
rect 1756 591 1768 625
rect 1710 553 1768 591
rect 1710 519 1722 553
rect 1756 519 1768 553
rect 1710 506 1768 519
<< ndiffc >>
rect 50 1013 84 1047
rect 50 941 84 975
rect 138 1012 172 1046
rect 138 941 172 975
rect 254 858 288 892
rect 322 858 356 892
rect 390 858 424 892
rect 246 770 280 804
rect 314 770 348 804
rect 382 770 416 804
rect 230 312 264 346
rect 318 312 352 346
rect 430 312 464 346
rect 518 312 552 346
rect 630 312 664 346
rect 718 312 752 346
rect 830 312 864 346
rect 918 312 952 346
rect 1030 312 1064 346
rect 1118 312 1152 346
rect 1230 312 1264 346
rect 1318 312 1352 346
rect 1430 312 1464 346
rect 1430 244 1464 278
rect 1430 176 1464 210
rect 1518 312 1552 346
rect 1518 244 1552 278
rect 1634 300 1668 334
rect 1722 300 1756 334
rect 1518 176 1552 210
<< pdiffc >>
rect 1094 1040 1128 1074
rect 1094 972 1128 1006
rect 1182 1048 1216 1082
rect 1326 1078 1360 1112
rect 1422 1078 1456 1112
rect 1182 980 1216 1014
rect 802 848 836 882
rect 870 848 904 882
rect 938 848 972 882
rect 1430 868 1464 902
rect 802 760 836 794
rect 870 760 904 794
rect 938 760 972 794
rect 1430 784 1464 818
rect 1430 700 1464 734
rect 1430 616 1464 650
rect 230 532 264 566
rect 318 532 352 566
rect 430 532 464 566
rect 518 532 552 566
rect 630 532 664 566
rect 718 532 752 566
rect 830 532 864 566
rect 918 532 952 566
rect 1030 532 1064 566
rect 1118 532 1152 566
rect 1230 532 1264 566
rect 1318 532 1352 566
rect 1430 532 1464 566
rect 1518 868 1552 902
rect 1518 784 1552 818
rect 1518 700 1552 734
rect 1518 616 1552 650
rect 1518 532 1552 566
rect 1634 675 1668 709
rect 1634 603 1668 637
rect 1634 532 1668 566
rect 1722 662 1756 696
rect 1722 591 1756 625
rect 1722 519 1756 553
<< psubdiff >>
rect 564 884 650 886
rect 564 850 590 884
rect 624 850 650 884
rect 564 848 650 850
rect 564 790 650 792
rect 564 756 590 790
rect 624 756 650 790
rect 564 754 650 756
<< nsubdiff >>
rect 816 1210 847 1244
rect 881 1210 942 1244
rect 1008 1210 1039 1244
rect 1073 1210 1104 1244
rect 1200 1210 1231 1244
rect 1265 1210 1296 1244
rect 1392 1210 1423 1244
rect 1457 1210 1488 1244
rect 1584 1210 1615 1244
rect 1649 1210 1680 1244
<< psubdiffcont >>
rect 590 850 624 884
rect 590 756 624 790
<< nsubdiffcont >>
rect 847 1210 881 1244
rect 1039 1210 1073 1244
rect 1231 1210 1265 1244
rect 1423 1210 1457 1244
rect 1615 1210 1649 1244
<< poly >>
rect 96 1092 126 1118
rect 922 1110 1170 1150
rect 1376 1138 1406 1164
rect 922 1090 968 1110
rect 1140 1090 1170 1110
rect 902 1068 968 1090
rect 902 1034 918 1068
rect 952 1034 968 1068
rect 902 1024 968 1034
rect 96 896 126 924
rect 1376 1034 1406 1054
rect 1294 1004 1406 1034
rect 1294 980 1368 1004
rect 1476 986 1506 1012
rect 1294 946 1311 980
rect 1345 946 1368 980
rect 1294 934 1368 946
rect 96 894 164 896
rect 94 874 164 894
rect 94 840 110 874
rect 144 846 164 874
rect 144 840 238 846
rect 94 816 238 840
rect 454 816 480 846
rect 1140 836 1170 922
rect 760 806 786 836
rect 1002 806 1170 836
rect 276 590 306 616
rect 476 590 506 616
rect 676 590 706 616
rect 876 590 906 616
rect 1076 590 1106 616
rect 1276 590 1306 616
rect 1680 722 1710 748
rect 276 490 306 506
rect 476 490 506 506
rect 676 490 706 506
rect 876 490 906 506
rect 1076 490 1106 506
rect 1276 490 1306 506
rect 1476 490 1506 506
rect 262 470 306 490
rect 462 470 506 490
rect 662 470 706 490
rect 862 470 906 490
rect 1062 470 1106 490
rect 1262 470 1306 490
rect 1462 470 1506 490
rect 218 456 306 470
rect 218 422 234 456
rect 268 422 306 456
rect 218 410 306 422
rect 418 456 506 470
rect 418 422 434 456
rect 468 422 506 456
rect 418 410 506 422
rect 618 456 706 470
rect 618 422 634 456
rect 668 422 706 456
rect 618 410 706 422
rect 818 456 906 470
rect 818 422 834 456
rect 868 422 906 456
rect 818 410 906 422
rect 1018 456 1106 470
rect 1018 422 1034 456
rect 1068 422 1106 456
rect 1018 410 1106 422
rect 1218 456 1306 470
rect 1218 422 1234 456
rect 1268 422 1306 456
rect 1218 410 1306 422
rect 1418 456 1506 470
rect 1680 468 1710 506
rect 1418 422 1434 456
rect 1468 422 1506 456
rect 1418 410 1506 422
rect 1620 456 1710 468
rect 1620 422 1636 456
rect 1670 422 1710 456
rect 1620 410 1710 422
rect 262 388 306 410
rect 462 388 506 410
rect 662 388 706 410
rect 862 388 906 410
rect 1062 388 1106 410
rect 1262 388 1306 410
rect 1462 388 1506 410
rect 276 372 306 388
rect 476 372 506 388
rect 676 372 706 388
rect 876 372 906 388
rect 1076 372 1106 388
rect 1276 372 1306 388
rect 1476 372 1506 388
rect 1680 374 1710 410
rect 276 262 306 288
rect 476 262 506 288
rect 676 262 706 288
rect 876 262 906 288
rect 1076 262 1106 288
rect 1276 262 1306 288
rect 1680 240 1710 266
rect 1476 106 1506 132
<< polycont >>
rect 918 1034 952 1068
rect 1311 946 1345 980
rect 110 840 144 874
rect 234 422 268 456
rect 434 422 468 456
rect 634 422 668 456
rect 834 422 868 456
rect 1034 422 1068 456
rect 1234 422 1268 456
rect 1434 422 1468 456
rect 1636 422 1670 456
<< locali >>
rect 0 1210 24 1244
rect 58 1210 160 1244
rect 194 1210 296 1244
rect 330 1210 432 1244
rect 466 1210 568 1244
rect 602 1210 704 1244
rect 738 1210 840 1244
rect 881 1210 976 1244
rect 1010 1210 1039 1244
rect 1073 1210 1112 1244
rect 1146 1210 1231 1244
rect 1282 1210 1384 1244
rect 1418 1210 1423 1244
rect 1457 1210 1520 1244
rect 1554 1210 1615 1244
rect 1649 1210 1656 1244
rect 1690 1210 1804 1244
rect 1292 1112 1360 1210
rect 50 1047 84 1092
rect 50 975 84 1012
rect 50 924 84 941
rect 138 1046 172 1092
rect 1094 1074 1128 1090
rect 860 1068 1094 1072
rect 860 1057 918 1068
rect 860 1023 877 1057
rect 911 1034 918 1057
rect 952 1040 1094 1068
rect 952 1034 1128 1040
rect 911 1023 1128 1034
rect 138 975 674 1012
rect 172 956 674 975
rect 860 1006 1128 1023
rect 860 972 1094 1006
rect 860 968 1128 972
rect 138 924 172 941
rect 278 948 674 956
rect 278 892 418 948
rect 542 898 674 948
rect 1094 922 1128 968
rect 1182 1082 1222 1098
rect 1216 1024 1222 1082
rect 1292 1078 1326 1112
rect 1292 1054 1360 1078
rect 1420 1112 1668 1138
rect 1420 1078 1422 1112
rect 1456 1078 1668 1112
rect 1420 1054 1668 1078
rect 1182 1014 1222 1024
rect 1216 980 1222 1014
rect 14 874 160 878
rect 14 840 110 874
rect 144 840 160 874
rect 238 858 254 892
rect 288 858 322 892
rect 356 858 390 892
rect 424 858 454 892
rect 542 884 676 898
rect 14 838 160 840
rect 542 850 590 884
rect 624 850 676 884
rect 1182 882 1222 980
rect 1292 960 1311 980
rect 1292 926 1310 960
rect 1345 946 1362 980
rect 1344 926 1362 946
rect 1292 912 1362 926
rect 42 770 246 804
rect 280 770 314 804
rect 348 770 382 804
rect 416 770 456 804
rect 542 798 676 850
rect 786 848 802 882
rect 836 848 870 882
rect 904 848 938 882
rect 972 848 1222 882
rect 1430 902 1464 952
rect 1430 818 1464 868
rect 42 754 456 770
rect 544 790 674 798
rect 544 756 590 790
rect 624 756 674 790
rect 786 760 802 794
rect 836 760 870 794
rect 904 760 938 794
rect 972 760 1002 794
rect 1430 766 1464 784
rect 42 254 116 754
rect 544 740 674 756
rect 830 688 948 760
rect 1234 734 1464 766
rect 1234 700 1430 734
rect 1234 688 1464 700
rect 230 650 1464 688
rect 230 624 1430 650
rect 230 566 264 624
rect 230 506 264 532
rect 318 566 352 590
rect 318 456 352 532
rect 430 566 464 624
rect 430 506 464 532
rect 518 566 552 590
rect 518 456 552 532
rect 630 566 664 624
rect 630 506 664 532
rect 718 566 752 590
rect 718 456 752 532
rect 830 566 864 624
rect 830 506 864 532
rect 918 566 952 590
rect 918 456 952 532
rect 1030 566 1064 624
rect 1030 506 1064 532
rect 1118 566 1152 590
rect 1118 456 1152 532
rect 1230 566 1264 624
rect 1230 506 1264 532
rect 1318 566 1352 590
rect 1318 456 1352 532
rect 1430 566 1464 616
rect 1430 506 1464 532
rect 1518 902 1552 952
rect 1518 818 1552 868
rect 1518 734 1552 784
rect 1518 650 1552 700
rect 1518 566 1552 616
rect 1518 468 1552 532
rect 1634 709 1668 1054
rect 1634 637 1668 675
rect 1634 566 1668 603
rect 1634 506 1668 532
rect 1722 696 1756 722
rect 1722 625 1756 662
rect 1722 553 1756 591
rect 1518 456 1686 468
rect 198 422 234 456
rect 268 422 284 456
rect 318 422 434 456
rect 468 422 484 456
rect 518 422 634 456
rect 668 422 684 456
rect 718 422 834 456
rect 868 422 884 456
rect 918 422 1034 456
rect 1068 422 1084 456
rect 1118 422 1234 456
rect 1268 422 1284 456
rect 1318 422 1434 456
rect 1468 422 1484 456
rect 1518 422 1584 456
rect 1618 422 1636 456
rect 1670 422 1686 456
rect 230 346 264 372
rect 230 254 264 312
rect 318 346 352 422
rect 318 288 352 312
rect 430 346 464 372
rect 430 254 464 312
rect 518 346 552 422
rect 518 288 552 312
rect 630 346 664 372
rect 630 254 664 312
rect 718 346 752 422
rect 718 288 752 312
rect 830 346 864 372
rect 830 254 864 312
rect 918 346 952 422
rect 918 288 952 312
rect 1030 346 1064 372
rect 1030 254 1064 312
rect 1118 346 1152 422
rect 1118 288 1152 312
rect 1230 346 1264 372
rect 1230 254 1264 312
rect 1318 346 1352 422
rect 1518 410 1686 422
rect 1722 462 1756 519
rect 1722 416 1804 462
rect 1318 288 1352 312
rect 1430 346 1464 372
rect 1430 278 1464 312
rect 1400 254 1430 266
rect 42 244 1430 254
rect 42 210 1464 244
rect 42 190 1430 210
rect 1400 180 1430 190
rect 1430 154 1464 176
rect 1518 346 1552 410
rect 1518 278 1552 312
rect 1634 334 1668 374
rect 1634 266 1668 300
rect 1722 334 1756 416
rect 1722 266 1756 300
rect 1518 210 1552 244
rect 1518 154 1552 176
rect 0 30 24 64
rect 58 30 160 64
rect 194 30 296 64
rect 330 30 432 64
rect 466 30 568 64
rect 602 30 704 64
rect 738 30 840 64
rect 874 30 976 64
rect 1010 30 1112 64
rect 1146 30 1248 64
rect 1282 30 1384 64
rect 1418 30 1520 64
rect 1554 30 1656 64
rect 1690 30 1804 64
<< viali >>
rect 24 1210 58 1244
rect 160 1210 194 1244
rect 296 1210 330 1244
rect 432 1210 466 1244
rect 568 1210 602 1244
rect 704 1210 738 1244
rect 840 1210 847 1244
rect 847 1210 874 1244
rect 976 1210 1010 1244
rect 1112 1210 1146 1244
rect 1248 1210 1265 1244
rect 1265 1210 1282 1244
rect 1384 1210 1418 1244
rect 1520 1210 1554 1244
rect 1656 1210 1690 1244
rect 50 1013 84 1046
rect 50 1012 84 1013
rect 877 1023 911 1057
rect 1182 1048 1216 1058
rect 1182 1024 1216 1048
rect 1422 1078 1456 1112
rect 590 850 624 884
rect 1310 946 1311 960
rect 1311 946 1344 960
rect 1310 926 1344 946
rect 590 756 624 790
rect 164 422 198 456
rect 1584 422 1618 456
rect 1634 300 1668 334
rect 24 30 58 64
rect 160 30 194 64
rect 296 30 330 64
rect 432 30 466 64
rect 568 30 602 64
rect 704 30 738 64
rect 840 30 874 64
rect 976 30 1010 64
rect 1112 30 1146 64
rect 1248 30 1282 64
rect 1384 30 1418 64
rect 1520 30 1554 64
rect 1656 30 1690 64
<< metal1 >>
rect 0 1244 1804 1280
rect 0 1210 24 1244
rect 58 1210 160 1244
rect 194 1210 296 1244
rect 330 1210 432 1244
rect 466 1210 568 1244
rect 602 1210 704 1244
rect 738 1210 840 1244
rect 874 1210 976 1244
rect 1010 1210 1112 1244
rect 1146 1210 1248 1244
rect 1282 1210 1384 1244
rect 1418 1210 1520 1244
rect 1554 1210 1656 1244
rect 1690 1210 1804 1244
rect 0 1184 1804 1210
rect 1410 1112 1468 1124
rect 1410 1078 1422 1112
rect 1456 1078 1468 1112
rect 38 1057 928 1072
rect 1410 1068 1468 1078
rect 38 1046 877 1057
rect 38 1012 50 1046
rect 84 1023 877 1046
rect 911 1023 928 1057
rect 84 1012 928 1023
rect 1170 1058 1470 1068
rect 1170 1024 1182 1058
rect 1216 1024 1470 1058
rect 1170 1014 1470 1024
rect 38 1000 928 1012
rect 1298 960 1780 976
rect 1298 926 1310 960
rect 1344 926 1780 960
rect 1298 914 1780 926
rect 544 898 674 900
rect 542 884 676 898
rect 542 850 590 884
rect 624 850 676 884
rect 542 790 676 850
rect 542 756 590 790
rect 624 756 676 790
rect 542 690 676 756
rect 10 594 1804 690
rect 152 456 1626 468
rect 152 422 164 456
rect 198 422 1584 456
rect 1618 422 1626 456
rect 152 412 1626 422
rect 152 410 1624 412
rect 1742 346 1782 594
rect 1622 334 1782 346
rect 1622 300 1634 334
rect 1668 300 1782 334
rect 1622 288 1782 300
rect 0 64 1804 96
rect 0 30 24 64
rect 58 30 160 64
rect 194 30 296 64
rect 330 30 432 64
rect 466 30 568 64
rect 602 30 704 64
rect 738 30 840 64
rect 874 30 976 64
rect 1010 30 1112 64
rect 1146 30 1248 64
rect 1282 30 1384 64
rect 1418 30 1520 64
rect 1554 30 1656 64
rect 1690 30 1804 64
rect 0 0 1804 30
<< labels >>
rlabel locali s 14 858 14 858 4 VCtrl
port 1 nsew
rlabel metal1 s 0 48 0 48 4 VDD
port 2 nsew
rlabel metal1 s 0 1232 0 1232 4 VDD
port 2 nsew
rlabel metal1 s 10 642 10 642 4 GND
port 3 nsew
rlabel locali s 1804 438 1804 438 4 Clk_Out
port 4 nsew
rlabel metal1 s 1780 944 1780 944 4 ENb
port 5 nsew
<< end >>
