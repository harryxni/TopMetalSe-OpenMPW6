magic
tech sky130A
magscale 1 2
timestamp 1608330103
<< error_p >>
rect -29 231 29 237
rect -29 197 -17 231
rect -29 191 29 197
<< nwell >>
rect -211 -242 211 369
<< pmos >>
rect -15 -150 15 150
<< pdiff >>
rect -73 138 -15 150
rect -73 -138 -61 138
rect -27 -138 -15 138
rect -73 -150 -15 -138
rect 15 138 73 150
rect 15 -138 27 138
rect 61 -138 73 138
rect 15 -150 73 -138
<< pdiffc >>
rect -61 -138 -27 138
rect 27 -138 61 138
<< nsubdiff >>
rect -120 299 -79 333
rect 79 299 128 333
<< nsubdiffcont >>
rect -79 299 79 333
<< poly >>
rect -33 231 33 247
rect -33 197 -17 231
rect 17 197 33 231
rect -33 181 33 197
rect -15 150 15 181
rect -15 -187 15 -150
<< polycont >>
rect -17 197 17 231
<< locali >>
rect -120 299 -79 333
rect 79 299 128 333
rect -33 197 -17 231
rect 17 197 33 231
rect -61 138 -27 154
rect -61 -154 -27 -138
rect 27 138 61 154
rect 27 -154 61 -138
<< viali >>
rect -17 197 17 231
rect -61 -138 -27 138
rect 27 -138 61 138
<< metal1 >>
rect -29 231 29 237
rect -29 197 -17 231
rect 17 197 29 231
rect -29 191 29 197
rect -67 138 -21 150
rect -67 -138 -61 138
rect -27 -138 -21 138
rect -67 -150 -21 -138
rect 21 138 67 150
rect 21 -138 27 138
rect 61 -138 67 138
rect 21 -150 67 -138
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -158 -316 158 316
string parameters w 1.5 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
