magic
tech sky130A
magscale 1 2
timestamp 1654643737
<< nwell >>
rect 1010 -1030 1930 -510
<< pwell >>
rect 3204 -1074 4856 -764
rect 2334 -1506 2586 -1074
rect 2844 -1486 4856 -1074
rect 2844 -1506 3096 -1486
rect 5204 -1626 6856 -764
<< pmoslvt >>
rect 1280 -960 1480 -760
<< nmoslvt >>
rect 2360 -1410 2560 -1170
rect 2870 -1410 3070 -1170
rect 3230 -1330 4830 -930
rect 5230 -1330 6830 -930
<< ndiff >>
rect 3230 -843 4830 -790
rect 3230 -877 3265 -843
rect 3299 -877 3333 -843
rect 3367 -877 3401 -843
rect 3435 -877 3469 -843
rect 3503 -877 3537 -843
rect 3571 -877 3605 -843
rect 3639 -877 3673 -843
rect 3707 -877 3741 -843
rect 3775 -877 3809 -843
rect 3843 -877 3877 -843
rect 3911 -877 3945 -843
rect 3979 -877 4013 -843
rect 4047 -877 4081 -843
rect 4115 -877 4149 -843
rect 4183 -877 4217 -843
rect 4251 -877 4285 -843
rect 4319 -877 4353 -843
rect 4387 -877 4421 -843
rect 4455 -877 4489 -843
rect 4523 -877 4557 -843
rect 4591 -877 4625 -843
rect 4659 -877 4693 -843
rect 4727 -877 4761 -843
rect 4795 -877 4830 -843
rect 3230 -930 4830 -877
rect 5230 -843 6830 -790
rect 5230 -877 5265 -843
rect 5299 -877 5333 -843
rect 5367 -877 5401 -843
rect 5435 -877 5469 -843
rect 5503 -877 5537 -843
rect 5571 -877 5605 -843
rect 5639 -877 5673 -843
rect 5707 -877 5741 -843
rect 5775 -877 5809 -843
rect 5843 -877 5877 -843
rect 5911 -877 5945 -843
rect 5979 -877 6013 -843
rect 6047 -877 6081 -843
rect 6115 -877 6149 -843
rect 6183 -877 6217 -843
rect 6251 -877 6285 -843
rect 6319 -877 6353 -843
rect 6387 -877 6421 -843
rect 6455 -877 6489 -843
rect 6523 -877 6557 -843
rect 6591 -877 6625 -843
rect 6659 -877 6693 -843
rect 6727 -877 6761 -843
rect 6795 -877 6830 -843
rect 5230 -930 6830 -877
rect 2360 -1113 2560 -1100
rect 2360 -1147 2409 -1113
rect 2443 -1147 2477 -1113
rect 2511 -1147 2560 -1113
rect 2360 -1170 2560 -1147
rect 2870 -1113 3070 -1100
rect 2870 -1147 2919 -1113
rect 2953 -1147 2987 -1113
rect 3021 -1147 3070 -1113
rect 2870 -1170 3070 -1147
rect 3230 -1383 4830 -1330
rect 2360 -1433 2560 -1410
rect 2360 -1467 2409 -1433
rect 2443 -1467 2477 -1433
rect 2511 -1467 2560 -1433
rect 2360 -1480 2560 -1467
rect 2870 -1433 3070 -1410
rect 2870 -1467 2919 -1433
rect 2953 -1467 2987 -1433
rect 3021 -1467 3070 -1433
rect 3230 -1417 3265 -1383
rect 3299 -1417 3333 -1383
rect 3367 -1417 3401 -1383
rect 3435 -1417 3469 -1383
rect 3503 -1417 3537 -1383
rect 3571 -1417 3605 -1383
rect 3639 -1417 3673 -1383
rect 3707 -1417 3741 -1383
rect 3775 -1417 3809 -1383
rect 3843 -1417 3877 -1383
rect 3911 -1417 3945 -1383
rect 3979 -1417 4013 -1383
rect 4047 -1417 4081 -1383
rect 4115 -1417 4149 -1383
rect 4183 -1417 4217 -1383
rect 4251 -1417 4285 -1383
rect 4319 -1417 4353 -1383
rect 4387 -1417 4421 -1383
rect 4455 -1417 4489 -1383
rect 4523 -1417 4557 -1383
rect 4591 -1417 4625 -1383
rect 4659 -1417 4693 -1383
rect 4727 -1417 4761 -1383
rect 4795 -1417 4830 -1383
rect 3230 -1460 4830 -1417
rect 5230 -1383 6830 -1330
rect 5230 -1417 5265 -1383
rect 5299 -1417 5333 -1383
rect 5367 -1417 5401 -1383
rect 5435 -1417 5469 -1383
rect 5503 -1417 5537 -1383
rect 5571 -1417 5605 -1383
rect 5639 -1417 5673 -1383
rect 5707 -1417 5741 -1383
rect 5775 -1417 5809 -1383
rect 5843 -1417 5877 -1383
rect 5911 -1417 5945 -1383
rect 5979 -1417 6013 -1383
rect 6047 -1417 6081 -1383
rect 6115 -1417 6149 -1383
rect 6183 -1417 6217 -1383
rect 6251 -1417 6285 -1383
rect 6319 -1417 6353 -1383
rect 6387 -1417 6421 -1383
rect 6455 -1417 6489 -1383
rect 6523 -1417 6557 -1383
rect 6591 -1417 6625 -1383
rect 6659 -1417 6693 -1383
rect 6727 -1417 6761 -1383
rect 6795 -1417 6830 -1383
rect 5230 -1460 6830 -1417
rect 2870 -1480 3070 -1467
<< pdiff >>
rect 1190 -809 1280 -760
rect 1190 -843 1213 -809
rect 1247 -843 1280 -809
rect 1190 -877 1280 -843
rect 1190 -911 1213 -877
rect 1247 -911 1280 -877
rect 1190 -960 1280 -911
rect 1480 -809 1590 -760
rect 1480 -843 1513 -809
rect 1547 -843 1590 -809
rect 1480 -877 1590 -843
rect 1480 -911 1513 -877
rect 1547 -911 1590 -877
rect 1480 -960 1590 -911
<< ndiffc >>
rect 3265 -877 3299 -843
rect 3333 -877 3367 -843
rect 3401 -877 3435 -843
rect 3469 -877 3503 -843
rect 3537 -877 3571 -843
rect 3605 -877 3639 -843
rect 3673 -877 3707 -843
rect 3741 -877 3775 -843
rect 3809 -877 3843 -843
rect 3877 -877 3911 -843
rect 3945 -877 3979 -843
rect 4013 -877 4047 -843
rect 4081 -877 4115 -843
rect 4149 -877 4183 -843
rect 4217 -877 4251 -843
rect 4285 -877 4319 -843
rect 4353 -877 4387 -843
rect 4421 -877 4455 -843
rect 4489 -877 4523 -843
rect 4557 -877 4591 -843
rect 4625 -877 4659 -843
rect 4693 -877 4727 -843
rect 4761 -877 4795 -843
rect 5265 -877 5299 -843
rect 5333 -877 5367 -843
rect 5401 -877 5435 -843
rect 5469 -877 5503 -843
rect 5537 -877 5571 -843
rect 5605 -877 5639 -843
rect 5673 -877 5707 -843
rect 5741 -877 5775 -843
rect 5809 -877 5843 -843
rect 5877 -877 5911 -843
rect 5945 -877 5979 -843
rect 6013 -877 6047 -843
rect 6081 -877 6115 -843
rect 6149 -877 6183 -843
rect 6217 -877 6251 -843
rect 6285 -877 6319 -843
rect 6353 -877 6387 -843
rect 6421 -877 6455 -843
rect 6489 -877 6523 -843
rect 6557 -877 6591 -843
rect 6625 -877 6659 -843
rect 6693 -877 6727 -843
rect 6761 -877 6795 -843
rect 2409 -1147 2443 -1113
rect 2477 -1147 2511 -1113
rect 2919 -1147 2953 -1113
rect 2987 -1147 3021 -1113
rect 2409 -1467 2443 -1433
rect 2477 -1467 2511 -1433
rect 2919 -1467 2953 -1433
rect 2987 -1467 3021 -1433
rect 3265 -1417 3299 -1383
rect 3333 -1417 3367 -1383
rect 3401 -1417 3435 -1383
rect 3469 -1417 3503 -1383
rect 3537 -1417 3571 -1383
rect 3605 -1417 3639 -1383
rect 3673 -1417 3707 -1383
rect 3741 -1417 3775 -1383
rect 3809 -1417 3843 -1383
rect 3877 -1417 3911 -1383
rect 3945 -1417 3979 -1383
rect 4013 -1417 4047 -1383
rect 4081 -1417 4115 -1383
rect 4149 -1417 4183 -1383
rect 4217 -1417 4251 -1383
rect 4285 -1417 4319 -1383
rect 4353 -1417 4387 -1383
rect 4421 -1417 4455 -1383
rect 4489 -1417 4523 -1383
rect 4557 -1417 4591 -1383
rect 4625 -1417 4659 -1383
rect 4693 -1417 4727 -1383
rect 4761 -1417 4795 -1383
rect 5265 -1417 5299 -1383
rect 5333 -1417 5367 -1383
rect 5401 -1417 5435 -1383
rect 5469 -1417 5503 -1383
rect 5537 -1417 5571 -1383
rect 5605 -1417 5639 -1383
rect 5673 -1417 5707 -1383
rect 5741 -1417 5775 -1383
rect 5809 -1417 5843 -1383
rect 5877 -1417 5911 -1383
rect 5945 -1417 5979 -1383
rect 6013 -1417 6047 -1383
rect 6081 -1417 6115 -1383
rect 6149 -1417 6183 -1383
rect 6217 -1417 6251 -1383
rect 6285 -1417 6319 -1383
rect 6353 -1417 6387 -1383
rect 6421 -1417 6455 -1383
rect 6489 -1417 6523 -1383
rect 6557 -1417 6591 -1383
rect 6625 -1417 6659 -1383
rect 6693 -1417 6727 -1383
rect 6761 -1417 6795 -1383
<< pdiffc >>
rect 1213 -843 1247 -809
rect 1213 -911 1247 -877
rect 1513 -843 1547 -809
rect 1513 -911 1547 -877
<< psubdiff >>
rect 5230 -1518 6830 -1460
rect 5230 -1552 5265 -1518
rect 5299 -1552 5333 -1518
rect 5367 -1552 5401 -1518
rect 5435 -1552 5469 -1518
rect 5503 -1552 5537 -1518
rect 5571 -1552 5605 -1518
rect 5639 -1552 5673 -1518
rect 5707 -1552 5741 -1518
rect 5775 -1552 5809 -1518
rect 5843 -1552 5877 -1518
rect 5911 -1552 5945 -1518
rect 5979 -1552 6013 -1518
rect 6047 -1552 6081 -1518
rect 6115 -1552 6149 -1518
rect 6183 -1552 6217 -1518
rect 6251 -1552 6285 -1518
rect 6319 -1552 6353 -1518
rect 6387 -1552 6421 -1518
rect 6455 -1552 6489 -1518
rect 6523 -1552 6557 -1518
rect 6591 -1552 6625 -1518
rect 6659 -1552 6693 -1518
rect 6727 -1552 6761 -1518
rect 6795 -1552 6830 -1518
rect 5230 -1600 6830 -1552
<< nsubdiff >>
rect 1090 -809 1190 -760
rect 1090 -843 1118 -809
rect 1152 -843 1190 -809
rect 1090 -877 1190 -843
rect 1090 -911 1118 -877
rect 1152 -911 1190 -877
rect 1090 -960 1190 -911
<< psubdiffcont >>
rect 5265 -1552 5299 -1518
rect 5333 -1552 5367 -1518
rect 5401 -1552 5435 -1518
rect 5469 -1552 5503 -1518
rect 5537 -1552 5571 -1518
rect 5605 -1552 5639 -1518
rect 5673 -1552 5707 -1518
rect 5741 -1552 5775 -1518
rect 5809 -1552 5843 -1518
rect 5877 -1552 5911 -1518
rect 5945 -1552 5979 -1518
rect 6013 -1552 6047 -1518
rect 6081 -1552 6115 -1518
rect 6149 -1552 6183 -1518
rect 6217 -1552 6251 -1518
rect 6285 -1552 6319 -1518
rect 6353 -1552 6387 -1518
rect 6421 -1552 6455 -1518
rect 6489 -1552 6523 -1518
rect 6557 -1552 6591 -1518
rect 6625 -1552 6659 -1518
rect 6693 -1552 6727 -1518
rect 6761 -1552 6795 -1518
<< nsubdiffcont >>
rect 1118 -843 1152 -809
rect 1118 -911 1152 -877
<< poly >>
rect 1280 -760 1480 -730
rect 1280 -990 1480 -960
rect 1280 -1063 1360 -990
rect 1280 -1097 1303 -1063
rect 1337 -1097 1360 -1063
rect 1280 -1130 1360 -1097
rect 2330 -1330 2360 -1170
rect 2230 -1353 2360 -1330
rect 2230 -1387 2263 -1353
rect 2297 -1387 2360 -1353
rect 2230 -1410 2360 -1387
rect 2560 -1410 2590 -1170
rect 2840 -1330 2870 -1170
rect 2740 -1353 2870 -1330
rect 2740 -1387 2773 -1353
rect 2807 -1387 2870 -1353
rect 2740 -1410 2870 -1387
rect 3070 -1410 3100 -1170
rect 3200 -1330 3230 -930
rect 4830 -1180 4860 -930
rect 4830 -1204 5020 -1180
rect 4830 -1306 4894 -1204
rect 4996 -1306 5020 -1204
rect 4830 -1330 5020 -1306
rect 5200 -1330 5230 -930
rect 6830 -1180 6860 -930
rect 6830 -1204 7020 -1180
rect 6830 -1306 6894 -1204
rect 6996 -1306 7020 -1204
rect 6830 -1330 7020 -1306
<< polycont >>
rect 1303 -1097 1337 -1063
rect 2263 -1387 2297 -1353
rect 2773 -1387 2807 -1353
rect 4894 -1306 4996 -1204
rect 6894 -1306 6996 -1204
<< locali >>
rect 1090 -622 1190 -600
rect 1090 -656 1123 -622
rect 1157 -656 1190 -622
rect 1090 -694 1190 -656
rect 1090 -728 1123 -694
rect 1157 -728 1190 -694
rect 1090 -770 1190 -728
rect 1090 -809 1280 -770
rect 1090 -843 1118 -809
rect 1152 -843 1213 -809
rect 1247 -843 1280 -809
rect 1090 -877 1280 -843
rect 1090 -911 1118 -877
rect 1152 -911 1213 -877
rect 1247 -911 1280 -877
rect 1090 -950 1280 -911
rect 1480 -809 1580 -770
rect 1480 -843 1513 -809
rect 1547 -843 1580 -809
rect 1480 -877 1580 -843
rect 1480 -911 1513 -877
rect 1547 -911 1580 -877
rect 3230 -838 5150 -790
rect 3230 -872 3257 -838
rect 3291 -843 3329 -838
rect 3363 -843 3401 -838
rect 3435 -843 3473 -838
rect 3507 -843 3545 -838
rect 3579 -843 3617 -838
rect 3651 -843 3689 -838
rect 3723 -843 3761 -838
rect 3795 -843 3833 -838
rect 3867 -843 3905 -838
rect 3939 -843 3977 -838
rect 4011 -843 4049 -838
rect 4083 -843 4121 -838
rect 4155 -843 4193 -838
rect 4227 -843 4265 -838
rect 4299 -843 4337 -838
rect 4371 -843 4409 -838
rect 4443 -843 4481 -838
rect 4515 -843 4553 -838
rect 4587 -843 4625 -838
rect 4659 -843 4697 -838
rect 4731 -843 4769 -838
rect 3299 -872 3329 -843
rect 3230 -877 3265 -872
rect 3299 -877 3333 -872
rect 3367 -877 3401 -843
rect 3435 -877 3469 -843
rect 3507 -872 3537 -843
rect 3579 -872 3605 -843
rect 3651 -872 3673 -843
rect 3723 -872 3741 -843
rect 3795 -872 3809 -843
rect 3867 -872 3877 -843
rect 3939 -872 3945 -843
rect 4011 -872 4013 -843
rect 3503 -877 3537 -872
rect 3571 -877 3605 -872
rect 3639 -877 3673 -872
rect 3707 -877 3741 -872
rect 3775 -877 3809 -872
rect 3843 -877 3877 -872
rect 3911 -877 3945 -872
rect 3979 -877 4013 -872
rect 4047 -872 4049 -843
rect 4115 -872 4121 -843
rect 4183 -872 4193 -843
rect 4251 -872 4265 -843
rect 4319 -872 4337 -843
rect 4387 -872 4409 -843
rect 4455 -872 4481 -843
rect 4523 -872 4553 -843
rect 4047 -877 4081 -872
rect 4115 -877 4149 -872
rect 4183 -877 4217 -872
rect 4251 -877 4285 -872
rect 4319 -877 4353 -872
rect 4387 -877 4421 -872
rect 4455 -877 4489 -872
rect 4523 -877 4557 -872
rect 4591 -877 4625 -843
rect 4659 -877 4693 -843
rect 4731 -872 4761 -843
rect 4803 -872 5150 -838
rect 4727 -877 4761 -872
rect 4795 -877 5150 -872
rect 3230 -910 5150 -877
rect 5230 -838 7150 -790
rect 5230 -872 5257 -838
rect 5291 -843 5329 -838
rect 5363 -843 5401 -838
rect 5435 -843 5473 -838
rect 5507 -843 5545 -838
rect 5579 -843 5617 -838
rect 5651 -843 5689 -838
rect 5723 -843 5761 -838
rect 5795 -843 5833 -838
rect 5867 -843 5905 -838
rect 5939 -843 5977 -838
rect 6011 -843 6049 -838
rect 6083 -843 6121 -838
rect 6155 -843 6193 -838
rect 6227 -843 6265 -838
rect 6299 -843 6337 -838
rect 6371 -843 6409 -838
rect 6443 -843 6481 -838
rect 6515 -843 6553 -838
rect 6587 -843 6625 -838
rect 6659 -843 6697 -838
rect 6731 -843 6769 -838
rect 5299 -872 5329 -843
rect 5230 -877 5265 -872
rect 5299 -877 5333 -872
rect 5367 -877 5401 -843
rect 5435 -877 5469 -843
rect 5507 -872 5537 -843
rect 5579 -872 5605 -843
rect 5651 -872 5673 -843
rect 5723 -872 5741 -843
rect 5795 -872 5809 -843
rect 5867 -872 5877 -843
rect 5939 -872 5945 -843
rect 6011 -872 6013 -843
rect 5503 -877 5537 -872
rect 5571 -877 5605 -872
rect 5639 -877 5673 -872
rect 5707 -877 5741 -872
rect 5775 -877 5809 -872
rect 5843 -877 5877 -872
rect 5911 -877 5945 -872
rect 5979 -877 6013 -872
rect 6047 -872 6049 -843
rect 6115 -872 6121 -843
rect 6183 -872 6193 -843
rect 6251 -872 6265 -843
rect 6319 -872 6337 -843
rect 6387 -872 6409 -843
rect 6455 -872 6481 -843
rect 6523 -872 6553 -843
rect 6047 -877 6081 -872
rect 6115 -877 6149 -872
rect 6183 -877 6217 -872
rect 6251 -877 6285 -872
rect 6319 -877 6353 -872
rect 6387 -877 6421 -872
rect 6455 -877 6489 -872
rect 6523 -877 6557 -872
rect 6591 -877 6625 -843
rect 6659 -877 6693 -843
rect 6731 -872 6761 -843
rect 6803 -872 7150 -838
rect 6727 -877 6761 -872
rect 6795 -877 7150 -872
rect 5230 -910 7150 -877
rect 1480 -950 1580 -911
rect 1500 -1040 1580 -950
rect 1090 -1063 1580 -1040
rect 1090 -1068 1303 -1063
rect 1090 -1102 1138 -1068
rect 1172 -1097 1303 -1068
rect 1337 -1068 1580 -1063
rect 1337 -1097 1472 -1068
rect 1172 -1102 1472 -1097
rect 1506 -1102 1544 -1068
rect 1578 -1102 1580 -1068
rect 1090 -1130 1580 -1102
rect 2250 -1093 2560 -1090
rect 2250 -1127 2407 -1093
rect 2441 -1113 2479 -1093
rect 2250 -1147 2409 -1127
rect 2443 -1147 2477 -1113
rect 2513 -1127 2560 -1093
rect 2511 -1147 2560 -1127
rect 2250 -1150 2560 -1147
rect 2760 -1098 3070 -1090
rect 2760 -1132 2917 -1098
rect 2951 -1113 2989 -1098
rect 2760 -1147 2919 -1132
rect 2953 -1147 2987 -1113
rect 3023 -1132 3070 -1098
rect 3021 -1147 3070 -1132
rect 2760 -1150 3070 -1147
rect 2250 -1330 2310 -1150
rect 2760 -1330 2820 -1150
rect 5040 -1200 5150 -910
rect 7040 -1200 7150 -910
rect 4860 -1204 5150 -1200
rect 4860 -1306 4894 -1204
rect 4996 -1238 5150 -1204
rect 5022 -1272 5060 -1238
rect 5094 -1272 5150 -1238
rect 4996 -1306 5150 -1272
rect 4860 -1310 5150 -1306
rect 6860 -1204 7150 -1200
rect 6860 -1306 6894 -1204
rect 6996 -1238 7150 -1204
rect 7022 -1272 7060 -1238
rect 7094 -1272 7150 -1238
rect 6996 -1306 7150 -1272
rect 6860 -1310 7150 -1306
rect 2180 -1340 2310 -1330
rect 2110 -1353 2310 -1340
rect 2110 -1387 2112 -1353
rect 2146 -1387 2184 -1353
rect 2218 -1387 2263 -1353
rect 2297 -1387 2310 -1353
rect 2110 -1400 2310 -1387
rect 2180 -1410 2310 -1400
rect 2600 -1353 2820 -1330
rect 2600 -1387 2622 -1353
rect 2656 -1387 2694 -1353
rect 2728 -1387 2773 -1353
rect 2807 -1387 2820 -1353
rect 2600 -1410 2820 -1387
rect 3230 -1383 4820 -1330
rect 2250 -1420 2310 -1410
rect 2360 -1433 2560 -1410
rect 2760 -1420 2820 -1410
rect 2360 -1467 2409 -1433
rect 2443 -1467 2477 -1433
rect 2511 -1467 2560 -1433
rect 2360 -1562 2560 -1467
rect 2360 -1668 2371 -1562
rect 2549 -1668 2560 -1562
rect 2360 -1690 2560 -1668
rect 2870 -1433 3070 -1410
rect 2870 -1467 2919 -1433
rect 2953 -1467 2987 -1433
rect 3021 -1467 3070 -1433
rect 2870 -1562 3070 -1467
rect 2870 -1668 2881 -1562
rect 3059 -1668 3070 -1562
rect 2870 -1690 3070 -1668
rect 3230 -1417 3265 -1383
rect 3299 -1417 3333 -1383
rect 3367 -1417 3401 -1383
rect 3435 -1417 3469 -1383
rect 3503 -1417 3537 -1383
rect 3571 -1417 3605 -1383
rect 3639 -1417 3673 -1383
rect 3707 -1417 3741 -1383
rect 3775 -1417 3809 -1383
rect 3843 -1417 3877 -1383
rect 3911 -1417 3945 -1383
rect 3979 -1417 4013 -1383
rect 4047 -1417 4081 -1383
rect 4115 -1417 4149 -1383
rect 4183 -1417 4217 -1383
rect 4251 -1417 4285 -1383
rect 4319 -1417 4353 -1383
rect 4387 -1417 4421 -1383
rect 4455 -1417 4489 -1383
rect 4523 -1417 4557 -1383
rect 4591 -1417 4625 -1383
rect 4659 -1417 4693 -1383
rect 4727 -1417 4761 -1383
rect 4795 -1417 4820 -1383
rect 3230 -1460 4820 -1417
rect 5230 -1383 6820 -1330
rect 5230 -1417 5265 -1383
rect 5299 -1417 5333 -1383
rect 5367 -1417 5401 -1383
rect 5435 -1417 5469 -1383
rect 5503 -1417 5537 -1383
rect 5571 -1417 5605 -1383
rect 5639 -1417 5673 -1383
rect 5707 -1417 5741 -1383
rect 5775 -1417 5809 -1383
rect 5843 -1417 5877 -1383
rect 5911 -1417 5945 -1383
rect 5979 -1417 6013 -1383
rect 6047 -1417 6081 -1383
rect 6115 -1417 6149 -1383
rect 6183 -1417 6217 -1383
rect 6251 -1417 6285 -1383
rect 6319 -1417 6353 -1383
rect 6387 -1417 6421 -1383
rect 6455 -1417 6489 -1383
rect 6523 -1417 6557 -1383
rect 6591 -1417 6625 -1383
rect 6659 -1417 6693 -1383
rect 6727 -1417 6761 -1383
rect 6795 -1417 6820 -1383
rect 3230 -1574 4830 -1460
rect 3230 -1896 3257 -1574
rect 4803 -1896 4830 -1574
rect 3230 -1940 4830 -1896
rect 5230 -1476 6820 -1417
rect 5230 -1518 6830 -1476
rect 5230 -1552 5265 -1518
rect 5299 -1552 5333 -1518
rect 5367 -1552 5401 -1518
rect 5435 -1552 5469 -1518
rect 5503 -1552 5537 -1518
rect 5571 -1552 5605 -1518
rect 5639 -1552 5673 -1518
rect 5707 -1552 5741 -1518
rect 5775 -1552 5809 -1518
rect 5843 -1552 5877 -1518
rect 5911 -1552 5945 -1518
rect 5979 -1552 6013 -1518
rect 6047 -1552 6081 -1518
rect 6115 -1552 6149 -1518
rect 6183 -1552 6217 -1518
rect 6251 -1552 6285 -1518
rect 6319 -1552 6353 -1518
rect 6387 -1552 6421 -1518
rect 6455 -1552 6489 -1518
rect 6523 -1552 6557 -1518
rect 6591 -1552 6625 -1518
rect 6659 -1552 6693 -1518
rect 6727 -1552 6761 -1518
rect 6795 -1552 6830 -1518
rect 5230 -1574 6830 -1552
rect 5230 -1896 5257 -1574
rect 6803 -1896 6830 -1574
rect 5230 -1950 6830 -1896
<< viali >>
rect 1123 -656 1157 -622
rect 1123 -728 1157 -694
rect 3257 -843 3291 -838
rect 3329 -843 3363 -838
rect 3401 -843 3435 -838
rect 3473 -843 3507 -838
rect 3545 -843 3579 -838
rect 3617 -843 3651 -838
rect 3689 -843 3723 -838
rect 3761 -843 3795 -838
rect 3833 -843 3867 -838
rect 3905 -843 3939 -838
rect 3977 -843 4011 -838
rect 4049 -843 4083 -838
rect 4121 -843 4155 -838
rect 4193 -843 4227 -838
rect 4265 -843 4299 -838
rect 4337 -843 4371 -838
rect 4409 -843 4443 -838
rect 4481 -843 4515 -838
rect 4553 -843 4587 -838
rect 4625 -843 4659 -838
rect 4697 -843 4731 -838
rect 4769 -843 4803 -838
rect 3257 -872 3265 -843
rect 3265 -872 3291 -843
rect 3329 -872 3333 -843
rect 3333 -872 3363 -843
rect 3401 -872 3435 -843
rect 3473 -872 3503 -843
rect 3503 -872 3507 -843
rect 3545 -872 3571 -843
rect 3571 -872 3579 -843
rect 3617 -872 3639 -843
rect 3639 -872 3651 -843
rect 3689 -872 3707 -843
rect 3707 -872 3723 -843
rect 3761 -872 3775 -843
rect 3775 -872 3795 -843
rect 3833 -872 3843 -843
rect 3843 -872 3867 -843
rect 3905 -872 3911 -843
rect 3911 -872 3939 -843
rect 3977 -872 3979 -843
rect 3979 -872 4011 -843
rect 4049 -872 4081 -843
rect 4081 -872 4083 -843
rect 4121 -872 4149 -843
rect 4149 -872 4155 -843
rect 4193 -872 4217 -843
rect 4217 -872 4227 -843
rect 4265 -872 4285 -843
rect 4285 -872 4299 -843
rect 4337 -872 4353 -843
rect 4353 -872 4371 -843
rect 4409 -872 4421 -843
rect 4421 -872 4443 -843
rect 4481 -872 4489 -843
rect 4489 -872 4515 -843
rect 4553 -872 4557 -843
rect 4557 -872 4587 -843
rect 4625 -872 4659 -843
rect 4697 -872 4727 -843
rect 4727 -872 4731 -843
rect 4769 -872 4795 -843
rect 4795 -872 4803 -843
rect 5257 -843 5291 -838
rect 5329 -843 5363 -838
rect 5401 -843 5435 -838
rect 5473 -843 5507 -838
rect 5545 -843 5579 -838
rect 5617 -843 5651 -838
rect 5689 -843 5723 -838
rect 5761 -843 5795 -838
rect 5833 -843 5867 -838
rect 5905 -843 5939 -838
rect 5977 -843 6011 -838
rect 6049 -843 6083 -838
rect 6121 -843 6155 -838
rect 6193 -843 6227 -838
rect 6265 -843 6299 -838
rect 6337 -843 6371 -838
rect 6409 -843 6443 -838
rect 6481 -843 6515 -838
rect 6553 -843 6587 -838
rect 6625 -843 6659 -838
rect 6697 -843 6731 -838
rect 6769 -843 6803 -838
rect 5257 -872 5265 -843
rect 5265 -872 5291 -843
rect 5329 -872 5333 -843
rect 5333 -872 5363 -843
rect 5401 -872 5435 -843
rect 5473 -872 5503 -843
rect 5503 -872 5507 -843
rect 5545 -872 5571 -843
rect 5571 -872 5579 -843
rect 5617 -872 5639 -843
rect 5639 -872 5651 -843
rect 5689 -872 5707 -843
rect 5707 -872 5723 -843
rect 5761 -872 5775 -843
rect 5775 -872 5795 -843
rect 5833 -872 5843 -843
rect 5843 -872 5867 -843
rect 5905 -872 5911 -843
rect 5911 -872 5939 -843
rect 5977 -872 5979 -843
rect 5979 -872 6011 -843
rect 6049 -872 6081 -843
rect 6081 -872 6083 -843
rect 6121 -872 6149 -843
rect 6149 -872 6155 -843
rect 6193 -872 6217 -843
rect 6217 -872 6227 -843
rect 6265 -872 6285 -843
rect 6285 -872 6299 -843
rect 6337 -872 6353 -843
rect 6353 -872 6371 -843
rect 6409 -872 6421 -843
rect 6421 -872 6443 -843
rect 6481 -872 6489 -843
rect 6489 -872 6515 -843
rect 6553 -872 6557 -843
rect 6557 -872 6587 -843
rect 6625 -872 6659 -843
rect 6697 -872 6727 -843
rect 6727 -872 6731 -843
rect 6769 -872 6795 -843
rect 6795 -872 6803 -843
rect 1138 -1102 1172 -1068
rect 1472 -1102 1506 -1068
rect 1544 -1102 1578 -1068
rect 2407 -1113 2441 -1093
rect 2479 -1113 2513 -1093
rect 2407 -1127 2409 -1113
rect 2409 -1127 2441 -1113
rect 2479 -1127 2511 -1113
rect 2511 -1127 2513 -1113
rect 2917 -1113 2951 -1098
rect 2989 -1113 3023 -1098
rect 2917 -1132 2919 -1113
rect 2919 -1132 2951 -1113
rect 2989 -1132 3021 -1113
rect 3021 -1132 3023 -1113
rect 4916 -1272 4950 -1238
rect 4988 -1272 4996 -1238
rect 4996 -1272 5022 -1238
rect 5060 -1272 5094 -1238
rect 6916 -1272 6950 -1238
rect 6988 -1272 6996 -1238
rect 6996 -1272 7022 -1238
rect 7060 -1272 7094 -1238
rect 2112 -1387 2146 -1353
rect 2184 -1387 2218 -1353
rect 2622 -1387 2656 -1353
rect 2694 -1387 2728 -1353
rect 2371 -1668 2549 -1562
rect 2881 -1668 3059 -1562
rect 3257 -1896 4803 -1574
rect 5257 -1896 6803 -1574
<< metal1 >>
rect 860 -622 1930 -220
rect 860 -656 1123 -622
rect 1157 -656 1930 -622
rect 860 -694 1930 -656
rect 860 -728 1123 -694
rect 1157 -728 1930 -694
rect 860 -750 1930 -728
rect 2360 -690 2560 -674
rect 2360 -870 2370 -690
rect 2550 -870 2560 -690
rect 820 -1059 1220 -1040
rect 820 -1111 866 -1059
rect 918 -1111 930 -1059
rect 982 -1111 994 -1059
rect 1046 -1111 1058 -1059
rect 1110 -1111 1122 -1059
rect 1174 -1111 1220 -1059
rect 820 -1130 1220 -1111
rect 1450 -1059 1930 -1040
rect 1450 -1111 1467 -1059
rect 1519 -1111 1531 -1059
rect 1583 -1111 1595 -1059
rect 1647 -1111 1659 -1059
rect 1711 -1111 1723 -1059
rect 1775 -1111 1787 -1059
rect 1839 -1111 1851 -1059
rect 1903 -1111 1930 -1059
rect 1450 -1130 1930 -1111
rect 2360 -1093 2560 -870
rect 2360 -1127 2407 -1093
rect 2441 -1127 2479 -1093
rect 2513 -1127 2560 -1093
rect 2360 -1150 2560 -1127
rect 2870 -690 3070 -674
rect 2870 -870 2880 -690
rect 3060 -870 3070 -690
rect 2870 -1098 3070 -870
rect 3230 -824 4830 -790
rect 3230 -838 3268 -824
rect 3320 -838 3332 -824
rect 3230 -872 3257 -838
rect 3320 -872 3329 -838
rect 3230 -876 3268 -872
rect 3320 -876 3332 -872
rect 3384 -876 3396 -824
rect 3448 -876 3460 -824
rect 3512 -876 3524 -824
rect 3576 -838 3588 -824
rect 3640 -838 3652 -824
rect 3704 -838 3716 -824
rect 3768 -838 3780 -824
rect 3832 -838 3844 -824
rect 3896 -838 3908 -824
rect 3579 -872 3588 -838
rect 3651 -872 3652 -838
rect 3832 -872 3833 -838
rect 3896 -872 3905 -838
rect 3576 -876 3588 -872
rect 3640 -876 3652 -872
rect 3704 -876 3716 -872
rect 3768 -876 3780 -872
rect 3832 -876 3844 -872
rect 3896 -876 3908 -872
rect 3960 -876 3972 -824
rect 4024 -876 4036 -824
rect 4088 -876 4100 -824
rect 4152 -838 4164 -824
rect 4216 -838 4228 -824
rect 4280 -838 4292 -824
rect 4344 -838 4356 -824
rect 4408 -838 4420 -824
rect 4472 -838 4484 -824
rect 4155 -872 4164 -838
rect 4227 -872 4228 -838
rect 4408 -872 4409 -838
rect 4472 -872 4481 -838
rect 4152 -876 4164 -872
rect 4216 -876 4228 -872
rect 4280 -876 4292 -872
rect 4344 -876 4356 -872
rect 4408 -876 4420 -872
rect 4472 -876 4484 -872
rect 4536 -876 4548 -824
rect 4600 -876 4612 -824
rect 4664 -876 4676 -824
rect 4728 -838 4740 -824
rect 4792 -838 4830 -824
rect 4731 -872 4740 -838
rect 4803 -872 4830 -838
rect 4728 -876 4740 -872
rect 4792 -876 4830 -872
rect 3230 -910 4830 -876
rect 5230 -824 6830 -790
rect 5230 -838 5268 -824
rect 5320 -838 5332 -824
rect 5230 -872 5257 -838
rect 5320 -872 5329 -838
rect 5230 -876 5268 -872
rect 5320 -876 5332 -872
rect 5384 -876 5396 -824
rect 5448 -876 5460 -824
rect 5512 -876 5524 -824
rect 5576 -838 5588 -824
rect 5640 -838 5652 -824
rect 5704 -838 5716 -824
rect 5768 -838 5780 -824
rect 5832 -838 5844 -824
rect 5896 -838 5908 -824
rect 5579 -872 5588 -838
rect 5651 -872 5652 -838
rect 5832 -872 5833 -838
rect 5896 -872 5905 -838
rect 5576 -876 5588 -872
rect 5640 -876 5652 -872
rect 5704 -876 5716 -872
rect 5768 -876 5780 -872
rect 5832 -876 5844 -872
rect 5896 -876 5908 -872
rect 5960 -876 5972 -824
rect 6024 -876 6036 -824
rect 6088 -876 6100 -824
rect 6152 -838 6164 -824
rect 6216 -838 6228 -824
rect 6280 -838 6292 -824
rect 6344 -838 6356 -824
rect 6408 -838 6420 -824
rect 6472 -838 6484 -824
rect 6155 -872 6164 -838
rect 6227 -872 6228 -838
rect 6408 -872 6409 -838
rect 6472 -872 6481 -838
rect 6152 -876 6164 -872
rect 6216 -876 6228 -872
rect 6280 -876 6292 -872
rect 6344 -876 6356 -872
rect 6408 -876 6420 -872
rect 6472 -876 6484 -872
rect 6536 -876 6548 -824
rect 6600 -876 6612 -824
rect 6664 -876 6676 -824
rect 6728 -838 6740 -824
rect 6792 -838 6830 -824
rect 6731 -872 6740 -838
rect 6803 -872 6830 -838
rect 6728 -876 6740 -872
rect 6792 -876 6830 -872
rect 5230 -910 6830 -876
rect 2870 -1132 2917 -1098
rect 2951 -1132 2989 -1098
rect 3023 -1132 3070 -1098
rect 2870 -1150 3070 -1132
rect 4860 -1229 5150 -1200
rect 4860 -1238 4920 -1229
rect 4860 -1272 4916 -1238
rect 4860 -1281 4920 -1272
rect 4972 -1281 4984 -1229
rect 5036 -1281 5048 -1229
rect 5100 -1281 5150 -1229
rect 4860 -1310 5150 -1281
rect 6860 -1229 7150 -1200
rect 6860 -1238 6920 -1229
rect 6860 -1272 6916 -1238
rect 6860 -1281 6920 -1272
rect 6972 -1281 6984 -1229
rect 7036 -1281 7048 -1229
rect 7100 -1281 7150 -1229
rect 6860 -1310 7150 -1281
rect 2090 -1344 2310 -1330
rect 2090 -1396 2100 -1344
rect 2152 -1396 2164 -1344
rect 2216 -1353 2228 -1344
rect 2218 -1387 2228 -1353
rect 2216 -1396 2228 -1387
rect 2280 -1396 2310 -1344
rect 2090 -1410 2310 -1396
rect 2600 -1344 2820 -1330
rect 2600 -1396 2610 -1344
rect 2662 -1396 2674 -1344
rect 2726 -1353 2738 -1344
rect 2728 -1387 2738 -1353
rect 2726 -1396 2738 -1387
rect 2790 -1396 2820 -1344
rect 2600 -1410 2820 -1396
rect 1530 -1562 7180 -1530
rect 1530 -1668 2371 -1562
rect 2549 -1668 2881 -1562
rect 3059 -1574 7180 -1562
rect 3059 -1668 3257 -1574
rect 1530 -1896 3257 -1668
rect 4803 -1896 5257 -1574
rect 6803 -1896 7180 -1574
rect 1530 -2170 7180 -1896
<< via1 >>
rect 2370 -870 2550 -690
rect 866 -1111 918 -1059
rect 930 -1111 982 -1059
rect 994 -1111 1046 -1059
rect 1058 -1111 1110 -1059
rect 1122 -1068 1174 -1059
rect 1122 -1102 1138 -1068
rect 1138 -1102 1172 -1068
rect 1172 -1102 1174 -1068
rect 1122 -1111 1174 -1102
rect 1467 -1068 1519 -1059
rect 1467 -1102 1472 -1068
rect 1472 -1102 1506 -1068
rect 1506 -1102 1519 -1068
rect 1467 -1111 1519 -1102
rect 1531 -1068 1583 -1059
rect 1531 -1102 1544 -1068
rect 1544 -1102 1578 -1068
rect 1578 -1102 1583 -1068
rect 1531 -1111 1583 -1102
rect 1595 -1111 1647 -1059
rect 1659 -1111 1711 -1059
rect 1723 -1111 1775 -1059
rect 1787 -1111 1839 -1059
rect 1851 -1111 1903 -1059
rect 2880 -870 3060 -690
rect 3268 -838 3320 -824
rect 3332 -838 3384 -824
rect 3268 -872 3291 -838
rect 3291 -872 3320 -838
rect 3332 -872 3363 -838
rect 3363 -872 3384 -838
rect 3268 -876 3320 -872
rect 3332 -876 3384 -872
rect 3396 -838 3448 -824
rect 3396 -872 3401 -838
rect 3401 -872 3435 -838
rect 3435 -872 3448 -838
rect 3396 -876 3448 -872
rect 3460 -838 3512 -824
rect 3460 -872 3473 -838
rect 3473 -872 3507 -838
rect 3507 -872 3512 -838
rect 3460 -876 3512 -872
rect 3524 -838 3576 -824
rect 3588 -838 3640 -824
rect 3652 -838 3704 -824
rect 3716 -838 3768 -824
rect 3780 -838 3832 -824
rect 3844 -838 3896 -824
rect 3908 -838 3960 -824
rect 3524 -872 3545 -838
rect 3545 -872 3576 -838
rect 3588 -872 3617 -838
rect 3617 -872 3640 -838
rect 3652 -872 3689 -838
rect 3689 -872 3704 -838
rect 3716 -872 3723 -838
rect 3723 -872 3761 -838
rect 3761 -872 3768 -838
rect 3780 -872 3795 -838
rect 3795 -872 3832 -838
rect 3844 -872 3867 -838
rect 3867 -872 3896 -838
rect 3908 -872 3939 -838
rect 3939 -872 3960 -838
rect 3524 -876 3576 -872
rect 3588 -876 3640 -872
rect 3652 -876 3704 -872
rect 3716 -876 3768 -872
rect 3780 -876 3832 -872
rect 3844 -876 3896 -872
rect 3908 -876 3960 -872
rect 3972 -838 4024 -824
rect 3972 -872 3977 -838
rect 3977 -872 4011 -838
rect 4011 -872 4024 -838
rect 3972 -876 4024 -872
rect 4036 -838 4088 -824
rect 4036 -872 4049 -838
rect 4049 -872 4083 -838
rect 4083 -872 4088 -838
rect 4036 -876 4088 -872
rect 4100 -838 4152 -824
rect 4164 -838 4216 -824
rect 4228 -838 4280 -824
rect 4292 -838 4344 -824
rect 4356 -838 4408 -824
rect 4420 -838 4472 -824
rect 4484 -838 4536 -824
rect 4100 -872 4121 -838
rect 4121 -872 4152 -838
rect 4164 -872 4193 -838
rect 4193 -872 4216 -838
rect 4228 -872 4265 -838
rect 4265 -872 4280 -838
rect 4292 -872 4299 -838
rect 4299 -872 4337 -838
rect 4337 -872 4344 -838
rect 4356 -872 4371 -838
rect 4371 -872 4408 -838
rect 4420 -872 4443 -838
rect 4443 -872 4472 -838
rect 4484 -872 4515 -838
rect 4515 -872 4536 -838
rect 4100 -876 4152 -872
rect 4164 -876 4216 -872
rect 4228 -876 4280 -872
rect 4292 -876 4344 -872
rect 4356 -876 4408 -872
rect 4420 -876 4472 -872
rect 4484 -876 4536 -872
rect 4548 -838 4600 -824
rect 4548 -872 4553 -838
rect 4553 -872 4587 -838
rect 4587 -872 4600 -838
rect 4548 -876 4600 -872
rect 4612 -838 4664 -824
rect 4612 -872 4625 -838
rect 4625 -872 4659 -838
rect 4659 -872 4664 -838
rect 4612 -876 4664 -872
rect 4676 -838 4728 -824
rect 4740 -838 4792 -824
rect 4676 -872 4697 -838
rect 4697 -872 4728 -838
rect 4740 -872 4769 -838
rect 4769 -872 4792 -838
rect 4676 -876 4728 -872
rect 4740 -876 4792 -872
rect 5268 -838 5320 -824
rect 5332 -838 5384 -824
rect 5268 -872 5291 -838
rect 5291 -872 5320 -838
rect 5332 -872 5363 -838
rect 5363 -872 5384 -838
rect 5268 -876 5320 -872
rect 5332 -876 5384 -872
rect 5396 -838 5448 -824
rect 5396 -872 5401 -838
rect 5401 -872 5435 -838
rect 5435 -872 5448 -838
rect 5396 -876 5448 -872
rect 5460 -838 5512 -824
rect 5460 -872 5473 -838
rect 5473 -872 5507 -838
rect 5507 -872 5512 -838
rect 5460 -876 5512 -872
rect 5524 -838 5576 -824
rect 5588 -838 5640 -824
rect 5652 -838 5704 -824
rect 5716 -838 5768 -824
rect 5780 -838 5832 -824
rect 5844 -838 5896 -824
rect 5908 -838 5960 -824
rect 5524 -872 5545 -838
rect 5545 -872 5576 -838
rect 5588 -872 5617 -838
rect 5617 -872 5640 -838
rect 5652 -872 5689 -838
rect 5689 -872 5704 -838
rect 5716 -872 5723 -838
rect 5723 -872 5761 -838
rect 5761 -872 5768 -838
rect 5780 -872 5795 -838
rect 5795 -872 5832 -838
rect 5844 -872 5867 -838
rect 5867 -872 5896 -838
rect 5908 -872 5939 -838
rect 5939 -872 5960 -838
rect 5524 -876 5576 -872
rect 5588 -876 5640 -872
rect 5652 -876 5704 -872
rect 5716 -876 5768 -872
rect 5780 -876 5832 -872
rect 5844 -876 5896 -872
rect 5908 -876 5960 -872
rect 5972 -838 6024 -824
rect 5972 -872 5977 -838
rect 5977 -872 6011 -838
rect 6011 -872 6024 -838
rect 5972 -876 6024 -872
rect 6036 -838 6088 -824
rect 6036 -872 6049 -838
rect 6049 -872 6083 -838
rect 6083 -872 6088 -838
rect 6036 -876 6088 -872
rect 6100 -838 6152 -824
rect 6164 -838 6216 -824
rect 6228 -838 6280 -824
rect 6292 -838 6344 -824
rect 6356 -838 6408 -824
rect 6420 -838 6472 -824
rect 6484 -838 6536 -824
rect 6100 -872 6121 -838
rect 6121 -872 6152 -838
rect 6164 -872 6193 -838
rect 6193 -872 6216 -838
rect 6228 -872 6265 -838
rect 6265 -872 6280 -838
rect 6292 -872 6299 -838
rect 6299 -872 6337 -838
rect 6337 -872 6344 -838
rect 6356 -872 6371 -838
rect 6371 -872 6408 -838
rect 6420 -872 6443 -838
rect 6443 -872 6472 -838
rect 6484 -872 6515 -838
rect 6515 -872 6536 -838
rect 6100 -876 6152 -872
rect 6164 -876 6216 -872
rect 6228 -876 6280 -872
rect 6292 -876 6344 -872
rect 6356 -876 6408 -872
rect 6420 -876 6472 -872
rect 6484 -876 6536 -872
rect 6548 -838 6600 -824
rect 6548 -872 6553 -838
rect 6553 -872 6587 -838
rect 6587 -872 6600 -838
rect 6548 -876 6600 -872
rect 6612 -838 6664 -824
rect 6612 -872 6625 -838
rect 6625 -872 6659 -838
rect 6659 -872 6664 -838
rect 6612 -876 6664 -872
rect 6676 -838 6728 -824
rect 6740 -838 6792 -824
rect 6676 -872 6697 -838
rect 6697 -872 6728 -838
rect 6740 -872 6769 -838
rect 6769 -872 6792 -838
rect 6676 -876 6728 -872
rect 6740 -876 6792 -872
rect 4920 -1238 4972 -1229
rect 4920 -1272 4950 -1238
rect 4950 -1272 4972 -1238
rect 4920 -1281 4972 -1272
rect 4984 -1238 5036 -1229
rect 4984 -1272 4988 -1238
rect 4988 -1272 5022 -1238
rect 5022 -1272 5036 -1238
rect 4984 -1281 5036 -1272
rect 5048 -1238 5100 -1229
rect 5048 -1272 5060 -1238
rect 5060 -1272 5094 -1238
rect 5094 -1272 5100 -1238
rect 5048 -1281 5100 -1272
rect 6920 -1238 6972 -1229
rect 6920 -1272 6950 -1238
rect 6950 -1272 6972 -1238
rect 6920 -1281 6972 -1272
rect 6984 -1238 7036 -1229
rect 6984 -1272 6988 -1238
rect 6988 -1272 7022 -1238
rect 7022 -1272 7036 -1238
rect 6984 -1281 7036 -1272
rect 7048 -1238 7100 -1229
rect 7048 -1272 7060 -1238
rect 7060 -1272 7094 -1238
rect 7094 -1272 7100 -1238
rect 7048 -1281 7100 -1272
rect 2100 -1353 2152 -1344
rect 2100 -1387 2112 -1353
rect 2112 -1387 2146 -1353
rect 2146 -1387 2152 -1353
rect 2100 -1396 2152 -1387
rect 2164 -1353 2216 -1344
rect 2164 -1387 2184 -1353
rect 2184 -1387 2216 -1353
rect 2164 -1396 2216 -1387
rect 2228 -1396 2280 -1344
rect 2610 -1353 2662 -1344
rect 2610 -1387 2622 -1353
rect 2622 -1387 2656 -1353
rect 2656 -1387 2662 -1353
rect 2610 -1396 2662 -1387
rect 2674 -1353 2726 -1344
rect 2674 -1387 2694 -1353
rect 2694 -1387 2726 -1353
rect 2674 -1396 2726 -1387
rect 2738 -1396 2790 -1344
<< metal2 >>
rect 2350 -690 2570 -670
rect 2350 -870 2370 -690
rect 2550 -870 2570 -690
rect 2350 -890 2570 -870
rect 2860 -690 3080 -670
rect 2860 -870 2880 -690
rect 3060 -870 3080 -690
rect 2860 -890 3080 -870
rect 3230 -822 4830 -790
rect 3230 -824 3282 -822
rect 3338 -824 3362 -822
rect 3418 -824 3442 -822
rect 3498 -824 3522 -822
rect 3578 -824 3602 -822
rect 3658 -824 3682 -822
rect 3738 -824 3762 -822
rect 3818 -824 3842 -822
rect 3898 -824 3922 -822
rect 3978 -824 4002 -822
rect 4058 -824 4082 -822
rect 4138 -824 4162 -822
rect 4218 -824 4242 -822
rect 4298 -824 4322 -822
rect 4378 -824 4402 -822
rect 4458 -824 4482 -822
rect 4538 -824 4562 -822
rect 4618 -824 4642 -822
rect 4698 -824 4722 -822
rect 4778 -824 4830 -822
rect 3230 -876 3268 -824
rect 3512 -876 3522 -824
rect 3578 -876 3588 -824
rect 3832 -876 3842 -824
rect 3898 -876 3908 -824
rect 4152 -876 4162 -824
rect 4218 -876 4228 -824
rect 4472 -876 4482 -824
rect 4538 -876 4548 -824
rect 4792 -876 4830 -824
rect 3230 -878 3282 -876
rect 3338 -878 3362 -876
rect 3418 -878 3442 -876
rect 3498 -878 3522 -876
rect 3578 -878 3602 -876
rect 3658 -878 3682 -876
rect 3738 -878 3762 -876
rect 3818 -878 3842 -876
rect 3898 -878 3922 -876
rect 3978 -878 4002 -876
rect 4058 -878 4082 -876
rect 4138 -878 4162 -876
rect 4218 -878 4242 -876
rect 4298 -878 4322 -876
rect 4378 -878 4402 -876
rect 4458 -878 4482 -876
rect 4538 -878 4562 -876
rect 4618 -878 4642 -876
rect 4698 -878 4722 -876
rect 4778 -878 4830 -876
rect 3230 -910 4830 -878
rect 5230 -822 6830 -790
rect 5230 -824 5282 -822
rect 5338 -824 5362 -822
rect 5418 -824 5442 -822
rect 5498 -824 5522 -822
rect 5578 -824 5602 -822
rect 5658 -824 5682 -822
rect 5738 -824 5762 -822
rect 5818 -824 5842 -822
rect 5898 -824 5922 -822
rect 5978 -824 6002 -822
rect 6058 -824 6082 -822
rect 6138 -824 6162 -822
rect 6218 -824 6242 -822
rect 6298 -824 6322 -822
rect 6378 -824 6402 -822
rect 6458 -824 6482 -822
rect 6538 -824 6562 -822
rect 6618 -824 6642 -822
rect 6698 -824 6722 -822
rect 6778 -824 6830 -822
rect 5230 -876 5268 -824
rect 5512 -876 5522 -824
rect 5578 -876 5588 -824
rect 5832 -876 5842 -824
rect 5898 -876 5908 -824
rect 6152 -876 6162 -824
rect 6218 -876 6228 -824
rect 6472 -876 6482 -824
rect 6538 -876 6548 -824
rect 6792 -876 6830 -824
rect 5230 -878 5282 -876
rect 5338 -878 5362 -876
rect 5418 -878 5442 -876
rect 5498 -878 5522 -876
rect 5578 -878 5602 -876
rect 5658 -878 5682 -876
rect 5738 -878 5762 -876
rect 5818 -878 5842 -876
rect 5898 -878 5922 -876
rect 5978 -878 6002 -876
rect 6058 -878 6082 -876
rect 6138 -878 6162 -876
rect 6218 -878 6242 -876
rect 6298 -878 6322 -876
rect 6378 -878 6402 -876
rect 6458 -878 6482 -876
rect 6538 -878 6562 -876
rect 6618 -878 6642 -876
rect 6698 -878 6722 -876
rect 6778 -878 6830 -876
rect 5230 -910 6830 -878
rect 790 -1059 1220 -1040
rect 790 -1111 866 -1059
rect 918 -1111 930 -1059
rect 982 -1111 994 -1059
rect 1046 -1111 1058 -1059
rect 1110 -1111 1122 -1059
rect 1174 -1111 1220 -1059
rect 790 -1130 1220 -1111
rect 1450 -1057 1930 -1040
rect 1450 -1059 1502 -1057
rect 1558 -1059 1582 -1057
rect 1638 -1059 1662 -1057
rect 1718 -1059 1742 -1057
rect 1798 -1059 1822 -1057
rect 1878 -1059 1930 -1057
rect 1450 -1111 1467 -1059
rect 1647 -1111 1659 -1059
rect 1718 -1111 1723 -1059
rect 1903 -1111 1930 -1059
rect 1450 -1113 1502 -1111
rect 1558 -1113 1582 -1111
rect 1638 -1113 1662 -1111
rect 1718 -1113 1742 -1111
rect 1798 -1113 1822 -1111
rect 1878 -1113 1930 -1111
rect 1450 -1130 1930 -1113
rect 4860 -1229 5150 -1200
rect 4860 -1281 4920 -1229
rect 4972 -1281 4984 -1229
rect 5036 -1281 5048 -1229
rect 5100 -1281 5150 -1229
rect 4860 -1310 5150 -1281
rect 6860 -1229 7150 -1200
rect 6860 -1281 6920 -1229
rect 6972 -1281 6984 -1229
rect 7036 -1281 7048 -1229
rect 7100 -1281 7150 -1229
rect 6860 -1310 7150 -1281
rect 2090 -1344 2310 -1330
rect 2090 -1396 2100 -1344
rect 2152 -1396 2164 -1344
rect 2216 -1396 2228 -1344
rect 2280 -1396 2310 -1344
rect 2090 -1410 2310 -1396
rect 2600 -1344 2820 -1330
rect 2600 -1396 2610 -1344
rect 2662 -1396 2674 -1344
rect 2726 -1396 2738 -1344
rect 2790 -1396 2820 -1344
rect 2600 -1410 2820 -1396
rect 2090 -2235 2180 -1410
rect 2600 -2225 2690 -1410
rect 5040 -2205 5150 -1310
rect 7040 -2205 7150 -1310
<< via2 >>
rect 2392 -848 2528 -712
rect 2902 -848 3038 -712
rect 3282 -824 3338 -822
rect 3362 -824 3418 -822
rect 3442 -824 3498 -822
rect 3522 -824 3578 -822
rect 3602 -824 3658 -822
rect 3682 -824 3738 -822
rect 3762 -824 3818 -822
rect 3842 -824 3898 -822
rect 3922 -824 3978 -822
rect 4002 -824 4058 -822
rect 4082 -824 4138 -822
rect 4162 -824 4218 -822
rect 4242 -824 4298 -822
rect 4322 -824 4378 -822
rect 4402 -824 4458 -822
rect 4482 -824 4538 -822
rect 4562 -824 4618 -822
rect 4642 -824 4698 -822
rect 4722 -824 4778 -822
rect 3282 -876 3320 -824
rect 3320 -876 3332 -824
rect 3332 -876 3338 -824
rect 3362 -876 3384 -824
rect 3384 -876 3396 -824
rect 3396 -876 3418 -824
rect 3442 -876 3448 -824
rect 3448 -876 3460 -824
rect 3460 -876 3498 -824
rect 3522 -876 3524 -824
rect 3524 -876 3576 -824
rect 3576 -876 3578 -824
rect 3602 -876 3640 -824
rect 3640 -876 3652 -824
rect 3652 -876 3658 -824
rect 3682 -876 3704 -824
rect 3704 -876 3716 -824
rect 3716 -876 3738 -824
rect 3762 -876 3768 -824
rect 3768 -876 3780 -824
rect 3780 -876 3818 -824
rect 3842 -876 3844 -824
rect 3844 -876 3896 -824
rect 3896 -876 3898 -824
rect 3922 -876 3960 -824
rect 3960 -876 3972 -824
rect 3972 -876 3978 -824
rect 4002 -876 4024 -824
rect 4024 -876 4036 -824
rect 4036 -876 4058 -824
rect 4082 -876 4088 -824
rect 4088 -876 4100 -824
rect 4100 -876 4138 -824
rect 4162 -876 4164 -824
rect 4164 -876 4216 -824
rect 4216 -876 4218 -824
rect 4242 -876 4280 -824
rect 4280 -876 4292 -824
rect 4292 -876 4298 -824
rect 4322 -876 4344 -824
rect 4344 -876 4356 -824
rect 4356 -876 4378 -824
rect 4402 -876 4408 -824
rect 4408 -876 4420 -824
rect 4420 -876 4458 -824
rect 4482 -876 4484 -824
rect 4484 -876 4536 -824
rect 4536 -876 4538 -824
rect 4562 -876 4600 -824
rect 4600 -876 4612 -824
rect 4612 -876 4618 -824
rect 4642 -876 4664 -824
rect 4664 -876 4676 -824
rect 4676 -876 4698 -824
rect 4722 -876 4728 -824
rect 4728 -876 4740 -824
rect 4740 -876 4778 -824
rect 3282 -878 3338 -876
rect 3362 -878 3418 -876
rect 3442 -878 3498 -876
rect 3522 -878 3578 -876
rect 3602 -878 3658 -876
rect 3682 -878 3738 -876
rect 3762 -878 3818 -876
rect 3842 -878 3898 -876
rect 3922 -878 3978 -876
rect 4002 -878 4058 -876
rect 4082 -878 4138 -876
rect 4162 -878 4218 -876
rect 4242 -878 4298 -876
rect 4322 -878 4378 -876
rect 4402 -878 4458 -876
rect 4482 -878 4538 -876
rect 4562 -878 4618 -876
rect 4642 -878 4698 -876
rect 4722 -878 4778 -876
rect 5282 -824 5338 -822
rect 5362 -824 5418 -822
rect 5442 -824 5498 -822
rect 5522 -824 5578 -822
rect 5602 -824 5658 -822
rect 5682 -824 5738 -822
rect 5762 -824 5818 -822
rect 5842 -824 5898 -822
rect 5922 -824 5978 -822
rect 6002 -824 6058 -822
rect 6082 -824 6138 -822
rect 6162 -824 6218 -822
rect 6242 -824 6298 -822
rect 6322 -824 6378 -822
rect 6402 -824 6458 -822
rect 6482 -824 6538 -822
rect 6562 -824 6618 -822
rect 6642 -824 6698 -822
rect 6722 -824 6778 -822
rect 5282 -876 5320 -824
rect 5320 -876 5332 -824
rect 5332 -876 5338 -824
rect 5362 -876 5384 -824
rect 5384 -876 5396 -824
rect 5396 -876 5418 -824
rect 5442 -876 5448 -824
rect 5448 -876 5460 -824
rect 5460 -876 5498 -824
rect 5522 -876 5524 -824
rect 5524 -876 5576 -824
rect 5576 -876 5578 -824
rect 5602 -876 5640 -824
rect 5640 -876 5652 -824
rect 5652 -876 5658 -824
rect 5682 -876 5704 -824
rect 5704 -876 5716 -824
rect 5716 -876 5738 -824
rect 5762 -876 5768 -824
rect 5768 -876 5780 -824
rect 5780 -876 5818 -824
rect 5842 -876 5844 -824
rect 5844 -876 5896 -824
rect 5896 -876 5898 -824
rect 5922 -876 5960 -824
rect 5960 -876 5972 -824
rect 5972 -876 5978 -824
rect 6002 -876 6024 -824
rect 6024 -876 6036 -824
rect 6036 -876 6058 -824
rect 6082 -876 6088 -824
rect 6088 -876 6100 -824
rect 6100 -876 6138 -824
rect 6162 -876 6164 -824
rect 6164 -876 6216 -824
rect 6216 -876 6218 -824
rect 6242 -876 6280 -824
rect 6280 -876 6292 -824
rect 6292 -876 6298 -824
rect 6322 -876 6344 -824
rect 6344 -876 6356 -824
rect 6356 -876 6378 -824
rect 6402 -876 6408 -824
rect 6408 -876 6420 -824
rect 6420 -876 6458 -824
rect 6482 -876 6484 -824
rect 6484 -876 6536 -824
rect 6536 -876 6538 -824
rect 6562 -876 6600 -824
rect 6600 -876 6612 -824
rect 6612 -876 6618 -824
rect 6642 -876 6664 -824
rect 6664 -876 6676 -824
rect 6676 -876 6698 -824
rect 6722 -876 6728 -824
rect 6728 -876 6740 -824
rect 6740 -876 6778 -824
rect 5282 -878 5338 -876
rect 5362 -878 5418 -876
rect 5442 -878 5498 -876
rect 5522 -878 5578 -876
rect 5602 -878 5658 -876
rect 5682 -878 5738 -876
rect 5762 -878 5818 -876
rect 5842 -878 5898 -876
rect 5922 -878 5978 -876
rect 6002 -878 6058 -876
rect 6082 -878 6138 -876
rect 6162 -878 6218 -876
rect 6242 -878 6298 -876
rect 6322 -878 6378 -876
rect 6402 -878 6458 -876
rect 6482 -878 6538 -876
rect 6562 -878 6618 -876
rect 6642 -878 6698 -876
rect 6722 -878 6778 -876
rect 1502 -1059 1558 -1057
rect 1582 -1059 1638 -1057
rect 1662 -1059 1718 -1057
rect 1742 -1059 1798 -1057
rect 1822 -1059 1878 -1057
rect 1502 -1111 1519 -1059
rect 1519 -1111 1531 -1059
rect 1531 -1111 1558 -1059
rect 1582 -1111 1583 -1059
rect 1583 -1111 1595 -1059
rect 1595 -1111 1638 -1059
rect 1662 -1111 1711 -1059
rect 1711 -1111 1718 -1059
rect 1742 -1111 1775 -1059
rect 1775 -1111 1787 -1059
rect 1787 -1111 1798 -1059
rect 1822 -1111 1839 -1059
rect 1839 -1111 1851 -1059
rect 1851 -1111 1878 -1059
rect 1502 -1113 1558 -1111
rect 1582 -1113 1638 -1111
rect 1662 -1113 1718 -1111
rect 1742 -1113 1798 -1111
rect 1822 -1113 1878 -1111
<< metal3 >>
rect 2360 -670 2560 -370
rect 2870 -670 3070 -370
rect 2350 -712 2570 -670
rect 2350 -848 2392 -712
rect 2528 -848 2570 -712
rect 2350 -890 2570 -848
rect 2860 -712 3080 -670
rect 2860 -848 2902 -712
rect 3038 -848 3080 -712
rect 2860 -890 3080 -848
rect 3230 -822 4830 -680
rect 3230 -878 3282 -822
rect 3338 -878 3362 -822
rect 3418 -878 3442 -822
rect 3498 -878 3522 -822
rect 3578 -878 3602 -822
rect 3658 -878 3682 -822
rect 3738 -878 3762 -822
rect 3818 -878 3842 -822
rect 3898 -878 3922 -822
rect 3978 -878 4002 -822
rect 4058 -878 4082 -822
rect 4138 -878 4162 -822
rect 4218 -878 4242 -822
rect 4298 -878 4322 -822
rect 4378 -878 4402 -822
rect 4458 -878 4482 -822
rect 4538 -878 4562 -822
rect 4618 -878 4642 -822
rect 4698 -878 4722 -822
rect 4778 -878 4830 -822
rect 3230 -910 4830 -878
rect 5230 -822 6830 -680
rect 5230 -878 5282 -822
rect 5338 -878 5362 -822
rect 5418 -878 5442 -822
rect 5498 -878 5522 -822
rect 5578 -878 5602 -822
rect 5658 -878 5682 -822
rect 5738 -878 5762 -822
rect 5818 -878 5842 -822
rect 5898 -878 5922 -822
rect 5978 -878 6002 -822
rect 6058 -878 6082 -822
rect 6138 -878 6162 -822
rect 6218 -878 6242 -822
rect 6298 -878 6322 -822
rect 6378 -878 6402 -822
rect 6458 -878 6482 -822
rect 6538 -878 6562 -822
rect 6618 -878 6642 -822
rect 6698 -878 6722 -822
rect 6778 -878 6830 -822
rect 5230 -910 6830 -878
rect 1450 -1057 1930 -1040
rect 1450 -1113 1502 -1057
rect 1558 -1113 1582 -1057
rect 1638 -1113 1662 -1057
rect 1718 -1113 1742 -1057
rect 1798 -1113 1822 -1057
rect 1878 -1113 1930 -1057
rect 1450 -1130 1930 -1113
rect 1840 -2236 1930 -1130
<< labels >>
rlabel metal1 s 870 -670 870 -670 4 VDD
port 1 nsew
rlabel metal2 s 2130 -1630 2130 -1630 4 NB1
port 2 nsew
rlabel metal2 s 2640 -1630 2640 -1630 4 NB2
port 3 nsew
rlabel metal2 s 5090 -1630 5090 -1630 4 OUT_IB
port 4 nsew
rlabel metal2 s 7100 -1630 7100 -1630 4 AMP_IB
port 5 nsew
rlabel metal1 s 1650 -1540 1650 -1540 4 GND
port 6 nsew
rlabel metal3 s 1840 -2236 1930 -2200 4 SF_IB
port 7 nsew
<< end >>
