magic
tech sky130A
magscale 1 2
timestamp 1654768983
<< metal1 >>
rect 401167 675692 401537 675698
rect 143673 675270 146631 675660
rect 173157 675322 401167 675692
rect 143673 670736 144063 675270
rect 173157 674103 173527 675322
rect 401167 675316 401537 675322
rect 152191 673733 173527 674103
rect 154966 673475 154972 673585
rect 155082 673475 155088 673585
rect 154972 672526 155082 673475
rect 364863 673430 365033 673460
rect 177593 673260 365033 673430
rect 178695 672526 178865 673260
rect 154972 672416 178922 672526
rect 143673 670340 144063 670346
rect 13647 669652 50982 669972
rect 13647 657326 13967 669652
rect 50662 664728 50982 669652
rect 53663 664728 53983 664734
rect 50662 664408 53663 664728
rect 53663 664402 53983 664408
rect 13647 657000 13967 657006
rect 364863 369194 365033 673260
rect 397829 665127 398129 665133
rect 380003 553714 380293 553720
rect 380003 428041 380293 553424
rect 380003 427751 396461 428041
rect 396171 370414 396461 427751
rect 364863 369024 367371 369194
rect 397829 357864 398129 664827
rect 395827 357564 398129 357864
<< via1 >>
rect 401167 675322 401537 675692
rect 154972 673475 155082 673585
rect 143673 670346 144063 670736
rect 53663 664408 53983 664728
rect 13647 657006 13967 657326
rect 397829 664827 398129 665127
rect 380003 553424 380293 553714
<< metal2 >>
rect 178455 689116 178515 689125
rect 145941 689061 178455 689111
rect 69665 676370 69775 676379
rect 46334 676260 69665 676370
rect 46334 669571 46444 676260
rect 69665 676251 69775 676260
rect 145941 674802 145991 689061
rect 178455 689047 178515 689056
rect 401167 675692 401537 675701
rect 401161 675322 401167 675692
rect 401537 675322 401543 675692
rect 401167 675313 401537 675322
rect 145941 674752 146221 674802
rect 147471 671904 147561 673735
rect 55827 671823 147561 671904
rect 55827 671794 147548 671823
rect 55827 671030 55937 671794
rect 147981 671172 148071 673745
rect 150421 673079 150531 673785
rect 152421 673585 152531 673785
rect 154972 673585 155082 673591
rect 231029 673585 231038 673684
rect 152412 673475 152421 673585
rect 152531 673475 154972 673585
rect 155082 673475 155098 673585
rect 155830 673475 231038 673585
rect 152431 673466 152531 673475
rect 154972 673469 155082 673475
rect 155846 673079 155956 673475
rect 231029 673374 231038 673475
rect 231348 673585 231357 673684
rect 231348 673475 241562 673585
rect 231348 673374 231357 673475
rect 150242 672969 155956 673079
rect 56588 671062 148395 671172
rect 147981 671023 148071 671062
rect 143673 670736 144063 670745
rect 143667 670346 143673 670736
rect 144063 670346 144069 670736
rect 143673 670337 144063 670346
rect 397829 665127 398129 665136
rect 397823 664827 397829 665127
rect 398129 664827 398135 665127
rect 397829 664818 398129 664827
rect 53668 664728 53978 664732
rect 53657 664408 53663 664728
rect 53983 664408 53989 664728
rect 53668 664404 53978 664408
rect 13638 657006 13647 657326
rect 13967 657006 13976 657326
rect 358400 639678 358710 639687
rect 358400 639359 358710 639368
rect 380003 553714 380293 553723
rect 379997 553424 380003 553714
rect 380293 553424 380299 553714
rect 380003 553415 380293 553424
rect 361653 363482 362756 363662
rect 362576 362993 362756 363482
rect 362389 362745 368047 362993
rect 365000 358894 365170 358903
rect 365170 358724 368461 358894
rect 365000 358715 365170 358724
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 69665 676260 69775 676370
rect 178455 689056 178515 689116
rect 401167 675322 401537 675692
rect 152421 673475 152531 673585
rect 231038 673374 231348 673684
rect 143673 670346 144063 670736
rect 397829 664827 398129 665127
rect 53668 664413 53978 664723
rect 13647 657006 13967 657326
rect 358400 639368 358710 639678
rect 380003 553424 380293 553714
rect 365000 358724 365170 358894
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 703390 418394 704800
rect 413394 703190 427730 703390
rect 413394 702300 418394 703190
rect 18694 692120 21194 702300
rect 68940 693513 71440 702300
rect 122330 696788 124830 702300
rect 122330 696678 126146 696788
rect 122330 693513 124830 696678
rect 18694 692119 22220 692120
rect 18694 692011 22111 692119
rect 22219 692011 22225 692119
rect 18694 692010 22220 692011
rect 18694 687950 21194 692010
rect -800 682742 1700 685242
rect -800 680242 8830 682742
rect 6330 658270 8830 680242
rect 69665 676375 69775 693513
rect 69660 676370 69780 676375
rect 69660 676260 69665 676370
rect 69775 676260 69780 676370
rect 69660 676255 69780 676260
rect 126036 674594 126146 696678
rect 177230 693513 179730 702300
rect 228438 698529 229478 698530
rect 228433 697491 228439 698529
rect 229477 697491 229483 698529
rect 331191 698285 332129 698286
rect 178455 689121 178515 693513
rect 178450 689116 178520 689121
rect 178450 689056 178455 689116
rect 178515 689056 178520 689116
rect 178450 689051 178520 689056
rect 228438 686295 229478 697491
rect 331186 697349 331192 698285
rect 332128 697349 332134 698285
rect 147741 686095 233572 686295
rect 147741 675242 147941 686095
rect 228438 685734 229478 686095
rect 331191 685196 332129 697349
rect 148251 684996 334616 685196
rect 148251 675274 148451 684996
rect 331191 684805 332129 684996
rect 427530 683959 427730 703190
rect 465394 702300 470394 704800
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 150041 683839 433994 683959
rect 150041 675080 150161 683839
rect 427530 683735 427730 683839
rect 152091 683277 152211 683401
rect 466776 683277 469276 702300
rect 152091 683157 471789 683277
rect 152091 675080 152211 683157
rect 466776 681546 469276 683157
rect 401162 675692 401542 675697
rect 401162 675322 401167 675692
rect 401537 675322 401542 675692
rect 401162 675317 401542 675322
rect 126031 674486 126037 674594
rect 126145 674486 126151 674594
rect 126036 674485 126146 674486
rect 231033 673996 231353 673997
rect 147221 672916 147311 673734
rect 231028 673678 231034 673996
rect 231352 673678 231358 673996
rect 152416 673585 152536 673590
rect 152416 673475 152421 673585
rect 152531 673475 152536 673585
rect 152416 673470 152536 673475
rect 231033 673374 231038 673678
rect 231348 673374 231353 673678
rect 231033 673369 231353 673374
rect 55254 672826 147311 672916
rect 55377 671464 55467 672826
rect 401167 670886 401537 675317
rect 510594 670886 513054 702340
rect 566594 702300 571594 704800
rect 574600 682984 582176 683000
rect 574600 682800 584800 682984
rect 574440 682402 584800 682800
rect 574440 678818 575238 682402
rect 582000 678818 584800 682402
rect 574440 678370 584800 678818
rect 582300 677984 584800 678370
rect 143668 670736 144068 670741
rect 143668 670731 143673 670736
rect 144063 670731 144068 670736
rect 143668 670335 144068 670341
rect 386054 668426 513054 670886
rect 53664 664728 53982 664733
rect 53663 664727 53983 664728
rect 53663 664409 53664 664727
rect 53982 664409 53983 664727
rect 53663 664408 53983 664409
rect 53664 664403 53982 664408
rect 6330 657331 14285 658270
rect 6330 657326 13652 657331
rect 6330 657006 13647 657326
rect 6330 657001 13652 657006
rect 13972 657001 14285 657331
rect 6330 655770 14285 657001
rect -800 643842 1660 648642
rect 386054 640879 388514 668426
rect 397829 665132 398129 668426
rect 397824 665127 398134 665132
rect 397824 664827 397829 665127
rect 398129 664827 398134 665127
rect 397824 664822 398134 664827
rect 582340 642244 584800 644584
rect 372543 640427 388514 640879
rect 358442 639688 388514 640427
rect 558429 639784 584800 642244
rect 358396 639683 388514 639688
rect 358395 639682 388514 639683
rect 358395 639364 358396 639682
rect 358714 639364 388514 639682
rect 358395 639363 388514 639364
rect 358396 639358 388514 639363
rect 358442 638872 388514 639358
rect -800 633842 1660 638642
rect 372543 638419 388514 638872
rect 582340 629784 584800 634584
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 558429 583562 584800 583674
rect -800 559442 1660 564242
rect 582340 555352 584800 555362
rect -800 549442 1660 554242
rect 359769 553719 584800 555352
rect 359769 553429 379998 553719
rect 380298 553429 584800 553719
rect 359769 553424 380003 553429
rect 380293 553424 584800 553429
rect 359769 553237 584800 553424
rect 359769 552919 359907 553237
rect 360225 552919 584800 553237
rect 359769 552892 584800 552919
rect 582340 550562 584800 552892
rect 582340 540562 584800 545362
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 504833 494140 584800 494252
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 504833 449718 584800 449830
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect 24171 420470 24291 426309
rect -800 420358 24407 420470
rect -800 419176 480 419288
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 23023 377248
rect -800 375954 480 376066
rect 22911 357975 23023 377136
rect 24171 359517 24291 420358
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 492062 362420 584800 362532
rect 365000 362221 365170 362227
rect 35309 359517 35429 361429
rect 24171 359397 35429 359517
rect 39253 357975 39373 361409
rect 22911 357863 40458 357975
rect 43333 357427 43453 361455
rect 14606 357307 43453 357427
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect 14606 335208 14726 357307
rect -800 335096 15405 335208
rect 14606 335072 14726 335096
rect -800 333914 480 334026
rect -800 332732 480 332844
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 9839 290804
rect -800 289510 480 289622
rect 9727 289082 9839 290692
rect 47277 289082 47397 361377
rect 365000 358899 365170 362051
rect 364995 358894 365175 358899
rect 361284 358660 363551 358780
rect 364995 358724 365000 358894
rect 365170 358724 365175 358894
rect 364995 358719 365175 358724
rect 363431 355489 363551 358660
rect 492062 355489 492174 362420
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 504833 358874 584800 358986
rect 363431 355369 493623 355489
rect 361279 354716 444537 354836
rect 361369 350636 441316 350756
rect 361381 346692 435926 346812
rect 435806 318609 435926 346692
rect 441196 337264 441316 350636
rect 444417 344507 444537 354716
rect 492062 354703 492174 355369
rect 444417 344387 570754 344507
rect 441196 337144 454512 337264
rect 435806 318489 448006 318609
rect 9482 288962 47397 289082
rect 9727 288921 9839 288962
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 447886 112941 448006 318489
rect 454392 276364 454512 337144
rect 570634 317310 570754 344387
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 570463 317198 584800 317310
rect 570634 315026 570754 317198
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 504833 313652 584800 313764
rect 454392 276244 580683 276364
rect 580563 272888 580683 276244
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 580563 272776 584800 272888
rect 580563 272105 580683 272776
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 504833 269230 584800 269342
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect 447886 112821 571679 112941
rect 571559 92866 571679 112821
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 570398 92754 584800 92866
rect 571559 89505 571679 92754
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 22111 692011 22219 692119
rect 228439 697491 229477 698529
rect 331192 697349 332128 698285
rect 126037 674486 126145 674594
rect 231034 673684 231352 673996
rect 231034 673678 231038 673684
rect 231038 673678 231348 673684
rect 231348 673678 231352 673684
rect 575238 678818 582000 682402
rect 143668 670346 143673 670731
rect 143673 670346 144063 670731
rect 144063 670346 144068 670731
rect 143668 670341 144068 670346
rect 53664 664723 53982 664727
rect 53664 664413 53668 664723
rect 53668 664413 53978 664723
rect 53978 664413 53982 664723
rect 53664 664409 53982 664413
rect 13652 657326 13972 657331
rect 13652 657006 13967 657326
rect 13967 657006 13972 657326
rect 13652 657001 13972 657006
rect 358396 639678 358714 639682
rect 358396 639368 358400 639678
rect 358400 639368 358710 639678
rect 358710 639368 358714 639678
rect 358396 639364 358714 639368
rect 379998 553714 380298 553719
rect 379998 553429 380003 553714
rect 380003 553429 380293 553714
rect 380293 553429 380298 553714
rect 359907 552919 360225 553237
rect 365000 362051 365170 362221
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 703788 334294 704800
rect 329294 702300 329837 703788
rect 329590 700672 329837 702300
rect 333913 702300 334294 703788
rect 333913 700672 334190 702300
rect 329590 700390 334190 700672
rect 229190 699708 231180 699960
rect 229190 698530 229597 699708
rect 228350 698529 229597 698530
rect 228350 697491 228439 698529
rect 229477 697552 229597 698529
rect 229477 697491 231180 697552
rect 228350 697490 231180 697491
rect 229190 697460 231180 697490
rect 331191 698285 332129 700390
rect 331191 697349 331192 698285
rect 332128 697349 332129 698285
rect 331191 697042 332129 697349
rect 22110 692119 31923 692120
rect 22110 692011 22111 692119
rect 22219 692011 31923 692119
rect 22110 692010 31923 692011
rect 13651 657331 13973 657332
rect 13651 657001 13652 657331
rect 13972 657001 13973 657331
rect 13651 657000 13973 657001
rect 31813 358331 31923 692010
rect 574553 682650 577887 682687
rect 574553 682402 582200 682650
rect 574553 678818 575238 682402
rect 582000 678818 582200 682402
rect 574553 678570 582200 678818
rect 46878 674594 126146 674595
rect 46878 674486 126037 674594
rect 126145 674486 126146 674594
rect 46878 674485 126146 674486
rect 46878 670057 46988 674485
rect 231033 673996 231353 673997
rect 231033 673678 231034 673996
rect 231352 673678 231353 673996
rect 231033 673677 231353 673678
rect 143667 670731 144069 670732
rect 143667 670730 143668 670731
rect 144068 670730 144069 670731
rect 408464 665164 409289 666667
rect 574553 665164 577887 678570
rect 53663 664727 53983 664728
rect 53663 664409 53664 664727
rect 53982 664409 53983 664727
rect 53663 664408 53983 664409
rect 408150 661830 577887 665164
rect 358395 639682 358715 639683
rect 358395 639364 358396 639682
rect 358714 639364 358715 639682
rect 358395 639363 358715 639364
rect 379997 553719 380299 553720
rect 379997 553429 379998 553719
rect 380298 553429 380299 553719
rect 379997 553428 380299 553429
rect 359906 553237 360226 553238
rect 359906 552919 359907 553237
rect 360225 552919 360226 553237
rect 359906 552918 360226 552919
rect 408464 367222 409289 661830
rect 395276 366397 409289 367222
rect 31813 358221 50244 358331
<< via4 >>
rect 329837 700672 333913 703788
rect 229597 697552 231180 699708
rect 231057 673701 231329 673973
rect 143667 670341 143668 670730
rect 143668 670341 144068 670730
rect 144068 670341 144069 670730
rect 143667 670340 144069 670341
rect 53687 664432 53959 664704
rect 358419 639387 358691 639659
rect 359930 552942 360202 553214
rect 364925 362221 365245 362296
rect 364925 362051 365000 362221
rect 365000 362051 365170 362221
rect 365170 362051 365245 362221
rect 364925 361976 365245 362051
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 703788 334294 704800
rect 329294 702300 329837 703788
rect 229160 699708 231660 702300
rect 329590 700672 329837 702300
rect 333913 702300 334294 703788
rect 333913 700672 334230 702300
rect 329590 700360 334230 700672
rect 229160 697552 229597 699708
rect 231180 697552 231660 699708
rect 229160 697490 231660 697552
rect 230913 679619 374371 679939
rect 231033 673973 231353 679619
rect 231033 673701 231057 673973
rect 231329 673701 231353 673973
rect 231033 673677 231353 673701
rect 143643 670730 144093 670754
rect 143643 670340 143667 670730
rect 144069 670340 144093 670730
rect 143643 670316 144093 670340
rect 53663 664704 54897 664728
rect 53663 664432 53687 664704
rect 53959 664432 54897 664704
rect 53663 664408 54897 664432
rect 374051 655260 374371 679619
rect 362730 654940 374371 655260
rect 358395 639659 358715 639683
rect 358395 639387 358419 639659
rect 358691 639387 358715 639659
rect 358395 639363 358715 639387
rect 359906 553214 360226 553238
rect 359906 552942 359930 553214
rect 360202 552942 360226 553214
rect 359906 552918 360226 552942
rect 362730 366160 363050 654940
rect 362730 365840 365245 366160
rect 364925 362320 365245 365840
rect 364901 362296 365269 362320
rect 364901 361976 364925 362296
rect 365245 361976 365269 362296
rect 364901 361952 365269 361976
use array_SR  array_SR_0
timestamp 1654762130
transform 1 0 54469 0 1 344190
box -21076 586 311448 327367
use bias  bias_0
timestamp 1654639008
transform 1 0 145381 0 1 675880
box 790 -2236 7180 -220
use opamp_wrapper  opamp_wrapper_0
timestamp 1654750071
transform 1 0 369481 0 1 359134
box -2280 -1640 26995 13665
<< labels >>
flabel metal3 s -800 381864 480 381976 0 FreeSans 1400 0 0 0 gpio_analog[10]
port 2 nsew
flabel metal3 s -800 338642 480 338754 0 FreeSans 1400 0 0 0 gpio_analog[11]
port 3 nsew
flabel metal3 s -800 295420 480 295532 0 FreeSans 1400 0 0 0 gpio_analog[12]
port 4 nsew
flabel metal3 s -800 252398 480 252510 0 FreeSans 1400 0 0 0 gpio_analog[13]
port 5 nsew
flabel metal3 s -800 124776 480 124888 0 FreeSans 1400 0 0 0 gpio_analog[14]
port 6 nsew
flabel metal3 s -800 81554 480 81666 0 FreeSans 1400 0 0 0 gpio_analog[15]
port 7 nsew
flabel metal3 s -800 38332 480 38444 0 FreeSans 1400 0 0 0 gpio_analog[16]
port 8 nsew
flabel metal3 s -800 16910 480 17022 0 FreeSans 1400 0 0 0 gpio_analog[17]
port 9 nsew
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1400 0 0 0 gpio_analog[3]
port 12 nsew
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1400 0 0 0 gpio_analog[4]
port 13 nsew
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1400 0 0 0 gpio_analog[5]
port 14 nsew
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1400 0 0 0 gpio_analog[6]
port 15 nsew
flabel metal3 s -800 511530 480 511642 0 FreeSans 1400 0 0 0 gpio_analog[7]
port 16 nsew
flabel metal3 s -800 468308 480 468420 0 FreeSans 1400 0 0 0 gpio_analog[8]
port 17 nsew
flabel metal3 s -800 425086 480 425198 0 FreeSans 1400 0 0 0 gpio_analog[9]
port 18 nsew
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1400 0 0 0 gpio_noesd[0]
port 19 nsew
flabel metal3 s -800 380682 480 380794 0 FreeSans 1400 0 0 0 gpio_noesd[10]
port 20 nsew
flabel metal3 s -800 337460 480 337572 0 FreeSans 1400 0 0 0 gpio_noesd[11]
port 21 nsew
flabel metal3 s -800 294238 480 294350 0 FreeSans 1400 0 0 0 gpio_noesd[12]
port 22 nsew
flabel metal3 s -800 251216 480 251328 0 FreeSans 1400 0 0 0 gpio_noesd[13]
port 23 nsew
flabel metal3 s -800 123594 480 123706 0 FreeSans 1400 0 0 0 gpio_noesd[14]
port 24 nsew
flabel metal3 s -800 80372 480 80484 0 FreeSans 1400 0 0 0 gpio_noesd[15]
port 25 nsew
flabel metal3 s -800 37150 480 37262 0 FreeSans 1400 0 0 0 gpio_noesd[16]
port 26 nsew
flabel metal3 s -800 15728 480 15840 0 FreeSans 1400 0 0 0 gpio_noesd[17]
port 27 nsew
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1400 0 0 0 gpio_noesd[1]
port 28 nsew
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1400 0 0 0 gpio_noesd[2]
port 29 nsew
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1400 0 0 0 gpio_noesd[3]
port 30 nsew
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1400 0 0 0 gpio_noesd[4]
port 31 nsew
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1400 0 0 0 gpio_noesd[5]
port 32 nsew
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1400 0 0 0 gpio_noesd[6]
port 33 nsew
flabel metal3 s -800 510348 480 510460 0 FreeSans 1400 0 0 0 gpio_noesd[7]
port 34 nsew
flabel metal3 s -800 467126 480 467238 0 FreeSans 1400 0 0 0 gpio_noesd[8]
port 35 nsew
flabel metal3 s -800 423904 480 424016 0 FreeSans 1400 0 0 0 gpio_noesd[9]
port 36 nsew
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1400 0 0 0 io_analog[0]
port 37 nsew
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1400 0 0 0 io_analog[10]
port 38 nsew
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 2400 180 0 0 io_analog[1]
port 39 nsew
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 2400 180 0 0 io_analog[2]
port 40 nsew
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 2400 180 0 0 io_analog[3]
port 41 nsew
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 2400 180 0 0 io_analog[7]
port 45 nsew
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 2400 180 0 0 io_analog[8]
port 46 nsew
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 2400 180 0 0 io_analog[9]
port 47 nsew
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 2400 180 0 0 io_clamp_high[0]
port 48 nsew
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 2400 180 0 0 io_clamp_high[1]
port 49 nsew
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 2400 180 0 0 io_clamp_high[2]
port 50 nsew
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 2400 180 0 0 io_clamp_low[0]
port 51 nsew
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 2400 180 0 0 io_clamp_low[1]
port 52 nsew
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 2400 180 0 0 io_clamp_low[2]
port 53 nsew
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1400 0 0 0 io_in[0]
port 54 nsew
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1400 0 0 0 io_in[10]
port 55 nsew
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1400 0 0 0 io_in[11]
port 56 nsew
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1400 0 0 0 io_in[12]
port 57 nsew
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1400 0 0 0 io_in[13]
port 58 nsew
flabel metal3 s -800 507984 480 508096 0 FreeSans 1400 0 0 0 io_in[14]
port 59 nsew
flabel metal3 s -800 464762 480 464874 0 FreeSans 1400 0 0 0 io_in[15]
port 60 nsew
flabel metal3 s -800 421540 480 421652 0 FreeSans 1400 0 0 0 io_in[16]
port 61 nsew
flabel metal3 s -800 378318 480 378430 0 FreeSans 1400 0 0 0 io_in[17]
port 62 nsew
flabel metal3 s -800 335096 480 335208 0 FreeSans 1400 0 0 0 io_in[18]
port 63 nsew
flabel metal3 s -800 291874 480 291986 0 FreeSans 1400 0 0 0 io_in[19]
port 64 nsew
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1400 0 0 0 io_in[1]
port 65 nsew
flabel metal3 s -800 248852 480 248964 0 FreeSans 1400 0 0 0 io_in[20]
port 66 nsew
flabel metal3 s -800 121230 480 121342 0 FreeSans 1400 0 0 0 io_in[21]
port 67 nsew
flabel metal3 s -800 78008 480 78120 0 FreeSans 1400 0 0 0 io_in[22]
port 68 nsew
flabel metal3 s -800 34786 480 34898 0 FreeSans 1400 0 0 0 io_in[23]
port 69 nsew
flabel metal3 s -800 13364 480 13476 0 FreeSans 1400 0 0 0 io_in[24]
port 70 nsew
flabel metal3 s -800 8636 480 8748 0 FreeSans 1400 0 0 0 io_in[25]
port 71 nsew
flabel metal3 s -800 3908 480 4020 0 FreeSans 1400 0 0 0 io_in[26]
port 72 nsew
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1400 0 0 0 io_in[2]
port 73 nsew
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1400 0 0 0 io_in[3]
port 74 nsew
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1400 0 0 0 io_in[4]
port 75 nsew
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1400 0 0 0 io_in[5]
port 76 nsew
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1400 0 0 0 io_in[6]
port 77 nsew
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1400 0 0 0 io_in[7]
port 78 nsew
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1400 0 0 0 io_in[8]
port 79 nsew
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1400 0 0 0 io_in[9]
port 80 nsew
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1400 0 0 0 io_in_3v3[0]
port 81 nsew
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1400 0 0 0 io_in_3v3[10]
port 82 nsew
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1400 0 0 0 io_in_3v3[11]
port 83 nsew
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1400 0 0 0 io_in_3v3[12]
port 84 nsew
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1400 0 0 0 io_in_3v3[13]
port 85 nsew
flabel metal3 s -800 509166 480 509278 0 FreeSans 1400 0 0 0 io_in_3v3[14]
port 86 nsew
flabel metal3 s -800 465944 480 466056 0 FreeSans 1400 0 0 0 io_in_3v3[15]
port 87 nsew
flabel metal3 s -800 422722 480 422834 0 FreeSans 1400 0 0 0 io_in_3v3[16]
port 88 nsew
flabel metal3 s -800 379500 480 379612 0 FreeSans 1400 0 0 0 io_in_3v3[17]
port 89 nsew
flabel metal3 s -800 336278 480 336390 0 FreeSans 1400 0 0 0 io_in_3v3[18]
port 90 nsew
flabel metal3 s -800 293056 480 293168 0 FreeSans 1400 0 0 0 io_in_3v3[19]
port 91 nsew
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1400 0 0 0 io_in_3v3[1]
port 92 nsew
flabel metal3 s -800 250034 480 250146 0 FreeSans 1400 0 0 0 io_in_3v3[20]
port 93 nsew
flabel metal3 s -800 122412 480 122524 0 FreeSans 1400 0 0 0 io_in_3v3[21]
port 94 nsew
flabel metal3 s -800 79190 480 79302 0 FreeSans 1400 0 0 0 io_in_3v3[22]
port 95 nsew
flabel metal3 s -800 35968 480 36080 0 FreeSans 1400 0 0 0 io_in_3v3[23]
port 96 nsew
flabel metal3 s -800 14546 480 14658 0 FreeSans 1400 0 0 0 io_in_3v3[24]
port 97 nsew
flabel metal3 s -800 9818 480 9930 0 FreeSans 1400 0 0 0 io_in_3v3[25]
port 98 nsew
flabel metal3 s -800 5090 480 5202 0 FreeSans 1400 0 0 0 io_in_3v3[26]
port 99 nsew
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1400 0 0 0 io_in_3v3[2]
port 100 nsew
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1400 0 0 0 io_in_3v3[3]
port 101 nsew
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1400 0 0 0 io_in_3v3[4]
port 102 nsew
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1400 0 0 0 io_in_3v3[5]
port 103 nsew
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1400 0 0 0 io_in_3v3[6]
port 104 nsew
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1400 0 0 0 io_in_3v3[7]
port 105 nsew
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1400 0 0 0 io_in_3v3[8]
port 106 nsew
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1400 0 0 0 io_in_3v3[9]
port 107 nsew
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1400 0 0 0 io_oeb[0]
port 108 nsew
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1400 0 0 0 io_oeb[10]
port 109 nsew
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1400 0 0 0 io_oeb[11]
port 110 nsew
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1400 0 0 0 io_oeb[12]
port 111 nsew
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1400 0 0 0 io_oeb[13]
port 112 nsew
flabel metal3 s -800 505620 480 505732 0 FreeSans 1400 0 0 0 io_oeb[14]
port 113 nsew
flabel metal3 s -800 462398 480 462510 0 FreeSans 1400 0 0 0 io_oeb[15]
port 114 nsew
flabel metal3 s -800 419176 480 419288 0 FreeSans 1400 0 0 0 io_oeb[16]
port 115 nsew
flabel metal3 s -800 375954 480 376066 0 FreeSans 1400 0 0 0 io_oeb[17]
port 116 nsew
flabel metal3 s -800 332732 480 332844 0 FreeSans 1400 0 0 0 io_oeb[18]
port 117 nsew
flabel metal3 s -800 289510 480 289622 0 FreeSans 1400 0 0 0 io_oeb[19]
port 118 nsew
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1400 0 0 0 io_oeb[1]
port 119 nsew
flabel metal3 s -800 246488 480 246600 0 FreeSans 1400 0 0 0 io_oeb[20]
port 120 nsew
flabel metal3 s -800 118866 480 118978 0 FreeSans 1400 0 0 0 io_oeb[21]
port 121 nsew
flabel metal3 s -800 75644 480 75756 0 FreeSans 1400 0 0 0 io_oeb[22]
port 122 nsew
flabel metal3 s -800 32422 480 32534 0 FreeSans 1400 0 0 0 io_oeb[23]
port 123 nsew
flabel metal3 s -800 11000 480 11112 0 FreeSans 1400 0 0 0 io_oeb[24]
port 124 nsew
flabel metal3 s -800 6272 480 6384 0 FreeSans 1400 0 0 0 io_oeb[25]
port 125 nsew
flabel metal3 s -800 1544 480 1656 0 FreeSans 1400 0 0 0 io_oeb[26]
port 126 nsew
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1400 0 0 0 io_oeb[2]
port 127 nsew
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1400 0 0 0 io_oeb[3]
port 128 nsew
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1400 0 0 0 io_oeb[4]
port 129 nsew
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1400 0 0 0 io_oeb[5]
port 130 nsew
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1400 0 0 0 io_oeb[6]
port 131 nsew
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1400 0 0 0 io_oeb[7]
port 132 nsew
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1400 0 0 0 io_oeb[8]
port 133 nsew
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1400 0 0 0 io_oeb[9]
port 134 nsew
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1400 0 0 0 io_out[0]
port 135 nsew
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1400 0 0 0 io_out[10]
port 136 nsew
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1400 0 0 0 io_out[11]
port 137 nsew
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1400 0 0 0 io_out[12]
port 138 nsew
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1400 0 0 0 io_out[13]
port 139 nsew
flabel metal3 s -800 506802 480 506914 0 FreeSans 1400 0 0 0 io_out[14]
port 140 nsew
flabel metal3 s -800 463580 480 463692 0 FreeSans 1400 0 0 0 io_out[15]
port 141 nsew
flabel metal3 s -800 420358 480 420470 0 FreeSans 1400 0 0 0 io_out[16]
port 142 nsew
flabel metal3 s -800 377136 480 377248 0 FreeSans 1400 0 0 0 io_out[17]
port 143 nsew
flabel metal3 s -800 333914 480 334026 0 FreeSans 1400 0 0 0 io_out[18]
port 144 nsew
flabel metal3 s -800 290692 480 290804 0 FreeSans 1400 0 0 0 io_out[19]
port 145 nsew
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1400 0 0 0 io_out[1]
port 146 nsew
flabel metal3 s -800 247670 480 247782 0 FreeSans 1400 0 0 0 io_out[20]
port 147 nsew
flabel metal3 s -800 120048 480 120160 0 FreeSans 1400 0 0 0 io_out[21]
port 148 nsew
flabel metal3 s -800 76826 480 76938 0 FreeSans 1400 0 0 0 io_out[22]
port 149 nsew
flabel metal3 s -800 33604 480 33716 0 FreeSans 1400 0 0 0 io_out[23]
port 150 nsew
flabel metal3 s -800 12182 480 12294 0 FreeSans 1400 0 0 0 io_out[24]
port 151 nsew
flabel metal3 s -800 7454 480 7566 0 FreeSans 1400 0 0 0 io_out[25]
port 152 nsew
flabel metal3 s -800 2726 480 2838 0 FreeSans 1400 0 0 0 io_out[26]
port 153 nsew
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1400 0 0 0 io_out[2]
port 154 nsew
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1400 0 0 0 io_out[3]
port 155 nsew
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1400 0 0 0 io_out[4]
port 156 nsew
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1400 0 0 0 io_out[5]
port 157 nsew
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1400 0 0 0 io_out[6]
port 158 nsew
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1400 0 0 0 io_out[7]
port 159 nsew
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1400 0 0 0 io_out[8]
port 160 nsew
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1400 0 0 0 io_out[9]
port 161 nsew
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1400 90 0 0 la_data_in[0]
port 162 nsew
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1400 90 0 0 la_data_in[100]
port 163 nsew
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1400 90 0 0 la_data_in[101]
port 164 nsew
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1400 90 0 0 la_data_in[102]
port 165 nsew
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1400 90 0 0 la_data_in[103]
port 166 nsew
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1400 90 0 0 la_data_in[104]
port 167 nsew
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1400 90 0 0 la_data_in[105]
port 168 nsew
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1400 90 0 0 la_data_in[106]
port 169 nsew
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1400 90 0 0 la_data_in[107]
port 170 nsew
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1400 90 0 0 la_data_in[108]
port 171 nsew
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1400 90 0 0 la_data_in[109]
port 172 nsew
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1400 90 0 0 la_data_in[10]
port 173 nsew
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1400 90 0 0 la_data_in[110]
port 174 nsew
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1400 90 0 0 la_data_in[111]
port 175 nsew
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1400 90 0 0 la_data_in[112]
port 176 nsew
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1400 90 0 0 la_data_in[113]
port 177 nsew
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1400 90 0 0 la_data_in[114]
port 178 nsew
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1400 90 0 0 la_data_in[115]
port 179 nsew
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1400 90 0 0 la_data_in[116]
port 180 nsew
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1400 90 0 0 la_data_in[117]
port 181 nsew
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1400 90 0 0 la_data_in[118]
port 182 nsew
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1400 90 0 0 la_data_in[119]
port 183 nsew
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1400 90 0 0 la_data_in[11]
port 184 nsew
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1400 90 0 0 la_data_in[120]
port 185 nsew
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1400 90 0 0 la_data_in[121]
port 186 nsew
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1400 90 0 0 la_data_in[122]
port 187 nsew
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1400 90 0 0 la_data_in[123]
port 188 nsew
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1400 90 0 0 la_data_in[124]
port 189 nsew
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1400 90 0 0 la_data_in[125]
port 190 nsew
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1400 90 0 0 la_data_in[126]
port 191 nsew
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1400 90 0 0 la_data_in[127]
port 192 nsew
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1400 90 0 0 la_data_in[12]
port 193 nsew
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1400 90 0 0 la_data_in[13]
port 194 nsew
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1400 90 0 0 la_data_in[14]
port 195 nsew
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1400 90 0 0 la_data_in[15]
port 196 nsew
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1400 90 0 0 la_data_in[16]
port 197 nsew
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1400 90 0 0 la_data_in[17]
port 198 nsew
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1400 90 0 0 la_data_in[18]
port 199 nsew
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1400 90 0 0 la_data_in[19]
port 200 nsew
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1400 90 0 0 la_data_in[1]
port 201 nsew
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1400 90 0 0 la_data_in[20]
port 202 nsew
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1400 90 0 0 la_data_in[21]
port 203 nsew
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1400 90 0 0 la_data_in[22]
port 204 nsew
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1400 90 0 0 la_data_in[23]
port 205 nsew
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1400 90 0 0 la_data_in[24]
port 206 nsew
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1400 90 0 0 la_data_in[25]
port 207 nsew
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1400 90 0 0 la_data_in[26]
port 208 nsew
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1400 90 0 0 la_data_in[27]
port 209 nsew
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1400 90 0 0 la_data_in[28]
port 210 nsew
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1400 90 0 0 la_data_in[29]
port 211 nsew
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1400 90 0 0 la_data_in[2]
port 212 nsew
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1400 90 0 0 la_data_in[30]
port 213 nsew
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1400 90 0 0 la_data_in[31]
port 214 nsew
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1400 90 0 0 la_data_in[32]
port 215 nsew
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1400 90 0 0 la_data_in[33]
port 216 nsew
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1400 90 0 0 la_data_in[34]
port 217 nsew
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1400 90 0 0 la_data_in[35]
port 218 nsew
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1400 90 0 0 la_data_in[36]
port 219 nsew
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1400 90 0 0 la_data_in[37]
port 220 nsew
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1400 90 0 0 la_data_in[38]
port 221 nsew
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1400 90 0 0 la_data_in[39]
port 222 nsew
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1400 90 0 0 la_data_in[3]
port 223 nsew
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1400 90 0 0 la_data_in[40]
port 224 nsew
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1400 90 0 0 la_data_in[41]
port 225 nsew
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1400 90 0 0 la_data_in[42]
port 226 nsew
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1400 90 0 0 la_data_in[43]
port 227 nsew
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1400 90 0 0 la_data_in[44]
port 228 nsew
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1400 90 0 0 la_data_in[45]
port 229 nsew
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1400 90 0 0 la_data_in[46]
port 230 nsew
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1400 90 0 0 la_data_in[47]
port 231 nsew
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1400 90 0 0 la_data_in[48]
port 232 nsew
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1400 90 0 0 la_data_in[49]
port 233 nsew
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1400 90 0 0 la_data_in[4]
port 234 nsew
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1400 90 0 0 la_data_in[50]
port 235 nsew
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1400 90 0 0 la_data_in[51]
port 236 nsew
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1400 90 0 0 la_data_in[52]
port 237 nsew
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1400 90 0 0 la_data_in[53]
port 238 nsew
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1400 90 0 0 la_data_in[54]
port 239 nsew
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1400 90 0 0 la_data_in[55]
port 240 nsew
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1400 90 0 0 la_data_in[56]
port 241 nsew
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1400 90 0 0 la_data_in[57]
port 242 nsew
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1400 90 0 0 la_data_in[58]
port 243 nsew
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1400 90 0 0 la_data_in[59]
port 244 nsew
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1400 90 0 0 la_data_in[5]
port 245 nsew
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1400 90 0 0 la_data_in[60]
port 246 nsew
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1400 90 0 0 la_data_in[61]
port 247 nsew
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1400 90 0 0 la_data_in[62]
port 248 nsew
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1400 90 0 0 la_data_in[63]
port 249 nsew
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1400 90 0 0 la_data_in[64]
port 250 nsew
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1400 90 0 0 la_data_in[65]
port 251 nsew
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1400 90 0 0 la_data_in[66]
port 252 nsew
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1400 90 0 0 la_data_in[67]
port 253 nsew
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1400 90 0 0 la_data_in[68]
port 254 nsew
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1400 90 0 0 la_data_in[69]
port 255 nsew
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1400 90 0 0 la_data_in[6]
port 256 nsew
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1400 90 0 0 la_data_in[70]
port 257 nsew
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1400 90 0 0 la_data_in[71]
port 258 nsew
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1400 90 0 0 la_data_in[72]
port 259 nsew
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1400 90 0 0 la_data_in[73]
port 260 nsew
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1400 90 0 0 la_data_in[74]
port 261 nsew
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1400 90 0 0 la_data_in[75]
port 262 nsew
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1400 90 0 0 la_data_in[76]
port 263 nsew
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1400 90 0 0 la_data_in[77]
port 264 nsew
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1400 90 0 0 la_data_in[78]
port 265 nsew
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1400 90 0 0 la_data_in[79]
port 266 nsew
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1400 90 0 0 la_data_in[7]
port 267 nsew
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1400 90 0 0 la_data_in[80]
port 268 nsew
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1400 90 0 0 la_data_in[81]
port 269 nsew
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1400 90 0 0 la_data_in[82]
port 270 nsew
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1400 90 0 0 la_data_in[83]
port 271 nsew
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1400 90 0 0 la_data_in[84]
port 272 nsew
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1400 90 0 0 la_data_in[85]
port 273 nsew
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1400 90 0 0 la_data_in[86]
port 274 nsew
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1400 90 0 0 la_data_in[87]
port 275 nsew
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1400 90 0 0 la_data_in[88]
port 276 nsew
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1400 90 0 0 la_data_in[89]
port 277 nsew
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1400 90 0 0 la_data_in[8]
port 278 nsew
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1400 90 0 0 la_data_in[90]
port 279 nsew
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1400 90 0 0 la_data_in[91]
port 280 nsew
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1400 90 0 0 la_data_in[92]
port 281 nsew
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1400 90 0 0 la_data_in[93]
port 282 nsew
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1400 90 0 0 la_data_in[94]
port 283 nsew
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1400 90 0 0 la_data_in[95]
port 284 nsew
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1400 90 0 0 la_data_in[96]
port 285 nsew
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1400 90 0 0 la_data_in[97]
port 286 nsew
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1400 90 0 0 la_data_in[98]
port 287 nsew
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1400 90 0 0 la_data_in[99]
port 288 nsew
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1400 90 0 0 la_data_in[9]
port 289 nsew
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1400 90 0 0 la_data_out[0]
port 290 nsew
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1400 90 0 0 la_data_out[100]
port 291 nsew
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1400 90 0 0 la_data_out[101]
port 292 nsew
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1400 90 0 0 la_data_out[102]
port 293 nsew
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1400 90 0 0 la_data_out[103]
port 294 nsew
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1400 90 0 0 la_data_out[104]
port 295 nsew
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1400 90 0 0 la_data_out[105]
port 296 nsew
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1400 90 0 0 la_data_out[106]
port 297 nsew
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1400 90 0 0 la_data_out[107]
port 298 nsew
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1400 90 0 0 la_data_out[108]
port 299 nsew
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1400 90 0 0 la_data_out[109]
port 300 nsew
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1400 90 0 0 la_data_out[10]
port 301 nsew
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1400 90 0 0 la_data_out[110]
port 302 nsew
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1400 90 0 0 la_data_out[111]
port 303 nsew
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1400 90 0 0 la_data_out[112]
port 304 nsew
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1400 90 0 0 la_data_out[113]
port 305 nsew
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1400 90 0 0 la_data_out[114]
port 306 nsew
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1400 90 0 0 la_data_out[115]
port 307 nsew
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1400 90 0 0 la_data_out[116]
port 308 nsew
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1400 90 0 0 la_data_out[117]
port 309 nsew
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1400 90 0 0 la_data_out[118]
port 310 nsew
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1400 90 0 0 la_data_out[119]
port 311 nsew
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1400 90 0 0 la_data_out[11]
port 312 nsew
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1400 90 0 0 la_data_out[120]
port 313 nsew
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1400 90 0 0 la_data_out[121]
port 314 nsew
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1400 90 0 0 la_data_out[122]
port 315 nsew
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1400 90 0 0 la_data_out[123]
port 316 nsew
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1400 90 0 0 la_data_out[124]
port 317 nsew
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1400 90 0 0 la_data_out[125]
port 318 nsew
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1400 90 0 0 la_data_out[126]
port 319 nsew
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1400 90 0 0 la_data_out[127]
port 320 nsew
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1400 90 0 0 la_data_out[12]
port 321 nsew
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1400 90 0 0 la_data_out[13]
port 322 nsew
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1400 90 0 0 la_data_out[14]
port 323 nsew
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1400 90 0 0 la_data_out[15]
port 324 nsew
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1400 90 0 0 la_data_out[16]
port 325 nsew
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1400 90 0 0 la_data_out[17]
port 326 nsew
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1400 90 0 0 la_data_out[18]
port 327 nsew
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1400 90 0 0 la_data_out[19]
port 328 nsew
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1400 90 0 0 la_data_out[1]
port 329 nsew
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1400 90 0 0 la_data_out[20]
port 330 nsew
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1400 90 0 0 la_data_out[21]
port 331 nsew
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1400 90 0 0 la_data_out[22]
port 332 nsew
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1400 90 0 0 la_data_out[23]
port 333 nsew
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1400 90 0 0 la_data_out[24]
port 334 nsew
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1400 90 0 0 la_data_out[25]
port 335 nsew
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1400 90 0 0 la_data_out[26]
port 336 nsew
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1400 90 0 0 la_data_out[27]
port 337 nsew
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1400 90 0 0 la_data_out[28]
port 338 nsew
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1400 90 0 0 la_data_out[29]
port 339 nsew
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1400 90 0 0 la_data_out[2]
port 340 nsew
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1400 90 0 0 la_data_out[30]
port 341 nsew
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1400 90 0 0 la_data_out[31]
port 342 nsew
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1400 90 0 0 la_data_out[32]
port 343 nsew
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1400 90 0 0 la_data_out[33]
port 344 nsew
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1400 90 0 0 la_data_out[34]
port 345 nsew
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1400 90 0 0 la_data_out[35]
port 346 nsew
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1400 90 0 0 la_data_out[36]
port 347 nsew
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1400 90 0 0 la_data_out[37]
port 348 nsew
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1400 90 0 0 la_data_out[38]
port 349 nsew
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1400 90 0 0 la_data_out[39]
port 350 nsew
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1400 90 0 0 la_data_out[3]
port 351 nsew
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1400 90 0 0 la_data_out[40]
port 352 nsew
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1400 90 0 0 la_data_out[41]
port 353 nsew
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1400 90 0 0 la_data_out[42]
port 354 nsew
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1400 90 0 0 la_data_out[43]
port 355 nsew
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1400 90 0 0 la_data_out[44]
port 356 nsew
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1400 90 0 0 la_data_out[45]
port 357 nsew
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1400 90 0 0 la_data_out[46]
port 358 nsew
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1400 90 0 0 la_data_out[47]
port 359 nsew
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1400 90 0 0 la_data_out[48]
port 360 nsew
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1400 90 0 0 la_data_out[49]
port 361 nsew
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1400 90 0 0 la_data_out[4]
port 362 nsew
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1400 90 0 0 la_data_out[50]
port 363 nsew
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1400 90 0 0 la_data_out[51]
port 364 nsew
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1400 90 0 0 la_data_out[52]
port 365 nsew
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1400 90 0 0 la_data_out[53]
port 366 nsew
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1400 90 0 0 la_data_out[54]
port 367 nsew
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1400 90 0 0 la_data_out[55]
port 368 nsew
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1400 90 0 0 la_data_out[56]
port 369 nsew
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1400 90 0 0 la_data_out[57]
port 370 nsew
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1400 90 0 0 la_data_out[58]
port 371 nsew
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1400 90 0 0 la_data_out[59]
port 372 nsew
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1400 90 0 0 la_data_out[5]
port 373 nsew
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1400 90 0 0 la_data_out[60]
port 374 nsew
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1400 90 0 0 la_data_out[61]
port 375 nsew
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1400 90 0 0 la_data_out[62]
port 376 nsew
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1400 90 0 0 la_data_out[63]
port 377 nsew
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1400 90 0 0 la_data_out[64]
port 378 nsew
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1400 90 0 0 la_data_out[65]
port 379 nsew
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1400 90 0 0 la_data_out[66]
port 380 nsew
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1400 90 0 0 la_data_out[67]
port 381 nsew
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1400 90 0 0 la_data_out[68]
port 382 nsew
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1400 90 0 0 la_data_out[69]
port 383 nsew
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1400 90 0 0 la_data_out[6]
port 384 nsew
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1400 90 0 0 la_data_out[70]
port 385 nsew
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1400 90 0 0 la_data_out[71]
port 386 nsew
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1400 90 0 0 la_data_out[72]
port 387 nsew
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1400 90 0 0 la_data_out[73]
port 388 nsew
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1400 90 0 0 la_data_out[74]
port 389 nsew
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1400 90 0 0 la_data_out[75]
port 390 nsew
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1400 90 0 0 la_data_out[76]
port 391 nsew
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1400 90 0 0 la_data_out[77]
port 392 nsew
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1400 90 0 0 la_data_out[78]
port 393 nsew
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1400 90 0 0 la_data_out[79]
port 394 nsew
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1400 90 0 0 la_data_out[7]
port 395 nsew
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1400 90 0 0 la_data_out[80]
port 396 nsew
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1400 90 0 0 la_data_out[81]
port 397 nsew
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1400 90 0 0 la_data_out[82]
port 398 nsew
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1400 90 0 0 la_data_out[83]
port 399 nsew
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1400 90 0 0 la_data_out[84]
port 400 nsew
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1400 90 0 0 la_data_out[85]
port 401 nsew
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1400 90 0 0 la_data_out[86]
port 402 nsew
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1400 90 0 0 la_data_out[87]
port 403 nsew
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1400 90 0 0 la_data_out[88]
port 404 nsew
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1400 90 0 0 la_data_out[89]
port 405 nsew
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1400 90 0 0 la_data_out[8]
port 406 nsew
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1400 90 0 0 la_data_out[90]
port 407 nsew
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1400 90 0 0 la_data_out[91]
port 408 nsew
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1400 90 0 0 la_data_out[92]
port 409 nsew
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1400 90 0 0 la_data_out[93]
port 410 nsew
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1400 90 0 0 la_data_out[94]
port 411 nsew
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1400 90 0 0 la_data_out[95]
port 412 nsew
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1400 90 0 0 la_data_out[96]
port 413 nsew
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1400 90 0 0 la_data_out[97]
port 414 nsew
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1400 90 0 0 la_data_out[98]
port 415 nsew
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1400 90 0 0 la_data_out[99]
port 416 nsew
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1400 90 0 0 la_data_out[9]
port 417 nsew
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1400 90 0 0 la_oenb[0]
port 418 nsew
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1400 90 0 0 la_oenb[100]
port 419 nsew
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1400 90 0 0 la_oenb[101]
port 420 nsew
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1400 90 0 0 la_oenb[102]
port 421 nsew
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1400 90 0 0 la_oenb[103]
port 422 nsew
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1400 90 0 0 la_oenb[104]
port 423 nsew
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1400 90 0 0 la_oenb[105]
port 424 nsew
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1400 90 0 0 la_oenb[106]
port 425 nsew
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1400 90 0 0 la_oenb[107]
port 426 nsew
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1400 90 0 0 la_oenb[108]
port 427 nsew
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1400 90 0 0 la_oenb[109]
port 428 nsew
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1400 90 0 0 la_oenb[10]
port 429 nsew
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1400 90 0 0 la_oenb[110]
port 430 nsew
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1400 90 0 0 la_oenb[111]
port 431 nsew
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1400 90 0 0 la_oenb[112]
port 432 nsew
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1400 90 0 0 la_oenb[113]
port 433 nsew
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1400 90 0 0 la_oenb[114]
port 434 nsew
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1400 90 0 0 la_oenb[115]
port 435 nsew
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1400 90 0 0 la_oenb[116]
port 436 nsew
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1400 90 0 0 la_oenb[117]
port 437 nsew
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1400 90 0 0 la_oenb[118]
port 438 nsew
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1400 90 0 0 la_oenb[119]
port 439 nsew
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1400 90 0 0 la_oenb[11]
port 440 nsew
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1400 90 0 0 la_oenb[120]
port 441 nsew
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1400 90 0 0 la_oenb[121]
port 442 nsew
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1400 90 0 0 la_oenb[122]
port 443 nsew
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1400 90 0 0 la_oenb[123]
port 444 nsew
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1400 90 0 0 la_oenb[124]
port 445 nsew
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1400 90 0 0 la_oenb[125]
port 446 nsew
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1400 90 0 0 la_oenb[126]
port 447 nsew
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1400 90 0 0 la_oenb[127]
port 448 nsew
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1400 90 0 0 la_oenb[12]
port 449 nsew
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1400 90 0 0 la_oenb[13]
port 450 nsew
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1400 90 0 0 la_oenb[14]
port 451 nsew
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1400 90 0 0 la_oenb[15]
port 452 nsew
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1400 90 0 0 la_oenb[16]
port 453 nsew
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1400 90 0 0 la_oenb[17]
port 454 nsew
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1400 90 0 0 la_oenb[18]
port 455 nsew
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1400 90 0 0 la_oenb[19]
port 456 nsew
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1400 90 0 0 la_oenb[1]
port 457 nsew
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1400 90 0 0 la_oenb[20]
port 458 nsew
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1400 90 0 0 la_oenb[21]
port 459 nsew
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1400 90 0 0 la_oenb[22]
port 460 nsew
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1400 90 0 0 la_oenb[23]
port 461 nsew
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1400 90 0 0 la_oenb[24]
port 462 nsew
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1400 90 0 0 la_oenb[25]
port 463 nsew
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1400 90 0 0 la_oenb[26]
port 464 nsew
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1400 90 0 0 la_oenb[27]
port 465 nsew
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1400 90 0 0 la_oenb[28]
port 466 nsew
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1400 90 0 0 la_oenb[29]
port 467 nsew
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1400 90 0 0 la_oenb[2]
port 468 nsew
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1400 90 0 0 la_oenb[30]
port 469 nsew
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1400 90 0 0 la_oenb[31]
port 470 nsew
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1400 90 0 0 la_oenb[32]
port 471 nsew
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1400 90 0 0 la_oenb[33]
port 472 nsew
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1400 90 0 0 la_oenb[34]
port 473 nsew
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1400 90 0 0 la_oenb[35]
port 474 nsew
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1400 90 0 0 la_oenb[36]
port 475 nsew
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1400 90 0 0 la_oenb[37]
port 476 nsew
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1400 90 0 0 la_oenb[38]
port 477 nsew
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1400 90 0 0 la_oenb[39]
port 478 nsew
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1400 90 0 0 la_oenb[3]
port 479 nsew
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1400 90 0 0 la_oenb[40]
port 480 nsew
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1400 90 0 0 la_oenb[41]
port 481 nsew
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1400 90 0 0 la_oenb[42]
port 482 nsew
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1400 90 0 0 la_oenb[43]
port 483 nsew
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1400 90 0 0 la_oenb[44]
port 484 nsew
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1400 90 0 0 la_oenb[45]
port 485 nsew
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1400 90 0 0 la_oenb[46]
port 486 nsew
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1400 90 0 0 la_oenb[47]
port 487 nsew
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1400 90 0 0 la_oenb[48]
port 488 nsew
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1400 90 0 0 la_oenb[49]
port 489 nsew
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1400 90 0 0 la_oenb[4]
port 490 nsew
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1400 90 0 0 la_oenb[50]
port 491 nsew
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1400 90 0 0 la_oenb[51]
port 492 nsew
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1400 90 0 0 la_oenb[52]
port 493 nsew
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1400 90 0 0 la_oenb[53]
port 494 nsew
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1400 90 0 0 la_oenb[54]
port 495 nsew
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1400 90 0 0 la_oenb[55]
port 496 nsew
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1400 90 0 0 la_oenb[56]
port 497 nsew
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1400 90 0 0 la_oenb[57]
port 498 nsew
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1400 90 0 0 la_oenb[58]
port 499 nsew
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1400 90 0 0 la_oenb[59]
port 500 nsew
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1400 90 0 0 la_oenb[5]
port 501 nsew
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1400 90 0 0 la_oenb[60]
port 502 nsew
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1400 90 0 0 la_oenb[61]
port 503 nsew
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1400 90 0 0 la_oenb[62]
port 504 nsew
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1400 90 0 0 la_oenb[63]
port 505 nsew
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1400 90 0 0 la_oenb[64]
port 506 nsew
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1400 90 0 0 la_oenb[65]
port 507 nsew
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1400 90 0 0 la_oenb[66]
port 508 nsew
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1400 90 0 0 la_oenb[67]
port 509 nsew
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1400 90 0 0 la_oenb[68]
port 510 nsew
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1400 90 0 0 la_oenb[69]
port 511 nsew
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1400 90 0 0 la_oenb[6]
port 512 nsew
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1400 90 0 0 la_oenb[70]
port 513 nsew
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1400 90 0 0 la_oenb[71]
port 514 nsew
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1400 90 0 0 la_oenb[72]
port 515 nsew
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1400 90 0 0 la_oenb[73]
port 516 nsew
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1400 90 0 0 la_oenb[74]
port 517 nsew
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1400 90 0 0 la_oenb[75]
port 518 nsew
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1400 90 0 0 la_oenb[76]
port 519 nsew
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1400 90 0 0 la_oenb[77]
port 520 nsew
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1400 90 0 0 la_oenb[78]
port 521 nsew
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1400 90 0 0 la_oenb[79]
port 522 nsew
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1400 90 0 0 la_oenb[7]
port 523 nsew
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1400 90 0 0 la_oenb[80]
port 524 nsew
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1400 90 0 0 la_oenb[81]
port 525 nsew
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1400 90 0 0 la_oenb[82]
port 526 nsew
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1400 90 0 0 la_oenb[83]
port 527 nsew
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1400 90 0 0 la_oenb[84]
port 528 nsew
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1400 90 0 0 la_oenb[85]
port 529 nsew
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1400 90 0 0 la_oenb[86]
port 530 nsew
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1400 90 0 0 la_oenb[87]
port 531 nsew
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1400 90 0 0 la_oenb[88]
port 532 nsew
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1400 90 0 0 la_oenb[89]
port 533 nsew
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1400 90 0 0 la_oenb[8]
port 534 nsew
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1400 90 0 0 la_oenb[90]
port 535 nsew
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1400 90 0 0 la_oenb[91]
port 536 nsew
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1400 90 0 0 la_oenb[92]
port 537 nsew
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1400 90 0 0 la_oenb[93]
port 538 nsew
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1400 90 0 0 la_oenb[94]
port 539 nsew
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1400 90 0 0 la_oenb[95]
port 540 nsew
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1400 90 0 0 la_oenb[96]
port 541 nsew
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1400 90 0 0 la_oenb[97]
port 542 nsew
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1400 90 0 0 la_oenb[98]
port 543 nsew
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1400 90 0 0 la_oenb[99]
port 544 nsew
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1400 90 0 0 la_oenb[9]
port 545 nsew
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1400 90 0 0 user_clock2
port 546 nsew
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1400 90 0 0 user_irq[0]
port 547 nsew
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1400 90 0 0 user_irq[1]
port 548 nsew
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1400 90 0 0 user_irq[2]
port 549 nsew
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1400 0 0 0 vccd1
port 550 nsew
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1400 0 0 0 vccd1
port 550 nsew
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1400 0 0 0 vccd2
port 551 nsew
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1400 0 0 0 vccd2
port 551 nsew
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1400 0 0 0 vdda2
port 553 nsew
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1400 0 0 0 vdda2
port 553 nsew
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 2400 180 0 0 vssa1
port 554 nsew
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 2400 180 0 0 vssa1
port 554 nsew
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1400 0 0 0 vssa1
port 554 nsew
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1400 0 0 0 vssa1
port 554 nsew
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1400 0 0 0 vssa2
port 555 nsew
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1400 0 0 0 vssa2
port 555 nsew
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1400 0 0 0 vssd1
port 556 nsew
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1400 0 0 0 vssd1
port 556 nsew
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1400 0 0 0 vssd2
port 557 nsew
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1400 0 0 0 vssd2
port 557 nsew
flabel metal2 s 524 -800 636 480 0 FreeSans 1400 90 0 0 wb_clk_i
port 558 nsew
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1400 90 0 0 wb_rst_i
port 559 nsew
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1400 90 0 0 wbs_ack_o
port 560 nsew
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1400 90 0 0 wbs_adr_i[0]
port 561 nsew
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1400 90 0 0 wbs_adr_i[10]
port 562 nsew
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1400 90 0 0 wbs_adr_i[11]
port 563 nsew
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1400 90 0 0 wbs_adr_i[12]
port 564 nsew
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1400 90 0 0 wbs_adr_i[13]
port 565 nsew
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1400 90 0 0 wbs_adr_i[14]
port 566 nsew
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1400 90 0 0 wbs_adr_i[15]
port 567 nsew
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1400 90 0 0 wbs_adr_i[16]
port 568 nsew
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1400 90 0 0 wbs_adr_i[17]
port 569 nsew
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1400 90 0 0 wbs_adr_i[18]
port 570 nsew
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1400 90 0 0 wbs_adr_i[19]
port 571 nsew
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1400 90 0 0 wbs_adr_i[1]
port 572 nsew
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1400 90 0 0 wbs_adr_i[20]
port 573 nsew
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1400 90 0 0 wbs_adr_i[21]
port 574 nsew
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1400 90 0 0 wbs_adr_i[22]
port 575 nsew
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1400 90 0 0 wbs_adr_i[23]
port 576 nsew
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1400 90 0 0 wbs_adr_i[24]
port 577 nsew
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1400 90 0 0 wbs_adr_i[25]
port 578 nsew
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1400 90 0 0 wbs_adr_i[26]
port 579 nsew
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1400 90 0 0 wbs_adr_i[27]
port 580 nsew
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1400 90 0 0 wbs_adr_i[28]
port 581 nsew
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1400 90 0 0 wbs_adr_i[29]
port 582 nsew
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1400 90 0 0 wbs_adr_i[2]
port 583 nsew
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1400 90 0 0 wbs_adr_i[30]
port 584 nsew
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1400 90 0 0 wbs_adr_i[31]
port 585 nsew
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1400 90 0 0 wbs_adr_i[3]
port 586 nsew
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1400 90 0 0 wbs_adr_i[4]
port 587 nsew
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1400 90 0 0 wbs_adr_i[5]
port 588 nsew
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1400 90 0 0 wbs_adr_i[6]
port 589 nsew
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1400 90 0 0 wbs_adr_i[7]
port 590 nsew
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1400 90 0 0 wbs_adr_i[8]
port 591 nsew
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1400 90 0 0 wbs_adr_i[9]
port 592 nsew
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1400 90 0 0 wbs_cyc_i
port 593 nsew
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1400 90 0 0 wbs_dat_i[0]
port 594 nsew
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1400 90 0 0 wbs_dat_i[10]
port 595 nsew
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1400 90 0 0 wbs_dat_i[11]
port 596 nsew
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1400 90 0 0 wbs_dat_i[12]
port 597 nsew
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1400 90 0 0 wbs_dat_i[13]
port 598 nsew
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1400 90 0 0 wbs_dat_i[14]
port 599 nsew
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1400 90 0 0 wbs_dat_i[15]
port 600 nsew
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1400 90 0 0 wbs_dat_i[16]
port 601 nsew
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1400 90 0 0 wbs_dat_i[17]
port 602 nsew
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1400 90 0 0 wbs_dat_i[18]
port 603 nsew
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1400 90 0 0 wbs_dat_i[19]
port 604 nsew
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1400 90 0 0 wbs_dat_i[1]
port 605 nsew
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1400 90 0 0 wbs_dat_i[20]
port 606 nsew
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1400 90 0 0 wbs_dat_i[21]
port 607 nsew
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1400 90 0 0 wbs_dat_i[22]
port 608 nsew
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1400 90 0 0 wbs_dat_i[23]
port 609 nsew
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1400 90 0 0 wbs_dat_i[24]
port 610 nsew
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1400 90 0 0 wbs_dat_i[25]
port 611 nsew
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1400 90 0 0 wbs_dat_i[26]
port 612 nsew
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1400 90 0 0 wbs_dat_i[27]
port 613 nsew
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1400 90 0 0 wbs_dat_i[28]
port 614 nsew
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1400 90 0 0 wbs_dat_i[29]
port 615 nsew
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1400 90 0 0 wbs_dat_i[2]
port 616 nsew
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1400 90 0 0 wbs_dat_i[30]
port 617 nsew
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1400 90 0 0 wbs_dat_i[31]
port 618 nsew
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1400 90 0 0 wbs_dat_i[3]
port 619 nsew
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1400 90 0 0 wbs_dat_i[4]
port 620 nsew
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1400 90 0 0 wbs_dat_i[5]
port 621 nsew
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1400 90 0 0 wbs_dat_i[6]
port 622 nsew
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1400 90 0 0 wbs_dat_i[7]
port 623 nsew
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1400 90 0 0 wbs_dat_i[8]
port 624 nsew
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1400 90 0 0 wbs_dat_i[9]
port 625 nsew
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1400 90 0 0 wbs_dat_o[0]
port 626 nsew
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1400 90 0 0 wbs_dat_o[10]
port 627 nsew
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1400 90 0 0 wbs_dat_o[11]
port 628 nsew
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1400 90 0 0 wbs_dat_o[12]
port 629 nsew
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1400 90 0 0 wbs_dat_o[13]
port 630 nsew
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1400 90 0 0 wbs_dat_o[14]
port 631 nsew
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1400 90 0 0 wbs_dat_o[15]
port 632 nsew
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1400 90 0 0 wbs_dat_o[16]
port 633 nsew
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1400 90 0 0 wbs_dat_o[17]
port 634 nsew
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1400 90 0 0 wbs_dat_o[18]
port 635 nsew
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1400 90 0 0 wbs_dat_o[19]
port 636 nsew
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1400 90 0 0 wbs_dat_o[1]
port 637 nsew
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1400 90 0 0 wbs_dat_o[20]
port 638 nsew
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1400 90 0 0 wbs_dat_o[21]
port 639 nsew
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1400 90 0 0 wbs_dat_o[22]
port 640 nsew
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1400 90 0 0 wbs_dat_o[23]
port 641 nsew
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1400 90 0 0 wbs_dat_o[24]
port 642 nsew
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1400 90 0 0 wbs_dat_o[25]
port 643 nsew
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1400 90 0 0 wbs_dat_o[26]
port 644 nsew
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1400 90 0 0 wbs_dat_o[27]
port 645 nsew
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1400 90 0 0 wbs_dat_o[28]
port 646 nsew
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1400 90 0 0 wbs_dat_o[29]
port 647 nsew
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1400 90 0 0 wbs_dat_o[2]
port 648 nsew
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1400 90 0 0 wbs_dat_o[30]
port 649 nsew
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1400 90 0 0 wbs_dat_o[31]
port 650 nsew
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1400 90 0 0 wbs_dat_o[3]
port 651 nsew
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1400 90 0 0 wbs_dat_o[4]
port 652 nsew
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1400 90 0 0 wbs_dat_o[5]
port 653 nsew
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1400 90 0 0 wbs_dat_o[6]
port 654 nsew
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1400 90 0 0 wbs_dat_o[7]
port 655 nsew
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1400 90 0 0 wbs_dat_o[8]
port 656 nsew
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1400 90 0 0 wbs_dat_o[9]
port 657 nsew
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1400 90 0 0 wbs_sel_i[0]
port 658 nsew
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1400 90 0 0 wbs_sel_i[1]
port 659 nsew
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1400 90 0 0 wbs_sel_i[2]
port 660 nsew
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1400 90 0 0 wbs_sel_i[3]
port 661 nsew
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1400 90 0 0 wbs_stb_i
port 662 nsew
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1400 90 0 0 wbs_we_i
port 663 nsew
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1400 0 0 0 gpio_analog[0]
port 1 nsew
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1400 0 0 0 gpio_analog[1]
port 10 nsew
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1400 0 0 0 gpio_analog[2]
port 11 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
