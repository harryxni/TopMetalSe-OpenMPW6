* SPICE3 file created from pixel.ext - technology: sky130A

.subckt pixel gring test_net VREF ROW_SEL NB1 VBIAS NB2 AMP_IN SF_IB PIX_OUT CSA_VREF
+ VDD GND
X0 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt ad=25.3 pd=56.2 as=0 ps=0 w=2 l=2
X1 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.57 pd=12.3 as=0 ps=0 w=0.65 l=0.65
X2 a_4120_n520# VBIAS a_4120_n750# GND sky130_fd_pr__nfet_01v8_lvt ad=0.35 pd=2.7 as=3.99 ps=17.6 w=1 l=0.8
X3 test_net a_4600_n810# GND VDD sky130_fd_pr__pfet_01v8_lvt ad=0.5 pd=3 as=0.83 ps=5.9 w=1 l=1
X4 VDD SF_IB test_net VDD sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=1
X5 a_5460_10# a_4350_10# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0.35 pd=2.7 as=0 ps=0 w=1 l=2
X6 a_3860_n520# VBIAS a_3860_n1150# GND sky130_fd_pr__nfet_01v8_lvt ad=0.35 pd=2.7 as=3.52 ps=17.6 w=1 l=0.8
X7 VDD a_4120_n520# a_4600_n810# GND sky130_fd_pr__nfet_01v8_lvt ad=1.15 pd=8.3 as=0.5 ps=3 w=1 l=1
X8 a_4350_10# a_3860_n520# a_3860_n520# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.35 pd=2.7 as=0.35 ps=2.7 w=1 l=2
X9 a_4120_n750# AMP_IN a_4050_n2590# GND sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=3.22 ps=17.9 w=7 l=0.15
X10 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2 l=3.35
X11 a_4120_n520# a_3860_n520# a_5460_10# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.35 pd=2.7 as=0 ps=0 w=1 l=2
X12 GND NB1 a_4050_n2590# GND sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.2 l=1
X13 a_5750_n920# ROW_SEL PIX_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=1.2 pd=5.9 as=5.4 ps=9.4 w=2 l=1
X14 a_4050_n2590# VREF a_3860_n1150# GND sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=7 l=0.15
X15 a_4600_n810# NB2 GND GND sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=1.15
X16 AMP_IN a_4600_n810# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 VDD a_4350_10# a_4350_10# VDD sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=2
X18 VDD test_net a_5750_n920# GND sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X19 AMP_IN CSA_VREF a_4600_n810# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.294 pd=2.24 as=0.273 ps=2.14 w=0.42 l=8
X20 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.6 l=0.35
C0 gring SF_IB 0.249f
C1 test_net AMP_IN 0.125f
C2 a_4120_n520# a_3860_n520# 0.104f
C3 CSA_VREF AMP_IN 1.03f
C4 NB1 PIX_OUT 0.161f
C5 NB2 AMP_IN 0.328f
C6 test_net a_4600_n810# 0.149f
C7 VBIAS AMP_IN 0.263f
C8 SF_IB PIX_OUT 0.105f
C9 CSA_VREF a_4600_n810# 0.587f
C10 a_4600_n810# NB2 0.288f
C11 CSA_VREF gring 0.194f
C12 VDD AMP_IN 0.463f
C13 NB1 ROW_SEL 0.124f
C14 a_4600_n810# VDD 0.563f
C15 VDD gring 0.33f
C16 VDD a_4350_10# 0.613f
C17 CSA_VREF PIX_OUT 0.237f
C18 VREF VBIAS 0.259f
C19 VDD PIX_OUT 0.185f
C20 VREF VDD 0.14f
C21 a_4600_n810# AMP_IN 0.929f
C22 CSA_VREF ROW_SEL 0.21f
C23 VBIAS a_4120_n520# 0.204f
C24 CSA_VREF a_3860_n520# 0.204f
C25 NB2 ROW_SEL 0.143f
C26 gring AMP_IN 3.09f
C27 VDD a_4120_n520# 0.655f
C28 VDD ROW_SEL 0.197f
C29 VDD a_3860_n520# 1.01f
C30 PIX_OUT AMP_IN 0.534f
C31 VREF AMP_IN 0.12f
C32 CSA_VREF SF_IB 0.896f
C33 gring PIX_OUT 0.737f
C34 VREF gring 0.135f
C35 a_4120_n520# AMP_IN 0.125f
C36 ROW_SEL AMP_IN 0.785f
C37 test_net CSA_VREF 0.104f
C38 VDD SF_IB 0.633f
C39 a_4600_n810# a_4120_n520# 0.34f
C40 a_4600_n810# ROW_SEL 0.207f
C41 a_4120_n520# a_4350_10# 0.114f
C42 CSA_VREF NB2 0.109f
C43 ROW_SEL gring 0.152f
C44 a_4350_10# a_3860_n520# 0.417f
C45 VBIAS NB2 0.262f
C46 test_net VDD 0.146f
C47 NB1 AMP_IN 0.494f
C48 CSA_VREF VDD 0.815f
C49 VDD NB2 0.31f
C50 SF_IB AMP_IN 0.151f
C51 VBIAS VDD 0.229f
C52 ROW_SEL PIX_OUT 0.332f
C53 NB1 gring 0.27f
.ends

