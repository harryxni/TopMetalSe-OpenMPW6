magic
tech sky130A
magscale 1 2
timestamp 1654904798
<< metal1 >>
rect 302508 324533 302708 324539
rect 302508 321358 302708 324333
rect 303926 321358 304246 321364
rect 302508 321038 303926 321358
rect 108 319922 308 320311
rect 302508 320098 302708 321038
rect 303926 321032 304246 321038
rect 102 319722 108 319922
rect 308 319722 314 319922
rect 102 319700 314 319722
rect 108 319450 308 319700
rect 303926 318358 304246 318364
rect 302536 318038 303926 318358
rect 303926 318032 304246 318038
rect 108 316922 308 317311
rect 102 316722 108 316922
rect 308 316722 314 316922
rect 102 316700 314 316722
rect 108 316450 308 316700
rect 303926 315358 304246 315364
rect 302536 315038 303926 315358
rect 303926 315032 304246 315038
rect 108 313922 308 314311
rect 102 313722 108 313922
rect 308 313722 314 313922
rect 102 313700 314 313722
rect 108 313450 308 313700
rect 303926 312358 304246 312364
rect 302536 312038 303926 312358
rect 303926 312032 304246 312038
rect 108 310922 308 311311
rect 102 310722 108 310922
rect 308 310722 314 310922
rect 102 310700 314 310722
rect 108 310450 308 310700
rect 303926 309358 304246 309364
rect 302536 309038 303926 309358
rect 303926 309032 304246 309038
rect 108 307922 308 308311
rect 102 307722 108 307922
rect 308 307722 314 307922
rect 102 307700 314 307722
rect 108 307450 308 307700
rect 303926 306358 304246 306364
rect 302536 306038 303926 306358
rect 303926 306032 304246 306038
rect 108 304922 308 305311
rect 102 304722 108 304922
rect 308 304722 314 304922
rect 102 304700 314 304722
rect 108 304450 308 304700
rect 303926 303358 304246 303364
rect 302536 303038 303926 303358
rect 303926 303032 304246 303038
rect 108 301922 308 302311
rect 102 301722 108 301922
rect 308 301722 314 301922
rect 102 301700 314 301722
rect 108 301450 308 301700
rect 303926 300358 304246 300364
rect 302536 300038 303926 300358
rect 303926 300032 304246 300038
rect 108 298922 308 299311
rect 102 298722 108 298922
rect 308 298722 314 298922
rect 102 298700 314 298722
rect 108 298450 308 298700
rect 303926 297358 304246 297364
rect 302536 297038 303926 297358
rect 303926 297032 304246 297038
rect 108 295922 308 296311
rect 102 295722 108 295922
rect 308 295722 314 295922
rect 102 295700 314 295722
rect 108 295450 308 295700
rect 303926 294358 304246 294364
rect 302536 294038 303926 294358
rect 303926 294032 304246 294038
rect 108 292922 308 293311
rect 102 292722 108 292922
rect 308 292722 314 292922
rect 102 292700 314 292722
rect 108 292450 308 292700
rect 303926 291358 304246 291364
rect 302536 291038 303926 291358
rect 303926 291032 304246 291038
rect 108 289922 308 290311
rect 102 289722 108 289922
rect 308 289722 314 289922
rect 102 289700 314 289722
rect 108 289450 308 289700
rect 303926 288358 304246 288364
rect 302536 288038 303926 288358
rect 303926 288032 304246 288038
rect 108 286922 308 287311
rect 102 286722 108 286922
rect 308 286722 314 286922
rect 102 286700 314 286722
rect 108 286450 308 286700
rect 303926 285358 304246 285364
rect 302536 285038 303926 285358
rect 303926 285032 304246 285038
rect 108 283922 308 284311
rect 102 283722 108 283922
rect 308 283722 314 283922
rect 102 283700 314 283722
rect 108 283450 308 283700
rect 303926 282358 304246 282364
rect 302536 282038 303926 282358
rect 303926 282032 304246 282038
rect 108 280922 308 281311
rect 102 280722 108 280922
rect 308 280722 314 280922
rect 102 280700 314 280722
rect 108 280450 308 280700
rect 303926 279358 304246 279364
rect 302536 279038 303926 279358
rect 303926 279032 304246 279038
rect 108 277922 308 278311
rect 102 277722 108 277922
rect 308 277722 314 277922
rect 102 277700 314 277722
rect 108 277450 308 277700
rect 303926 276358 304246 276364
rect 302536 276038 303926 276358
rect 303926 276032 304246 276038
rect 108 274922 308 275311
rect 102 274722 108 274922
rect 308 274722 314 274922
rect 102 274700 314 274722
rect 108 274450 308 274700
rect 303926 273358 304246 273364
rect 302536 273038 303926 273358
rect 303926 273032 304246 273038
rect 108 271922 308 272311
rect 102 271722 108 271922
rect 308 271722 314 271922
rect 102 271700 314 271722
rect 108 271450 308 271700
rect 303926 270358 304246 270364
rect 302536 270038 303926 270358
rect 303926 270032 304246 270038
rect 108 268922 308 269311
rect 102 268722 108 268922
rect 308 268722 314 268922
rect 102 268700 314 268722
rect 108 268450 308 268700
rect 303926 267358 304246 267364
rect 302536 267038 303926 267358
rect 303926 267032 304246 267038
rect 108 265922 308 266311
rect 102 265722 108 265922
rect 308 265722 314 265922
rect 102 265700 314 265722
rect 108 265450 308 265700
rect 303926 264358 304246 264364
rect 302536 264038 303926 264358
rect 303926 264032 304246 264038
rect 108 262922 308 263311
rect 102 262722 108 262922
rect 308 262722 314 262922
rect 102 262700 314 262722
rect 108 262450 308 262700
rect 303926 261358 304246 261364
rect 302536 261038 303926 261358
rect 303926 261032 304246 261038
rect 108 259922 308 260311
rect 102 259722 108 259922
rect 308 259722 314 259922
rect 102 259700 314 259722
rect 108 259450 308 259700
rect 303926 258358 304246 258364
rect 302536 258038 303926 258358
rect 303926 258032 304246 258038
rect 108 256922 308 257311
rect 102 256722 108 256922
rect 308 256722 314 256922
rect 102 256700 314 256722
rect 108 256450 308 256700
rect 303926 255358 304246 255364
rect 302536 255038 303926 255358
rect 303926 255032 304246 255038
rect 108 253922 308 254311
rect 102 253722 108 253922
rect 308 253722 314 253922
rect 102 253700 314 253722
rect 108 253450 308 253700
rect 303926 252358 304246 252364
rect 302536 252038 303926 252358
rect 303926 252032 304246 252038
rect 108 250922 308 251311
rect 102 250722 108 250922
rect 308 250722 314 250922
rect 102 250700 314 250722
rect 108 250450 308 250700
rect 303926 249358 304246 249364
rect 302536 249038 303926 249358
rect 303926 249032 304246 249038
rect 108 247922 308 248311
rect 102 247722 108 247922
rect 308 247722 314 247922
rect 102 247700 314 247722
rect 108 247450 308 247700
rect 303926 246358 304246 246364
rect 302536 246038 303926 246358
rect 303926 246032 304246 246038
rect 108 244922 308 245311
rect 102 244722 108 244922
rect 308 244722 314 244922
rect 102 244700 314 244722
rect 108 244450 308 244700
rect 303926 243358 304246 243364
rect 302536 243038 303926 243358
rect 303926 243032 304246 243038
rect 108 241922 308 242311
rect 102 241722 108 241922
rect 308 241722 314 241922
rect 102 241700 314 241722
rect 108 241450 308 241700
rect 303926 240358 304246 240364
rect 302536 240038 303926 240358
rect 303926 240032 304246 240038
rect 108 238922 308 239311
rect 102 238722 108 238922
rect 308 238722 314 238922
rect 102 238700 314 238722
rect 108 238450 308 238700
rect 303926 237358 304246 237364
rect 302536 237038 303926 237358
rect 303926 237032 304246 237038
rect 108 235922 308 236311
rect 102 235722 108 235922
rect 308 235722 314 235922
rect 102 235700 314 235722
rect 108 235450 308 235700
rect 303926 234358 304246 234364
rect 302536 234038 303926 234358
rect 303926 234032 304246 234038
rect 108 232922 308 233311
rect 102 232722 108 232922
rect 308 232722 314 232922
rect 102 232700 314 232722
rect 108 232450 308 232700
rect 303926 231358 304246 231364
rect 302536 231038 303926 231358
rect 303926 231032 304246 231038
rect 108 229922 308 230311
rect 102 229722 108 229922
rect 308 229722 314 229922
rect 102 229700 314 229722
rect 108 229450 308 229700
rect 303926 228358 304246 228364
rect 302536 228038 303926 228358
rect 303926 228032 304246 228038
rect 108 226922 308 227311
rect 102 226722 108 226922
rect 308 226722 314 226922
rect 102 226700 314 226722
rect 108 226450 308 226700
rect 303926 225358 304246 225364
rect 302536 225038 303926 225358
rect 303926 225032 304246 225038
rect 108 223922 308 224311
rect 102 223722 108 223922
rect 308 223722 314 223922
rect 102 223700 314 223722
rect 108 223450 308 223700
rect 303926 222358 304246 222364
rect 302536 222038 303926 222358
rect 303926 222032 304246 222038
rect 108 220922 308 221311
rect 102 220722 108 220922
rect 308 220722 314 220922
rect 102 220700 314 220722
rect 108 220450 308 220700
rect 303926 219358 304246 219364
rect 302536 219038 303926 219358
rect 303926 219032 304246 219038
rect 108 217922 308 218311
rect 102 217722 108 217922
rect 308 217722 314 217922
rect 102 217700 314 217722
rect 108 217450 308 217700
rect 303926 216358 304246 216364
rect 302536 216038 303926 216358
rect 303926 216032 304246 216038
rect 108 214922 308 215311
rect 102 214722 108 214922
rect 308 214722 314 214922
rect 102 214700 314 214722
rect 108 214450 308 214700
rect 303926 213358 304246 213364
rect 302536 213038 303926 213358
rect 303926 213032 304246 213038
rect 108 211922 308 212311
rect 102 211722 108 211922
rect 308 211722 314 211922
rect 102 211700 314 211722
rect 108 211450 308 211700
rect 303926 210358 304246 210364
rect 302536 210038 303926 210358
rect 303926 210032 304246 210038
rect 108 208922 308 209311
rect 102 208722 108 208922
rect 308 208722 314 208922
rect 102 208700 314 208722
rect 108 208450 308 208700
rect 303926 207358 304246 207364
rect 302536 207038 303926 207358
rect 303926 207032 304246 207038
rect 108 205922 308 206311
rect 102 205722 108 205922
rect 308 205722 314 205922
rect 102 205700 314 205722
rect 108 205450 308 205700
rect 303926 204358 304246 204364
rect 302536 204038 303926 204358
rect 303926 204032 304246 204038
rect 108 202922 308 203311
rect 102 202722 108 202922
rect 308 202722 314 202922
rect 102 202700 314 202722
rect 108 202450 308 202700
rect 303926 201358 304246 201364
rect 302536 201038 303926 201358
rect 303926 201032 304246 201038
rect 108 199922 308 200311
rect 102 199722 108 199922
rect 308 199722 314 199922
rect 102 199700 314 199722
rect 108 199450 308 199700
rect 303926 198358 304246 198364
rect 302536 198038 303926 198358
rect 303926 198032 304246 198038
rect 108 196922 308 197311
rect 102 196722 108 196922
rect 308 196722 314 196922
rect 102 196700 314 196722
rect 108 196450 308 196700
rect 303926 195358 304246 195364
rect 302536 195038 303926 195358
rect 303926 195032 304246 195038
rect 108 193922 308 194311
rect 102 193722 108 193922
rect 308 193722 314 193922
rect 102 193700 314 193722
rect 108 193450 308 193700
rect 303926 192358 304246 192364
rect 302536 192038 303926 192358
rect 303926 192032 304246 192038
rect 108 190922 308 191311
rect 102 190722 108 190922
rect 308 190722 314 190922
rect 102 190700 314 190722
rect 108 190450 308 190700
rect 303926 189358 304246 189364
rect 302536 189038 303926 189358
rect 303926 189032 304246 189038
rect 108 187922 308 188311
rect 102 187722 108 187922
rect 308 187722 314 187922
rect 102 187700 314 187722
rect 108 187450 308 187700
rect 303926 186358 304246 186364
rect 302536 186038 303926 186358
rect 303926 186032 304246 186038
rect 108 184922 308 185311
rect 102 184722 108 184922
rect 308 184722 314 184922
rect 102 184700 314 184722
rect 108 184450 308 184700
rect 303926 183358 304246 183364
rect 302536 183038 303926 183358
rect 303926 183032 304246 183038
rect 108 181922 308 182311
rect 102 181722 108 181922
rect 308 181722 314 181922
rect 102 181700 314 181722
rect 108 181450 308 181700
rect 303926 180358 304246 180364
rect 302536 180038 303926 180358
rect 303926 180032 304246 180038
rect 108 178922 308 179311
rect 102 178722 108 178922
rect 308 178722 314 178922
rect 102 178700 314 178722
rect 108 178450 308 178700
rect 303926 177358 304246 177364
rect 302536 177038 303926 177358
rect 303926 177032 304246 177038
rect 108 175922 308 176311
rect 102 175722 108 175922
rect 308 175722 314 175922
rect 102 175700 314 175722
rect 108 175450 308 175700
rect 303926 174358 304246 174364
rect 302536 174038 303926 174358
rect 303926 174032 304246 174038
rect 108 172922 308 173311
rect 102 172722 108 172922
rect 308 172722 314 172922
rect 102 172700 314 172722
rect 108 172450 308 172700
rect 303926 171358 304246 171364
rect 302536 171038 303926 171358
rect 303926 171032 304246 171038
rect 108 169922 308 170311
rect 102 169722 108 169922
rect 308 169722 314 169922
rect 102 169700 314 169722
rect 108 169450 308 169700
rect 303926 168358 304246 168364
rect 302536 168038 303926 168358
rect 303926 168032 304246 168038
rect 108 166922 308 167311
rect 102 166722 108 166922
rect 308 166722 314 166922
rect 102 166700 314 166722
rect 108 166450 308 166700
rect 303926 165358 304246 165364
rect 302536 165038 303926 165358
rect 303926 165032 304246 165038
rect 108 163922 308 164311
rect 102 163722 108 163922
rect 308 163722 314 163922
rect 102 163700 314 163722
rect 108 163450 308 163700
rect 303926 162358 304246 162364
rect 302536 162038 303926 162358
rect 303926 162032 304246 162038
rect 108 160922 308 161311
rect 102 160722 108 160922
rect 308 160722 314 160922
rect 102 160700 314 160722
rect 108 160450 308 160700
rect 303926 159358 304246 159364
rect 302536 159038 303926 159358
rect 303926 159032 304246 159038
rect 108 157922 308 158311
rect 102 157722 108 157922
rect 308 157722 314 157922
rect 102 157700 314 157722
rect 108 157450 308 157700
rect 303926 156358 304246 156364
rect 302536 156038 303926 156358
rect 303926 156032 304246 156038
rect 108 154922 308 155311
rect 102 154722 108 154922
rect 308 154722 314 154922
rect 102 154700 314 154722
rect 108 154450 308 154700
rect 303926 153358 304246 153364
rect 302536 153038 303926 153358
rect 303926 153032 304246 153038
rect 108 151922 308 152311
rect 102 151722 108 151922
rect 308 151722 314 151922
rect 102 151700 314 151722
rect 108 151450 308 151700
rect 303926 150358 304246 150364
rect 302536 150038 303926 150358
rect 303926 150032 304246 150038
rect 108 148922 308 149311
rect 102 148722 108 148922
rect 308 148722 314 148922
rect 102 148700 314 148722
rect 108 148450 308 148700
rect 303926 147358 304246 147364
rect 302536 147038 303926 147358
rect 303926 147032 304246 147038
rect 108 145922 308 146311
rect 102 145722 108 145922
rect 308 145722 314 145922
rect 102 145700 314 145722
rect 108 145450 308 145700
rect 303926 144358 304246 144364
rect 302536 144038 303926 144358
rect 303926 144032 304246 144038
rect 108 142922 308 143311
rect 102 142722 108 142922
rect 308 142722 314 142922
rect 102 142700 314 142722
rect 108 142450 308 142700
rect 303926 141358 304246 141364
rect 302536 141038 303926 141358
rect 303926 141032 304246 141038
rect 108 139922 308 140311
rect 102 139722 108 139922
rect 308 139722 314 139922
rect 102 139700 314 139722
rect 108 139450 308 139700
rect 303926 138358 304246 138364
rect 302536 138038 303926 138358
rect 303926 138032 304246 138038
rect 108 136922 308 137311
rect 102 136722 108 136922
rect 308 136722 314 136922
rect 102 136700 314 136722
rect 108 136450 308 136700
rect 303926 135358 304246 135364
rect 302536 135038 303926 135358
rect 303926 135032 304246 135038
rect 108 133922 308 134311
rect 102 133722 108 133922
rect 308 133722 314 133922
rect 102 133700 314 133722
rect 108 133450 308 133700
rect 303926 132358 304246 132364
rect 302536 132038 303926 132358
rect 303926 132032 304246 132038
rect 108 130922 308 131311
rect 102 130722 108 130922
rect 308 130722 314 130922
rect 102 130700 314 130722
rect 108 130450 308 130700
rect 303926 129358 304246 129364
rect 302536 129038 303926 129358
rect 303926 129032 304246 129038
rect 108 127922 308 128311
rect 102 127722 108 127922
rect 308 127722 314 127922
rect 102 127700 314 127722
rect 108 127450 308 127700
rect 303926 126358 304246 126364
rect 302536 126038 303926 126358
rect 303926 126032 304246 126038
rect 108 124922 308 125311
rect 102 124722 108 124922
rect 308 124722 314 124922
rect 102 124700 314 124722
rect 108 124450 308 124700
rect 303926 123358 304246 123364
rect 302536 123038 303926 123358
rect 303926 123032 304246 123038
rect 108 121922 308 122311
rect 102 121722 108 121922
rect 308 121722 314 121922
rect 102 121700 314 121722
rect 108 121450 308 121700
rect 303926 120358 304246 120364
rect 302536 120038 303926 120358
rect 303926 120032 304246 120038
rect 108 118922 308 119311
rect 102 118722 108 118922
rect 308 118722 314 118922
rect 102 118700 314 118722
rect 108 118450 308 118700
rect 303926 117358 304246 117364
rect 302536 117038 303926 117358
rect 303926 117032 304246 117038
rect 108 115922 308 116311
rect 102 115722 108 115922
rect 308 115722 314 115922
rect 102 115700 314 115722
rect 108 115450 308 115700
rect 303926 114358 304246 114364
rect 302536 114038 303926 114358
rect 303926 114032 304246 114038
rect 108 112922 308 113311
rect 102 112722 108 112922
rect 308 112722 314 112922
rect 102 112700 314 112722
rect 108 112450 308 112700
rect 303926 111358 304246 111364
rect 302536 111038 303926 111358
rect 303926 111032 304246 111038
rect 108 109922 308 110311
rect 102 109722 108 109922
rect 308 109722 314 109922
rect 102 109700 314 109722
rect 108 109450 308 109700
rect 303926 108358 304246 108364
rect 302536 108038 303926 108358
rect 303926 108032 304246 108038
rect 108 106922 308 107311
rect 102 106722 108 106922
rect 308 106722 314 106922
rect 102 106700 314 106722
rect 108 106450 308 106700
rect 303926 105358 304246 105364
rect 302536 105038 303926 105358
rect 303926 105032 304246 105038
rect 108 103922 308 104311
rect 102 103722 108 103922
rect 308 103722 314 103922
rect 102 103700 314 103722
rect 108 103450 308 103700
rect 303926 102358 304246 102364
rect 302536 102038 303926 102358
rect 303926 102032 304246 102038
rect 108 100922 308 101311
rect 102 100722 108 100922
rect 308 100722 314 100922
rect 102 100700 314 100722
rect 108 100450 308 100700
rect 303926 99358 304246 99364
rect 302536 99038 303926 99358
rect 303926 99032 304246 99038
rect 108 97922 308 98311
rect 102 97722 108 97922
rect 308 97722 314 97922
rect 102 97700 314 97722
rect 108 97450 308 97700
rect 303926 96358 304246 96364
rect 302536 96038 303926 96358
rect 303926 96032 304246 96038
rect 108 94922 308 95311
rect 102 94722 108 94922
rect 308 94722 314 94922
rect 102 94700 314 94722
rect 108 94450 308 94700
rect 303926 93358 304246 93364
rect 302536 93038 303926 93358
rect 303926 93032 304246 93038
rect 108 91922 308 92311
rect 102 91722 108 91922
rect 308 91722 314 91922
rect 102 91700 314 91722
rect 108 91450 308 91700
rect 303926 90358 304246 90364
rect 302536 90038 303926 90358
rect 303926 90032 304246 90038
rect 108 88922 308 89311
rect 102 88722 108 88922
rect 308 88722 314 88922
rect 102 88700 314 88722
rect 108 88450 308 88700
rect 303926 87358 304246 87364
rect 302536 87038 303926 87358
rect 303926 87032 304246 87038
rect 108 85922 308 86311
rect 102 85722 108 85922
rect 308 85722 314 85922
rect 102 85700 314 85722
rect 108 85450 308 85700
rect 303926 84358 304246 84364
rect 302536 84038 303926 84358
rect 303926 84032 304246 84038
rect 108 82922 308 83311
rect 102 82722 108 82922
rect 308 82722 314 82922
rect 102 82700 314 82722
rect 108 82450 308 82700
rect 303926 81358 304246 81364
rect 302536 81038 303926 81358
rect 303926 81032 304246 81038
rect 108 79922 308 80311
rect 102 79722 108 79922
rect 308 79722 314 79922
rect 102 79700 314 79722
rect 108 79450 308 79700
rect 303926 78358 304246 78364
rect 302536 78038 303926 78358
rect 303926 78032 304246 78038
rect 108 76922 308 77311
rect 102 76722 108 76922
rect 308 76722 314 76922
rect 102 76700 314 76722
rect 108 76450 308 76700
rect 303926 75358 304246 75364
rect 302536 75038 303926 75358
rect 303926 75032 304246 75038
rect 108 73922 308 74311
rect 102 73722 108 73922
rect 308 73722 314 73922
rect 102 73700 314 73722
rect 108 73450 308 73700
rect 303926 72358 304246 72364
rect 302536 72038 303926 72358
rect 303926 72032 304246 72038
rect 108 70922 308 71311
rect 102 70722 108 70922
rect 308 70722 314 70922
rect 102 70700 314 70722
rect 108 70450 308 70700
rect 303926 69358 304246 69364
rect 302536 69038 303926 69358
rect 303926 69032 304246 69038
rect 108 67922 308 68311
rect 102 67722 108 67922
rect 308 67722 314 67922
rect 102 67700 314 67722
rect 108 67450 308 67700
rect 303926 66358 304246 66364
rect 302536 66038 303926 66358
rect 303926 66032 304246 66038
rect 108 64922 308 65311
rect 102 64722 108 64922
rect 308 64722 314 64922
rect 102 64700 314 64722
rect 108 64450 308 64700
rect 303926 63358 304246 63364
rect 302536 63038 303926 63358
rect 303926 63032 304246 63038
rect 108 61922 308 62311
rect 102 61722 108 61922
rect 308 61722 314 61922
rect 102 61700 314 61722
rect 108 61450 308 61700
rect 303926 60358 304246 60364
rect 302536 60038 303926 60358
rect 303926 60032 304246 60038
rect 108 58922 308 59311
rect 102 58722 108 58922
rect 308 58722 314 58922
rect 102 58700 314 58722
rect 108 58450 308 58700
rect 303926 57358 304246 57364
rect 302536 57038 303926 57358
rect 303926 57032 304246 57038
rect 108 55922 308 56311
rect 102 55722 108 55922
rect 308 55722 314 55922
rect 102 55700 314 55722
rect 108 55450 308 55700
rect 303926 54358 304246 54364
rect 302536 54038 303926 54358
rect 303926 54032 304246 54038
rect 108 52922 308 53311
rect 102 52722 108 52922
rect 308 52722 314 52922
rect 102 52700 314 52722
rect 108 52450 308 52700
rect 303926 51358 304246 51364
rect 302536 51038 303926 51358
rect 303926 51032 304246 51038
rect 108 49922 308 50311
rect 102 49722 108 49922
rect 308 49722 314 49922
rect 102 49700 314 49722
rect 108 49450 308 49700
rect 303926 48358 304246 48364
rect 302536 48038 303926 48358
rect 303926 48032 304246 48038
rect 108 46922 308 47311
rect 102 46722 108 46922
rect 308 46722 314 46922
rect 102 46700 314 46722
rect 108 46450 308 46700
rect 303926 45358 304246 45364
rect 302536 45038 303926 45358
rect 303926 45032 304246 45038
rect 108 43922 308 44311
rect 102 43722 108 43922
rect 308 43722 314 43922
rect 102 43700 314 43722
rect 108 43450 308 43700
rect 303926 42358 304246 42364
rect 302536 42038 303926 42358
rect 303926 42032 304246 42038
rect 108 40922 308 41311
rect 102 40722 108 40922
rect 308 40722 314 40922
rect 102 40700 314 40722
rect 108 40450 308 40700
rect 303926 39358 304246 39364
rect 302536 39038 303926 39358
rect 303926 39032 304246 39038
rect 108 37922 308 38311
rect 102 37722 108 37922
rect 308 37722 314 37922
rect 102 37700 314 37722
rect 108 37450 308 37700
rect 303926 36358 304246 36364
rect 302536 36038 303926 36358
rect 303926 36032 304246 36038
rect 108 34922 308 35311
rect 102 34722 108 34922
rect 308 34722 314 34922
rect 102 34700 314 34722
rect 108 34450 308 34700
rect 303926 33358 304246 33364
rect 302536 33038 303926 33358
rect 303926 33032 304246 33038
rect 108 31922 308 32311
rect 102 31722 108 31922
rect 308 31722 314 31922
rect 102 31700 314 31722
rect 108 31450 308 31700
rect 303926 30358 304246 30364
rect 302536 30038 303926 30358
rect 303926 30032 304246 30038
rect 108 28922 308 29311
rect 102 28722 108 28922
rect 308 28722 314 28922
rect 102 28700 314 28722
rect 108 28450 308 28700
rect 303926 27358 304246 27364
rect 302536 27038 303926 27358
rect 303926 27032 304246 27038
rect 108 25922 308 26311
rect 102 25722 108 25922
rect 308 25722 314 25922
rect 102 25700 314 25722
rect 108 25450 308 25700
rect 303926 24358 304246 24364
rect 302536 24038 303926 24358
rect 303926 24032 304246 24038
rect 108 22922 308 23311
rect 102 22722 108 22922
rect 308 22722 314 22922
rect 102 22700 314 22722
rect 108 22450 308 22700
rect 303926 21358 304246 21364
rect 302536 21038 303926 21358
rect 303926 21032 304246 21038
rect 108 19900 308 20808
rect 302508 20408 302828 20608
rect 102 19700 314 19900
rect 108 17947 308 19700
rect 3658 18440 3664 18760
rect 3984 18440 3990 18760
rect 18082 18440 18088 18760
rect 18408 18440 18414 18760
rect 32908 18440 32914 18760
rect 33234 18440 33240 18760
rect 64250 18440 64256 18760
rect 64576 18440 64582 18760
rect 121672 18440 121678 18760
rect 121998 18440 122004 18760
rect 167542 18440 167548 18760
rect 167868 18440 167874 18760
rect 180542 18440 180548 18760
rect 180868 18440 180874 18760
rect 189542 18440 189548 18760
rect 189868 18440 189874 18760
rect 198542 18440 198548 18760
rect 198868 18440 198874 18760
rect 204542 18440 204548 18760
rect 204868 18440 204874 18760
rect 211542 18440 211548 18760
rect 211868 18440 211874 18760
rect 223542 18440 223548 18760
rect 223868 18440 223874 18760
rect 232542 18440 232548 18760
rect 232868 18440 232874 18760
rect 238542 18440 238548 18760
rect 238868 18440 238874 18760
rect 250542 18440 250548 18760
rect 250868 18440 250874 18760
rect 263942 18440 263948 18760
rect 264268 18440 264274 18760
rect 269942 18440 269948 18760
rect 270268 18440 270274 18760
rect 272942 18440 272948 18760
rect 273268 18440 273274 18760
rect 275942 18440 275948 18760
rect 276268 18440 276274 18760
rect 281942 18440 281948 18760
rect 282268 18440 282274 18760
rect 285942 18440 285948 18760
rect 286268 18440 286274 18760
rect 293942 18440 293948 18760
rect 294268 18440 294274 18760
rect 296942 18440 296948 18760
rect 297268 18440 297274 18760
rect 299942 18440 299948 18760
rect 300268 18440 300274 18760
rect 302942 18440 302948 18760
rect 303268 18440 303274 18760
rect -6205 17747 -6199 17947
rect -5999 17747 308 17947
rect 3664 17938 3984 18440
rect 18088 17938 18408 18440
rect 32914 17938 33234 18440
rect 64256 17938 64576 18440
rect 121678 17938 121998 18440
rect 167548 17938 167868 18440
rect 180548 17938 180868 18440
rect 189548 17938 189868 18440
rect 198548 17938 198868 18440
rect 204548 17938 204868 18440
rect 211548 17938 211868 18440
rect 223548 17938 223868 18440
rect 232548 17938 232868 18440
rect 238548 17938 238868 18440
rect 250548 17938 250868 18440
rect 263948 17938 264268 18440
rect 269948 17938 270268 18440
rect 272948 17938 273268 18440
rect 275948 17938 276268 18440
rect 281948 17938 282268 18440
rect 285948 17938 286268 18440
rect 293948 17938 294268 18440
rect 296948 17938 297268 18440
rect 299948 17938 300268 18440
rect 302948 18259 303268 18440
rect 108 15588 308 17747
rect 302947 16416 303269 18259
rect 302947 16088 303269 16094
rect 108 15382 308 15388
<< via1 >>
rect 302508 324333 302708 324533
rect 303926 321038 304246 321358
rect 108 319722 308 319922
rect 303926 318038 304246 318358
rect 108 316722 308 316922
rect 303926 315038 304246 315358
rect 108 313722 308 313922
rect 303926 312038 304246 312358
rect 108 310722 308 310922
rect 303926 309038 304246 309358
rect 108 307722 308 307922
rect 303926 306038 304246 306358
rect 108 304722 308 304922
rect 303926 303038 304246 303358
rect 108 301722 308 301922
rect 303926 300038 304246 300358
rect 108 298722 308 298922
rect 303926 297038 304246 297358
rect 108 295722 308 295922
rect 303926 294038 304246 294358
rect 108 292722 308 292922
rect 303926 291038 304246 291358
rect 108 289722 308 289922
rect 303926 288038 304246 288358
rect 108 286722 308 286922
rect 303926 285038 304246 285358
rect 108 283722 308 283922
rect 303926 282038 304246 282358
rect 108 280722 308 280922
rect 303926 279038 304246 279358
rect 108 277722 308 277922
rect 303926 276038 304246 276358
rect 108 274722 308 274922
rect 303926 273038 304246 273358
rect 108 271722 308 271922
rect 303926 270038 304246 270358
rect 108 268722 308 268922
rect 303926 267038 304246 267358
rect 108 265722 308 265922
rect 303926 264038 304246 264358
rect 108 262722 308 262922
rect 303926 261038 304246 261358
rect 108 259722 308 259922
rect 303926 258038 304246 258358
rect 108 256722 308 256922
rect 303926 255038 304246 255358
rect 108 253722 308 253922
rect 303926 252038 304246 252358
rect 108 250722 308 250922
rect 303926 249038 304246 249358
rect 108 247722 308 247922
rect 303926 246038 304246 246358
rect 108 244722 308 244922
rect 303926 243038 304246 243358
rect 108 241722 308 241922
rect 303926 240038 304246 240358
rect 108 238722 308 238922
rect 303926 237038 304246 237358
rect 108 235722 308 235922
rect 303926 234038 304246 234358
rect 108 232722 308 232922
rect 303926 231038 304246 231358
rect 108 229722 308 229922
rect 303926 228038 304246 228358
rect 108 226722 308 226922
rect 303926 225038 304246 225358
rect 108 223722 308 223922
rect 303926 222038 304246 222358
rect 108 220722 308 220922
rect 303926 219038 304246 219358
rect 108 217722 308 217922
rect 303926 216038 304246 216358
rect 108 214722 308 214922
rect 303926 213038 304246 213358
rect 108 211722 308 211922
rect 303926 210038 304246 210358
rect 108 208722 308 208922
rect 303926 207038 304246 207358
rect 108 205722 308 205922
rect 303926 204038 304246 204358
rect 108 202722 308 202922
rect 303926 201038 304246 201358
rect 108 199722 308 199922
rect 303926 198038 304246 198358
rect 108 196722 308 196922
rect 303926 195038 304246 195358
rect 108 193722 308 193922
rect 303926 192038 304246 192358
rect 108 190722 308 190922
rect 303926 189038 304246 189358
rect 108 187722 308 187922
rect 303926 186038 304246 186358
rect 108 184722 308 184922
rect 303926 183038 304246 183358
rect 108 181722 308 181922
rect 303926 180038 304246 180358
rect 108 178722 308 178922
rect 303926 177038 304246 177358
rect 108 175722 308 175922
rect 303926 174038 304246 174358
rect 108 172722 308 172922
rect 303926 171038 304246 171358
rect 108 169722 308 169922
rect 303926 168038 304246 168358
rect 108 166722 308 166922
rect 303926 165038 304246 165358
rect 108 163722 308 163922
rect 303926 162038 304246 162358
rect 108 160722 308 160922
rect 303926 159038 304246 159358
rect 108 157722 308 157922
rect 303926 156038 304246 156358
rect 108 154722 308 154922
rect 303926 153038 304246 153358
rect 108 151722 308 151922
rect 303926 150038 304246 150358
rect 108 148722 308 148922
rect 303926 147038 304246 147358
rect 108 145722 308 145922
rect 303926 144038 304246 144358
rect 108 142722 308 142922
rect 303926 141038 304246 141358
rect 108 139722 308 139922
rect 303926 138038 304246 138358
rect 108 136722 308 136922
rect 303926 135038 304246 135358
rect 108 133722 308 133922
rect 303926 132038 304246 132358
rect 108 130722 308 130922
rect 303926 129038 304246 129358
rect 108 127722 308 127922
rect 303926 126038 304246 126358
rect 108 124722 308 124922
rect 303926 123038 304246 123358
rect 108 121722 308 121922
rect 303926 120038 304246 120358
rect 108 118722 308 118922
rect 303926 117038 304246 117358
rect 108 115722 308 115922
rect 303926 114038 304246 114358
rect 108 112722 308 112922
rect 303926 111038 304246 111358
rect 108 109722 308 109922
rect 303926 108038 304246 108358
rect 108 106722 308 106922
rect 303926 105038 304246 105358
rect 108 103722 308 103922
rect 303926 102038 304246 102358
rect 108 100722 308 100922
rect 303926 99038 304246 99358
rect 108 97722 308 97922
rect 303926 96038 304246 96358
rect 108 94722 308 94922
rect 303926 93038 304246 93358
rect 108 91722 308 91922
rect 303926 90038 304246 90358
rect 108 88722 308 88922
rect 303926 87038 304246 87358
rect 108 85722 308 85922
rect 303926 84038 304246 84358
rect 108 82722 308 82922
rect 303926 81038 304246 81358
rect 108 79722 308 79922
rect 303926 78038 304246 78358
rect 108 76722 308 76922
rect 303926 75038 304246 75358
rect 108 73722 308 73922
rect 303926 72038 304246 72358
rect 108 70722 308 70922
rect 303926 69038 304246 69358
rect 108 67722 308 67922
rect 303926 66038 304246 66358
rect 108 64722 308 64922
rect 303926 63038 304246 63358
rect 108 61722 308 61922
rect 303926 60038 304246 60358
rect 108 58722 308 58922
rect 303926 57038 304246 57358
rect 108 55722 308 55922
rect 303926 54038 304246 54358
rect 108 52722 308 52922
rect 303926 51038 304246 51358
rect 108 49722 308 49922
rect 303926 48038 304246 48358
rect 108 46722 308 46922
rect 303926 45038 304246 45358
rect 108 43722 308 43922
rect 303926 42038 304246 42358
rect 108 40722 308 40922
rect 303926 39038 304246 39358
rect 108 37722 308 37922
rect 303926 36038 304246 36358
rect 108 34722 308 34922
rect 303926 33038 304246 33358
rect 108 31722 308 31922
rect 303926 30038 304246 30358
rect 108 28722 308 28922
rect 303926 27038 304246 27358
rect 108 25722 308 25922
rect 303926 24038 304246 24358
rect 108 22722 308 22922
rect 303926 21038 304246 21358
rect 3664 18440 3984 18760
rect 18088 18440 18408 18760
rect 32914 18440 33234 18760
rect 64256 18440 64576 18760
rect 121678 18440 121998 18760
rect 167548 18440 167868 18760
rect 180548 18440 180868 18760
rect 189548 18440 189868 18760
rect 198548 18440 198868 18760
rect 204548 18440 204868 18760
rect 211548 18440 211868 18760
rect 223548 18440 223868 18760
rect 232548 18440 232868 18760
rect 238548 18440 238868 18760
rect 250548 18440 250868 18760
rect 263948 18440 264268 18760
rect 269948 18440 270268 18760
rect 272948 18440 273268 18760
rect 275948 18440 276268 18760
rect 281948 18440 282268 18760
rect 285948 18440 286268 18760
rect 293948 18440 294268 18760
rect 296948 18440 297268 18760
rect 299948 18440 300268 18760
rect 302948 18440 303268 18760
rect -6199 17747 -5999 17947
rect 302947 16094 303269 16416
rect 108 15388 308 15588
<< metal2 >>
rect -8167 325381 -1627 325491
rect -5180 322443 -2033 322533
rect -5132 319402 -2403 319458
rect -5168 316366 -2742 316422
rect -5148 313238 -3102 313294
rect -3535 310258 -3445 310275
rect -5148 310202 -3445 310258
rect -5138 307166 -3932 307222
rect -5158 304038 -4342 304094
rect -4398 302338 -4342 304038
rect -3988 303948 -3932 307166
rect -3535 306948 -3445 310202
rect -3158 309948 -3102 313238
rect -2798 312948 -2742 316366
rect -2459 315930 -2403 319402
rect -2123 318948 -2033 322443
rect -1737 320838 -1627 325381
rect 1358 321239 1468 327121
rect 2119 321418 2229 326997
rect 302508 324533 302708 324542
rect 302502 324333 302508 324533
rect 302708 324333 302714 324533
rect 302508 324324 302708 324333
rect 303931 321358 304241 321362
rect 303920 321038 303926 321358
rect 304246 321038 304252 321358
rect 303931 321034 304241 321038
rect -1737 320728 -782 320838
rect 108 319922 308 319928
rect 99 319722 108 319922
rect 308 319722 317 319922
rect 108 319716 308 319722
rect -2123 318858 -802 318948
rect 303931 318358 304241 318362
rect 303920 318038 303926 318358
rect 304246 318038 304252 318358
rect 303931 318034 304241 318038
rect 108 316922 308 316928
rect 99 316722 108 316922
rect 308 316722 317 316922
rect 108 316716 308 316722
rect -2459 315874 -579 315930
rect 303931 315358 304241 315362
rect 303920 315038 303926 315358
rect 304246 315038 304252 315358
rect 303931 315034 304241 315038
rect 108 313922 308 313928
rect 99 313722 108 313922
rect 308 313722 317 313922
rect 108 313716 308 313722
rect -2798 312892 -622 312948
rect 303931 312358 304241 312362
rect 303920 312038 303926 312358
rect 304246 312038 304252 312358
rect 303931 312034 304241 312038
rect 108 310922 308 310928
rect 99 310722 108 310922
rect 308 310722 317 310922
rect 108 310716 308 310722
rect -3165 309858 -755 309948
rect 303931 309358 304241 309362
rect 303920 309038 303926 309358
rect 304246 309038 304252 309358
rect 303931 309034 304241 309038
rect 108 307922 308 307928
rect 99 307722 108 307922
rect 308 307722 317 307922
rect 108 307716 308 307722
rect -3535 306858 -802 306948
rect 303931 306358 304241 306362
rect 303920 306038 303926 306358
rect 304246 306038 304252 306358
rect 303931 306034 304241 306038
rect 108 304922 308 304928
rect 99 304722 108 304922
rect 308 304722 317 304922
rect 108 304716 308 304722
rect -4005 303858 -775 303948
rect 303931 303358 304241 303362
rect 303920 303038 303926 303358
rect 304246 303038 304252 303358
rect 303931 303034 304241 303038
rect -4398 302282 -692 302338
rect -1485 301058 -1005 301065
rect -5128 301002 -1005 301058
rect -1485 300975 -1005 301002
rect -5148 297966 -1542 298022
rect -1635 294948 -1545 297966
rect -1095 297948 -1005 300975
rect -835 300858 -745 302282
rect 108 301922 308 301928
rect 99 301722 108 301922
rect 308 301722 317 301922
rect 108 301716 308 301722
rect 303931 300358 304241 300362
rect 303920 300038 303926 300358
rect 304246 300038 304252 300358
rect 303931 300034 304241 300038
rect 108 298922 308 298928
rect 99 298722 108 298922
rect 308 298722 317 298922
rect 108 298716 308 298722
rect -1095 297858 -745 297948
rect 303931 297358 304241 297362
rect 303920 297038 303926 297358
rect 304246 297038 304252 297358
rect 303931 297034 304241 297038
rect 108 295922 308 295928
rect 99 295722 108 295922
rect 308 295722 317 295922
rect 108 295716 308 295722
rect -5148 294838 -2152 294894
rect -1635 294858 -725 294948
rect -3095 291858 -3005 292055
rect -2208 291918 -2152 294838
rect 303931 294358 304241 294362
rect 303920 294038 303926 294358
rect 304246 294038 304252 294358
rect 303931 294034 304241 294038
rect 108 292922 308 292928
rect 99 292722 108 292922
rect 308 292722 317 292922
rect 108 292716 308 292722
rect -2208 291862 -452 291918
rect -5148 291802 -3005 291858
rect -3095 288948 -3005 291802
rect 303931 291358 304241 291362
rect 303920 291038 303926 291358
rect 304246 291038 304252 291358
rect 303931 291034 304241 291038
rect 108 289922 308 289928
rect 99 289722 108 289922
rect 308 289722 317 289922
rect 108 289716 308 289722
rect -3095 288858 -785 288948
rect -3915 288730 -3825 288815
rect -5148 288674 -3825 288730
rect -3915 285948 -3825 288674
rect 303931 288358 304241 288362
rect 303920 288038 303926 288358
rect 304246 288038 304252 288358
rect 303931 288034 304241 288038
rect 108 286922 308 286928
rect 99 286722 108 286922
rect 308 286722 317 286922
rect 108 286716 308 286722
rect -3915 285858 -765 285948
rect -5138 285638 -4232 285694
rect -4288 284088 -4232 285638
rect 303931 285358 304241 285362
rect 303920 285038 303926 285358
rect 304246 285038 304252 285358
rect 303931 285034 304241 285038
rect -1105 284088 -1015 284105
rect -4288 284032 -962 284088
rect -1105 282948 -1015 284032
rect 108 283922 308 283928
rect 99 283722 108 283922
rect 308 283722 317 283922
rect 108 283716 308 283722
rect -1105 282858 -802 282948
rect -2205 282658 -2115 282765
rect -5158 282602 -2115 282658
rect -2205 279948 -2115 282602
rect 303931 282358 304241 282362
rect 303920 282038 303926 282358
rect 304246 282038 304252 282358
rect 303931 282034 304241 282038
rect 108 280922 308 280928
rect 99 280722 108 280922
rect 308 280722 317 280922
rect 108 280716 308 280722
rect -2205 279858 -802 279948
rect -5218 279474 -1962 279530
rect -2055 276948 -1965 279474
rect 303931 279358 304241 279362
rect 303920 279038 303926 279358
rect 304246 279038 304252 279358
rect 303931 279034 304241 279038
rect 108 277922 308 277928
rect 99 277722 108 277922
rect 308 277722 317 277922
rect 108 277716 308 277722
rect -2055 276858 -785 276948
rect -892 276494 -802 276525
rect -5188 276438 -802 276494
rect -892 273858 -802 276438
rect 303931 276358 304241 276362
rect 303920 276038 303926 276358
rect 304246 276038 304252 276358
rect 303931 276034 304241 276038
rect 108 274922 308 274928
rect 99 274722 108 274922
rect 308 274722 317 274922
rect 108 274716 308 274722
rect -3965 273458 -3875 273585
rect -5228 273402 -3875 273458
rect -3965 270948 -3875 273402
rect 303931 273358 304241 273362
rect 303920 273038 303926 273358
rect 304246 273038 304252 273358
rect 303931 273034 304241 273038
rect 108 271922 308 271928
rect 99 271722 108 271922
rect 308 271722 317 271922
rect 108 271716 308 271722
rect -3965 270858 -802 270948
rect 303931 270358 304241 270362
rect -5168 270274 -4582 270330
rect -4638 267948 -4582 270274
rect 303920 270038 303926 270358
rect 304246 270038 304252 270358
rect 303931 270034 304241 270038
rect 108 268922 308 268928
rect 99 268722 108 268922
rect 308 268722 317 268922
rect 108 268716 308 268722
rect -4638 267882 -802 267948
rect -4615 267858 -802 267882
rect -4285 267294 -4195 267425
rect 303931 267358 304241 267362
rect -5148 267238 -4195 267294
rect -4285 264948 -4195 267238
rect 303920 267038 303926 267358
rect 304246 267038 304252 267358
rect 303931 267034 304241 267038
rect 108 265922 308 265928
rect 99 265722 108 265922
rect 308 265722 317 265922
rect 108 265716 308 265722
rect -4285 264858 -802 264948
rect 303931 264358 304241 264362
rect -5148 264110 -1932 264166
rect -1988 261948 -1932 264110
rect 303920 264038 303926 264358
rect 304246 264038 304252 264358
rect 303931 264034 304241 264038
rect 108 262922 308 262928
rect 99 262722 108 262922
rect 308 262722 317 262922
rect 108 262716 308 262722
rect -1988 261858 -802 261948
rect -1988 261812 -1932 261858
rect 303931 261358 304241 261362
rect -5178 261074 -1092 261130
rect -1148 258948 -1092 261074
rect 303920 261038 303926 261358
rect 304246 261038 304252 261358
rect 303931 261034 304241 261038
rect 108 259922 308 259928
rect 99 259722 108 259922
rect 308 259722 317 259922
rect 108 259716 308 259722
rect -1148 258858 -775 258948
rect -1148 258822 -1092 258858
rect 303931 258358 304241 258362
rect -5218 258038 -1112 258094
rect 303920 258038 303926 258358
rect 304246 258038 304252 258358
rect -1168 255948 -1112 258038
rect 303931 258034 304241 258038
rect 108 256922 308 256928
rect 99 256722 108 256922
rect 308 256722 317 256922
rect 108 256716 308 256722
rect -1168 255858 -802 255948
rect -1168 255842 -1112 255858
rect 303931 255358 304241 255362
rect 303920 255038 303926 255358
rect 304246 255038 304252 255358
rect 303931 255034 304241 255038
rect -5168 254910 -1172 254966
rect -1228 252948 -1172 254910
rect 108 253922 308 253928
rect 99 253722 108 253922
rect 308 253722 317 253922
rect 108 253716 308 253722
rect -1228 252858 -802 252948
rect -1228 252852 -1172 252858
rect 303931 252358 304241 252362
rect 303920 252038 303926 252358
rect 304246 252038 304252 252358
rect 303931 252034 304241 252038
rect -5208 251874 -1402 251930
rect -1458 249948 -1402 251874
rect 108 250922 308 250928
rect 99 250722 108 250922
rect 308 250722 317 250922
rect 108 250716 308 250722
rect -1458 249892 -795 249948
rect -1435 249858 -795 249892
rect 303931 249358 304241 249362
rect -885 248894 -795 249085
rect 303920 249038 303926 249358
rect 304246 249038 304252 249358
rect 303931 249034 304241 249038
rect -5128 248838 -792 248894
rect -885 246858 -795 248838
rect 108 247922 308 247928
rect 99 247722 108 247922
rect 308 247722 317 247922
rect 108 247716 308 247722
rect 303931 246358 304241 246362
rect 303920 246038 303926 246358
rect 304246 246038 304252 246358
rect 303931 246034 304241 246038
rect -892 245766 -802 245885
rect -5268 245710 -802 245766
rect -892 243858 -802 245710
rect 108 244922 308 244928
rect 99 244722 108 244922
rect 308 244722 317 244922
rect 108 244716 308 244722
rect 303931 243358 304241 243362
rect 303920 243038 303926 243358
rect 304246 243038 304252 243358
rect 303931 243034 304241 243038
rect -5228 242674 -832 242730
rect -888 240852 -832 242674
rect 108 241922 308 241928
rect 99 241722 108 241922
rect 308 241722 317 241922
rect 108 241716 308 241722
rect 303931 240358 304241 240362
rect 303920 240038 303926 240358
rect 304246 240038 304252 240358
rect 303931 240034 304241 240038
rect -5158 239638 -812 239694
rect -868 237892 -812 239638
rect 108 238922 308 238928
rect 99 238722 108 238922
rect 308 238722 317 238922
rect 108 238716 308 238722
rect 303931 237358 304241 237362
rect 303920 237038 303926 237358
rect 304246 237038 304252 237358
rect 303931 237034 304241 237038
rect -892 236566 -802 236725
rect -5188 236510 -802 236566
rect -892 234858 -802 236510
rect 108 235922 308 235928
rect 99 235722 108 235922
rect 308 235722 317 235922
rect 108 235716 308 235722
rect 303931 234358 304241 234362
rect 303920 234038 303926 234358
rect 304246 234038 304252 234358
rect 303931 234034 304241 234038
rect -5168 233474 -892 233530
rect -948 231852 -892 233474
rect 108 232922 308 232928
rect 99 232722 108 232922
rect 308 232722 317 232922
rect 108 232716 308 232722
rect 303931 231358 304241 231362
rect 303920 231038 303926 231358
rect 304246 231038 304252 231358
rect 303931 231034 304241 231038
rect -5168 228948 -5112 230402
rect 108 229922 308 229928
rect 99 229722 108 229922
rect 308 229722 317 229922
rect 108 229716 308 229722
rect -5168 228892 -785 228948
rect -5155 228858 -785 228892
rect 303931 228358 304241 228362
rect 303920 228038 303926 228358
rect 304246 228038 304252 228358
rect 303931 228034 304241 228038
rect -5138 227310 -612 227366
rect -835 225858 -745 227310
rect 108 226922 308 226928
rect 99 226722 108 226922
rect 308 226722 317 226922
rect 108 226716 308 226722
rect 303931 225358 304241 225362
rect 303920 225038 303926 225358
rect 304246 225038 304252 225358
rect 303931 225034 304241 225038
rect -5195 224265 -802 224355
rect -892 222858 -802 224265
rect 108 223922 308 223928
rect 99 223722 108 223922
rect 308 223722 317 223922
rect 108 223716 308 223722
rect 303931 222358 304241 222362
rect 303920 222038 303926 222358
rect 304246 222038 304252 222358
rect 303931 222034 304241 222038
rect -5148 221146 -808 221202
rect -864 219882 -808 221146
rect 108 220922 308 220928
rect 99 220722 108 220922
rect 308 220722 317 220922
rect 108 220716 308 220722
rect 303931 219358 304241 219362
rect 303920 219038 303926 219358
rect 304246 219038 304252 219358
rect 303931 219034 304241 219038
rect -808 218178 -752 218202
rect -5128 218122 -752 218178
rect -808 216872 -752 218122
rect 108 217922 308 217928
rect 99 217722 108 217922
rect 308 217722 317 217922
rect 108 217716 308 217722
rect 303931 216358 304241 216362
rect 303920 216038 303926 216358
rect 304246 216038 304252 216358
rect 303931 216034 304241 216038
rect -5128 215082 -752 215138
rect -808 213858 -752 215082
rect 108 214922 308 214928
rect 99 214722 108 214922
rect 308 214722 317 214922
rect 108 214716 308 214722
rect 303931 213358 304241 213362
rect 303920 213038 303926 213358
rect 304246 213038 304252 213358
rect 303931 213034 304241 213038
rect -5135 211915 -802 212005
rect 108 211922 308 211928
rect -892 210858 -802 211915
rect 99 211722 108 211922
rect 308 211722 317 211922
rect 108 211716 308 211722
rect 303931 210358 304241 210362
rect 303920 210038 303926 210358
rect 304246 210038 304252 210358
rect 303931 210034 304241 210038
rect -5128 208910 -732 208966
rect 108 208922 308 208928
rect -892 207872 -732 208910
rect 99 208722 108 208922
rect 308 208722 317 208922
rect 108 208716 308 208722
rect -892 207858 -765 207872
rect 303931 207358 304241 207362
rect 303920 207038 303926 207358
rect 304246 207038 304252 207358
rect 303931 207034 304241 207038
rect 108 205922 308 205928
rect -5168 205782 -802 205838
rect -858 204842 -802 205782
rect 99 205722 108 205922
rect 308 205722 317 205922
rect 108 205716 308 205722
rect 303931 204358 304241 204362
rect 303920 204038 303926 204358
rect 304246 204038 304252 204358
rect 303931 204034 304241 204038
rect 108 202922 308 202928
rect -5158 202746 -762 202802
rect -885 201858 -795 202746
rect 99 202722 108 202922
rect 308 202722 317 202922
rect 108 202716 308 202722
rect 303931 201358 304241 201362
rect 303920 201038 303926 201358
rect 304246 201038 304252 201358
rect 303931 201034 304241 201038
rect 108 199922 308 199928
rect -5208 199710 -722 199766
rect 99 199722 108 199922
rect 308 199722 317 199922
rect 108 199716 308 199722
rect -778 198852 -722 199710
rect 303931 198358 304241 198362
rect 303920 198038 303926 198358
rect 304246 198038 304252 198358
rect 303931 198034 304241 198038
rect 108 196922 308 196928
rect 99 196722 108 196922
rect 308 196722 317 196922
rect 108 196716 308 196722
rect -5145 196582 -1202 196638
rect -1258 195948 -1202 196582
rect -1258 195858 -793 195948
rect -1258 195805 -1202 195858
rect 303931 195358 304241 195362
rect 303920 195038 303926 195358
rect 304246 195038 304252 195358
rect 303931 195034 304241 195038
rect 108 193922 308 193928
rect 99 193722 108 193922
rect 308 193722 317 193922
rect 108 193716 308 193722
rect -5145 193552 -4891 193642
rect -4981 192948 -4891 193552
rect -4981 192858 -782 192948
rect 303931 192358 304241 192362
rect 303920 192038 303926 192358
rect 304246 192038 304252 192358
rect 303931 192034 304241 192038
rect 108 190922 308 190928
rect 99 190722 108 190922
rect 308 190722 317 190922
rect 108 190716 308 190722
rect -5134 190510 -737 190566
rect -793 189806 -737 190510
rect 303931 189358 304241 189362
rect 303920 189038 303926 189358
rect 304246 189038 304252 189358
rect 303931 189034 304241 189038
rect 108 187922 308 187928
rect 99 187722 108 187922
rect 308 187722 317 187922
rect 108 187716 308 187722
rect -5140 186948 -5050 187461
rect -5140 186858 -793 186948
rect 303931 186358 304241 186362
rect 303920 186038 303926 186358
rect 304246 186038 304252 186358
rect 303931 186034 304241 186038
rect 108 184922 308 184928
rect 99 184722 108 184922
rect 308 184722 317 184922
rect 108 184716 308 184722
rect -5140 183948 -5050 184425
rect -5140 183858 -578 183948
rect 303931 183358 304241 183362
rect 303920 183038 303926 183358
rect 304246 183038 304252 183358
rect 303931 183034 304241 183038
rect 108 181922 308 181928
rect 99 181722 108 181922
rect 308 181722 317 181922
rect 108 181716 308 181722
rect -5185 180948 -5095 181338
rect -5185 180858 -802 180948
rect 303931 180358 304241 180362
rect 303920 180038 303926 180358
rect 304246 180038 304252 180358
rect 303931 180034 304241 180038
rect 108 178922 308 178928
rect 99 178722 108 178922
rect 308 178722 317 178922
rect 108 178716 308 178722
rect -5168 177948 -5078 178234
rect -5168 177858 -572 177948
rect 303931 177358 304241 177362
rect 303920 177038 303926 177358
rect 304246 177038 304252 177358
rect 303931 177034 304241 177038
rect 108 175922 308 175928
rect 99 175722 108 175922
rect 308 175722 317 175922
rect 108 175716 308 175722
rect -5128 174948 -5072 175202
rect -5128 174858 -691 174948
rect -5128 174790 -5072 174858
rect 303931 174358 304241 174362
rect 303920 174038 303926 174358
rect 304246 174038 304252 174358
rect 303931 174034 304241 174038
rect 108 172922 308 172928
rect 99 172722 108 172922
rect 308 172722 317 172922
rect 108 172716 308 172722
rect -5208 171948 -5118 172065
rect -5208 171858 -782 171948
rect 303931 171358 304241 171362
rect 303920 171038 303926 171358
rect 304246 171038 304252 171358
rect 303931 171034 304241 171038
rect 108 169922 308 169928
rect 99 169722 108 169922
rect 308 169722 317 169922
rect 108 169716 308 169722
rect -5157 168948 -5067 169080
rect -5157 168858 -802 168948
rect 303931 168358 304241 168362
rect 303920 168038 303926 168358
rect 304246 168038 304252 168358
rect 303931 168034 304241 168038
rect 108 166922 308 166928
rect 99 166722 108 166922
rect 308 166722 317 166922
rect 108 166716 308 166722
rect -5145 165948 -5055 166032
rect -5145 165858 -731 165948
rect 303931 165358 304241 165362
rect 303920 165038 303926 165358
rect 304246 165038 304252 165358
rect 303931 165034 304241 165038
rect 108 163922 308 163928
rect 99 163722 108 163922
rect 308 163722 317 163922
rect 108 163716 308 163722
rect -5145 162858 -771 162948
rect 303931 162358 304241 162362
rect 303920 162038 303926 162358
rect 304246 162038 304252 162358
rect 303931 162034 304241 162038
rect 108 160922 308 160928
rect 99 160722 108 160922
rect 308 160722 317 160922
rect 108 160716 308 160722
rect -3852 159858 -799 159948
rect -5208 159782 -5202 159838
rect -3852 159779 -816 159858
rect 303931 159358 304241 159362
rect 303920 159038 303926 159358
rect 304246 159038 304252 159358
rect 303931 159034 304241 159038
rect 108 157922 308 157928
rect 99 157722 108 157922
rect 308 157722 317 157922
rect 108 157716 308 157722
rect -827 156901 -737 156948
rect -5162 156856 -737 156901
rect -5168 156743 -737 156856
rect 303931 156358 304241 156362
rect 303920 156038 303926 156358
rect 304246 156038 304252 156358
rect 303931 156034 304241 156038
rect 108 154922 308 154928
rect 99 154722 108 154922
rect 308 154722 317 154922
rect 108 154716 308 154722
rect -883 153678 -793 153948
rect -5134 153588 -793 153678
rect 303931 153358 304241 153362
rect 303920 153038 303926 153358
rect 304246 153038 304252 153358
rect 303931 153034 304241 153038
rect 108 151922 308 151928
rect 99 151722 108 151922
rect 308 151722 317 151922
rect 108 151716 308 151722
rect -5242 150585 -5010 150658
rect -892 150585 -802 150948
rect -5242 150568 -802 150585
rect -5100 150495 -802 150568
rect 303931 150358 304241 150362
rect 303920 150038 303926 150358
rect 304246 150038 304252 150358
rect 303931 150034 304241 150038
rect 108 148922 308 148928
rect 99 148722 108 148922
rect 308 148722 317 148922
rect 108 148716 308 148722
rect -5123 147429 -5033 147554
rect -883 147429 -793 147948
rect -5123 147339 -793 147429
rect 303931 147358 304241 147362
rect 303920 147038 303926 147358
rect 304246 147038 304252 147358
rect 303931 147034 304241 147038
rect 108 145922 308 145928
rect 99 145722 108 145922
rect 308 145722 317 145922
rect 108 145716 308 145722
rect -883 144569 -793 144948
rect -5179 144479 -793 144569
rect -5179 144417 -839 144479
rect 303931 144358 304241 144362
rect 303920 144038 303926 144358
rect 304246 144038 304252 144358
rect 303931 144034 304241 144038
rect 108 142922 308 142928
rect 99 142722 108 142922
rect 308 142722 317 142922
rect 108 142716 308 142722
rect -866 141505 -776 141948
rect -5140 141415 -776 141505
rect -5140 141352 -816 141415
rect 303931 141358 304241 141362
rect 303920 141038 303926 141358
rect 304246 141038 304252 141358
rect 303931 141034 304241 141038
rect 108 139922 308 139928
rect 99 139722 108 139922
rect 308 139722 317 139922
rect 108 139716 308 139722
rect -861 138338 -771 138948
rect 303931 138358 304241 138362
rect -5179 138248 -771 138338
rect 303920 138038 303926 138358
rect 304246 138038 304252 138358
rect 303931 138034 304241 138038
rect 108 136922 308 136928
rect 99 136722 108 136922
rect 308 136722 317 136922
rect 108 136716 308 136722
rect -892 135341 -802 135948
rect 303931 135358 304241 135362
rect -5191 135251 -802 135341
rect -5134 135183 -805 135251
rect 303920 135038 303926 135358
rect 304246 135038 304252 135358
rect 303931 135034 304241 135038
rect 108 133922 308 133928
rect 99 133722 108 133922
rect 308 133722 317 133922
rect 108 133716 308 133722
rect -849 132368 -759 132948
rect -5174 132278 -759 132368
rect 303931 132358 304241 132362
rect -5174 132187 -5084 132278
rect 303920 132038 303926 132358
rect 304246 132038 304252 132358
rect 303931 132034 304241 132038
rect 108 130922 308 130928
rect 99 130722 108 130922
rect 308 130722 317 130922
rect 108 130716 308 130722
rect -881 129085 -791 129948
rect 303931 129358 304241 129362
rect -5186 128937 -791 129085
rect 303920 129038 303926 129358
rect 304246 129038 304252 129358
rect 303931 129034 304241 129038
rect 108 127922 308 127928
rect 99 127722 108 127922
rect 308 127722 317 127922
rect 108 127716 308 127722
rect -853 126085 -763 126948
rect 303931 126358 304241 126362
rect -5198 125938 -763 126085
rect 303920 126038 303926 126358
rect 304246 126038 304252 126358
rect 303931 126034 304241 126038
rect 108 124922 308 124928
rect 99 124722 108 124922
rect 308 124722 317 124922
rect 108 124716 308 124722
rect -892 122977 -802 123948
rect 303931 123358 304241 123362
rect 303920 123038 303926 123358
rect 304246 123038 304252 123358
rect 303931 123034 304241 123038
rect -5141 122790 -802 122977
rect 108 121922 308 121928
rect 99 121722 108 121922
rect 308 121722 317 121922
rect 108 121716 308 121722
rect -5128 120948 -5072 121158
rect -5141 120858 -763 120948
rect -5128 119854 -5072 120858
rect 303931 120358 304241 120362
rect 303920 120038 303926 120358
rect 304246 120038 304252 120358
rect 303931 120034 304241 120038
rect 108 118922 308 118928
rect 99 118722 108 118922
rect 308 118722 317 118922
rect 108 118716 308 118722
rect -5186 117858 -802 117948
rect -5186 116775 -5096 117858
rect 303931 117358 304241 117362
rect 303920 117038 303926 117358
rect 304246 117038 304252 117358
rect 303931 117034 304241 117038
rect 108 115922 308 115928
rect 99 115722 108 115922
rect 308 115722 317 115922
rect 108 115716 308 115722
rect -5158 114858 -614 114948
rect -5158 113650 -5068 114858
rect 303931 114358 304241 114362
rect 303920 114038 303926 114358
rect 304246 114038 304252 114358
rect 303931 114034 304241 114038
rect 108 112922 308 112928
rect 99 112722 108 112922
rect 308 112722 317 112922
rect 108 112716 308 112722
rect -5192 111858 -768 111948
rect -5192 110633 -5102 111858
rect 303931 111358 304241 111362
rect 303920 111038 303926 111358
rect 304246 111038 304252 111358
rect 303931 111034 304241 111038
rect 108 109922 308 109928
rect 99 109722 108 109922
rect 308 109722 317 109922
rect 108 109716 308 109722
rect -5124 108858 -802 108948
rect -5124 107622 -5034 108858
rect 303931 108358 304241 108362
rect 303920 108038 303926 108358
rect 304246 108038 304252 108358
rect 303931 108034 304241 108038
rect 108 106922 308 106928
rect 99 106722 108 106922
rect 308 106722 317 106922
rect 108 106716 308 106722
rect -836 104588 -746 105948
rect 303931 105358 304241 105362
rect 303920 105038 303926 105358
rect 304246 105038 304252 105358
rect 303931 105034 304241 105038
rect -5164 104498 -746 104588
rect -5164 104490 -768 104498
rect 108 103922 308 103928
rect 99 103722 108 103922
rect 308 103722 317 103922
rect 108 103716 308 103722
rect -892 101548 -802 102948
rect 303931 102358 304241 102362
rect 303920 102038 303926 102358
rect 304246 102038 304252 102358
rect 303931 102034 304241 102038
rect -5175 101458 -802 101548
rect -892 101259 -802 101458
rect 108 100922 308 100928
rect 99 100722 108 100922
rect 308 100722 317 100922
rect 108 100716 308 100722
rect -892 98429 -802 99948
rect 303931 99358 304241 99362
rect 303920 99038 303926 99358
rect 304246 99038 304252 99358
rect 303931 99034 304241 99038
rect -5209 98339 -802 98429
rect -892 98077 -802 98339
rect 108 97922 308 97928
rect 99 97722 108 97922
rect 308 97722 317 97922
rect 108 97716 308 97722
rect -881 95396 -791 96948
rect 303931 96358 304241 96362
rect 303920 96038 303926 96358
rect 304246 96038 304252 96358
rect 303931 96034 304241 96038
rect -5181 95306 -791 95396
rect -881 95009 -791 95306
rect 108 94922 308 94928
rect 99 94722 108 94922
rect 308 94722 317 94922
rect 108 94716 308 94722
rect -870 92316 -780 93948
rect 303931 93358 304241 93362
rect 303920 93038 303926 93358
rect 304246 93038 304252 93358
rect 303931 93034 304241 93038
rect -5232 92226 -780 92316
rect -870 91913 -780 92226
rect 108 91922 308 91928
rect 99 91722 108 91922
rect 308 91722 317 91922
rect 108 91716 308 91722
rect -853 89209 -763 90948
rect 303931 90358 304241 90362
rect 303920 90038 303926 90358
rect 304246 90038 304252 90358
rect 303931 90034 304241 90038
rect -5192 89119 -763 89209
rect -853 89016 -763 89119
rect 108 88922 308 88928
rect 99 88722 108 88922
rect 308 88722 317 88922
rect 108 88716 308 88722
rect -836 86198 -746 87948
rect 303931 87358 304241 87362
rect 303920 87038 303926 87358
rect 304246 87038 304252 87358
rect 303931 87034 304241 87038
rect -5129 86108 -746 86198
rect -836 85977 -746 86108
rect 108 85922 308 85928
rect 99 85722 108 85922
rect 308 85722 317 85922
rect 108 85716 308 85722
rect -796 83153 -706 84948
rect 303931 84358 304241 84362
rect 303920 84038 303926 84358
rect 304246 84038 304252 84358
rect 303931 84034 304241 84038
rect -5221 83063 -706 83153
rect -796 82721 -706 83063
rect 108 82922 308 82928
rect 99 82722 108 82922
rect 308 82722 317 82922
rect 108 82716 308 82722
rect -881 80022 -791 81948
rect 303931 81358 304241 81362
rect 303920 81038 303926 81358
rect 304246 81038 304252 81358
rect 303931 81034 304241 81038
rect -5203 79932 -791 80022
rect -881 79527 -791 79932
rect 108 79922 308 79928
rect 99 79722 108 79922
rect 308 79722 317 79922
rect 108 79716 308 79722
rect -858 76949 -768 78948
rect 303931 78358 304241 78362
rect 303920 78038 303926 78358
rect 304246 78038 304252 78358
rect 303931 78034 304241 78038
rect -5209 76859 -768 76949
rect 108 76922 308 76928
rect -858 76391 -768 76859
rect 99 76722 108 76922
rect 308 76722 317 76922
rect 108 76716 308 76722
rect -5164 73773 -5074 74058
rect -790 73773 -700 75948
rect 303931 75358 304241 75362
rect 303920 75038 303926 75358
rect 304246 75038 304252 75358
rect 303931 75034 304241 75038
rect 108 73922 308 73928
rect -5164 73683 -700 73773
rect 99 73722 108 73922
rect 308 73722 317 73922
rect 108 73716 308 73722
rect -790 73477 -700 73683
rect -830 70796 -740 72948
rect 303931 72358 304241 72362
rect 303920 72038 303926 72358
rect 304246 72038 304252 72358
rect 303931 72034 304241 72038
rect 108 70922 308 70928
rect -5152 70706 -740 70796
rect 99 70722 108 70922
rect 308 70722 317 70922
rect 108 70716 308 70722
rect -830 70581 -740 70706
rect -5169 67654 -5079 67774
rect -892 67654 -802 69948
rect 303931 69358 304241 69362
rect 303920 69038 303926 69358
rect 304246 69038 304252 69358
rect 303931 69034 304241 69038
rect 108 67922 308 67928
rect 99 67722 108 67922
rect 308 67722 317 67922
rect 108 67716 308 67722
rect -5169 67564 -802 67654
rect -892 67370 -802 67564
rect -608 64618 -552 66924
rect 303931 66358 304241 66362
rect 303920 66038 303926 66358
rect 304246 66038 304252 66358
rect 303931 66034 304241 66038
rect 108 64922 308 64928
rect 99 64722 108 64922
rect 308 64722 317 64922
rect 108 64716 308 64722
rect -5226 64562 -552 64618
rect -5209 63858 -643 63948
rect -5209 61354 -5119 63858
rect 303931 63358 304241 63362
rect 303920 63038 303926 63358
rect 304246 63038 304252 63358
rect 303931 63034 304241 63038
rect 108 61922 308 61928
rect 99 61722 108 61922
rect 308 61722 317 61922
rect 108 61716 308 61722
rect -5243 60858 -700 60948
rect -5243 58378 -5153 60858
rect 303931 60358 304241 60362
rect 303920 60038 303926 60358
rect 304246 60038 304252 60358
rect 303931 60034 304241 60038
rect 108 58922 308 58928
rect 99 58722 108 58922
rect 308 58722 317 58922
rect 108 58716 308 58722
rect -5215 57858 -774 57948
rect -5215 55224 -5125 57858
rect 303931 57358 304241 57362
rect 303920 57038 303926 57358
rect 304246 57038 304252 57358
rect 303931 57034 304241 57038
rect 108 55922 308 55928
rect 99 55722 108 55922
rect 308 55722 317 55922
rect 108 55716 308 55722
rect -5243 54858 -774 54948
rect -5243 52316 -5153 54858
rect 303931 54358 304241 54362
rect 303920 54038 303926 54358
rect 304246 54038 304252 54358
rect 303931 54034 304241 54038
rect 108 52922 308 52928
rect 99 52722 108 52922
rect 308 52722 317 52922
rect 108 52716 308 52722
rect -322 49346 -266 52178
rect 303931 51358 304241 51362
rect 303920 51038 303926 51358
rect 304246 51038 304252 51358
rect 303931 51034 304241 51038
rect 108 49922 308 49928
rect 99 49722 108 49922
rect 308 49722 317 49922
rect 108 49716 308 49722
rect -5147 49290 -266 49346
rect -5226 48858 -489 48948
rect -5226 45970 -5136 48858
rect 303931 48358 304241 48362
rect 303920 48038 303926 48358
rect 304246 48038 304252 48358
rect 303931 48034 304241 48038
rect 108 46922 308 46928
rect 99 46722 108 46922
rect 308 46722 317 46922
rect 108 46716 308 46722
rect -3541 45858 -802 45948
rect -3541 43182 -3451 45858
rect 303931 45358 304241 45362
rect 303920 45038 303926 45358
rect 304246 45038 304252 45358
rect 303931 45034 304241 45038
rect 108 43922 308 43928
rect 99 43722 108 43922
rect 308 43722 317 43922
rect 108 43716 308 43722
rect -5188 43126 -3343 43182
rect -3541 42491 -3451 43126
rect -2360 42948 -2304 43190
rect -2459 42858 -802 42948
rect -2360 40054 -2304 42858
rect 303931 42358 304241 42362
rect 303920 42038 303926 42358
rect 304246 42038 304252 42358
rect 303931 42034 304241 42038
rect 108 40922 308 40928
rect 99 40722 108 40922
rect 308 40722 317 40922
rect 108 40716 308 40722
rect -5257 39998 -2304 40054
rect -751 38442 -661 39948
rect 303931 39358 304241 39362
rect 303920 39038 303926 39358
rect 304246 39038 304252 39358
rect 303931 39034 304241 39038
rect -1991 38386 -497 38442
rect -1991 37018 -1935 38386
rect -751 38281 -661 38386
rect 108 37922 308 37928
rect 99 37722 108 37922
rect 308 37722 317 37922
rect 108 37716 308 37722
rect -5131 36962 -1935 37018
rect -463 35565 -373 36948
rect 303931 36358 304241 36362
rect 303920 36038 303926 36358
rect 304246 36038 304252 36358
rect 303931 36034 304241 36038
rect -2435 35509 -373 35565
rect -2435 33982 -2379 35509
rect -463 35254 -373 35509
rect 108 34922 308 34928
rect 99 34722 108 34922
rect 308 34722 317 34922
rect 108 34716 308 34722
rect -5144 33926 -2379 33982
rect -772 32850 -716 34558
rect 303931 33358 304241 33362
rect 303920 33038 303926 33358
rect 304246 33038 304252 33358
rect 303931 33034 304241 33038
rect -3299 32794 -716 32850
rect -3299 30854 -3243 32794
rect 108 31922 308 31928
rect 99 31722 108 31922
rect 308 31722 317 31922
rect 108 31716 308 31722
rect -5175 30798 -3243 30854
rect -720 29741 -630 30948
rect 303931 30358 304241 30362
rect 303920 30038 303926 30358
rect 304246 30038 304252 30358
rect 303931 30034 304241 30038
rect -2905 29685 -584 29741
rect -2905 27818 -2849 29685
rect -720 29385 -584 29685
rect -720 29261 -630 29385
rect 108 28922 308 28928
rect 99 28722 108 28922
rect 308 28722 317 28922
rect 108 28716 308 28722
rect -5175 27762 -2849 27818
rect -757 26901 -667 27948
rect 303931 27358 304241 27362
rect 303920 27038 303926 27358
rect 304246 27038 304252 27358
rect 303931 27034 304241 27038
rect -2592 26845 -628 26901
rect -2592 24782 -2536 26845
rect -757 26590 -667 26845
rect 108 25922 308 25928
rect 99 25722 108 25922
rect 308 25722 317 25922
rect 108 25716 308 25722
rect -5188 24726 -2536 24782
rect -764 23911 -674 24948
rect 303931 24358 304241 24362
rect 303920 24038 303926 24358
rect 304246 24038 304252 24358
rect 303931 24034 304241 24038
rect -5244 23855 -459 23911
rect -5244 21598 -5188 23855
rect -764 23519 -674 23855
rect 108 22922 308 22928
rect 99 22722 108 22922
rect 308 22722 317 22922
rect 108 22716 308 22722
rect -4016 21858 -736 21948
rect -4016 18618 -3926 21858
rect 303931 21358 304241 21362
rect 303920 21038 303926 21358
rect 304246 21038 304252 21358
rect 303931 21034 304241 21038
rect 302848 19472 303028 19478
rect 302848 19292 307364 19472
rect 302848 19278 303028 19292
rect 38313 19214 38563 19226
rect 19851 19189 20101 19202
rect 19851 18979 19874 19189
rect 20084 18979 20101 19189
rect 29084 19062 29304 19071
rect 13790 18930 14040 18950
rect 19851 18944 20101 18979
rect 25909 19007 26226 19029
rect 13650 18925 14040 18930
rect 7470 18887 7720 18911
rect 5317 18785 5567 18810
rect 4518 18780 5567 18785
rect 3664 18760 3984 18766
rect -5180 18510 -3805 18618
rect -5180 18496 -3926 18510
rect 2316 18440 2566 18467
rect 3660 18445 3664 18755
rect 3984 18445 3988 18755
rect 4518 18570 5333 18780
rect 5543 18570 5567 18780
rect 7470 18677 7487 18887
rect 7697 18677 7720 18887
rect 7470 18653 7720 18677
rect 10692 18831 10942 18858
rect 4518 18565 5567 18570
rect 1499 18435 2566 18440
rect 1499 18225 2333 18435
rect 2543 18225 2566 18435
rect 3664 18434 3984 18440
rect 1499 18220 2566 18225
rect -6199 17947 -5999 17956
rect -6199 17738 -5999 17747
rect 1499 16557 1719 18220
rect 2316 18209 2566 18220
rect 4518 16431 4738 18565
rect 5317 18552 5567 18565
rect 7482 16457 7702 18653
rect 10692 18621 10716 18831
rect 10926 18621 10942 18831
rect 10692 18600 10942 18621
rect 13650 18715 13806 18925
rect 14016 18715 14040 18925
rect 13650 18692 14040 18715
rect 16900 18812 17150 18825
rect 10711 16526 10931 18600
rect 13650 16450 13870 18692
rect 16900 18602 16916 18812
rect 17126 18602 17150 18812
rect 18088 18760 18408 18766
rect 16900 18567 17150 18602
rect 16911 16695 17131 18567
rect 18084 18445 18088 18755
rect 18408 18445 18412 18755
rect 18088 18434 18408 18440
rect 16747 16475 17131 16695
rect 19869 16482 20089 18944
rect 25909 18797 25948 19007
rect 26158 18797 26226 19007
rect 29075 18842 29084 19052
rect 29304 18842 29313 19052
rect 35298 19051 35585 19066
rect 32333 18987 32543 18991
rect 32124 18982 32548 18987
rect 25909 18763 26226 18797
rect 22872 18654 23189 18673
rect 22872 18444 22902 18654
rect 23112 18444 23189 18654
rect 22872 18407 23189 18444
rect 22897 16457 23117 18407
rect 25943 16450 26163 18763
rect 29084 16482 29304 18842
rect 32124 18772 32333 18982
rect 32543 18772 32548 18982
rect 35298 18841 35333 19051
rect 35543 18841 35585 19051
rect 38313 19004 38333 19214
rect 38543 19004 38563 19214
rect 56594 19158 56844 19179
rect 38313 18968 38563 19004
rect 47318 19126 47568 19145
rect 35298 18828 35585 18841
rect 32124 18767 32548 18772
rect 32124 18763 32543 18767
rect 32124 16526 32344 18763
rect 32914 18760 33234 18766
rect 32910 18445 32914 18755
rect 33234 18445 33238 18755
rect 32914 18434 33234 18440
rect 35328 17249 35548 18828
rect 35196 17029 35548 17249
rect 35196 16482 35416 17029
rect 38328 16513 38548 18968
rect 44320 18919 44570 18936
rect 41318 18868 41568 18892
rect 41318 18658 41333 18868
rect 41543 18658 41568 18868
rect 44320 18709 44333 18919
rect 44543 18709 44570 18919
rect 47318 18916 47333 19126
rect 47543 18916 47568 19126
rect 53520 19038 53770 19065
rect 47318 18887 47568 18916
rect 50500 19007 50750 19023
rect 44320 18678 44570 18709
rect 41318 18634 41568 18658
rect 41328 16457 41548 18634
rect 44328 16425 44548 18678
rect 47328 17633 47548 18887
rect 50500 18797 50521 19007
rect 50731 18797 50750 19007
rect 53520 18828 53542 19038
rect 53752 18828 53770 19038
rect 56594 18948 56620 19158
rect 56830 18948 56844 19158
rect 174366 19131 174586 19136
rect 75052 19026 75347 19045
rect 108901 19028 109121 19033
rect 68555 18953 68765 18957
rect 56594 18921 56844 18948
rect 68550 18948 69258 18953
rect 53520 18807 53770 18828
rect 50500 18765 50750 18797
rect 47328 17413 47734 17633
rect 47514 16507 47734 17413
rect 50516 16475 50736 18765
rect 53537 17810 53757 18807
rect 53537 17590 53889 17810
rect 53669 16507 53889 17590
rect 56615 16444 56835 18921
rect 59609 18867 59859 18886
rect 65737 18877 66011 18893
rect 59609 18862 60001 18867
rect 59609 18652 59635 18862
rect 59845 18652 60001 18862
rect 59609 18628 60001 18652
rect 59781 16494 60001 18628
rect 62620 18791 62870 18803
rect 62620 18786 62997 18791
rect 62620 18576 62637 18786
rect 62847 18576 62997 18786
rect 64256 18760 64576 18766
rect 62620 18545 62997 18576
rect 62777 16469 62997 18545
rect 64252 18445 64256 18755
rect 64576 18445 64580 18755
rect 65737 18667 65747 18877
rect 65957 18667 66011 18877
rect 68550 18738 68555 18948
rect 68765 18738 69258 18948
rect 75052 18816 75083 19026
rect 75293 18816 75347 19026
rect 96453 18871 96673 18876
rect 90412 18833 90632 18838
rect 75052 18783 75347 18816
rect 68550 18733 69258 18738
rect 68555 18729 68765 18733
rect 65737 18611 66011 18667
rect 64256 18434 64576 18440
rect 65947 16499 66003 18611
rect 69038 16506 69258 18733
rect 71928 18520 72148 18525
rect 71924 18310 71933 18520
rect 72143 18310 72152 18520
rect 71928 17006 72148 18310
rect 71928 16786 72278 17006
rect 72058 16506 72278 16786
rect 75078 16417 75298 18783
rect 81190 18706 81410 18711
rect 81186 18496 81195 18706
rect 81405 18496 81414 18706
rect 90408 18623 90417 18833
rect 90627 18623 90636 18833
rect 93556 18789 93776 18794
rect 78103 18082 78313 18086
rect 78098 18077 78318 18082
rect 78098 17867 78103 18077
rect 78313 17867 78318 18077
rect 78098 17154 78318 17867
rect 78098 16934 78453 17154
rect 78233 16493 78453 16934
rect 81190 16478 81410 18496
rect 87335 18310 87555 18315
rect 87331 18100 87340 18310
rect 87550 18100 87559 18310
rect 84274 17980 84494 17985
rect 84270 17770 84279 17980
rect 84489 17770 84498 17980
rect 84274 16493 84494 17770
rect 87335 16380 87555 18100
rect 90412 16440 90632 18623
rect 93552 18579 93561 18789
rect 93771 18579 93780 18789
rect 96449 18661 96458 18871
rect 96668 18661 96677 18871
rect 108897 18818 108906 19028
rect 109116 18818 109125 19028
rect 157843 18993 158063 18998
rect 114953 18980 115173 18985
rect 111948 18931 112168 18936
rect 105675 18751 105895 18756
rect 102711 18736 102931 18741
rect 93556 16448 93776 18579
rect 96453 17027 96673 18661
rect 102707 18526 102716 18736
rect 102926 18526 102935 18736
rect 105671 18541 105680 18751
rect 105890 18541 105899 18751
rect 99602 18502 99812 18506
rect 99597 18497 99817 18502
rect 99597 18287 99602 18497
rect 99812 18287 99817 18497
rect 96453 16807 96815 17027
rect 96595 16478 96815 16807
rect 99597 16515 99817 18287
rect 102711 16410 102931 18526
rect 105675 16997 105895 18541
rect 105675 16777 106015 16997
rect 105795 16463 106015 16777
rect 108901 16455 109121 18818
rect 111944 18721 111953 18931
rect 112163 18721 112172 18931
rect 114949 18770 114958 18980
rect 115168 18770 115177 18980
rect 117961 18973 118202 18992
rect 111948 16515 112168 18721
rect 114953 16453 115173 18770
rect 117961 18763 117973 18973
rect 118183 18763 118202 18973
rect 127241 18938 127461 18943
rect 117961 18747 118202 18763
rect 121128 18860 121383 18878
rect 117968 17905 118188 18747
rect 121128 18650 121155 18860
rect 121365 18650 121383 18860
rect 124118 18852 124338 18861
rect 124114 18842 124118 18847
rect 121678 18760 121998 18766
rect 121128 18614 121383 18650
rect 117968 17685 118369 17905
rect 118149 16483 118369 17685
rect 121150 16461 121370 18614
rect 121674 18445 121678 18755
rect 121998 18445 122002 18755
rect 124109 18632 124118 18842
rect 124338 18842 124342 18847
rect 124338 18632 124347 18842
rect 127237 18728 127246 18938
rect 127456 18728 127465 18938
rect 133412 18867 133632 18876
rect 133408 18857 133412 18862
rect 130250 18809 130470 18814
rect 121678 18434 121998 18440
rect 124118 16552 124338 18632
rect 127241 16461 127461 18728
rect 130246 18599 130255 18809
rect 130465 18599 130474 18809
rect 133403 18647 133412 18857
rect 133632 18857 133636 18862
rect 133632 18647 133641 18857
rect 154792 18854 155012 18859
rect 145578 18839 145798 18844
rect 148754 18839 148974 18844
rect 142599 18664 142819 18669
rect 130250 16476 130470 18599
rect 133412 16461 133632 18647
rect 139552 18596 139772 18601
rect 139548 18386 139557 18596
rect 139767 18386 139776 18596
rect 142595 18454 142604 18664
rect 142814 18454 142823 18664
rect 145574 18629 145583 18839
rect 145793 18629 145802 18839
rect 148750 18629 148759 18839
rect 148969 18629 148978 18839
rect 151772 18770 151992 18775
rect 136467 18237 136687 18242
rect 136463 18027 136472 18237
rect 136682 18027 136691 18237
rect 136467 16400 136687 18027
rect 139552 16484 139772 18386
rect 142599 16468 142819 18454
rect 145578 16947 145798 18629
rect 145578 16727 145919 16947
rect 145699 16453 145919 16727
rect 148754 16407 148974 18629
rect 151768 18560 151777 18770
rect 151987 18560 151996 18770
rect 154788 18644 154797 18854
rect 155007 18644 155016 18854
rect 157839 18783 157848 18993
rect 158058 18783 158067 18993
rect 174362 18921 174371 19131
rect 174581 18921 174590 19131
rect 305385 19095 305605 19100
rect 290333 18956 290543 18960
rect 290328 18951 293619 18956
rect 229658 18935 229878 18940
rect 151772 16372 151992 18560
rect 154792 17614 155012 18644
rect 154792 17394 155166 17614
rect 154946 16464 155166 17394
rect 157843 17038 158063 18783
rect 167548 18760 167868 18766
rect 160886 18754 161106 18759
rect 160882 18544 160891 18754
rect 161101 18544 161110 18754
rect 160886 17192 161106 18544
rect 163243 18460 163453 18464
rect 163238 18455 164319 18460
rect 163238 18245 163243 18455
rect 163453 18245 164319 18455
rect 167544 18445 167548 18755
rect 167868 18445 167872 18755
rect 173066 18485 173336 18534
rect 167548 18434 167868 18440
rect 163238 18240 164319 18245
rect 163243 18236 163453 18240
rect 164099 17689 164319 18240
rect 173066 18275 173087 18485
rect 173297 18275 173336 18485
rect 173066 18238 173336 18275
rect 165933 18175 166143 18179
rect 165928 18170 167323 18175
rect 165928 17960 165933 18170
rect 166143 17960 167323 18170
rect 165928 17955 167323 17960
rect 165933 17951 166143 17955
rect 164053 17333 164319 17689
rect 157843 16818 158225 17038
rect 160886 16972 161245 17192
rect 158005 16495 158225 16818
rect 161025 16541 161245 16972
rect 164053 16441 164273 17333
rect 167103 16441 167323 17955
rect 173082 17607 173302 18238
rect 168868 17422 169078 17426
rect 168863 17417 170482 17422
rect 168863 17207 168868 17417
rect 169078 17207 170482 17417
rect 173082 17387 173510 17607
rect 168863 17202 170482 17207
rect 168868 17198 169078 17202
rect 170262 16503 170482 17202
rect 173290 16464 173510 17387
rect 174366 17560 174586 18921
rect 176311 18813 176564 18823
rect 176311 18808 179212 18813
rect 176311 18598 176333 18808
rect 176543 18598 179212 18808
rect 180548 18760 180868 18766
rect 189548 18760 189868 18766
rect 198548 18760 198868 18766
rect 204548 18760 204868 18766
rect 211548 18760 211868 18766
rect 223548 18760 223868 18766
rect 176311 18593 179212 18598
rect 176311 18578 176564 18593
rect 174366 17340 176668 17560
rect 176448 16457 176668 17340
rect 178992 17291 179212 18593
rect 180544 18445 180548 18755
rect 180868 18445 180872 18755
rect 189544 18445 189548 18755
rect 189868 18445 189872 18755
rect 198544 18445 198548 18755
rect 198868 18445 198872 18755
rect 204544 18445 204548 18755
rect 204868 18445 204872 18755
rect 206333 18456 206543 18460
rect 206328 18451 208700 18456
rect 180548 18434 180868 18440
rect 189548 18434 189868 18440
rect 198548 18434 198868 18440
rect 204548 18434 204868 18440
rect 206328 18241 206333 18451
rect 206543 18241 208700 18451
rect 211544 18445 211548 18755
rect 211868 18445 211872 18755
rect 215333 18564 215543 18568
rect 215328 18559 219617 18564
rect 211548 18434 211868 18440
rect 215328 18349 215333 18559
rect 215543 18349 219617 18559
rect 223544 18445 223548 18755
rect 223868 18445 223872 18755
rect 229654 18725 229663 18935
rect 229873 18725 229882 18935
rect 232548 18760 232868 18766
rect 238548 18760 238868 18766
rect 250548 18760 250868 18766
rect 263948 18760 264268 18766
rect 269948 18760 270268 18766
rect 272948 18760 273268 18766
rect 275948 18760 276268 18766
rect 281948 18760 282268 18766
rect 285948 18760 286268 18766
rect 223548 18434 223868 18440
rect 227194 18424 227414 18429
rect 215328 18344 219617 18349
rect 215333 18340 215543 18344
rect 206328 18236 208700 18241
rect 206333 18232 206543 18236
rect 185333 18037 185543 18041
rect 185328 18032 188126 18037
rect 182473 17855 182693 17860
rect 182469 17645 182478 17855
rect 182688 17645 182697 17855
rect 185328 17822 185333 18032
rect 185543 17822 188126 18032
rect 200915 17952 201135 17957
rect 196793 17925 197013 17930
rect 185328 17817 188126 17822
rect 185333 17813 185543 17817
rect 178992 17071 179704 17291
rect 179484 16495 179704 17071
rect 182473 16480 182693 17645
rect 184015 17153 184225 17157
rect 184010 17148 185875 17153
rect 184010 16938 184015 17148
rect 184225 16938 185875 17148
rect 184010 16933 185875 16938
rect 184015 16929 184225 16933
rect 185655 16457 185875 16933
rect 187906 16884 188126 17817
rect 196789 17715 196798 17925
rect 197008 17715 197017 17925
rect 200911 17742 200920 17952
rect 201130 17742 201139 17952
rect 206999 17747 207219 17752
rect 188333 17660 188543 17664
rect 188328 17655 191876 17660
rect 188328 17445 188333 17655
rect 188543 17445 191876 17655
rect 188328 17440 191876 17445
rect 188333 17436 188543 17440
rect 187906 16664 188841 16884
rect 188621 16449 188841 16664
rect 191656 16487 191876 17440
rect 193470 17020 193680 17024
rect 196793 17020 197013 17715
rect 193465 17015 195050 17020
rect 193465 16805 193470 17015
rect 193680 16805 195050 17015
rect 193465 16800 195050 16805
rect 196793 16800 198137 17020
rect 193470 16796 193680 16800
rect 194830 16452 195050 16800
rect 197917 16381 198137 16800
rect 200915 16470 201135 17742
rect 206995 17537 207004 17747
rect 207214 17537 207223 17747
rect 202008 16895 202218 16899
rect 202003 16890 204257 16895
rect 202003 16680 202008 16890
rect 202218 16680 204257 16890
rect 202003 16675 204257 16680
rect 202008 16671 202218 16675
rect 204037 16515 204257 16675
rect 206999 16523 207219 17537
rect 208480 17091 208700 18236
rect 213155 18094 213375 18099
rect 213151 17884 213160 18094
rect 213370 17884 213379 18094
rect 208480 16871 210431 17091
rect 210211 16506 210431 16871
rect 213155 16434 213375 17884
rect 213909 17270 214119 17274
rect 213904 17265 216497 17270
rect 213904 17055 213909 17265
rect 214119 17055 216497 17265
rect 213904 17050 216497 17055
rect 213909 17046 214119 17050
rect 216277 16372 216497 17050
rect 219397 16435 219617 18344
rect 227190 18214 227199 18424
rect 227409 18214 227418 18424
rect 221333 17712 221543 17716
rect 221328 17707 225720 17712
rect 221328 17497 221333 17707
rect 221543 17497 225720 17707
rect 221328 17492 225720 17497
rect 221333 17488 221543 17492
rect 220693 17229 220903 17233
rect 220688 17224 222682 17229
rect 220688 17014 220693 17224
rect 220903 17014 222682 17224
rect 220688 17009 222682 17014
rect 220693 17005 220903 17009
rect 222462 16426 222682 17009
rect 225500 16498 225720 17492
rect 227194 17524 227414 18214
rect 227194 17304 228839 17524
rect 228619 16480 228839 17304
rect 229658 17435 229878 18725
rect 232544 18445 232548 18755
rect 232868 18445 232872 18755
rect 233333 18690 233543 18694
rect 233328 18685 237602 18690
rect 233328 18475 233333 18685
rect 233543 18681 237602 18685
rect 233543 18475 237949 18681
rect 233328 18470 237949 18475
rect 233333 18466 233543 18470
rect 237356 18461 237949 18470
rect 232548 18434 232868 18440
rect 234650 18299 235040 18304
rect 234646 18089 234655 18299
rect 234865 18089 235040 18299
rect 234650 18084 235040 18089
rect 229658 17215 231877 17435
rect 231657 16542 231877 17215
rect 234820 16507 235040 18084
rect 237729 17961 237949 18461
rect 238544 18445 238548 18755
rect 238868 18445 238872 18755
rect 242333 18571 242543 18575
rect 242328 18566 245088 18571
rect 241672 18530 241892 18535
rect 238548 18434 238868 18440
rect 241668 18320 241677 18530
rect 241887 18320 241896 18530
rect 242328 18356 242333 18566
rect 242543 18356 245088 18566
rect 250544 18445 250548 18755
rect 250868 18445 250872 18755
rect 254333 18701 254543 18705
rect 254328 18696 257537 18701
rect 253925 18505 254145 18510
rect 250548 18434 250868 18440
rect 242328 18351 245088 18356
rect 242333 18347 242543 18351
rect 240916 18011 241136 18016
rect 237706 17778 237949 17961
rect 240912 17801 240921 18011
rect 241131 17801 241140 18011
rect 237706 16426 237926 17778
rect 240916 16485 241136 17801
rect 241672 17215 241892 18320
rect 241672 16995 244150 17215
rect 243930 16321 244150 16995
rect 244868 16987 245088 18351
rect 253921 18295 253930 18505
rect 254140 18295 254149 18505
rect 254328 18486 254333 18696
rect 254543 18486 257537 18696
rect 254328 18481 257537 18486
rect 254333 18477 254543 18481
rect 249644 17861 249924 17882
rect 249644 17856 253347 17861
rect 249644 17646 249672 17856
rect 249882 17646 253347 17856
rect 249644 17641 253347 17646
rect 249644 17623 249924 17641
rect 248716 17078 248926 17082
rect 248711 17073 250269 17078
rect 244868 16767 247273 16987
rect 248711 16863 248716 17073
rect 248926 16863 250269 17073
rect 248711 16858 250269 16863
rect 248716 16854 248926 16858
rect 247053 16521 247273 16767
rect 250049 16421 250269 16858
rect 253127 16521 253347 17641
rect 253925 17355 254145 18295
rect 257317 17358 257537 18481
rect 263944 18445 263948 18755
rect 264268 18445 264272 18755
rect 269032 18556 269252 18561
rect 263948 18434 264268 18440
rect 269028 18346 269037 18556
rect 269247 18346 269256 18556
rect 269944 18445 269948 18755
rect 270268 18445 270272 18755
rect 272944 18445 272948 18755
rect 273268 18445 273272 18755
rect 275944 18445 275948 18755
rect 276268 18445 276272 18755
rect 279676 18694 279896 18699
rect 279672 18484 279681 18694
rect 279891 18484 279900 18694
rect 269948 18434 270268 18440
rect 272948 18434 273268 18440
rect 275948 18434 276268 18440
rect 261049 18126 261259 18130
rect 261044 18121 265648 18126
rect 261044 17911 261049 18121
rect 261259 17911 265648 18121
rect 265875 17964 266085 17968
rect 261044 17906 265648 17911
rect 261049 17902 261259 17906
rect 259367 17358 259587 17386
rect 253925 17135 256417 17355
rect 257317 17138 259608 17358
rect 260058 17247 260268 17251
rect 260053 17242 262607 17247
rect 256197 16439 256417 17135
rect 259367 16507 259587 17138
rect 260053 17032 260058 17242
rect 260268 17032 262607 17242
rect 260053 17027 262607 17032
rect 260058 17023 260268 17027
rect 262387 16480 262607 17027
rect 265428 16438 265648 17906
rect 265870 17959 267379 17964
rect 265870 17749 265875 17959
rect 266085 17749 267379 17959
rect 265870 17744 267379 17749
rect 265875 17740 266085 17744
rect 267159 17371 267379 17744
rect 267159 17151 268752 17371
rect 267159 17148 267379 17151
rect 268532 16389 268752 17151
rect 269032 17090 269252 18346
rect 269333 18269 269543 18273
rect 269328 18264 274813 18269
rect 269328 18054 269333 18264
rect 269543 18054 274813 18264
rect 278878 18202 279098 18207
rect 269328 18049 274813 18054
rect 269333 18045 269543 18049
rect 269032 16870 271810 17090
rect 271590 16406 271810 16870
rect 274593 16503 274813 18049
rect 278874 17992 278883 18202
rect 279093 17992 279102 18202
rect 277693 17578 277913 17583
rect 277689 17368 277698 17578
rect 277908 17368 277917 17578
rect 277693 16482 277913 17368
rect 278878 17146 279098 17992
rect 279676 17916 279896 18484
rect 281944 18445 281948 18755
rect 282268 18445 282272 18755
rect 285944 18445 285948 18755
rect 286268 18445 286272 18755
rect 290328 18741 290333 18951
rect 290543 18741 293619 18951
rect 305381 18885 305390 19095
rect 305600 18885 305609 19095
rect 293948 18760 294268 18766
rect 296948 18760 297268 18766
rect 299948 18760 300268 18766
rect 302948 18760 303268 18766
rect 290328 18736 293619 18741
rect 290333 18732 290543 18736
rect 281948 18434 282268 18440
rect 285948 18434 286268 18440
rect 292407 18223 292627 18228
rect 284333 18138 284543 18142
rect 284328 18133 287822 18138
rect 284328 17923 284333 18133
rect 284543 17923 287822 18133
rect 292403 18013 292412 18223
rect 292622 18013 292631 18223
rect 284328 17918 287822 17923
rect 279676 17696 284112 17916
rect 284333 17914 284543 17918
rect 278878 16926 280971 17146
rect 280751 16364 280971 16926
rect 283892 16454 284112 17696
rect 286929 17508 287149 17513
rect 286925 17298 286934 17508
rect 287144 17298 287153 17508
rect 286929 16447 287149 17298
rect 287602 16980 287822 17918
rect 287602 16760 290186 16980
rect 289966 16489 290186 16760
rect 292407 16924 292627 18013
rect 293399 17354 293619 18736
rect 293944 18445 293948 18755
rect 294268 18445 294272 18755
rect 296944 18445 296948 18755
rect 297268 18445 297272 18755
rect 299944 18445 299948 18755
rect 300268 18445 300272 18755
rect 302944 18445 302948 18755
rect 303268 18445 303272 18755
rect 293948 18434 294268 18440
rect 296948 18434 297268 18440
rect 299948 18434 300268 18440
rect 302948 18434 303268 18440
rect 299258 17719 299478 17724
rect 299254 17509 299263 17719
rect 299473 17509 299482 17719
rect 293399 17134 296406 17354
rect 292407 16704 293307 16924
rect 293087 16447 293307 16704
rect 296186 16461 296406 17134
rect 299258 16890 299478 17509
rect 300256 17106 300466 17110
rect 299147 16670 299478 16890
rect 300251 17101 302500 17106
rect 300251 16891 300256 17101
rect 300466 16891 302500 17101
rect 300251 16886 302500 16891
rect 300256 16882 300466 16886
rect 299147 16399 299367 16670
rect 302280 16510 302500 16886
rect 305385 16504 305605 18885
rect 302947 16416 303269 16425
rect 302941 16094 302947 16416
rect 303269 16094 303275 16416
rect 302947 16085 303269 16094
rect 18088 15712 18408 15721
rect 3664 15694 3984 15703
rect 108 15588 308 15597
rect 102 15388 108 15588
rect 308 15388 314 15588
rect 108 15379 308 15388
rect 3658 15374 3664 15694
rect 3984 15374 3990 15694
rect 18082 15392 18088 15712
rect 18408 15392 18414 15712
rect 121678 15710 121998 15719
rect 167548 15712 167868 15721
rect 180548 15712 180868 15721
rect 189548 15712 189868 15721
rect 198548 15712 198868 15721
rect 204548 15712 204868 15721
rect 211548 15712 211868 15721
rect 223548 15712 223868 15721
rect 232548 15712 232868 15721
rect 238548 15712 238868 15721
rect 250548 15712 250868 15721
rect 263948 15712 264268 15721
rect 269948 15712 270268 15721
rect 272948 15712 273268 15721
rect 275948 15712 276268 15721
rect 281948 15712 282268 15721
rect 285948 15712 286268 15721
rect 293948 15712 294268 15721
rect 296948 15712 297268 15721
rect 299948 15712 300268 15721
rect 302948 15712 303268 15721
rect 32914 15688 33234 15697
rect 64256 15696 64576 15705
rect 18088 15383 18408 15392
rect 3664 15365 3984 15374
rect 32908 15368 32914 15688
rect 33234 15368 33240 15688
rect 64250 15376 64256 15696
rect 64576 15376 64582 15696
rect 121672 15390 121678 15710
rect 121998 15390 122004 15710
rect 167542 15392 167548 15712
rect 167868 15392 167874 15712
rect 180542 15392 180548 15712
rect 180868 15392 180874 15712
rect 189542 15392 189548 15712
rect 189868 15392 189874 15712
rect 198542 15392 198548 15712
rect 198868 15392 198874 15712
rect 204542 15392 204548 15712
rect 204868 15392 204874 15712
rect 211542 15392 211548 15712
rect 211868 15392 211874 15712
rect 223542 15392 223548 15712
rect 223868 15392 223874 15712
rect 232542 15392 232548 15712
rect 232868 15392 232874 15712
rect 238542 15392 238548 15712
rect 238868 15392 238874 15712
rect 250542 15392 250548 15712
rect 250868 15392 250874 15712
rect 263942 15392 263948 15712
rect 264268 15392 264274 15712
rect 269942 15392 269948 15712
rect 270268 15392 270274 15712
rect 272942 15392 272948 15712
rect 273268 15392 273274 15712
rect 275942 15392 275948 15712
rect 276268 15392 276274 15712
rect 281942 15392 281948 15712
rect 282268 15392 282274 15712
rect 285942 15392 285948 15712
rect 286268 15392 286274 15712
rect 293942 15392 293948 15712
rect 294268 15392 294274 15712
rect 296942 15392 296948 15712
rect 297268 15392 297274 15712
rect 299942 15392 299948 15712
rect 300268 15392 300274 15712
rect 302942 15392 302948 15712
rect 303268 15392 303274 15712
rect 121678 15381 121998 15390
rect 167548 15383 167868 15392
rect 180548 15383 180868 15392
rect 189548 15383 189868 15392
rect 198548 15383 198868 15392
rect 204548 15383 204868 15392
rect 211548 15383 211868 15392
rect 223548 15383 223868 15392
rect 232548 15383 232868 15392
rect 238548 15383 238868 15392
rect 250548 15383 250868 15392
rect 263948 15383 264268 15392
rect 269948 15383 270268 15392
rect 272948 15383 273268 15392
rect 275948 15383 276268 15392
rect 281948 15383 282268 15392
rect 285948 15383 286268 15392
rect 293948 15383 294268 15392
rect 296948 15383 297268 15392
rect 299948 15383 300268 15392
rect 302948 15383 303268 15392
rect 32914 15359 33234 15368
rect 64256 15367 64576 15376
<< via2 >>
rect 302508 324333 302708 324533
rect 303931 321043 304241 321353
rect 108 319722 308 319922
rect 303931 318043 304241 318353
rect 108 316722 308 316922
rect 303931 315043 304241 315353
rect 108 313722 308 313922
rect 303931 312043 304241 312353
rect 108 310722 308 310922
rect 303931 309043 304241 309353
rect 108 307722 308 307922
rect 303931 306043 304241 306353
rect 108 304722 308 304922
rect 303931 303043 304241 303353
rect 108 301722 308 301922
rect 303931 300043 304241 300353
rect 108 298722 308 298922
rect 303931 297043 304241 297353
rect 108 295722 308 295922
rect 303931 294043 304241 294353
rect 108 292722 308 292922
rect 303931 291043 304241 291353
rect 108 289722 308 289922
rect 303931 288043 304241 288353
rect 108 286722 308 286922
rect 303931 285043 304241 285353
rect 108 283722 308 283922
rect 303931 282043 304241 282353
rect 108 280722 308 280922
rect 303931 279043 304241 279353
rect 108 277722 308 277922
rect 303931 276043 304241 276353
rect 108 274722 308 274922
rect 303931 273043 304241 273353
rect 108 271722 308 271922
rect 303931 270043 304241 270353
rect 108 268722 308 268922
rect 303931 267043 304241 267353
rect 108 265722 308 265922
rect 303931 264043 304241 264353
rect 108 262722 308 262922
rect 303931 261043 304241 261353
rect 108 259722 308 259922
rect 303931 258043 304241 258353
rect 108 256722 308 256922
rect 303931 255043 304241 255353
rect 108 253722 308 253922
rect 303931 252043 304241 252353
rect 108 250722 308 250922
rect 303931 249043 304241 249353
rect 108 247722 308 247922
rect 303931 246043 304241 246353
rect 108 244722 308 244922
rect 303931 243043 304241 243353
rect 108 241722 308 241922
rect 303931 240043 304241 240353
rect 108 238722 308 238922
rect 303931 237043 304241 237353
rect 108 235722 308 235922
rect 303931 234043 304241 234353
rect 108 232722 308 232922
rect 303931 231043 304241 231353
rect 108 229722 308 229922
rect 303931 228043 304241 228353
rect 108 226722 308 226922
rect 303931 225043 304241 225353
rect 108 223722 308 223922
rect 303931 222043 304241 222353
rect 108 220722 308 220922
rect 303931 219043 304241 219353
rect 108 217722 308 217922
rect 303931 216043 304241 216353
rect 108 214722 308 214922
rect 303931 213043 304241 213353
rect 108 211722 308 211922
rect 303931 210043 304241 210353
rect 108 208722 308 208922
rect 303931 207043 304241 207353
rect 108 205722 308 205922
rect 303931 204043 304241 204353
rect 108 202722 308 202922
rect 303931 201043 304241 201353
rect 108 199722 308 199922
rect 303931 198043 304241 198353
rect 108 196722 308 196922
rect 303931 195043 304241 195353
rect 108 193722 308 193922
rect 303931 192043 304241 192353
rect 108 190722 308 190922
rect 303931 189043 304241 189353
rect 108 187722 308 187922
rect 303931 186043 304241 186353
rect 108 184722 308 184922
rect 303931 183043 304241 183353
rect 108 181722 308 181922
rect 303931 180043 304241 180353
rect 108 178722 308 178922
rect 303931 177043 304241 177353
rect 108 175722 308 175922
rect 303931 174043 304241 174353
rect 108 172722 308 172922
rect 303931 171043 304241 171353
rect 108 169722 308 169922
rect 303931 168043 304241 168353
rect 108 166722 308 166922
rect 303931 165043 304241 165353
rect 108 163722 308 163922
rect 303931 162043 304241 162353
rect 108 160722 308 160922
rect 303931 159043 304241 159353
rect 108 157722 308 157922
rect 303931 156043 304241 156353
rect 108 154722 308 154922
rect 303931 153043 304241 153353
rect 108 151722 308 151922
rect 303931 150043 304241 150353
rect 108 148722 308 148922
rect 303931 147043 304241 147353
rect 108 145722 308 145922
rect 303931 144043 304241 144353
rect 108 142722 308 142922
rect 303931 141043 304241 141353
rect 108 139722 308 139922
rect 303931 138043 304241 138353
rect 108 136722 308 136922
rect 303931 135043 304241 135353
rect 108 133722 308 133922
rect 303931 132043 304241 132353
rect 108 130722 308 130922
rect 303931 129043 304241 129353
rect 108 127722 308 127922
rect 303931 126043 304241 126353
rect 108 124722 308 124922
rect 303931 123043 304241 123353
rect 108 121722 308 121922
rect 303931 120043 304241 120353
rect 108 118722 308 118922
rect 303931 117043 304241 117353
rect 108 115722 308 115922
rect 303931 114043 304241 114353
rect 108 112722 308 112922
rect 303931 111043 304241 111353
rect 108 109722 308 109922
rect 303931 108043 304241 108353
rect 108 106722 308 106922
rect 303931 105043 304241 105353
rect 108 103722 308 103922
rect 303931 102043 304241 102353
rect 108 100722 308 100922
rect 303931 99043 304241 99353
rect 108 97722 308 97922
rect 303931 96043 304241 96353
rect 108 94722 308 94922
rect 303931 93043 304241 93353
rect 108 91722 308 91922
rect 303931 90043 304241 90353
rect 108 88722 308 88922
rect 303931 87043 304241 87353
rect 108 85722 308 85922
rect 303931 84043 304241 84353
rect 108 82722 308 82922
rect 303931 81043 304241 81353
rect 108 79722 308 79922
rect 303931 78043 304241 78353
rect 108 76722 308 76922
rect 303931 75043 304241 75353
rect 108 73722 308 73922
rect 303931 72043 304241 72353
rect 108 70722 308 70922
rect 303931 69043 304241 69353
rect 108 67722 308 67922
rect 303931 66043 304241 66353
rect 108 64722 308 64922
rect 303931 63043 304241 63353
rect 108 61722 308 61922
rect 303931 60043 304241 60353
rect 108 58722 308 58922
rect 303931 57043 304241 57353
rect 108 55722 308 55922
rect 303931 54043 304241 54353
rect 108 52722 308 52922
rect 303931 51043 304241 51353
rect 108 49722 308 49922
rect 303931 48043 304241 48353
rect 108 46722 308 46922
rect 303931 45043 304241 45353
rect 108 43722 308 43922
rect 303931 42043 304241 42353
rect 108 40722 308 40922
rect 303931 39043 304241 39353
rect 108 37722 308 37922
rect 303931 36043 304241 36353
rect 108 34722 308 34922
rect 303931 33043 304241 33353
rect 108 31722 308 31922
rect 303931 30043 304241 30353
rect 108 28722 308 28922
rect 303931 27043 304241 27353
rect 108 25722 308 25922
rect 303931 24043 304241 24353
rect 108 22722 308 22922
rect 303931 21043 304241 21353
rect 19874 18979 20084 19189
rect 3669 18445 3979 18755
rect 5333 18570 5543 18780
rect 7487 18677 7697 18887
rect 2333 18225 2543 18435
rect -6199 17747 -5999 17947
rect 10716 18621 10926 18831
rect 13806 18715 14016 18925
rect 16916 18602 17126 18812
rect 18093 18445 18403 18755
rect 25948 18797 26158 19007
rect 29084 18842 29304 19062
rect 22902 18444 23112 18654
rect 32333 18772 32543 18982
rect 35333 18841 35543 19051
rect 38333 19004 38543 19214
rect 32919 18445 33229 18755
rect 41333 18658 41543 18868
rect 44333 18709 44543 18919
rect 47333 18916 47543 19126
rect 50521 18797 50731 19007
rect 53542 18828 53752 19038
rect 56620 18948 56830 19158
rect 59635 18652 59845 18862
rect 62637 18576 62847 18786
rect 64261 18445 64571 18755
rect 65747 18667 65957 18877
rect 68555 18738 68765 18948
rect 75083 18816 75293 19026
rect 71933 18310 72143 18520
rect 81195 18496 81405 18706
rect 90417 18623 90627 18833
rect 78103 17867 78313 18077
rect 87340 18100 87550 18310
rect 84279 17770 84489 17980
rect 93561 18579 93771 18789
rect 96458 18661 96668 18871
rect 108906 18818 109116 19028
rect 102716 18526 102926 18736
rect 105680 18541 105890 18751
rect 99602 18287 99812 18497
rect 111953 18721 112163 18931
rect 114958 18770 115168 18980
rect 117973 18763 118183 18973
rect 121155 18650 121365 18860
rect 121683 18445 121993 18755
rect 124118 18632 124338 18852
rect 127246 18728 127456 18938
rect 130255 18599 130465 18809
rect 133412 18647 133632 18867
rect 139557 18386 139767 18596
rect 142604 18454 142814 18664
rect 145583 18629 145793 18839
rect 148759 18629 148969 18839
rect 136472 18027 136682 18237
rect 151777 18560 151987 18770
rect 154797 18644 155007 18854
rect 157848 18783 158058 18993
rect 174371 18921 174581 19131
rect 160891 18544 161101 18754
rect 163243 18245 163453 18455
rect 167553 18445 167863 18755
rect 173087 18275 173297 18485
rect 165933 17960 166143 18170
rect 168868 17207 169078 17417
rect 176333 18598 176543 18808
rect 180553 18445 180863 18755
rect 189553 18445 189863 18755
rect 198553 18445 198863 18755
rect 204553 18445 204863 18755
rect 206333 18241 206543 18451
rect 211553 18445 211863 18755
rect 215333 18349 215543 18559
rect 223553 18445 223863 18755
rect 229663 18725 229873 18935
rect 182478 17645 182688 17855
rect 185333 17822 185543 18032
rect 184015 16938 184225 17148
rect 196798 17715 197008 17925
rect 200920 17742 201130 17952
rect 188333 17445 188543 17655
rect 193470 16805 193680 17015
rect 207004 17537 207214 17747
rect 202008 16680 202218 16890
rect 213160 17884 213370 18094
rect 213909 17055 214119 17265
rect 227199 18214 227409 18424
rect 221333 17497 221543 17707
rect 220693 17014 220903 17224
rect 232553 18445 232863 18755
rect 233333 18475 233543 18685
rect 234655 18089 234865 18299
rect 238553 18445 238863 18755
rect 241677 18320 241887 18530
rect 242333 18356 242543 18566
rect 250553 18445 250863 18755
rect 240921 17801 241131 18011
rect 253930 18295 254140 18505
rect 254333 18486 254543 18696
rect 249672 17646 249882 17856
rect 248716 16863 248926 17073
rect 263953 18445 264263 18755
rect 269037 18346 269247 18556
rect 269953 18445 270263 18755
rect 272953 18445 273263 18755
rect 275953 18445 276263 18755
rect 279681 18484 279891 18694
rect 261049 17911 261259 18121
rect 260058 17032 260268 17242
rect 265875 17749 266085 17959
rect 269333 18054 269543 18264
rect 278883 17992 279093 18202
rect 277698 17368 277908 17578
rect 281953 18445 282263 18755
rect 285953 18445 286263 18755
rect 290333 18741 290543 18951
rect 305390 18885 305600 19095
rect 284333 17923 284543 18133
rect 292412 18013 292622 18223
rect 286934 17298 287144 17508
rect 293953 18445 294263 18755
rect 296953 18445 297263 18755
rect 299953 18445 300263 18755
rect 302953 18445 303263 18755
rect 299263 17509 299473 17719
rect 300256 16891 300466 17101
rect 302947 16094 303269 16416
rect 108 15388 308 15588
rect 3664 15374 3984 15694
rect 18088 15392 18408 15712
rect 32914 15368 33234 15688
rect 64256 15376 64576 15696
rect 121678 15390 121998 15710
rect 167548 15392 167868 15712
rect 180548 15392 180868 15712
rect 189548 15392 189868 15712
rect 198548 15392 198868 15712
rect 204548 15392 204868 15712
rect 211548 15392 211868 15712
rect 223548 15392 223868 15712
rect 232548 15392 232868 15712
rect 238548 15392 238868 15712
rect 250548 15392 250868 15712
rect 263948 15392 264268 15712
rect 269948 15392 270268 15712
rect 272948 15392 273268 15712
rect 275948 15392 276268 15712
rect 281948 15392 282268 15712
rect 285948 15392 286268 15712
rect 293948 15392 294268 15712
rect 296948 15392 297268 15712
rect 299948 15392 300268 15712
rect 302948 15392 303268 15712
<< metal3 >>
rect 908 322281 998 327367
rect 302503 324538 302713 324544
rect 302503 324333 302508 324338
rect 302708 324333 302713 324338
rect 302503 324328 302713 324333
rect 303927 321358 304245 321363
rect 303926 321357 304246 321358
rect 303926 321039 303927 321357
rect 304245 321039 304246 321357
rect 303926 321038 304246 321039
rect 303927 321033 304245 321038
rect 103 319922 313 319927
rect -2012 319722 -2006 319922
rect -1806 319722 108 319922
rect 308 319722 313 319922
rect 103 319717 313 319722
rect 303927 318358 304245 318363
rect 303926 318357 304246 318358
rect 303926 318039 303927 318357
rect 304245 318039 304246 318357
rect 303926 318038 304246 318039
rect 303927 318033 304245 318038
rect 103 316922 313 316927
rect -2012 316722 -2006 316922
rect -1806 316722 108 316922
rect 308 316722 313 316922
rect 103 316717 313 316722
rect 303927 315358 304245 315363
rect 303926 315357 304246 315358
rect 303926 315039 303927 315357
rect 304245 315039 304246 315357
rect 303926 315038 304246 315039
rect 303927 315033 304245 315038
rect 103 313922 313 313927
rect -2012 313722 -2006 313922
rect -1806 313722 108 313922
rect 308 313722 313 313922
rect 103 313717 313 313722
rect 303927 312358 304245 312363
rect 303926 312357 304246 312358
rect 303926 312039 303927 312357
rect 304245 312039 304246 312357
rect 303926 312038 304246 312039
rect 303927 312033 304245 312038
rect 103 310922 313 310927
rect -2012 310722 -2006 310922
rect -1806 310722 108 310922
rect 308 310722 313 310922
rect 103 310717 313 310722
rect 303927 309358 304245 309363
rect 303926 309357 304246 309358
rect 303926 309039 303927 309357
rect 304245 309039 304246 309357
rect 303926 309038 304246 309039
rect 303927 309033 304245 309038
rect 103 307922 313 307927
rect -2012 307722 -2006 307922
rect -1806 307722 108 307922
rect 308 307722 313 307922
rect 103 307717 313 307722
rect 303927 306358 304245 306363
rect 303926 306357 304246 306358
rect 303926 306039 303927 306357
rect 304245 306039 304246 306357
rect 303926 306038 304246 306039
rect 303927 306033 304245 306038
rect 103 304922 313 304927
rect -2012 304722 -2006 304922
rect -1806 304722 108 304922
rect 308 304722 313 304922
rect 103 304717 313 304722
rect 303927 303358 304245 303363
rect 303926 303357 304246 303358
rect 303926 303039 303927 303357
rect 304245 303039 304246 303357
rect 303926 303038 304246 303039
rect 303927 303033 304245 303038
rect 103 301922 313 301927
rect -2012 301722 -2006 301922
rect -1806 301722 108 301922
rect 308 301722 313 301922
rect 103 301717 313 301722
rect 303927 300358 304245 300363
rect 303926 300357 304246 300358
rect 303926 300039 303927 300357
rect 304245 300039 304246 300357
rect 303926 300038 304246 300039
rect 303927 300033 304245 300038
rect 103 298922 313 298927
rect -2012 298722 -2006 298922
rect -1806 298722 108 298922
rect 308 298722 313 298922
rect 103 298717 313 298722
rect 303927 297358 304245 297363
rect 303926 297357 304246 297358
rect 303926 297039 303927 297357
rect 304245 297039 304246 297357
rect 303926 297038 304246 297039
rect 303927 297033 304245 297038
rect 103 295922 313 295927
rect -2012 295722 -2006 295922
rect -1806 295722 108 295922
rect 308 295722 313 295922
rect 103 295717 313 295722
rect 303927 294358 304245 294363
rect 303926 294357 304246 294358
rect 303926 294039 303927 294357
rect 304245 294039 304246 294357
rect 303926 294038 304246 294039
rect 303927 294033 304245 294038
rect 103 292922 313 292927
rect -2012 292722 -2006 292922
rect -1806 292722 108 292922
rect 308 292722 313 292922
rect 103 292717 313 292722
rect 303927 291358 304245 291363
rect 303926 291357 304246 291358
rect 303926 291039 303927 291357
rect 304245 291039 304246 291357
rect 303926 291038 304246 291039
rect 303927 291033 304245 291038
rect 103 289922 313 289927
rect -2012 289722 -2006 289922
rect -1806 289722 108 289922
rect 308 289722 313 289922
rect 103 289717 313 289722
rect 303927 288358 304245 288363
rect 303926 288357 304246 288358
rect 303926 288039 303927 288357
rect 304245 288039 304246 288357
rect 303926 288038 304246 288039
rect 303927 288033 304245 288038
rect 103 286922 313 286927
rect -2012 286722 -2006 286922
rect -1806 286722 108 286922
rect 308 286722 313 286922
rect 103 286717 313 286722
rect 303927 285358 304245 285363
rect 303926 285357 304246 285358
rect 303926 285039 303927 285357
rect 304245 285039 304246 285357
rect 303926 285038 304246 285039
rect 303927 285033 304245 285038
rect 103 283922 313 283927
rect -2012 283722 -2006 283922
rect -1806 283722 108 283922
rect 308 283722 313 283922
rect 103 283717 313 283722
rect 303927 282358 304245 282363
rect 303926 282357 304246 282358
rect 303926 282039 303927 282357
rect 304245 282039 304246 282357
rect 303926 282038 304246 282039
rect 303927 282033 304245 282038
rect 103 280922 313 280927
rect -2012 280722 -2006 280922
rect -1806 280722 108 280922
rect 308 280722 313 280922
rect 103 280717 313 280722
rect 303927 279358 304245 279363
rect 303926 279357 304246 279358
rect 303926 279039 303927 279357
rect 304245 279039 304246 279357
rect 303926 279038 304246 279039
rect 303927 279033 304245 279038
rect 103 277922 313 277927
rect -2012 277722 -2006 277922
rect -1806 277722 108 277922
rect 308 277722 313 277922
rect 103 277717 313 277722
rect 303927 276358 304245 276363
rect 303926 276357 304246 276358
rect 303926 276039 303927 276357
rect 304245 276039 304246 276357
rect 303926 276038 304246 276039
rect 303927 276033 304245 276038
rect 103 274922 313 274927
rect -2012 274722 -2006 274922
rect -1806 274722 108 274922
rect 308 274722 313 274922
rect 103 274717 313 274722
rect 303927 273358 304245 273363
rect 303926 273357 304246 273358
rect 303926 273039 303927 273357
rect 304245 273039 304246 273357
rect 303926 273038 304246 273039
rect 303927 273033 304245 273038
rect 103 271922 313 271927
rect -2012 271722 -2006 271922
rect -1806 271722 108 271922
rect 308 271722 313 271922
rect 103 271717 313 271722
rect 303927 270358 304245 270363
rect 303926 270357 304246 270358
rect 303926 270039 303927 270357
rect 304245 270039 304246 270357
rect 303926 270038 304246 270039
rect 303927 270033 304245 270038
rect 103 268922 313 268927
rect -2012 268722 -2006 268922
rect -1806 268722 108 268922
rect 308 268722 313 268922
rect 103 268717 313 268722
rect 303927 267358 304245 267363
rect 303926 267357 304246 267358
rect 303926 267039 303927 267357
rect 304245 267039 304246 267357
rect 303926 267038 304246 267039
rect 303927 267033 304245 267038
rect 103 265922 313 265927
rect -2012 265722 -2006 265922
rect -1806 265722 108 265922
rect 308 265722 313 265922
rect 103 265717 313 265722
rect 303927 264358 304245 264363
rect 303926 264357 304246 264358
rect 303926 264039 303927 264357
rect 304245 264039 304246 264357
rect 303926 264038 304246 264039
rect 303927 264033 304245 264038
rect 103 262922 313 262927
rect -2012 262722 -2006 262922
rect -1806 262722 108 262922
rect 308 262722 313 262922
rect 103 262717 313 262722
rect 303927 261358 304245 261363
rect 303926 261357 304246 261358
rect 303926 261039 303927 261357
rect 304245 261039 304246 261357
rect 303926 261038 304246 261039
rect 303927 261033 304245 261038
rect 103 259922 313 259927
rect -2012 259722 -2006 259922
rect -1806 259722 108 259922
rect 308 259722 313 259922
rect 103 259717 313 259722
rect 303927 258358 304245 258363
rect 303926 258357 304246 258358
rect 303926 258039 303927 258357
rect 304245 258039 304246 258357
rect 303926 258038 304246 258039
rect 303927 258033 304245 258038
rect 103 256922 313 256927
rect -2012 256722 -2006 256922
rect -1806 256722 108 256922
rect 308 256722 313 256922
rect 103 256717 313 256722
rect 303927 255358 304245 255363
rect 303926 255357 304246 255358
rect 303926 255039 303927 255357
rect 304245 255039 304246 255357
rect 303926 255038 304246 255039
rect 303927 255033 304245 255038
rect 103 253922 313 253927
rect -2012 253722 -2006 253922
rect -1806 253722 108 253922
rect 308 253722 313 253922
rect 103 253717 313 253722
rect 303927 252358 304245 252363
rect 303926 252357 304246 252358
rect 303926 252039 303927 252357
rect 304245 252039 304246 252357
rect 303926 252038 304246 252039
rect 303927 252033 304245 252038
rect 103 250922 313 250927
rect -2012 250722 -2006 250922
rect -1806 250722 108 250922
rect 308 250722 313 250922
rect 103 250717 313 250722
rect 303927 249358 304245 249363
rect 303926 249357 304246 249358
rect 303926 249039 303927 249357
rect 304245 249039 304246 249357
rect 303926 249038 304246 249039
rect 303927 249033 304245 249038
rect 103 247922 313 247927
rect -2012 247722 -2006 247922
rect -1806 247722 108 247922
rect 308 247722 313 247922
rect 103 247717 313 247722
rect 303927 246358 304245 246363
rect 303926 246357 304246 246358
rect 303926 246039 303927 246357
rect 304245 246039 304246 246357
rect 303926 246038 304246 246039
rect 303927 246033 304245 246038
rect 103 244922 313 244927
rect -2012 244722 -2006 244922
rect -1806 244722 108 244922
rect 308 244722 313 244922
rect 103 244717 313 244722
rect 303927 243358 304245 243363
rect 303926 243357 304246 243358
rect 303926 243039 303927 243357
rect 304245 243039 304246 243357
rect 303926 243038 304246 243039
rect 303927 243033 304245 243038
rect 103 241922 313 241927
rect -2012 241722 -2006 241922
rect -1806 241722 108 241922
rect 308 241722 313 241922
rect 103 241717 313 241722
rect 303927 240358 304245 240363
rect 303926 240357 304246 240358
rect 303926 240039 303927 240357
rect 304245 240039 304246 240357
rect 303926 240038 304246 240039
rect 303927 240033 304245 240038
rect 103 238922 313 238927
rect -2012 238722 -2006 238922
rect -1806 238722 108 238922
rect 308 238722 313 238922
rect 103 238717 313 238722
rect 303927 237358 304245 237363
rect 303926 237357 304246 237358
rect 303926 237039 303927 237357
rect 304245 237039 304246 237357
rect 303926 237038 304246 237039
rect 303927 237033 304245 237038
rect 103 235922 313 235927
rect -2012 235722 -2006 235922
rect -1806 235722 108 235922
rect 308 235722 313 235922
rect 103 235717 313 235722
rect 303927 234358 304245 234363
rect 303926 234357 304246 234358
rect 303926 234039 303927 234357
rect 304245 234039 304246 234357
rect 303926 234038 304246 234039
rect 303927 234033 304245 234038
rect 103 232922 313 232927
rect -2012 232722 -2006 232922
rect -1806 232722 108 232922
rect 308 232722 313 232922
rect 103 232717 313 232722
rect 303927 231358 304245 231363
rect 303926 231357 304246 231358
rect 303926 231039 303927 231357
rect 304245 231039 304246 231357
rect 303926 231038 304246 231039
rect 303927 231033 304245 231038
rect 103 229922 313 229927
rect -2012 229722 -2006 229922
rect -1806 229722 108 229922
rect 308 229722 313 229922
rect 103 229717 313 229722
rect 303927 228358 304245 228363
rect 303926 228357 304246 228358
rect 303926 228039 303927 228357
rect 304245 228039 304246 228357
rect 303926 228038 304246 228039
rect 303927 228033 304245 228038
rect 103 226922 313 226927
rect -2012 226722 -2006 226922
rect -1806 226722 108 226922
rect 308 226722 313 226922
rect 103 226717 313 226722
rect 303927 225358 304245 225363
rect 303926 225357 304246 225358
rect 303926 225039 303927 225357
rect 304245 225039 304246 225357
rect 303926 225038 304246 225039
rect 303927 225033 304245 225038
rect 103 223922 313 223927
rect -2012 223722 -2006 223922
rect -1806 223722 108 223922
rect 308 223722 313 223922
rect 103 223717 313 223722
rect 303927 222358 304245 222363
rect 303926 222357 304246 222358
rect 303926 222039 303927 222357
rect 304245 222039 304246 222357
rect 303926 222038 304246 222039
rect 303927 222033 304245 222038
rect 103 220922 313 220927
rect -2012 220722 -2006 220922
rect -1806 220722 108 220922
rect 308 220722 313 220922
rect 103 220717 313 220722
rect 303927 219358 304245 219363
rect 303926 219357 304246 219358
rect 303926 219039 303927 219357
rect 304245 219039 304246 219357
rect 303926 219038 304246 219039
rect 303927 219033 304245 219038
rect 103 217922 313 217927
rect -2012 217722 -2006 217922
rect -1806 217722 108 217922
rect 308 217722 313 217922
rect 103 217717 313 217722
rect 303927 216358 304245 216363
rect 303926 216357 304246 216358
rect 303926 216039 303927 216357
rect 304245 216039 304246 216357
rect 303926 216038 304246 216039
rect 303927 216033 304245 216038
rect 103 214922 313 214927
rect -2012 214722 -2006 214922
rect -1806 214722 108 214922
rect 308 214722 313 214922
rect 103 214717 313 214722
rect 303927 213358 304245 213363
rect 303926 213357 304246 213358
rect 303926 213039 303927 213357
rect 304245 213039 304246 213357
rect 303926 213038 304246 213039
rect 303927 213033 304245 213038
rect 103 211922 313 211927
rect -2012 211722 -2006 211922
rect -1806 211722 108 211922
rect 308 211722 313 211922
rect 103 211717 313 211722
rect 303927 210358 304245 210363
rect 303926 210357 304246 210358
rect 303926 210039 303927 210357
rect 304245 210039 304246 210357
rect 303926 210038 304246 210039
rect 303927 210033 304245 210038
rect 103 208922 313 208927
rect -2012 208722 -2006 208922
rect -1806 208722 108 208922
rect 308 208722 313 208922
rect 103 208717 313 208722
rect 303927 207358 304245 207363
rect 303926 207357 304246 207358
rect 303926 207039 303927 207357
rect 304245 207039 304246 207357
rect 303926 207038 304246 207039
rect 303927 207033 304245 207038
rect 103 205922 313 205927
rect -2012 205722 -2006 205922
rect -1806 205722 108 205922
rect 308 205722 313 205922
rect 103 205717 313 205722
rect 303927 204358 304245 204363
rect 303926 204357 304246 204358
rect 303926 204039 303927 204357
rect 304245 204039 304246 204357
rect 303926 204038 304246 204039
rect 303927 204033 304245 204038
rect 103 202922 313 202927
rect -2012 202722 -2006 202922
rect -1806 202722 108 202922
rect 308 202722 313 202922
rect 103 202717 313 202722
rect 303927 201358 304245 201363
rect 303926 201357 304246 201358
rect 303926 201039 303927 201357
rect 304245 201039 304246 201357
rect 303926 201038 304246 201039
rect 303927 201033 304245 201038
rect 103 199922 313 199927
rect -2012 199722 -2006 199922
rect -1806 199722 108 199922
rect 308 199722 313 199922
rect 103 199717 313 199722
rect 303927 198358 304245 198363
rect 303926 198357 304246 198358
rect 303926 198039 303927 198357
rect 304245 198039 304246 198357
rect 303926 198038 304246 198039
rect 303927 198033 304245 198038
rect 103 196922 313 196927
rect -2012 196722 -2006 196922
rect -1806 196722 108 196922
rect 308 196722 313 196922
rect 103 196717 313 196722
rect 303927 195358 304245 195363
rect 303926 195357 304246 195358
rect 303926 195039 303927 195357
rect 304245 195039 304246 195357
rect 303926 195038 304246 195039
rect 303927 195033 304245 195038
rect 103 193922 313 193927
rect -2012 193722 -2006 193922
rect -1806 193722 108 193922
rect 308 193722 313 193922
rect 103 193717 313 193722
rect 303927 192358 304245 192363
rect 303926 192357 304246 192358
rect 303926 192039 303927 192357
rect 304245 192039 304246 192357
rect 303926 192038 304246 192039
rect 303927 192033 304245 192038
rect 103 190922 313 190927
rect -2012 190722 -2006 190922
rect -1806 190722 108 190922
rect 308 190722 313 190922
rect 103 190717 313 190722
rect 303927 189358 304245 189363
rect 303926 189357 304246 189358
rect 303926 189039 303927 189357
rect 304245 189039 304246 189357
rect 303926 189038 304246 189039
rect 303927 189033 304245 189038
rect 103 187922 313 187927
rect -2012 187722 -2006 187922
rect -1806 187722 108 187922
rect 308 187722 313 187922
rect 103 187717 313 187722
rect 303927 186358 304245 186363
rect 303926 186357 304246 186358
rect 303926 186039 303927 186357
rect 304245 186039 304246 186357
rect 303926 186038 304246 186039
rect 303927 186033 304245 186038
rect 103 184922 313 184927
rect -2012 184722 -2006 184922
rect -1806 184722 108 184922
rect 308 184722 313 184922
rect 103 184717 313 184722
rect 303927 183358 304245 183363
rect 303926 183357 304246 183358
rect 303926 183039 303927 183357
rect 304245 183039 304246 183357
rect 303926 183038 304246 183039
rect 303927 183033 304245 183038
rect 103 181922 313 181927
rect -2012 181722 -2006 181922
rect -1806 181722 108 181922
rect 308 181722 313 181922
rect 103 181717 313 181722
rect 303927 180358 304245 180363
rect 303926 180357 304246 180358
rect 303926 180039 303927 180357
rect 304245 180039 304246 180357
rect 303926 180038 304246 180039
rect 303927 180033 304245 180038
rect 103 178922 313 178927
rect -2012 178722 -2006 178922
rect -1806 178722 108 178922
rect 308 178722 313 178922
rect 103 178717 313 178722
rect 303927 177358 304245 177363
rect 303926 177357 304246 177358
rect 303926 177039 303927 177357
rect 304245 177039 304246 177357
rect 303926 177038 304246 177039
rect 303927 177033 304245 177038
rect 103 175922 313 175927
rect -2012 175722 -2006 175922
rect -1806 175722 108 175922
rect 308 175722 313 175922
rect 103 175717 313 175722
rect 303927 174358 304245 174363
rect 303926 174357 304246 174358
rect 303926 174039 303927 174357
rect 304245 174039 304246 174357
rect 303926 174038 304246 174039
rect 303927 174033 304245 174038
rect 103 172922 313 172927
rect -2012 172722 -2006 172922
rect -1806 172722 108 172922
rect 308 172722 313 172922
rect 103 172717 313 172722
rect 303927 171358 304245 171363
rect 303926 171357 304246 171358
rect 303926 171039 303927 171357
rect 304245 171039 304246 171357
rect 303926 171038 304246 171039
rect 303927 171033 304245 171038
rect 103 169922 313 169927
rect -2012 169722 -2006 169922
rect -1806 169722 108 169922
rect 308 169722 313 169922
rect 103 169717 313 169722
rect 303927 168358 304245 168363
rect 303926 168357 304246 168358
rect 303926 168039 303927 168357
rect 304245 168039 304246 168357
rect 303926 168038 304246 168039
rect 303927 168033 304245 168038
rect 103 166922 313 166927
rect -2012 166722 -2006 166922
rect -1806 166722 108 166922
rect 308 166722 313 166922
rect 103 166717 313 166722
rect 303927 165358 304245 165363
rect 303926 165357 304246 165358
rect 303926 165039 303927 165357
rect 304245 165039 304246 165357
rect 303926 165038 304246 165039
rect 303927 165033 304245 165038
rect 103 163922 313 163927
rect -2012 163722 -2006 163922
rect -1806 163722 108 163922
rect 308 163722 313 163922
rect 103 163717 313 163722
rect 303927 162358 304245 162363
rect 303926 162357 304246 162358
rect 303926 162039 303927 162357
rect 304245 162039 304246 162357
rect 303926 162038 304246 162039
rect 303927 162033 304245 162038
rect 103 160922 313 160927
rect -2012 160722 -2006 160922
rect -1806 160722 108 160922
rect 308 160722 313 160922
rect 103 160717 313 160722
rect 303927 159358 304245 159363
rect 303926 159357 304246 159358
rect 303926 159039 303927 159357
rect 304245 159039 304246 159357
rect 303926 159038 304246 159039
rect 303927 159033 304245 159038
rect 103 157922 313 157927
rect -2012 157722 -2006 157922
rect -1806 157722 108 157922
rect 308 157722 313 157922
rect 103 157717 313 157722
rect 303927 156358 304245 156363
rect 303926 156357 304246 156358
rect 303926 156039 303927 156357
rect 304245 156039 304246 156357
rect 303926 156038 304246 156039
rect 303927 156033 304245 156038
rect 103 154922 313 154927
rect -2012 154722 -2006 154922
rect -1806 154722 108 154922
rect 308 154722 313 154922
rect 103 154717 313 154722
rect 303927 153358 304245 153363
rect 303926 153357 304246 153358
rect 303926 153039 303927 153357
rect 304245 153039 304246 153357
rect 303926 153038 304246 153039
rect 303927 153033 304245 153038
rect 103 151922 313 151927
rect -2012 151722 -2006 151922
rect -1806 151722 108 151922
rect 308 151722 313 151922
rect 103 151717 313 151722
rect 303927 150358 304245 150363
rect 303926 150357 304246 150358
rect 303926 150039 303927 150357
rect 304245 150039 304246 150357
rect 303926 150038 304246 150039
rect 303927 150033 304245 150038
rect 103 148922 313 148927
rect -2012 148722 -2006 148922
rect -1806 148722 108 148922
rect 308 148722 313 148922
rect 103 148717 313 148722
rect 303927 147358 304245 147363
rect 303926 147357 304246 147358
rect 303926 147039 303927 147357
rect 304245 147039 304246 147357
rect 303926 147038 304246 147039
rect 303927 147033 304245 147038
rect 103 145922 313 145927
rect -2012 145722 -2006 145922
rect -1806 145722 108 145922
rect 308 145722 313 145922
rect 103 145717 313 145722
rect 303927 144358 304245 144363
rect 303926 144357 304246 144358
rect 303926 144039 303927 144357
rect 304245 144039 304246 144357
rect 303926 144038 304246 144039
rect 303927 144033 304245 144038
rect 103 142922 313 142927
rect -2012 142722 -2006 142922
rect -1806 142722 108 142922
rect 308 142722 313 142922
rect 103 142717 313 142722
rect 303927 141358 304245 141363
rect 303926 141357 304246 141358
rect 303926 141039 303927 141357
rect 304245 141039 304246 141357
rect 303926 141038 304246 141039
rect 303927 141033 304245 141038
rect 103 139922 313 139927
rect -2012 139722 -2006 139922
rect -1806 139722 108 139922
rect 308 139722 313 139922
rect 103 139717 313 139722
rect 303927 138358 304245 138363
rect 303926 138357 304246 138358
rect 303926 138039 303927 138357
rect 304245 138039 304246 138357
rect 303926 138038 304246 138039
rect 303927 138033 304245 138038
rect 103 136922 313 136927
rect -2012 136722 -2006 136922
rect -1806 136722 108 136922
rect 308 136722 313 136922
rect 103 136717 313 136722
rect 303927 135358 304245 135363
rect 303926 135357 304246 135358
rect 303926 135039 303927 135357
rect 304245 135039 304246 135357
rect 303926 135038 304246 135039
rect 303927 135033 304245 135038
rect 103 133922 313 133927
rect -2012 133722 -2006 133922
rect -1806 133722 108 133922
rect 308 133722 313 133922
rect 103 133717 313 133722
rect 303927 132358 304245 132363
rect 303926 132357 304246 132358
rect 303926 132039 303927 132357
rect 304245 132039 304246 132357
rect 303926 132038 304246 132039
rect 303927 132033 304245 132038
rect 103 130922 313 130927
rect -2012 130722 -2006 130922
rect -1806 130722 108 130922
rect 308 130722 313 130922
rect 103 130717 313 130722
rect 303927 129358 304245 129363
rect 303926 129357 304246 129358
rect 303926 129039 303927 129357
rect 304245 129039 304246 129357
rect 303926 129038 304246 129039
rect 303927 129033 304245 129038
rect 103 127922 313 127927
rect -2012 127722 -2006 127922
rect -1806 127722 108 127922
rect 308 127722 313 127922
rect 103 127717 313 127722
rect 303927 126358 304245 126363
rect 303926 126357 304246 126358
rect 303926 126039 303927 126357
rect 304245 126039 304246 126357
rect 303926 126038 304246 126039
rect 303927 126033 304245 126038
rect 103 124922 313 124927
rect -2012 124722 -2006 124922
rect -1806 124722 108 124922
rect 308 124722 313 124922
rect 103 124717 313 124722
rect 303927 123358 304245 123363
rect 303926 123357 304246 123358
rect 303926 123039 303927 123357
rect 304245 123039 304246 123357
rect 303926 123038 304246 123039
rect 303927 123033 304245 123038
rect 103 121922 313 121927
rect -2012 121722 -2006 121922
rect -1806 121722 108 121922
rect 308 121722 313 121922
rect 103 121717 313 121722
rect 303927 120358 304245 120363
rect 303926 120357 304246 120358
rect 303926 120039 303927 120357
rect 304245 120039 304246 120357
rect 303926 120038 304246 120039
rect 303927 120033 304245 120038
rect 103 118922 313 118927
rect -2012 118722 -2006 118922
rect -1806 118722 108 118922
rect 308 118722 313 118922
rect 103 118717 313 118722
rect 303927 117358 304245 117363
rect 303926 117357 304246 117358
rect 303926 117039 303927 117357
rect 304245 117039 304246 117357
rect 303926 117038 304246 117039
rect 303927 117033 304245 117038
rect 103 115922 313 115927
rect -2012 115722 -2006 115922
rect -1806 115722 108 115922
rect 308 115722 313 115922
rect 103 115717 313 115722
rect 303927 114358 304245 114363
rect 303926 114357 304246 114358
rect 303926 114039 303927 114357
rect 304245 114039 304246 114357
rect 303926 114038 304246 114039
rect 303927 114033 304245 114038
rect 103 112922 313 112927
rect -2012 112722 -2006 112922
rect -1806 112722 108 112922
rect 308 112722 313 112922
rect 103 112717 313 112722
rect 303927 111358 304245 111363
rect 303926 111357 304246 111358
rect 303926 111039 303927 111357
rect 304245 111039 304246 111357
rect 303926 111038 304246 111039
rect 303927 111033 304245 111038
rect 103 109922 313 109927
rect -2012 109722 -2006 109922
rect -1806 109722 108 109922
rect 308 109722 313 109922
rect 103 109717 313 109722
rect 303927 108358 304245 108363
rect 303926 108357 304246 108358
rect 303926 108039 303927 108357
rect 304245 108039 304246 108357
rect 303926 108038 304246 108039
rect 303927 108033 304245 108038
rect 103 106922 313 106927
rect -2012 106722 -2006 106922
rect -1806 106722 108 106922
rect 308 106722 313 106922
rect 103 106717 313 106722
rect 303927 105358 304245 105363
rect 303926 105357 304246 105358
rect 303926 105039 303927 105357
rect 304245 105039 304246 105357
rect 303926 105038 304246 105039
rect 303927 105033 304245 105038
rect 103 103922 313 103927
rect -2012 103722 -2006 103922
rect -1806 103722 108 103922
rect 308 103722 313 103922
rect 103 103717 313 103722
rect 303927 102358 304245 102363
rect 303926 102357 304246 102358
rect 303926 102039 303927 102357
rect 304245 102039 304246 102357
rect 303926 102038 304246 102039
rect 303927 102033 304245 102038
rect 103 100922 313 100927
rect -2012 100722 -2006 100922
rect -1806 100722 108 100922
rect 308 100722 313 100922
rect 103 100717 313 100722
rect 303927 99358 304245 99363
rect 303926 99357 304246 99358
rect 303926 99039 303927 99357
rect 304245 99039 304246 99357
rect 303926 99038 304246 99039
rect 303927 99033 304245 99038
rect 103 97922 313 97927
rect -2012 97722 -2006 97922
rect -1806 97722 108 97922
rect 308 97722 313 97922
rect 103 97717 313 97722
rect 303927 96358 304245 96363
rect 303926 96357 304246 96358
rect 303926 96039 303927 96357
rect 304245 96039 304246 96357
rect 303926 96038 304246 96039
rect 303927 96033 304245 96038
rect 103 94922 313 94927
rect -2012 94722 -2006 94922
rect -1806 94722 108 94922
rect 308 94722 313 94922
rect 103 94717 313 94722
rect 303927 93358 304245 93363
rect 303926 93357 304246 93358
rect 303926 93039 303927 93357
rect 304245 93039 304246 93357
rect 303926 93038 304246 93039
rect 303927 93033 304245 93038
rect 103 91922 313 91927
rect -2012 91722 -2006 91922
rect -1806 91722 108 91922
rect 308 91722 313 91922
rect 103 91717 313 91722
rect 303927 90358 304245 90363
rect 303926 90357 304246 90358
rect 303926 90039 303927 90357
rect 304245 90039 304246 90357
rect 303926 90038 304246 90039
rect 303927 90033 304245 90038
rect 103 88922 313 88927
rect -2012 88722 -2006 88922
rect -1806 88722 108 88922
rect 308 88722 313 88922
rect 103 88717 313 88722
rect 303927 87358 304245 87363
rect 303926 87357 304246 87358
rect 303926 87039 303927 87357
rect 304245 87039 304246 87357
rect 303926 87038 304246 87039
rect 303927 87033 304245 87038
rect 103 85922 313 85927
rect -2012 85722 -2006 85922
rect -1806 85722 108 85922
rect 308 85722 313 85922
rect 103 85717 313 85722
rect 303927 84358 304245 84363
rect 303926 84357 304246 84358
rect 303926 84039 303927 84357
rect 304245 84039 304246 84357
rect 303926 84038 304246 84039
rect 303927 84033 304245 84038
rect 103 82922 313 82927
rect -2012 82722 -2006 82922
rect -1806 82722 108 82922
rect 308 82722 313 82922
rect 103 82717 313 82722
rect 303927 81358 304245 81363
rect 303926 81357 304246 81358
rect 303926 81039 303927 81357
rect 304245 81039 304246 81357
rect 303926 81038 304246 81039
rect 303927 81033 304245 81038
rect 103 79922 313 79927
rect -2012 79722 -2006 79922
rect -1806 79722 108 79922
rect 308 79722 313 79922
rect 103 79717 313 79722
rect 303927 78358 304245 78363
rect 303926 78357 304246 78358
rect 303926 78039 303927 78357
rect 304245 78039 304246 78357
rect 303926 78038 304246 78039
rect 303927 78033 304245 78038
rect 103 76922 313 76927
rect -2012 76722 -2006 76922
rect -1806 76722 108 76922
rect 308 76722 313 76922
rect 103 76717 313 76722
rect 303927 75358 304245 75363
rect 303926 75357 304246 75358
rect 303926 75039 303927 75357
rect 304245 75039 304246 75357
rect 303926 75038 304246 75039
rect 303927 75033 304245 75038
rect 103 73922 313 73927
rect -2012 73722 -2006 73922
rect -1806 73722 108 73922
rect 308 73722 313 73922
rect 103 73717 313 73722
rect 303927 72358 304245 72363
rect 303926 72357 304246 72358
rect 303926 72039 303927 72357
rect 304245 72039 304246 72357
rect 303926 72038 304246 72039
rect 303927 72033 304245 72038
rect 103 70922 313 70927
rect -2012 70722 -2006 70922
rect -1806 70722 108 70922
rect 308 70722 313 70922
rect 103 70717 313 70722
rect 303927 69358 304245 69363
rect 303926 69357 304246 69358
rect 303926 69039 303927 69357
rect 304245 69039 304246 69357
rect 303926 69038 304246 69039
rect 303927 69033 304245 69038
rect 103 67922 313 67927
rect -2012 67722 -2006 67922
rect -1806 67722 108 67922
rect 308 67722 313 67922
rect 103 67717 313 67722
rect 303927 66358 304245 66363
rect 303926 66357 304246 66358
rect 303926 66039 303927 66357
rect 304245 66039 304246 66357
rect 303926 66038 304246 66039
rect 303927 66033 304245 66038
rect 103 64922 313 64927
rect -2012 64722 -2006 64922
rect -1806 64722 108 64922
rect 308 64722 313 64922
rect 103 64717 313 64722
rect 303927 63358 304245 63363
rect 303926 63357 304246 63358
rect 303926 63039 303927 63357
rect 304245 63039 304246 63357
rect 303926 63038 304246 63039
rect 303927 63033 304245 63038
rect 103 61922 313 61927
rect -2012 61722 -2006 61922
rect -1806 61722 108 61922
rect 308 61722 313 61922
rect 103 61717 313 61722
rect 303927 60358 304245 60363
rect 303926 60357 304246 60358
rect 303926 60039 303927 60357
rect 304245 60039 304246 60357
rect 303926 60038 304246 60039
rect 303927 60033 304245 60038
rect 103 58922 313 58927
rect -2012 58722 -2006 58922
rect -1806 58722 108 58922
rect 308 58722 313 58922
rect 103 58717 313 58722
rect 303927 57358 304245 57363
rect 303926 57357 304246 57358
rect 303926 57039 303927 57357
rect 304245 57039 304246 57357
rect 303926 57038 304246 57039
rect 303927 57033 304245 57038
rect 103 55922 313 55927
rect -2012 55722 -2006 55922
rect -1806 55722 108 55922
rect 308 55722 313 55922
rect 103 55717 313 55722
rect 303927 54358 304245 54363
rect 303926 54357 304246 54358
rect 303926 54039 303927 54357
rect 304245 54039 304246 54357
rect 303926 54038 304246 54039
rect 303927 54033 304245 54038
rect 103 52922 313 52927
rect -2012 52722 -2006 52922
rect -1806 52722 108 52922
rect 308 52722 313 52922
rect 103 52717 313 52722
rect 303927 51358 304245 51363
rect 303926 51357 304246 51358
rect 303926 51039 303927 51357
rect 304245 51039 304246 51357
rect 303926 51038 304246 51039
rect 303927 51033 304245 51038
rect 103 49922 313 49927
rect -2012 49722 -2006 49922
rect -1806 49722 108 49922
rect 308 49722 313 49922
rect 103 49717 313 49722
rect 303927 48358 304245 48363
rect 303926 48357 304246 48358
rect 303926 48039 303927 48357
rect 304245 48039 304246 48357
rect 303926 48038 304246 48039
rect 303927 48033 304245 48038
rect 103 46922 313 46927
rect -2012 46722 -2006 46922
rect -1806 46722 108 46922
rect 308 46722 313 46922
rect 103 46717 313 46722
rect 303927 45358 304245 45363
rect 303926 45357 304246 45358
rect 303926 45039 303927 45357
rect 304245 45039 304246 45357
rect 303926 45038 304246 45039
rect 303927 45033 304245 45038
rect 103 43922 313 43927
rect -2012 43722 -2006 43922
rect -1806 43722 108 43922
rect 308 43722 313 43922
rect 103 43717 313 43722
rect 303927 42358 304245 42363
rect 303926 42357 304246 42358
rect 303926 42039 303927 42357
rect 304245 42039 304246 42357
rect 303926 42038 304246 42039
rect 303927 42033 304245 42038
rect 103 40922 313 40927
rect -2012 40722 -2006 40922
rect -1806 40722 108 40922
rect 308 40722 313 40922
rect 103 40717 313 40722
rect 303927 39358 304245 39363
rect 303926 39357 304246 39358
rect 303926 39039 303927 39357
rect 304245 39039 304246 39357
rect 303926 39038 304246 39039
rect 303927 39033 304245 39038
rect 103 37922 313 37927
rect -2012 37722 -2006 37922
rect -1806 37722 108 37922
rect 308 37722 313 37922
rect 103 37717 313 37722
rect 303927 36358 304245 36363
rect 303926 36357 304246 36358
rect 303926 36039 303927 36357
rect 304245 36039 304246 36357
rect 303926 36038 304246 36039
rect 303927 36033 304245 36038
rect 103 34922 313 34927
rect -2012 34722 -2006 34922
rect -1806 34722 108 34922
rect 308 34722 313 34922
rect 103 34717 313 34722
rect 303927 33358 304245 33363
rect 303926 33357 304246 33358
rect 303926 33039 303927 33357
rect 304245 33039 304246 33357
rect 303926 33038 304246 33039
rect 303927 33033 304245 33038
rect 103 31922 313 31927
rect -2012 31722 -2006 31922
rect -1806 31722 108 31922
rect 308 31722 313 31922
rect 103 31717 313 31722
rect 303927 30358 304245 30363
rect 303926 30357 304246 30358
rect 303926 30039 303927 30357
rect 304245 30039 304246 30357
rect 303926 30038 304246 30039
rect 303927 30033 304245 30038
rect 103 28922 313 28927
rect -2012 28722 -2006 28922
rect -1806 28722 108 28922
rect 308 28722 313 28922
rect 103 28717 313 28722
rect 303927 27358 304245 27363
rect 303926 27357 304246 27358
rect 303926 27039 303927 27357
rect 304245 27039 304246 27357
rect 303926 27038 304246 27039
rect 303927 27033 304245 27038
rect 103 25922 313 25927
rect -2012 25722 -2006 25922
rect -1806 25722 108 25922
rect 308 25722 313 25922
rect 103 25717 313 25722
rect 303927 24358 304245 24363
rect 303926 24357 304246 24358
rect 303926 24039 303927 24357
rect 304245 24039 304246 24357
rect 303926 24038 304246 24039
rect 303927 24033 304245 24038
rect 103 22922 313 22927
rect -2012 22722 -2006 22922
rect -1806 22722 108 22922
rect 308 22722 313 22922
rect 103 22717 313 22722
rect 303927 21358 304245 21363
rect 303926 21357 304246 21358
rect 303926 21039 303927 21357
rect 304245 21039 304246 21357
rect 303926 21038 304246 21039
rect 303927 21033 304245 21038
rect 38328 19218 38548 19219
rect 19870 19194 20088 19199
rect 19869 19193 20089 19194
rect 19869 18975 19870 19193
rect 20088 18975 20089 19193
rect 29079 19062 29309 19067
rect 25944 19012 26162 19017
rect 19869 18974 20089 18975
rect 25943 19011 26163 19012
rect 19870 18969 20088 18974
rect 13802 18930 14020 18935
rect 13801 18929 14021 18930
rect 7482 18891 7702 18892
rect 5329 18785 5547 18790
rect 5328 18784 5548 18785
rect 3664 18759 3984 18760
rect 3659 18441 3665 18759
rect 3983 18441 3989 18759
rect 5328 18566 5329 18784
rect 5547 18566 5548 18784
rect 7477 18673 7483 18891
rect 7701 18673 7707 18891
rect 10712 18836 10930 18841
rect 10711 18835 10931 18836
rect 7482 18672 7702 18673
rect 10711 18617 10712 18835
rect 10930 18617 10931 18835
rect 13801 18711 13802 18929
rect 14020 18711 14021 18929
rect 16912 18817 17130 18822
rect 13801 18710 14021 18711
rect 16911 18816 17131 18817
rect 13802 18705 14020 18710
rect 10711 18616 10931 18617
rect 10712 18611 10930 18616
rect 16911 18598 16912 18816
rect 17130 18598 17131 18816
rect 25943 18793 25944 19011
rect 26162 18793 26163 19011
rect 29079 18842 29084 19062
rect 29304 18842 29309 19062
rect 35328 19055 35548 19056
rect 32329 18987 32547 18992
rect 29079 18837 29309 18842
rect 32328 18986 32548 18987
rect 25943 18792 26163 18793
rect 25944 18787 26162 18792
rect 32328 18768 32329 18986
rect 32547 18768 32548 18986
rect 35323 18837 35329 19055
rect 35547 18837 35553 19055
rect 38323 19000 38329 19218
rect 38547 19000 38553 19218
rect 56616 19163 56834 19168
rect 56615 19162 56835 19163
rect 47328 19130 47548 19131
rect 38328 18999 38548 19000
rect 44328 18923 44548 18924
rect 41328 18872 41548 18873
rect 35328 18836 35548 18837
rect 32328 18767 32548 18768
rect 32329 18762 32547 18767
rect 18088 18759 18408 18760
rect 32914 18759 33234 18760
rect 16911 18597 17131 18598
rect 16912 18592 17130 18597
rect 5328 18565 5548 18566
rect 5329 18560 5547 18565
rect 18083 18441 18089 18759
rect 18407 18441 18413 18759
rect 22898 18659 23116 18664
rect 22897 18658 23117 18659
rect 3664 18440 3984 18441
rect 18088 18440 18408 18441
rect 22897 18440 22898 18658
rect 23116 18440 23117 18658
rect 32909 18441 32915 18759
rect 33233 18441 33239 18759
rect 41323 18654 41329 18872
rect 41547 18654 41553 18872
rect 44323 18705 44329 18923
rect 44547 18705 44553 18923
rect 47323 18912 47329 19130
rect 47547 18912 47553 19130
rect 53538 19043 53756 19048
rect 53537 19042 53757 19043
rect 50517 19012 50735 19017
rect 50516 19011 50736 19012
rect 47328 18911 47548 18912
rect 50516 18793 50517 19011
rect 50735 18793 50736 19011
rect 53537 18824 53538 19042
rect 53756 18824 53757 19042
rect 56615 18944 56616 19162
rect 56834 18944 56835 19162
rect 174366 19135 174586 19136
rect 71929 19061 72147 19066
rect 71928 19060 72148 19061
rect 68328 18952 68770 18953
rect 56615 18943 56835 18944
rect 56616 18938 56834 18943
rect 65743 18882 65961 18887
rect 65742 18881 65962 18882
rect 59631 18867 59849 18872
rect 53537 18823 53757 18824
rect 59630 18866 59850 18867
rect 53538 18818 53756 18823
rect 50516 18792 50736 18793
rect 50517 18787 50735 18792
rect 44328 18704 44548 18705
rect 41328 18653 41548 18654
rect 59630 18648 59631 18866
rect 59849 18648 59850 18866
rect 62633 18791 62851 18796
rect 59630 18647 59850 18648
rect 62632 18790 62852 18791
rect 59631 18642 59849 18647
rect 62632 18572 62633 18790
rect 62851 18572 62852 18790
rect 64256 18759 64576 18760
rect 62632 18571 62852 18572
rect 62633 18566 62851 18571
rect 64251 18441 64257 18759
rect 64575 18441 64581 18759
rect 65742 18663 65743 18881
rect 65961 18663 65962 18881
rect 68323 18734 68329 18952
rect 68547 18948 68770 18952
rect 68547 18738 68555 18948
rect 68765 18738 68770 18948
rect 68547 18734 68770 18738
rect 68328 18733 68770 18734
rect 71928 18842 71929 19060
rect 72147 18842 72148 19060
rect 75079 19031 75297 19036
rect 108902 19033 109120 19038
rect 108901 19032 109121 19033
rect 65742 18662 65962 18663
rect 65743 18657 65961 18662
rect 71928 18520 72148 18842
rect 75078 19030 75298 19031
rect 75078 18812 75079 19030
rect 75297 18812 75298 19030
rect 81190 18905 81410 18906
rect 75078 18811 75298 18812
rect 75079 18806 75297 18811
rect 81185 18687 81191 18905
rect 81409 18687 81415 18905
rect 96453 18875 96673 18876
rect 90412 18837 90632 18838
rect 32914 18440 33234 18441
rect 64256 18440 64576 18441
rect 2328 18439 2548 18440
rect 22897 18439 23117 18440
rect 2323 18221 2329 18439
rect 2547 18221 2553 18439
rect 22898 18434 23116 18439
rect 71928 18310 71933 18520
rect 72143 18310 72148 18520
rect 81190 18496 81195 18687
rect 81405 18496 81410 18687
rect 90407 18619 90413 18837
rect 90631 18619 90637 18837
rect 93556 18793 93776 18794
rect 90412 18618 90632 18619
rect 93551 18575 93557 18793
rect 93775 18575 93781 18793
rect 96448 18657 96454 18875
rect 96672 18657 96678 18875
rect 108901 18814 108902 19032
rect 109120 18814 109121 19032
rect 157844 18998 158062 19003
rect 157843 18997 158063 18998
rect 114954 18985 115172 18990
rect 114953 18984 115173 18985
rect 111949 18936 112167 18941
rect 108901 18813 109121 18814
rect 111948 18935 112168 18936
rect 108902 18808 109120 18813
rect 105675 18755 105895 18756
rect 102712 18741 102930 18746
rect 102711 18740 102931 18741
rect 96453 18656 96673 18657
rect 93556 18574 93776 18575
rect 102711 18522 102712 18740
rect 102930 18522 102931 18740
rect 105670 18537 105676 18755
rect 105894 18537 105900 18755
rect 111948 18717 111949 18935
rect 112167 18717 112168 18935
rect 114953 18766 114954 18984
rect 115172 18766 115173 18984
rect 117969 18978 118187 18983
rect 114953 18765 115173 18766
rect 117968 18977 118188 18978
rect 114954 18760 115172 18765
rect 117968 18759 117969 18977
rect 118187 18759 118188 18977
rect 127242 18943 127460 18948
rect 127241 18942 127461 18943
rect 121151 18865 121369 18870
rect 117968 18758 118188 18759
rect 121150 18864 121370 18865
rect 117969 18753 118187 18758
rect 111948 18716 112168 18717
rect 111949 18711 112167 18716
rect 121150 18646 121151 18864
rect 121369 18646 121370 18864
rect 124113 18852 124343 18857
rect 121678 18759 121998 18760
rect 121150 18645 121370 18646
rect 121151 18640 121369 18645
rect 105675 18536 105895 18537
rect 102711 18521 102931 18522
rect 102712 18516 102930 18521
rect 99598 18502 99816 18507
rect 81190 18491 81410 18496
rect 99597 18501 99817 18502
rect 84275 18404 84493 18409
rect 84274 18403 84494 18404
rect 71928 18305 72148 18310
rect 78099 18307 78317 18312
rect 78098 18306 78318 18307
rect 2328 18220 2548 18221
rect 78098 18088 78099 18306
rect 78317 18088 78318 18306
rect 78098 18077 78318 18088
rect -6204 17947 -5994 17952
rect -6204 17942 -6199 17947
rect -5999 17942 -5994 17947
rect 78098 17867 78103 18077
rect 78313 17867 78318 18077
rect 78098 17862 78318 17867
rect 84274 18185 84275 18403
rect 84493 18185 84494 18403
rect 87336 18315 87554 18320
rect 84274 17980 84494 18185
rect 87335 18314 87555 18315
rect 87335 18096 87336 18314
rect 87554 18096 87555 18314
rect 99597 18283 99598 18501
rect 99816 18283 99817 18501
rect 121673 18441 121679 18759
rect 121997 18441 122003 18759
rect 124113 18632 124118 18852
rect 124338 18632 124343 18852
rect 127241 18724 127242 18942
rect 127460 18724 127461 18942
rect 133407 18867 133637 18872
rect 130251 18814 130469 18819
rect 127241 18723 127461 18724
rect 130250 18813 130470 18814
rect 127242 18718 127460 18723
rect 124113 18627 124343 18632
rect 130250 18595 130251 18813
rect 130469 18595 130470 18813
rect 133407 18647 133412 18867
rect 133632 18647 133637 18867
rect 154793 18859 155011 18864
rect 154792 18858 155012 18859
rect 145579 18844 145797 18849
rect 148755 18844 148973 18849
rect 145578 18843 145798 18844
rect 142600 18669 142818 18674
rect 133407 18642 133637 18647
rect 142599 18668 142819 18669
rect 139553 18601 139771 18606
rect 130250 18594 130470 18595
rect 139552 18600 139772 18601
rect 130251 18589 130469 18594
rect 121678 18440 121998 18441
rect 139552 18382 139553 18600
rect 139771 18382 139772 18600
rect 142599 18450 142600 18668
rect 142818 18450 142819 18668
rect 145578 18625 145579 18843
rect 145797 18625 145798 18843
rect 145578 18624 145798 18625
rect 148754 18843 148974 18844
rect 148754 18625 148755 18843
rect 148973 18625 148974 18843
rect 151773 18775 151991 18780
rect 148754 18624 148974 18625
rect 151772 18774 151992 18775
rect 145579 18619 145797 18624
rect 148755 18619 148973 18624
rect 151772 18556 151773 18774
rect 151991 18556 151992 18774
rect 154792 18640 154793 18858
rect 155011 18640 155012 18858
rect 157843 18779 157844 18997
rect 158062 18779 158063 18997
rect 174361 18917 174367 19135
rect 174585 18917 174591 19135
rect 305386 19100 305604 19105
rect 305385 19099 305605 19100
rect 290329 18956 290547 18961
rect 290328 18955 290548 18956
rect 229658 18939 229878 18940
rect 174366 18916 174586 18917
rect 176328 18812 176548 18813
rect 157843 18778 158063 18779
rect 157844 18773 158062 18778
rect 167548 18759 167868 18760
rect 160886 18758 161106 18759
rect 154792 18639 155012 18640
rect 154793 18634 155011 18639
rect 151772 18555 151992 18556
rect 151773 18550 151991 18555
rect 160881 18540 160887 18758
rect 161105 18540 161111 18758
rect 160886 18539 161106 18540
rect 163238 18459 163458 18460
rect 142599 18449 142819 18450
rect 142600 18444 142818 18449
rect 139552 18381 139772 18382
rect 139553 18376 139771 18381
rect 99597 18282 99817 18283
rect 99598 18277 99816 18282
rect 136467 18241 136687 18242
rect 163233 18241 163239 18459
rect 163457 18241 163463 18459
rect 167543 18441 167549 18759
rect 167867 18441 167873 18759
rect 176323 18594 176329 18812
rect 176547 18594 176553 18812
rect 180548 18759 180868 18760
rect 189548 18759 189868 18760
rect 198548 18759 198868 18760
rect 204548 18759 204868 18760
rect 211548 18759 211868 18760
rect 223548 18759 223868 18760
rect 176328 18593 176548 18594
rect 173083 18490 173301 18495
rect 173082 18489 173302 18490
rect 167548 18440 167868 18441
rect 173082 18271 173083 18489
rect 173301 18271 173302 18489
rect 180543 18441 180549 18759
rect 180867 18441 180873 18759
rect 189543 18441 189549 18759
rect 189867 18441 189873 18759
rect 198543 18441 198549 18759
rect 198867 18441 198873 18759
rect 204543 18441 204549 18759
rect 204867 18441 204873 18759
rect 206329 18456 206547 18461
rect 206328 18455 206548 18456
rect 180548 18440 180868 18441
rect 189548 18440 189868 18441
rect 198548 18440 198868 18441
rect 204548 18440 204868 18441
rect 173082 18270 173302 18271
rect 173083 18265 173301 18270
rect 87335 18095 87555 18096
rect 87336 18090 87554 18095
rect 136462 18023 136468 18241
rect 136686 18023 136692 18241
rect 163238 18240 163458 18241
rect 206328 18237 206329 18455
rect 206547 18237 206548 18455
rect 211543 18441 211549 18759
rect 211867 18441 211873 18759
rect 215329 18564 215547 18569
rect 215328 18563 215548 18564
rect 211548 18440 211868 18441
rect 215328 18345 215329 18563
rect 215547 18345 215548 18563
rect 223543 18441 223549 18759
rect 223867 18441 223873 18759
rect 229653 18721 229659 18939
rect 229877 18721 229883 18939
rect 232548 18759 232868 18760
rect 238548 18759 238868 18760
rect 250548 18759 250868 18760
rect 263948 18759 264268 18760
rect 269948 18759 270268 18760
rect 272948 18759 273268 18760
rect 275948 18759 276268 18760
rect 281948 18759 282268 18760
rect 285948 18759 286268 18760
rect 229658 18720 229878 18721
rect 232543 18441 232549 18759
rect 232867 18441 232873 18759
rect 233329 18690 233547 18695
rect 233328 18689 233548 18690
rect 233328 18471 233329 18689
rect 233547 18471 233548 18689
rect 233328 18470 233548 18471
rect 233329 18465 233547 18470
rect 238543 18441 238549 18759
rect 238867 18441 238873 18759
rect 242329 18571 242547 18576
rect 242328 18570 242548 18571
rect 241673 18535 241891 18540
rect 241672 18534 241892 18535
rect 223548 18440 223868 18441
rect 232548 18440 232868 18441
rect 238548 18440 238868 18441
rect 227194 18428 227414 18429
rect 215328 18344 215548 18345
rect 215329 18339 215547 18344
rect 206328 18236 206548 18237
rect 206329 18231 206547 18236
rect 227189 18210 227195 18428
rect 227413 18210 227419 18428
rect 241672 18316 241673 18534
rect 241891 18316 241892 18534
rect 242328 18352 242329 18570
rect 242547 18352 242548 18570
rect 250543 18441 250549 18759
rect 250867 18441 250873 18759
rect 254329 18701 254547 18706
rect 254328 18700 254548 18701
rect 253925 18509 254145 18510
rect 250548 18440 250868 18441
rect 242328 18351 242548 18352
rect 242329 18346 242547 18351
rect 241672 18315 241892 18316
rect 241673 18310 241891 18315
rect 234650 18303 234870 18304
rect 227194 18209 227414 18210
rect 165929 18175 166147 18180
rect 165928 18174 166148 18175
rect 136467 18022 136687 18023
rect 84274 17770 84279 17980
rect 84489 17770 84494 17980
rect 165928 17956 165929 18174
rect 166147 17956 166148 18174
rect 213156 18099 213374 18104
rect 213155 18098 213375 18099
rect 185329 18037 185547 18042
rect 165928 17955 166148 17956
rect 185328 18036 185548 18037
rect 165929 17950 166147 17955
rect 182473 17859 182693 17860
rect 84274 17765 84494 17770
rect -6204 17736 -5994 17742
rect 182468 17641 182474 17859
rect 182692 17641 182698 17859
rect 185328 17818 185329 18036
rect 185547 17818 185548 18036
rect 200916 17957 201134 17962
rect 200915 17956 201135 17957
rect 196793 17929 197013 17930
rect 185328 17817 185548 17818
rect 185329 17812 185547 17817
rect 196788 17711 196794 17929
rect 197012 17711 197018 17929
rect 200915 17738 200916 17956
rect 201134 17738 201135 17956
rect 213155 17880 213156 18098
rect 213374 17880 213375 18098
rect 234645 18085 234651 18303
rect 234869 18085 234875 18303
rect 253920 18291 253926 18509
rect 254144 18291 254150 18509
rect 254328 18482 254329 18700
rect 254547 18482 254548 18700
rect 254328 18481 254548 18482
rect 254329 18476 254547 18481
rect 263943 18441 263949 18759
rect 264267 18441 264273 18759
rect 269032 18560 269252 18561
rect 263948 18440 264268 18441
rect 269027 18342 269033 18560
rect 269251 18342 269257 18560
rect 269943 18441 269949 18759
rect 270267 18441 270273 18759
rect 272943 18441 272949 18759
rect 273267 18441 273273 18759
rect 275943 18441 275949 18759
rect 276267 18441 276273 18759
rect 279676 18698 279896 18699
rect 279671 18480 279677 18698
rect 279895 18480 279901 18698
rect 279676 18479 279896 18480
rect 281943 18441 281949 18759
rect 282267 18441 282273 18759
rect 285943 18441 285949 18759
rect 286267 18441 286273 18759
rect 290328 18737 290329 18955
rect 290547 18737 290548 18955
rect 305385 18881 305386 19099
rect 305604 18881 305605 19099
rect 305385 18880 305605 18881
rect 305386 18875 305604 18880
rect 293948 18759 294268 18760
rect 296948 18759 297268 18760
rect 299948 18759 300268 18760
rect 302948 18759 303268 18760
rect 290328 18736 290548 18737
rect 290329 18731 290547 18736
rect 293943 18441 293949 18759
rect 294267 18441 294273 18759
rect 296943 18441 296949 18759
rect 297267 18441 297273 18759
rect 299943 18441 299949 18759
rect 300267 18441 300273 18759
rect 302943 18441 302949 18759
rect 303267 18441 303273 18759
rect 269948 18440 270268 18441
rect 272948 18440 273268 18441
rect 275948 18440 276268 18441
rect 281948 18440 282268 18441
rect 285948 18440 286268 18441
rect 293948 18440 294268 18441
rect 296948 18440 297268 18441
rect 299948 18440 300268 18441
rect 302948 18440 303268 18441
rect 269032 18341 269252 18342
rect 253925 18290 254145 18291
rect 269329 18269 269547 18274
rect 269328 18268 269548 18269
rect 261045 18126 261263 18131
rect 261044 18125 261264 18126
rect 234650 18084 234870 18085
rect 240917 18016 241135 18021
rect 213155 17879 213375 17880
rect 240916 18015 241136 18016
rect 213156 17874 213374 17879
rect 240916 17797 240917 18015
rect 241135 17797 241136 18015
rect 261044 17907 261045 18125
rect 261263 17907 261264 18125
rect 269328 18050 269329 18268
rect 269547 18050 269548 18268
rect 292407 18227 292627 18228
rect 278878 18206 279098 18207
rect 269328 18049 269548 18050
rect 269329 18044 269547 18049
rect 278873 17988 278879 18206
rect 279097 17988 279103 18206
rect 284329 18138 284547 18143
rect 284328 18137 284548 18138
rect 278878 17987 279098 17988
rect 265871 17964 266089 17969
rect 261044 17906 261264 17907
rect 265870 17963 266090 17964
rect 261045 17901 261263 17906
rect 249667 17860 249887 17861
rect 240916 17796 241136 17797
rect 240917 17791 241135 17796
rect 207000 17752 207218 17757
rect 200915 17737 201135 17738
rect 206999 17751 207219 17752
rect 200916 17732 201134 17737
rect 196793 17710 197013 17711
rect 188329 17660 188547 17665
rect 188328 17659 188548 17660
rect 182473 17640 182693 17641
rect 188328 17441 188329 17659
rect 188547 17441 188548 17659
rect 206999 17533 207000 17751
rect 207218 17533 207219 17751
rect 221329 17712 221547 17717
rect 206999 17532 207219 17533
rect 221328 17711 221548 17712
rect 207000 17527 207218 17532
rect 221328 17493 221329 17711
rect 221547 17493 221548 17711
rect 249662 17642 249668 17860
rect 249886 17642 249892 17860
rect 265870 17745 265871 17963
rect 266089 17745 266090 17963
rect 284328 17919 284329 18137
rect 284547 17919 284548 18137
rect 292402 18009 292408 18227
rect 292626 18009 292632 18227
rect 292407 18008 292627 18009
rect 284328 17918 284548 17919
rect 284329 17913 284547 17918
rect 265870 17744 266090 17745
rect 265871 17739 266089 17744
rect 299259 17724 299477 17729
rect 299258 17723 299478 17724
rect 249667 17641 249887 17642
rect 277693 17582 277913 17583
rect 221328 17492 221548 17493
rect 221329 17487 221547 17492
rect 188328 17440 188548 17441
rect 188329 17435 188547 17440
rect 168864 17422 169082 17427
rect 168863 17421 169083 17422
rect 168863 17203 168864 17421
rect 169082 17203 169083 17421
rect 277688 17364 277694 17582
rect 277912 17364 277918 17582
rect 286930 17513 287148 17518
rect 286929 17512 287149 17513
rect 277693 17363 277913 17364
rect 286929 17294 286930 17512
rect 287148 17294 287149 17512
rect 299258 17505 299259 17723
rect 299477 17505 299478 17723
rect 299258 17504 299478 17505
rect 299259 17499 299477 17504
rect 286929 17293 287149 17294
rect 286930 17288 287148 17293
rect 213905 17270 214123 17275
rect 168863 17202 169083 17203
rect 213904 17269 214124 17270
rect 168864 17197 169082 17202
rect 184011 17153 184229 17158
rect 184010 17152 184230 17153
rect 184010 16934 184011 17152
rect 184229 16934 184230 17152
rect 213904 17051 213905 17269
rect 214123 17051 214124 17269
rect 260054 17247 260272 17252
rect 260053 17246 260273 17247
rect 220689 17229 220907 17234
rect 213904 17050 214124 17051
rect 220688 17228 220908 17229
rect 213905 17045 214123 17050
rect 193466 17020 193684 17025
rect 184010 16933 184230 16934
rect 193465 17019 193685 17020
rect 184011 16928 184229 16933
rect 193465 16801 193466 17019
rect 193684 16801 193685 17019
rect 220688 17010 220689 17228
rect 220907 17010 220908 17228
rect 248712 17078 248930 17083
rect 220688 17009 220908 17010
rect 248711 17077 248931 17078
rect 220689 17004 220907 17009
rect 202004 16895 202222 16900
rect 193465 16800 193685 16801
rect 202003 16894 202223 16895
rect 193466 16795 193684 16800
rect 202003 16676 202004 16894
rect 202222 16676 202223 16894
rect 248711 16859 248712 17077
rect 248930 16859 248931 17077
rect 260053 17028 260054 17246
rect 260272 17028 260273 17246
rect 300252 17106 300470 17111
rect 260053 17027 260273 17028
rect 300251 17105 300471 17106
rect 260054 17022 260272 17027
rect 300251 16887 300252 17105
rect 300470 16887 300471 17105
rect 300251 16886 300471 16887
rect 300252 16881 300470 16886
rect 248711 16858 248931 16859
rect 248712 16853 248930 16858
rect 202003 16675 202223 16676
rect 202004 16670 202222 16675
rect 302942 16416 303274 16421
rect 302942 16411 302947 16416
rect 303269 16411 303274 16416
rect 302942 16083 303274 16089
rect 18083 15712 18413 15717
rect 18083 15707 18088 15712
rect 18408 15707 18413 15712
rect 3659 15694 3989 15699
rect 3659 15689 3664 15694
rect 3984 15689 3989 15694
rect 103 15588 313 15593
rect 103 15583 108 15588
rect 308 15583 313 15588
rect 103 15377 313 15383
rect 121673 15710 122003 15715
rect 121673 15705 121678 15710
rect 121998 15705 122003 15710
rect 64251 15696 64581 15701
rect 18083 15381 18413 15387
rect 32909 15688 33239 15693
rect 32909 15683 32914 15688
rect 33234 15683 33239 15688
rect 3659 15363 3989 15369
rect 64251 15691 64256 15696
rect 64576 15691 64581 15696
rect 121673 15379 122003 15385
rect 167543 15712 167873 15717
rect 167543 15707 167548 15712
rect 167868 15707 167873 15712
rect 167543 15381 167873 15387
rect 180543 15712 180873 15717
rect 180543 15707 180548 15712
rect 180868 15707 180873 15712
rect 180543 15381 180873 15387
rect 189543 15712 189873 15717
rect 189543 15707 189548 15712
rect 189868 15707 189873 15712
rect 189543 15381 189873 15387
rect 198543 15712 198873 15717
rect 198543 15707 198548 15712
rect 198868 15707 198873 15712
rect 198543 15381 198873 15387
rect 204543 15712 204873 15717
rect 204543 15707 204548 15712
rect 204868 15707 204873 15712
rect 204543 15381 204873 15387
rect 211543 15712 211873 15717
rect 211543 15707 211548 15712
rect 211868 15707 211873 15712
rect 211543 15381 211873 15387
rect 223543 15712 223873 15717
rect 223543 15707 223548 15712
rect 223868 15707 223873 15712
rect 223543 15381 223873 15387
rect 232543 15712 232873 15717
rect 232543 15707 232548 15712
rect 232868 15707 232873 15712
rect 232543 15381 232873 15387
rect 238543 15712 238873 15717
rect 238543 15707 238548 15712
rect 238868 15707 238873 15712
rect 238543 15381 238873 15387
rect 250543 15712 250873 15717
rect 250543 15707 250548 15712
rect 250868 15707 250873 15712
rect 250543 15381 250873 15387
rect 263943 15712 264273 15717
rect 263943 15707 263948 15712
rect 264268 15707 264273 15712
rect 263943 15381 264273 15387
rect 269943 15712 270273 15717
rect 269943 15707 269948 15712
rect 270268 15707 270273 15712
rect 269943 15381 270273 15387
rect 272943 15712 273273 15717
rect 272943 15707 272948 15712
rect 273268 15707 273273 15712
rect 272943 15381 273273 15387
rect 275943 15712 276273 15717
rect 275943 15707 275948 15712
rect 276268 15707 276273 15712
rect 275943 15381 276273 15387
rect 281943 15712 282273 15717
rect 281943 15707 281948 15712
rect 282268 15707 282273 15712
rect 281943 15381 282273 15387
rect 285943 15712 286273 15717
rect 285943 15707 285948 15712
rect 286268 15707 286273 15712
rect 285943 15381 286273 15387
rect 293943 15712 294273 15717
rect 293943 15707 293948 15712
rect 294268 15707 294273 15712
rect 293943 15381 294273 15387
rect 296943 15712 297273 15717
rect 296943 15707 296948 15712
rect 297268 15707 297273 15712
rect 296943 15381 297273 15387
rect 299943 15712 300273 15717
rect 299943 15707 299948 15712
rect 300268 15707 300273 15712
rect 299943 15381 300273 15387
rect 302943 15712 303273 15717
rect 302943 15707 302948 15712
rect 303268 15707 303273 15712
rect 302943 15381 303273 15387
rect 64251 15365 64581 15371
rect 32909 15357 33239 15363
<< via3 >>
rect 302503 324533 302713 324538
rect 302503 324338 302508 324533
rect 302508 324338 302708 324533
rect 302708 324338 302713 324533
rect 303927 321353 304245 321357
rect 303927 321043 303931 321353
rect 303931 321043 304241 321353
rect 304241 321043 304245 321353
rect 303927 321039 304245 321043
rect -2006 319722 -1806 319922
rect 303927 318353 304245 318357
rect 303927 318043 303931 318353
rect 303931 318043 304241 318353
rect 304241 318043 304245 318353
rect 303927 318039 304245 318043
rect -2006 316722 -1806 316922
rect 303927 315353 304245 315357
rect 303927 315043 303931 315353
rect 303931 315043 304241 315353
rect 304241 315043 304245 315353
rect 303927 315039 304245 315043
rect -2006 313722 -1806 313922
rect 303927 312353 304245 312357
rect 303927 312043 303931 312353
rect 303931 312043 304241 312353
rect 304241 312043 304245 312353
rect 303927 312039 304245 312043
rect -2006 310722 -1806 310922
rect 303927 309353 304245 309357
rect 303927 309043 303931 309353
rect 303931 309043 304241 309353
rect 304241 309043 304245 309353
rect 303927 309039 304245 309043
rect -2006 307722 -1806 307922
rect 303927 306353 304245 306357
rect 303927 306043 303931 306353
rect 303931 306043 304241 306353
rect 304241 306043 304245 306353
rect 303927 306039 304245 306043
rect -2006 304722 -1806 304922
rect 303927 303353 304245 303357
rect 303927 303043 303931 303353
rect 303931 303043 304241 303353
rect 304241 303043 304245 303353
rect 303927 303039 304245 303043
rect -2006 301722 -1806 301922
rect 303927 300353 304245 300357
rect 303927 300043 303931 300353
rect 303931 300043 304241 300353
rect 304241 300043 304245 300353
rect 303927 300039 304245 300043
rect -2006 298722 -1806 298922
rect 303927 297353 304245 297357
rect 303927 297043 303931 297353
rect 303931 297043 304241 297353
rect 304241 297043 304245 297353
rect 303927 297039 304245 297043
rect -2006 295722 -1806 295922
rect 303927 294353 304245 294357
rect 303927 294043 303931 294353
rect 303931 294043 304241 294353
rect 304241 294043 304245 294353
rect 303927 294039 304245 294043
rect -2006 292722 -1806 292922
rect 303927 291353 304245 291357
rect 303927 291043 303931 291353
rect 303931 291043 304241 291353
rect 304241 291043 304245 291353
rect 303927 291039 304245 291043
rect -2006 289722 -1806 289922
rect 303927 288353 304245 288357
rect 303927 288043 303931 288353
rect 303931 288043 304241 288353
rect 304241 288043 304245 288353
rect 303927 288039 304245 288043
rect -2006 286722 -1806 286922
rect 303927 285353 304245 285357
rect 303927 285043 303931 285353
rect 303931 285043 304241 285353
rect 304241 285043 304245 285353
rect 303927 285039 304245 285043
rect -2006 283722 -1806 283922
rect 303927 282353 304245 282357
rect 303927 282043 303931 282353
rect 303931 282043 304241 282353
rect 304241 282043 304245 282353
rect 303927 282039 304245 282043
rect -2006 280722 -1806 280922
rect 303927 279353 304245 279357
rect 303927 279043 303931 279353
rect 303931 279043 304241 279353
rect 304241 279043 304245 279353
rect 303927 279039 304245 279043
rect -2006 277722 -1806 277922
rect 303927 276353 304245 276357
rect 303927 276043 303931 276353
rect 303931 276043 304241 276353
rect 304241 276043 304245 276353
rect 303927 276039 304245 276043
rect -2006 274722 -1806 274922
rect 303927 273353 304245 273357
rect 303927 273043 303931 273353
rect 303931 273043 304241 273353
rect 304241 273043 304245 273353
rect 303927 273039 304245 273043
rect -2006 271722 -1806 271922
rect 303927 270353 304245 270357
rect 303927 270043 303931 270353
rect 303931 270043 304241 270353
rect 304241 270043 304245 270353
rect 303927 270039 304245 270043
rect -2006 268722 -1806 268922
rect 303927 267353 304245 267357
rect 303927 267043 303931 267353
rect 303931 267043 304241 267353
rect 304241 267043 304245 267353
rect 303927 267039 304245 267043
rect -2006 265722 -1806 265922
rect 303927 264353 304245 264357
rect 303927 264043 303931 264353
rect 303931 264043 304241 264353
rect 304241 264043 304245 264353
rect 303927 264039 304245 264043
rect -2006 262722 -1806 262922
rect 303927 261353 304245 261357
rect 303927 261043 303931 261353
rect 303931 261043 304241 261353
rect 304241 261043 304245 261353
rect 303927 261039 304245 261043
rect -2006 259722 -1806 259922
rect 303927 258353 304245 258357
rect 303927 258043 303931 258353
rect 303931 258043 304241 258353
rect 304241 258043 304245 258353
rect 303927 258039 304245 258043
rect -2006 256722 -1806 256922
rect 303927 255353 304245 255357
rect 303927 255043 303931 255353
rect 303931 255043 304241 255353
rect 304241 255043 304245 255353
rect 303927 255039 304245 255043
rect -2006 253722 -1806 253922
rect 303927 252353 304245 252357
rect 303927 252043 303931 252353
rect 303931 252043 304241 252353
rect 304241 252043 304245 252353
rect 303927 252039 304245 252043
rect -2006 250722 -1806 250922
rect 303927 249353 304245 249357
rect 303927 249043 303931 249353
rect 303931 249043 304241 249353
rect 304241 249043 304245 249353
rect 303927 249039 304245 249043
rect -2006 247722 -1806 247922
rect 303927 246353 304245 246357
rect 303927 246043 303931 246353
rect 303931 246043 304241 246353
rect 304241 246043 304245 246353
rect 303927 246039 304245 246043
rect -2006 244722 -1806 244922
rect 303927 243353 304245 243357
rect 303927 243043 303931 243353
rect 303931 243043 304241 243353
rect 304241 243043 304245 243353
rect 303927 243039 304245 243043
rect -2006 241722 -1806 241922
rect 303927 240353 304245 240357
rect 303927 240043 303931 240353
rect 303931 240043 304241 240353
rect 304241 240043 304245 240353
rect 303927 240039 304245 240043
rect -2006 238722 -1806 238922
rect 303927 237353 304245 237357
rect 303927 237043 303931 237353
rect 303931 237043 304241 237353
rect 304241 237043 304245 237353
rect 303927 237039 304245 237043
rect -2006 235722 -1806 235922
rect 303927 234353 304245 234357
rect 303927 234043 303931 234353
rect 303931 234043 304241 234353
rect 304241 234043 304245 234353
rect 303927 234039 304245 234043
rect -2006 232722 -1806 232922
rect 303927 231353 304245 231357
rect 303927 231043 303931 231353
rect 303931 231043 304241 231353
rect 304241 231043 304245 231353
rect 303927 231039 304245 231043
rect -2006 229722 -1806 229922
rect 303927 228353 304245 228357
rect 303927 228043 303931 228353
rect 303931 228043 304241 228353
rect 304241 228043 304245 228353
rect 303927 228039 304245 228043
rect -2006 226722 -1806 226922
rect 303927 225353 304245 225357
rect 303927 225043 303931 225353
rect 303931 225043 304241 225353
rect 304241 225043 304245 225353
rect 303927 225039 304245 225043
rect -2006 223722 -1806 223922
rect 303927 222353 304245 222357
rect 303927 222043 303931 222353
rect 303931 222043 304241 222353
rect 304241 222043 304245 222353
rect 303927 222039 304245 222043
rect -2006 220722 -1806 220922
rect 303927 219353 304245 219357
rect 303927 219043 303931 219353
rect 303931 219043 304241 219353
rect 304241 219043 304245 219353
rect 303927 219039 304245 219043
rect -2006 217722 -1806 217922
rect 303927 216353 304245 216357
rect 303927 216043 303931 216353
rect 303931 216043 304241 216353
rect 304241 216043 304245 216353
rect 303927 216039 304245 216043
rect -2006 214722 -1806 214922
rect 303927 213353 304245 213357
rect 303927 213043 303931 213353
rect 303931 213043 304241 213353
rect 304241 213043 304245 213353
rect 303927 213039 304245 213043
rect -2006 211722 -1806 211922
rect 303927 210353 304245 210357
rect 303927 210043 303931 210353
rect 303931 210043 304241 210353
rect 304241 210043 304245 210353
rect 303927 210039 304245 210043
rect -2006 208722 -1806 208922
rect 303927 207353 304245 207357
rect 303927 207043 303931 207353
rect 303931 207043 304241 207353
rect 304241 207043 304245 207353
rect 303927 207039 304245 207043
rect -2006 205722 -1806 205922
rect 303927 204353 304245 204357
rect 303927 204043 303931 204353
rect 303931 204043 304241 204353
rect 304241 204043 304245 204353
rect 303927 204039 304245 204043
rect -2006 202722 -1806 202922
rect 303927 201353 304245 201357
rect 303927 201043 303931 201353
rect 303931 201043 304241 201353
rect 304241 201043 304245 201353
rect 303927 201039 304245 201043
rect -2006 199722 -1806 199922
rect 303927 198353 304245 198357
rect 303927 198043 303931 198353
rect 303931 198043 304241 198353
rect 304241 198043 304245 198353
rect 303927 198039 304245 198043
rect -2006 196722 -1806 196922
rect 303927 195353 304245 195357
rect 303927 195043 303931 195353
rect 303931 195043 304241 195353
rect 304241 195043 304245 195353
rect 303927 195039 304245 195043
rect -2006 193722 -1806 193922
rect 303927 192353 304245 192357
rect 303927 192043 303931 192353
rect 303931 192043 304241 192353
rect 304241 192043 304245 192353
rect 303927 192039 304245 192043
rect -2006 190722 -1806 190922
rect 303927 189353 304245 189357
rect 303927 189043 303931 189353
rect 303931 189043 304241 189353
rect 304241 189043 304245 189353
rect 303927 189039 304245 189043
rect -2006 187722 -1806 187922
rect 303927 186353 304245 186357
rect 303927 186043 303931 186353
rect 303931 186043 304241 186353
rect 304241 186043 304245 186353
rect 303927 186039 304245 186043
rect -2006 184722 -1806 184922
rect 303927 183353 304245 183357
rect 303927 183043 303931 183353
rect 303931 183043 304241 183353
rect 304241 183043 304245 183353
rect 303927 183039 304245 183043
rect -2006 181722 -1806 181922
rect 303927 180353 304245 180357
rect 303927 180043 303931 180353
rect 303931 180043 304241 180353
rect 304241 180043 304245 180353
rect 303927 180039 304245 180043
rect -2006 178722 -1806 178922
rect 303927 177353 304245 177357
rect 303927 177043 303931 177353
rect 303931 177043 304241 177353
rect 304241 177043 304245 177353
rect 303927 177039 304245 177043
rect -2006 175722 -1806 175922
rect 303927 174353 304245 174357
rect 303927 174043 303931 174353
rect 303931 174043 304241 174353
rect 304241 174043 304245 174353
rect 303927 174039 304245 174043
rect -2006 172722 -1806 172922
rect 303927 171353 304245 171357
rect 303927 171043 303931 171353
rect 303931 171043 304241 171353
rect 304241 171043 304245 171353
rect 303927 171039 304245 171043
rect -2006 169722 -1806 169922
rect 303927 168353 304245 168357
rect 303927 168043 303931 168353
rect 303931 168043 304241 168353
rect 304241 168043 304245 168353
rect 303927 168039 304245 168043
rect -2006 166722 -1806 166922
rect 303927 165353 304245 165357
rect 303927 165043 303931 165353
rect 303931 165043 304241 165353
rect 304241 165043 304245 165353
rect 303927 165039 304245 165043
rect -2006 163722 -1806 163922
rect 303927 162353 304245 162357
rect 303927 162043 303931 162353
rect 303931 162043 304241 162353
rect 304241 162043 304245 162353
rect 303927 162039 304245 162043
rect -2006 160722 -1806 160922
rect 303927 159353 304245 159357
rect 303927 159043 303931 159353
rect 303931 159043 304241 159353
rect 304241 159043 304245 159353
rect 303927 159039 304245 159043
rect -2006 157722 -1806 157922
rect 303927 156353 304245 156357
rect 303927 156043 303931 156353
rect 303931 156043 304241 156353
rect 304241 156043 304245 156353
rect 303927 156039 304245 156043
rect -2006 154722 -1806 154922
rect 303927 153353 304245 153357
rect 303927 153043 303931 153353
rect 303931 153043 304241 153353
rect 304241 153043 304245 153353
rect 303927 153039 304245 153043
rect -2006 151722 -1806 151922
rect 303927 150353 304245 150357
rect 303927 150043 303931 150353
rect 303931 150043 304241 150353
rect 304241 150043 304245 150353
rect 303927 150039 304245 150043
rect -2006 148722 -1806 148922
rect 303927 147353 304245 147357
rect 303927 147043 303931 147353
rect 303931 147043 304241 147353
rect 304241 147043 304245 147353
rect 303927 147039 304245 147043
rect -2006 145722 -1806 145922
rect 303927 144353 304245 144357
rect 303927 144043 303931 144353
rect 303931 144043 304241 144353
rect 304241 144043 304245 144353
rect 303927 144039 304245 144043
rect -2006 142722 -1806 142922
rect 303927 141353 304245 141357
rect 303927 141043 303931 141353
rect 303931 141043 304241 141353
rect 304241 141043 304245 141353
rect 303927 141039 304245 141043
rect -2006 139722 -1806 139922
rect 303927 138353 304245 138357
rect 303927 138043 303931 138353
rect 303931 138043 304241 138353
rect 304241 138043 304245 138353
rect 303927 138039 304245 138043
rect -2006 136722 -1806 136922
rect 303927 135353 304245 135357
rect 303927 135043 303931 135353
rect 303931 135043 304241 135353
rect 304241 135043 304245 135353
rect 303927 135039 304245 135043
rect -2006 133722 -1806 133922
rect 303927 132353 304245 132357
rect 303927 132043 303931 132353
rect 303931 132043 304241 132353
rect 304241 132043 304245 132353
rect 303927 132039 304245 132043
rect -2006 130722 -1806 130922
rect 303927 129353 304245 129357
rect 303927 129043 303931 129353
rect 303931 129043 304241 129353
rect 304241 129043 304245 129353
rect 303927 129039 304245 129043
rect -2006 127722 -1806 127922
rect 303927 126353 304245 126357
rect 303927 126043 303931 126353
rect 303931 126043 304241 126353
rect 304241 126043 304245 126353
rect 303927 126039 304245 126043
rect -2006 124722 -1806 124922
rect 303927 123353 304245 123357
rect 303927 123043 303931 123353
rect 303931 123043 304241 123353
rect 304241 123043 304245 123353
rect 303927 123039 304245 123043
rect -2006 121722 -1806 121922
rect 303927 120353 304245 120357
rect 303927 120043 303931 120353
rect 303931 120043 304241 120353
rect 304241 120043 304245 120353
rect 303927 120039 304245 120043
rect -2006 118722 -1806 118922
rect 303927 117353 304245 117357
rect 303927 117043 303931 117353
rect 303931 117043 304241 117353
rect 304241 117043 304245 117353
rect 303927 117039 304245 117043
rect -2006 115722 -1806 115922
rect 303927 114353 304245 114357
rect 303927 114043 303931 114353
rect 303931 114043 304241 114353
rect 304241 114043 304245 114353
rect 303927 114039 304245 114043
rect -2006 112722 -1806 112922
rect 303927 111353 304245 111357
rect 303927 111043 303931 111353
rect 303931 111043 304241 111353
rect 304241 111043 304245 111353
rect 303927 111039 304245 111043
rect -2006 109722 -1806 109922
rect 303927 108353 304245 108357
rect 303927 108043 303931 108353
rect 303931 108043 304241 108353
rect 304241 108043 304245 108353
rect 303927 108039 304245 108043
rect -2006 106722 -1806 106922
rect 303927 105353 304245 105357
rect 303927 105043 303931 105353
rect 303931 105043 304241 105353
rect 304241 105043 304245 105353
rect 303927 105039 304245 105043
rect -2006 103722 -1806 103922
rect 303927 102353 304245 102357
rect 303927 102043 303931 102353
rect 303931 102043 304241 102353
rect 304241 102043 304245 102353
rect 303927 102039 304245 102043
rect -2006 100722 -1806 100922
rect 303927 99353 304245 99357
rect 303927 99043 303931 99353
rect 303931 99043 304241 99353
rect 304241 99043 304245 99353
rect 303927 99039 304245 99043
rect -2006 97722 -1806 97922
rect 303927 96353 304245 96357
rect 303927 96043 303931 96353
rect 303931 96043 304241 96353
rect 304241 96043 304245 96353
rect 303927 96039 304245 96043
rect -2006 94722 -1806 94922
rect 303927 93353 304245 93357
rect 303927 93043 303931 93353
rect 303931 93043 304241 93353
rect 304241 93043 304245 93353
rect 303927 93039 304245 93043
rect -2006 91722 -1806 91922
rect 303927 90353 304245 90357
rect 303927 90043 303931 90353
rect 303931 90043 304241 90353
rect 304241 90043 304245 90353
rect 303927 90039 304245 90043
rect -2006 88722 -1806 88922
rect 303927 87353 304245 87357
rect 303927 87043 303931 87353
rect 303931 87043 304241 87353
rect 304241 87043 304245 87353
rect 303927 87039 304245 87043
rect -2006 85722 -1806 85922
rect 303927 84353 304245 84357
rect 303927 84043 303931 84353
rect 303931 84043 304241 84353
rect 304241 84043 304245 84353
rect 303927 84039 304245 84043
rect -2006 82722 -1806 82922
rect 303927 81353 304245 81357
rect 303927 81043 303931 81353
rect 303931 81043 304241 81353
rect 304241 81043 304245 81353
rect 303927 81039 304245 81043
rect -2006 79722 -1806 79922
rect 303927 78353 304245 78357
rect 303927 78043 303931 78353
rect 303931 78043 304241 78353
rect 304241 78043 304245 78353
rect 303927 78039 304245 78043
rect -2006 76722 -1806 76922
rect 303927 75353 304245 75357
rect 303927 75043 303931 75353
rect 303931 75043 304241 75353
rect 304241 75043 304245 75353
rect 303927 75039 304245 75043
rect -2006 73722 -1806 73922
rect 303927 72353 304245 72357
rect 303927 72043 303931 72353
rect 303931 72043 304241 72353
rect 304241 72043 304245 72353
rect 303927 72039 304245 72043
rect -2006 70722 -1806 70922
rect 303927 69353 304245 69357
rect 303927 69043 303931 69353
rect 303931 69043 304241 69353
rect 304241 69043 304245 69353
rect 303927 69039 304245 69043
rect -2006 67722 -1806 67922
rect 303927 66353 304245 66357
rect 303927 66043 303931 66353
rect 303931 66043 304241 66353
rect 304241 66043 304245 66353
rect 303927 66039 304245 66043
rect -2006 64722 -1806 64922
rect 303927 63353 304245 63357
rect 303927 63043 303931 63353
rect 303931 63043 304241 63353
rect 304241 63043 304245 63353
rect 303927 63039 304245 63043
rect -2006 61722 -1806 61922
rect 303927 60353 304245 60357
rect 303927 60043 303931 60353
rect 303931 60043 304241 60353
rect 304241 60043 304245 60353
rect 303927 60039 304245 60043
rect -2006 58722 -1806 58922
rect 303927 57353 304245 57357
rect 303927 57043 303931 57353
rect 303931 57043 304241 57353
rect 304241 57043 304245 57353
rect 303927 57039 304245 57043
rect -2006 55722 -1806 55922
rect 303927 54353 304245 54357
rect 303927 54043 303931 54353
rect 303931 54043 304241 54353
rect 304241 54043 304245 54353
rect 303927 54039 304245 54043
rect -2006 52722 -1806 52922
rect 303927 51353 304245 51357
rect 303927 51043 303931 51353
rect 303931 51043 304241 51353
rect 304241 51043 304245 51353
rect 303927 51039 304245 51043
rect -2006 49722 -1806 49922
rect 303927 48353 304245 48357
rect 303927 48043 303931 48353
rect 303931 48043 304241 48353
rect 304241 48043 304245 48353
rect 303927 48039 304245 48043
rect -2006 46722 -1806 46922
rect 303927 45353 304245 45357
rect 303927 45043 303931 45353
rect 303931 45043 304241 45353
rect 304241 45043 304245 45353
rect 303927 45039 304245 45043
rect -2006 43722 -1806 43922
rect 303927 42353 304245 42357
rect 303927 42043 303931 42353
rect 303931 42043 304241 42353
rect 304241 42043 304245 42353
rect 303927 42039 304245 42043
rect -2006 40722 -1806 40922
rect 303927 39353 304245 39357
rect 303927 39043 303931 39353
rect 303931 39043 304241 39353
rect 304241 39043 304245 39353
rect 303927 39039 304245 39043
rect -2006 37722 -1806 37922
rect 303927 36353 304245 36357
rect 303927 36043 303931 36353
rect 303931 36043 304241 36353
rect 304241 36043 304245 36353
rect 303927 36039 304245 36043
rect -2006 34722 -1806 34922
rect 303927 33353 304245 33357
rect 303927 33043 303931 33353
rect 303931 33043 304241 33353
rect 304241 33043 304245 33353
rect 303927 33039 304245 33043
rect -2006 31722 -1806 31922
rect 303927 30353 304245 30357
rect 303927 30043 303931 30353
rect 303931 30043 304241 30353
rect 304241 30043 304245 30353
rect 303927 30039 304245 30043
rect -2006 28722 -1806 28922
rect 303927 27353 304245 27357
rect 303927 27043 303931 27353
rect 303931 27043 304241 27353
rect 304241 27043 304245 27353
rect 303927 27039 304245 27043
rect -2006 25722 -1806 25922
rect 303927 24353 304245 24357
rect 303927 24043 303931 24353
rect 303931 24043 304241 24353
rect 304241 24043 304245 24353
rect 303927 24039 304245 24043
rect -2006 22722 -1806 22922
rect 303927 21353 304245 21357
rect 303927 21043 303931 21353
rect 303931 21043 304241 21353
rect 304241 21043 304245 21353
rect 303927 21039 304245 21043
rect 19870 19189 20088 19193
rect 19870 18979 19874 19189
rect 19874 18979 20084 19189
rect 20084 18979 20088 19189
rect 19870 18975 20088 18979
rect 3665 18755 3983 18759
rect 3665 18445 3669 18755
rect 3669 18445 3979 18755
rect 3979 18445 3983 18755
rect 3665 18441 3983 18445
rect 5329 18780 5547 18784
rect 5329 18570 5333 18780
rect 5333 18570 5543 18780
rect 5543 18570 5547 18780
rect 5329 18566 5547 18570
rect 7483 18887 7701 18891
rect 7483 18677 7487 18887
rect 7487 18677 7697 18887
rect 7697 18677 7701 18887
rect 7483 18673 7701 18677
rect 10712 18831 10930 18835
rect 10712 18621 10716 18831
rect 10716 18621 10926 18831
rect 10926 18621 10930 18831
rect 10712 18617 10930 18621
rect 13802 18925 14020 18929
rect 13802 18715 13806 18925
rect 13806 18715 14016 18925
rect 14016 18715 14020 18925
rect 13802 18711 14020 18715
rect 16912 18812 17130 18816
rect 16912 18602 16916 18812
rect 16916 18602 17126 18812
rect 17126 18602 17130 18812
rect 16912 18598 17130 18602
rect 25944 19007 26162 19011
rect 25944 18797 25948 19007
rect 25948 18797 26158 19007
rect 26158 18797 26162 19007
rect 25944 18793 26162 18797
rect 29085 18843 29303 19061
rect 32329 18982 32547 18986
rect 32329 18772 32333 18982
rect 32333 18772 32543 18982
rect 32543 18772 32547 18982
rect 32329 18768 32547 18772
rect 35329 19051 35547 19055
rect 35329 18841 35333 19051
rect 35333 18841 35543 19051
rect 35543 18841 35547 19051
rect 35329 18837 35547 18841
rect 38329 19214 38547 19218
rect 38329 19004 38333 19214
rect 38333 19004 38543 19214
rect 38543 19004 38547 19214
rect 38329 19000 38547 19004
rect 18089 18755 18407 18759
rect 18089 18445 18093 18755
rect 18093 18445 18403 18755
rect 18403 18445 18407 18755
rect 18089 18441 18407 18445
rect 22898 18654 23116 18658
rect 22898 18444 22902 18654
rect 22902 18444 23112 18654
rect 23112 18444 23116 18654
rect 22898 18440 23116 18444
rect 32915 18755 33233 18759
rect 32915 18445 32919 18755
rect 32919 18445 33229 18755
rect 33229 18445 33233 18755
rect 32915 18441 33233 18445
rect 41329 18868 41547 18872
rect 41329 18658 41333 18868
rect 41333 18658 41543 18868
rect 41543 18658 41547 18868
rect 41329 18654 41547 18658
rect 44329 18919 44547 18923
rect 44329 18709 44333 18919
rect 44333 18709 44543 18919
rect 44543 18709 44547 18919
rect 44329 18705 44547 18709
rect 47329 19126 47547 19130
rect 47329 18916 47333 19126
rect 47333 18916 47543 19126
rect 47543 18916 47547 19126
rect 47329 18912 47547 18916
rect 50517 19007 50735 19011
rect 50517 18797 50521 19007
rect 50521 18797 50731 19007
rect 50731 18797 50735 19007
rect 50517 18793 50735 18797
rect 53538 19038 53756 19042
rect 53538 18828 53542 19038
rect 53542 18828 53752 19038
rect 53752 18828 53756 19038
rect 53538 18824 53756 18828
rect 56616 19158 56834 19162
rect 56616 18948 56620 19158
rect 56620 18948 56830 19158
rect 56830 18948 56834 19158
rect 56616 18944 56834 18948
rect 59631 18862 59849 18866
rect 59631 18652 59635 18862
rect 59635 18652 59845 18862
rect 59845 18652 59849 18862
rect 59631 18648 59849 18652
rect 62633 18786 62851 18790
rect 62633 18576 62637 18786
rect 62637 18576 62847 18786
rect 62847 18576 62851 18786
rect 62633 18572 62851 18576
rect 64257 18755 64575 18759
rect 64257 18445 64261 18755
rect 64261 18445 64571 18755
rect 64571 18445 64575 18755
rect 64257 18441 64575 18445
rect 65743 18877 65961 18881
rect 65743 18667 65747 18877
rect 65747 18667 65957 18877
rect 65957 18667 65961 18877
rect 65743 18663 65961 18667
rect 68329 18734 68547 18952
rect 71929 18842 72147 19060
rect 75079 19026 75297 19030
rect 75079 18816 75083 19026
rect 75083 18816 75293 19026
rect 75293 18816 75297 19026
rect 75079 18812 75297 18816
rect 81191 18706 81409 18905
rect 81191 18687 81195 18706
rect 81195 18687 81405 18706
rect 81405 18687 81409 18706
rect 2329 18435 2547 18439
rect 2329 18225 2333 18435
rect 2333 18225 2543 18435
rect 2543 18225 2547 18435
rect 2329 18221 2547 18225
rect 90413 18833 90631 18837
rect 90413 18623 90417 18833
rect 90417 18623 90627 18833
rect 90627 18623 90631 18833
rect 90413 18619 90631 18623
rect 93557 18789 93775 18793
rect 93557 18579 93561 18789
rect 93561 18579 93771 18789
rect 93771 18579 93775 18789
rect 93557 18575 93775 18579
rect 96454 18871 96672 18875
rect 96454 18661 96458 18871
rect 96458 18661 96668 18871
rect 96668 18661 96672 18871
rect 96454 18657 96672 18661
rect 108902 19028 109120 19032
rect 108902 18818 108906 19028
rect 108906 18818 109116 19028
rect 109116 18818 109120 19028
rect 108902 18814 109120 18818
rect 102712 18736 102930 18740
rect 102712 18526 102716 18736
rect 102716 18526 102926 18736
rect 102926 18526 102930 18736
rect 102712 18522 102930 18526
rect 105676 18751 105894 18755
rect 105676 18541 105680 18751
rect 105680 18541 105890 18751
rect 105890 18541 105894 18751
rect 105676 18537 105894 18541
rect 111949 18931 112167 18935
rect 111949 18721 111953 18931
rect 111953 18721 112163 18931
rect 112163 18721 112167 18931
rect 111949 18717 112167 18721
rect 114954 18980 115172 18984
rect 114954 18770 114958 18980
rect 114958 18770 115168 18980
rect 115168 18770 115172 18980
rect 114954 18766 115172 18770
rect 117969 18973 118187 18977
rect 117969 18763 117973 18973
rect 117973 18763 118183 18973
rect 118183 18763 118187 18973
rect 117969 18759 118187 18763
rect 121151 18860 121369 18864
rect 121151 18650 121155 18860
rect 121155 18650 121365 18860
rect 121365 18650 121369 18860
rect 121151 18646 121369 18650
rect 78099 18088 78317 18306
rect -6204 17747 -6199 17942
rect -6199 17747 -5999 17942
rect -5999 17747 -5994 17942
rect 84275 18185 84493 18403
rect 87336 18310 87554 18314
rect 87336 18100 87340 18310
rect 87340 18100 87550 18310
rect 87550 18100 87554 18310
rect 87336 18096 87554 18100
rect 99598 18497 99816 18501
rect 99598 18287 99602 18497
rect 99602 18287 99812 18497
rect 99812 18287 99816 18497
rect 99598 18283 99816 18287
rect 121679 18755 121997 18759
rect 121679 18445 121683 18755
rect 121683 18445 121993 18755
rect 121993 18445 121997 18755
rect 121679 18441 121997 18445
rect 124119 18633 124337 18851
rect 127242 18938 127460 18942
rect 127242 18728 127246 18938
rect 127246 18728 127456 18938
rect 127456 18728 127460 18938
rect 127242 18724 127460 18728
rect 130251 18809 130469 18813
rect 130251 18599 130255 18809
rect 130255 18599 130465 18809
rect 130465 18599 130469 18809
rect 130251 18595 130469 18599
rect 133413 18648 133631 18866
rect 139553 18596 139771 18600
rect 139553 18386 139557 18596
rect 139557 18386 139767 18596
rect 139767 18386 139771 18596
rect 139553 18382 139771 18386
rect 142600 18664 142818 18668
rect 142600 18454 142604 18664
rect 142604 18454 142814 18664
rect 142814 18454 142818 18664
rect 142600 18450 142818 18454
rect 145579 18839 145797 18843
rect 145579 18629 145583 18839
rect 145583 18629 145793 18839
rect 145793 18629 145797 18839
rect 145579 18625 145797 18629
rect 148755 18839 148973 18843
rect 148755 18629 148759 18839
rect 148759 18629 148969 18839
rect 148969 18629 148973 18839
rect 148755 18625 148973 18629
rect 151773 18770 151991 18774
rect 151773 18560 151777 18770
rect 151777 18560 151987 18770
rect 151987 18560 151991 18770
rect 151773 18556 151991 18560
rect 154793 18854 155011 18858
rect 154793 18644 154797 18854
rect 154797 18644 155007 18854
rect 155007 18644 155011 18854
rect 154793 18640 155011 18644
rect 157844 18993 158062 18997
rect 157844 18783 157848 18993
rect 157848 18783 158058 18993
rect 158058 18783 158062 18993
rect 157844 18779 158062 18783
rect 174367 19131 174585 19135
rect 174367 18921 174371 19131
rect 174371 18921 174581 19131
rect 174581 18921 174585 19131
rect 174367 18917 174585 18921
rect 160887 18754 161105 18758
rect 160887 18544 160891 18754
rect 160891 18544 161101 18754
rect 161101 18544 161105 18754
rect 160887 18540 161105 18544
rect 163239 18455 163457 18459
rect 163239 18245 163243 18455
rect 163243 18245 163453 18455
rect 163453 18245 163457 18455
rect 163239 18241 163457 18245
rect 167549 18755 167867 18759
rect 167549 18445 167553 18755
rect 167553 18445 167863 18755
rect 167863 18445 167867 18755
rect 167549 18441 167867 18445
rect 176329 18808 176547 18812
rect 176329 18598 176333 18808
rect 176333 18598 176543 18808
rect 176543 18598 176547 18808
rect 176329 18594 176547 18598
rect 173083 18485 173301 18489
rect 173083 18275 173087 18485
rect 173087 18275 173297 18485
rect 173297 18275 173301 18485
rect 173083 18271 173301 18275
rect 180549 18755 180867 18759
rect 180549 18445 180553 18755
rect 180553 18445 180863 18755
rect 180863 18445 180867 18755
rect 180549 18441 180867 18445
rect 189549 18755 189867 18759
rect 189549 18445 189553 18755
rect 189553 18445 189863 18755
rect 189863 18445 189867 18755
rect 189549 18441 189867 18445
rect 198549 18755 198867 18759
rect 198549 18445 198553 18755
rect 198553 18445 198863 18755
rect 198863 18445 198867 18755
rect 198549 18441 198867 18445
rect 204549 18755 204867 18759
rect 204549 18445 204553 18755
rect 204553 18445 204863 18755
rect 204863 18445 204867 18755
rect 204549 18441 204867 18445
rect 136468 18237 136686 18241
rect 136468 18027 136472 18237
rect 136472 18027 136682 18237
rect 136682 18027 136686 18237
rect 136468 18023 136686 18027
rect 206329 18451 206547 18455
rect 206329 18241 206333 18451
rect 206333 18241 206543 18451
rect 206543 18241 206547 18451
rect 206329 18237 206547 18241
rect 211549 18755 211867 18759
rect 211549 18445 211553 18755
rect 211553 18445 211863 18755
rect 211863 18445 211867 18755
rect 211549 18441 211867 18445
rect 215329 18559 215547 18563
rect 215329 18349 215333 18559
rect 215333 18349 215543 18559
rect 215543 18349 215547 18559
rect 215329 18345 215547 18349
rect 223549 18755 223867 18759
rect 223549 18445 223553 18755
rect 223553 18445 223863 18755
rect 223863 18445 223867 18755
rect 223549 18441 223867 18445
rect 229659 18935 229877 18939
rect 229659 18725 229663 18935
rect 229663 18725 229873 18935
rect 229873 18725 229877 18935
rect 229659 18721 229877 18725
rect 232549 18755 232867 18759
rect 232549 18445 232553 18755
rect 232553 18445 232863 18755
rect 232863 18445 232867 18755
rect 232549 18441 232867 18445
rect 233329 18685 233547 18689
rect 233329 18475 233333 18685
rect 233333 18475 233543 18685
rect 233543 18475 233547 18685
rect 233329 18471 233547 18475
rect 238549 18755 238867 18759
rect 238549 18445 238553 18755
rect 238553 18445 238863 18755
rect 238863 18445 238867 18755
rect 238549 18441 238867 18445
rect 227195 18424 227413 18428
rect 227195 18214 227199 18424
rect 227199 18214 227409 18424
rect 227409 18214 227413 18424
rect 227195 18210 227413 18214
rect 241673 18530 241891 18534
rect 241673 18320 241677 18530
rect 241677 18320 241887 18530
rect 241887 18320 241891 18530
rect 241673 18316 241891 18320
rect 242329 18566 242547 18570
rect 242329 18356 242333 18566
rect 242333 18356 242543 18566
rect 242543 18356 242547 18566
rect 242329 18352 242547 18356
rect 250549 18755 250867 18759
rect 250549 18445 250553 18755
rect 250553 18445 250863 18755
rect 250863 18445 250867 18755
rect 250549 18441 250867 18445
rect 165929 18170 166147 18174
rect 165929 17960 165933 18170
rect 165933 17960 166143 18170
rect 166143 17960 166147 18170
rect 165929 17956 166147 17960
rect -6204 17742 -5994 17747
rect 182474 17855 182692 17859
rect 182474 17645 182478 17855
rect 182478 17645 182688 17855
rect 182688 17645 182692 17855
rect 182474 17641 182692 17645
rect 185329 18032 185547 18036
rect 185329 17822 185333 18032
rect 185333 17822 185543 18032
rect 185543 17822 185547 18032
rect 185329 17818 185547 17822
rect 196794 17925 197012 17929
rect 196794 17715 196798 17925
rect 196798 17715 197008 17925
rect 197008 17715 197012 17925
rect 196794 17711 197012 17715
rect 200916 17952 201134 17956
rect 200916 17742 200920 17952
rect 200920 17742 201130 17952
rect 201130 17742 201134 17952
rect 200916 17738 201134 17742
rect 213156 18094 213374 18098
rect 213156 17884 213160 18094
rect 213160 17884 213370 18094
rect 213370 17884 213374 18094
rect 213156 17880 213374 17884
rect 234651 18299 234869 18303
rect 234651 18089 234655 18299
rect 234655 18089 234865 18299
rect 234865 18089 234869 18299
rect 234651 18085 234869 18089
rect 253926 18505 254144 18509
rect 253926 18295 253930 18505
rect 253930 18295 254140 18505
rect 254140 18295 254144 18505
rect 253926 18291 254144 18295
rect 254329 18696 254547 18700
rect 254329 18486 254333 18696
rect 254333 18486 254543 18696
rect 254543 18486 254547 18696
rect 254329 18482 254547 18486
rect 263949 18755 264267 18759
rect 263949 18445 263953 18755
rect 263953 18445 264263 18755
rect 264263 18445 264267 18755
rect 263949 18441 264267 18445
rect 269033 18556 269251 18560
rect 269033 18346 269037 18556
rect 269037 18346 269247 18556
rect 269247 18346 269251 18556
rect 269033 18342 269251 18346
rect 269949 18755 270267 18759
rect 269949 18445 269953 18755
rect 269953 18445 270263 18755
rect 270263 18445 270267 18755
rect 269949 18441 270267 18445
rect 272949 18755 273267 18759
rect 272949 18445 272953 18755
rect 272953 18445 273263 18755
rect 273263 18445 273267 18755
rect 272949 18441 273267 18445
rect 275949 18755 276267 18759
rect 275949 18445 275953 18755
rect 275953 18445 276263 18755
rect 276263 18445 276267 18755
rect 275949 18441 276267 18445
rect 279677 18694 279895 18698
rect 279677 18484 279681 18694
rect 279681 18484 279891 18694
rect 279891 18484 279895 18694
rect 279677 18480 279895 18484
rect 281949 18755 282267 18759
rect 281949 18445 281953 18755
rect 281953 18445 282263 18755
rect 282263 18445 282267 18755
rect 281949 18441 282267 18445
rect 285949 18755 286267 18759
rect 285949 18445 285953 18755
rect 285953 18445 286263 18755
rect 286263 18445 286267 18755
rect 285949 18441 286267 18445
rect 290329 18951 290547 18955
rect 290329 18741 290333 18951
rect 290333 18741 290543 18951
rect 290543 18741 290547 18951
rect 290329 18737 290547 18741
rect 305386 19095 305604 19099
rect 305386 18885 305390 19095
rect 305390 18885 305600 19095
rect 305600 18885 305604 19095
rect 305386 18881 305604 18885
rect 293949 18755 294267 18759
rect 293949 18445 293953 18755
rect 293953 18445 294263 18755
rect 294263 18445 294267 18755
rect 293949 18441 294267 18445
rect 296949 18755 297267 18759
rect 296949 18445 296953 18755
rect 296953 18445 297263 18755
rect 297263 18445 297267 18755
rect 296949 18441 297267 18445
rect 299949 18755 300267 18759
rect 299949 18445 299953 18755
rect 299953 18445 300263 18755
rect 300263 18445 300267 18755
rect 299949 18441 300267 18445
rect 302949 18755 303267 18759
rect 302949 18445 302953 18755
rect 302953 18445 303263 18755
rect 303263 18445 303267 18755
rect 302949 18441 303267 18445
rect 240917 18011 241135 18015
rect 240917 17801 240921 18011
rect 240921 17801 241131 18011
rect 241131 17801 241135 18011
rect 240917 17797 241135 17801
rect 261045 18121 261263 18125
rect 261045 17911 261049 18121
rect 261049 17911 261259 18121
rect 261259 17911 261263 18121
rect 261045 17907 261263 17911
rect 269329 18264 269547 18268
rect 269329 18054 269333 18264
rect 269333 18054 269543 18264
rect 269543 18054 269547 18264
rect 269329 18050 269547 18054
rect 278879 18202 279097 18206
rect 278879 17992 278883 18202
rect 278883 17992 279093 18202
rect 279093 17992 279097 18202
rect 278879 17988 279097 17992
rect 188329 17655 188547 17659
rect 188329 17445 188333 17655
rect 188333 17445 188543 17655
rect 188543 17445 188547 17655
rect 188329 17441 188547 17445
rect 207000 17747 207218 17751
rect 207000 17537 207004 17747
rect 207004 17537 207214 17747
rect 207214 17537 207218 17747
rect 207000 17533 207218 17537
rect 221329 17707 221547 17711
rect 221329 17497 221333 17707
rect 221333 17497 221543 17707
rect 221543 17497 221547 17707
rect 221329 17493 221547 17497
rect 249668 17856 249886 17860
rect 249668 17646 249672 17856
rect 249672 17646 249882 17856
rect 249882 17646 249886 17856
rect 249668 17642 249886 17646
rect 265871 17959 266089 17963
rect 265871 17749 265875 17959
rect 265875 17749 266085 17959
rect 266085 17749 266089 17959
rect 265871 17745 266089 17749
rect 284329 18133 284547 18137
rect 284329 17923 284333 18133
rect 284333 17923 284543 18133
rect 284543 17923 284547 18133
rect 284329 17919 284547 17923
rect 292408 18223 292626 18227
rect 292408 18013 292412 18223
rect 292412 18013 292622 18223
rect 292622 18013 292626 18223
rect 292408 18009 292626 18013
rect 168864 17417 169082 17421
rect 168864 17207 168868 17417
rect 168868 17207 169078 17417
rect 169078 17207 169082 17417
rect 168864 17203 169082 17207
rect 277694 17578 277912 17582
rect 277694 17368 277698 17578
rect 277698 17368 277908 17578
rect 277908 17368 277912 17578
rect 277694 17364 277912 17368
rect 286930 17508 287148 17512
rect 286930 17298 286934 17508
rect 286934 17298 287144 17508
rect 287144 17298 287148 17508
rect 286930 17294 287148 17298
rect 299259 17719 299477 17723
rect 299259 17509 299263 17719
rect 299263 17509 299473 17719
rect 299473 17509 299477 17719
rect 299259 17505 299477 17509
rect 184011 17148 184229 17152
rect 184011 16938 184015 17148
rect 184015 16938 184225 17148
rect 184225 16938 184229 17148
rect 184011 16934 184229 16938
rect 213905 17265 214123 17269
rect 213905 17055 213909 17265
rect 213909 17055 214119 17265
rect 214119 17055 214123 17265
rect 213905 17051 214123 17055
rect 193466 17015 193684 17019
rect 193466 16805 193470 17015
rect 193470 16805 193680 17015
rect 193680 16805 193684 17015
rect 193466 16801 193684 16805
rect 220689 17224 220907 17228
rect 220689 17014 220693 17224
rect 220693 17014 220903 17224
rect 220903 17014 220907 17224
rect 220689 17010 220907 17014
rect 202004 16890 202222 16894
rect 202004 16680 202008 16890
rect 202008 16680 202218 16890
rect 202218 16680 202222 16890
rect 202004 16676 202222 16680
rect 248712 17073 248930 17077
rect 248712 16863 248716 17073
rect 248716 16863 248926 17073
rect 248926 16863 248930 17073
rect 248712 16859 248930 16863
rect 260054 17242 260272 17246
rect 260054 17032 260058 17242
rect 260058 17032 260268 17242
rect 260268 17032 260272 17242
rect 260054 17028 260272 17032
rect 300252 17101 300470 17105
rect 300252 16891 300256 17101
rect 300256 16891 300466 17101
rect 300466 16891 300470 17101
rect 300252 16887 300470 16891
rect 302942 16094 302947 16411
rect 302947 16094 303269 16411
rect 303269 16094 303274 16411
rect 302942 16089 303274 16094
rect 103 15388 108 15583
rect 108 15388 308 15583
rect 308 15388 313 15583
rect 103 15383 313 15388
rect 3659 15374 3664 15689
rect 3664 15374 3984 15689
rect 3984 15374 3989 15689
rect 18083 15392 18088 15707
rect 18088 15392 18408 15707
rect 18408 15392 18413 15707
rect 18083 15387 18413 15392
rect 3659 15369 3989 15374
rect 32909 15368 32914 15683
rect 32914 15368 33234 15683
rect 33234 15368 33239 15683
rect 32909 15363 33239 15368
rect 64251 15376 64256 15691
rect 64256 15376 64576 15691
rect 64576 15376 64581 15691
rect 121673 15390 121678 15705
rect 121678 15390 121998 15705
rect 121998 15390 122003 15705
rect 121673 15385 122003 15390
rect 167543 15392 167548 15707
rect 167548 15392 167868 15707
rect 167868 15392 167873 15707
rect 167543 15387 167873 15392
rect 180543 15392 180548 15707
rect 180548 15392 180868 15707
rect 180868 15392 180873 15707
rect 180543 15387 180873 15392
rect 189543 15392 189548 15707
rect 189548 15392 189868 15707
rect 189868 15392 189873 15707
rect 189543 15387 189873 15392
rect 198543 15392 198548 15707
rect 198548 15392 198868 15707
rect 198868 15392 198873 15707
rect 198543 15387 198873 15392
rect 204543 15392 204548 15707
rect 204548 15392 204868 15707
rect 204868 15392 204873 15707
rect 204543 15387 204873 15392
rect 211543 15392 211548 15707
rect 211548 15392 211868 15707
rect 211868 15392 211873 15707
rect 211543 15387 211873 15392
rect 223543 15392 223548 15707
rect 223548 15392 223868 15707
rect 223868 15392 223873 15707
rect 223543 15387 223873 15392
rect 232543 15392 232548 15707
rect 232548 15392 232868 15707
rect 232868 15392 232873 15707
rect 232543 15387 232873 15392
rect 238543 15392 238548 15707
rect 238548 15392 238868 15707
rect 238868 15392 238873 15707
rect 238543 15387 238873 15392
rect 250543 15392 250548 15707
rect 250548 15392 250868 15707
rect 250868 15392 250873 15707
rect 250543 15387 250873 15392
rect 263943 15392 263948 15707
rect 263948 15392 264268 15707
rect 264268 15392 264273 15707
rect 263943 15387 264273 15392
rect 269943 15392 269948 15707
rect 269948 15392 270268 15707
rect 270268 15392 270273 15707
rect 269943 15387 270273 15392
rect 272943 15392 272948 15707
rect 272948 15392 273268 15707
rect 273268 15392 273273 15707
rect 272943 15387 273273 15392
rect 275943 15392 275948 15707
rect 275948 15392 276268 15707
rect 276268 15392 276273 15707
rect 275943 15387 276273 15392
rect 281943 15392 281948 15707
rect 281948 15392 282268 15707
rect 282268 15392 282273 15707
rect 281943 15387 282273 15392
rect 285943 15392 285948 15707
rect 285948 15392 286268 15707
rect 286268 15392 286273 15707
rect 285943 15387 286273 15392
rect 293943 15392 293948 15707
rect 293948 15392 294268 15707
rect 294268 15392 294273 15707
rect 293943 15387 294273 15392
rect 296943 15392 296948 15707
rect 296948 15392 297268 15707
rect 297268 15392 297273 15707
rect 296943 15387 297273 15392
rect 299943 15392 299948 15707
rect 299948 15392 300268 15707
rect 300268 15392 300273 15707
rect 299943 15387 300273 15392
rect 302943 15392 302948 15707
rect 302948 15392 303268 15707
rect 303268 15392 303273 15707
rect 302943 15387 303273 15392
rect 64251 15371 64581 15376
<< metal4 >>
rect -7597 325867 -763 325977
rect -5203 322052 -1206 322076
rect -5203 321780 -1502 322052
rect -1230 321780 -1206 322052
rect -5203 321760 -1206 321780
rect -5203 321756 -1526 321760
rect -873 320928 -763 325867
rect 303926 321357 304246 321358
rect 303926 321039 303927 321357
rect 304245 321039 304246 321357
rect 303926 321038 304246 321039
rect -5974 319800 -3762 320120
rect -2007 319922 -1805 319923
rect -2674 319722 -2006 319922
rect -1806 319722 -1805 319922
rect -2007 319721 -1805 319722
rect -5203 319052 -1206 319076
rect -5203 318780 -1502 319052
rect -1230 318780 -1206 319052
rect -5203 318760 -1206 318780
rect -5203 318756 -1526 318760
rect 303926 318357 304246 318358
rect 303926 318039 303927 318357
rect 304245 318039 304246 318357
rect 303926 318038 304246 318039
rect -5974 316800 -3762 317120
rect -2007 316922 -1805 316923
rect -2674 316722 -2006 316922
rect -1806 316722 -1805 316922
rect -2007 316721 -1805 316722
rect -5203 316052 -1206 316076
rect -5203 315780 -1502 316052
rect -1230 315780 -1206 316052
rect -5203 315760 -1206 315780
rect -5203 315756 -1526 315760
rect 303926 315357 304246 315358
rect 303926 315039 303927 315357
rect 304245 315039 304246 315357
rect 303926 315038 304246 315039
rect -5974 313800 -3762 314120
rect -2007 313922 -1805 313923
rect -2674 313722 -2006 313922
rect -1806 313722 -1805 313922
rect -2007 313721 -1805 313722
rect -5203 313052 -1206 313076
rect -5203 312780 -1502 313052
rect -1230 312780 -1206 313052
rect -5203 312760 -1206 312780
rect -5203 312756 -1526 312760
rect 303926 312357 304246 312358
rect 303926 312039 303927 312357
rect 304245 312039 304246 312357
rect 303926 312038 304246 312039
rect -5974 310800 -3762 311120
rect -2007 310922 -1805 310923
rect -2674 310722 -2006 310922
rect -1806 310722 -1805 310922
rect -2007 310721 -1805 310722
rect -5203 310052 -1206 310076
rect -5203 309780 -1502 310052
rect -1230 309780 -1206 310052
rect -5203 309760 -1206 309780
rect -5203 309756 -1526 309760
rect 303926 309357 304246 309358
rect 303926 309039 303927 309357
rect 304245 309039 304246 309357
rect 303926 309038 304246 309039
rect -5974 307800 -3762 308120
rect -2007 307922 -1805 307923
rect -2674 307722 -2006 307922
rect -1806 307722 -1805 307922
rect -2007 307721 -1805 307722
rect -5203 307052 -1206 307076
rect -5203 306780 -1502 307052
rect -1230 306780 -1206 307052
rect -5203 306760 -1206 306780
rect -5203 306756 -1526 306760
rect 303926 306357 304246 306358
rect 303926 306039 303927 306357
rect 304245 306039 304246 306357
rect 303926 306038 304246 306039
rect -5974 304800 -3762 305120
rect -2007 304922 -1805 304923
rect -2674 304722 -2006 304922
rect -1806 304722 -1805 304922
rect -2007 304721 -1805 304722
rect -5203 304052 -1206 304076
rect -5203 303780 -1502 304052
rect -1230 303780 -1206 304052
rect -5203 303760 -1206 303780
rect -5203 303756 -1526 303760
rect 303926 303357 304246 303358
rect 303926 303039 303927 303357
rect 304245 303039 304246 303357
rect 303926 303038 304246 303039
rect -5974 301800 -3762 302120
rect -2007 301922 -1805 301923
rect -2674 301722 -2006 301922
rect -1806 301722 -1805 301922
rect -2007 301721 -1805 301722
rect -5203 301052 -1206 301076
rect -5203 300780 -1502 301052
rect -1230 300780 -1206 301052
rect -5203 300760 -1206 300780
rect -5203 300756 -1526 300760
rect 303926 300357 304246 300358
rect 303926 300039 303927 300357
rect 304245 300039 304246 300357
rect 303926 300038 304246 300039
rect -5974 298800 -3762 299120
rect -2007 298922 -1805 298923
rect -2674 298722 -2006 298922
rect -1806 298722 -1805 298922
rect -2007 298721 -1805 298722
rect -5203 298052 -1206 298076
rect -5203 297780 -1502 298052
rect -1230 297780 -1206 298052
rect -5203 297760 -1206 297780
rect -5203 297756 -1526 297760
rect 303926 297357 304246 297358
rect 303926 297039 303927 297357
rect 304245 297039 304246 297357
rect 303926 297038 304246 297039
rect -5974 295800 -3762 296120
rect -2007 295922 -1805 295923
rect -2674 295722 -2006 295922
rect -1806 295722 -1805 295922
rect -2007 295721 -1805 295722
rect -5203 295052 -1206 295076
rect -5203 294780 -1502 295052
rect -1230 294780 -1206 295052
rect -5203 294760 -1206 294780
rect -5203 294756 -1526 294760
rect 303926 294357 304246 294358
rect 303926 294039 303927 294357
rect 304245 294039 304246 294357
rect 303926 294038 304246 294039
rect -5974 292800 -3762 293120
rect -2007 292922 -1805 292923
rect -2674 292722 -2006 292922
rect -1806 292722 -1805 292922
rect -2007 292721 -1805 292722
rect -5203 292052 -1206 292076
rect -5203 291780 -1502 292052
rect -1230 291780 -1206 292052
rect -5203 291760 -1206 291780
rect -5203 291756 -1526 291760
rect 303926 291357 304246 291358
rect 303926 291039 303927 291357
rect 304245 291039 304246 291357
rect 303926 291038 304246 291039
rect -5974 289800 -3762 290120
rect -2007 289922 -1805 289923
rect -2674 289722 -2006 289922
rect -1806 289722 -1805 289922
rect -2007 289721 -1805 289722
rect -5203 289052 -1206 289076
rect -5203 288780 -1502 289052
rect -1230 288780 -1206 289052
rect -5203 288760 -1206 288780
rect -5203 288756 -1526 288760
rect 303926 288357 304246 288358
rect 303926 288039 303927 288357
rect 304245 288039 304246 288357
rect 303926 288038 304246 288039
rect -5974 286800 -3762 287120
rect -2007 286922 -1805 286923
rect -2674 286722 -2006 286922
rect -1806 286722 -1805 286922
rect -2007 286721 -1805 286722
rect -5203 286052 -1206 286076
rect -5203 285780 -1502 286052
rect -1230 285780 -1206 286052
rect -5203 285760 -1206 285780
rect -5203 285756 -1526 285760
rect 303926 285357 304246 285358
rect 303926 285039 303927 285357
rect 304245 285039 304246 285357
rect 303926 285038 304246 285039
rect -5974 283800 -3762 284120
rect -2007 283922 -1805 283923
rect -2674 283722 -2006 283922
rect -1806 283722 -1805 283922
rect -2007 283721 -1805 283722
rect -5203 283052 -1206 283076
rect -5203 282780 -1502 283052
rect -1230 282780 -1206 283052
rect -5203 282760 -1206 282780
rect -5203 282756 -1526 282760
rect 303926 282357 304246 282358
rect 303926 282039 303927 282357
rect 304245 282039 304246 282357
rect 303926 282038 304246 282039
rect -5974 280800 -3762 281120
rect -2007 280922 -1805 280923
rect -2674 280722 -2006 280922
rect -1806 280722 -1805 280922
rect -2007 280721 -1805 280722
rect -5203 280052 -1206 280076
rect -5203 279780 -1502 280052
rect -1230 279780 -1206 280052
rect -5203 279760 -1206 279780
rect -5203 279756 -1526 279760
rect 303926 279357 304246 279358
rect 303926 279039 303927 279357
rect 304245 279039 304246 279357
rect 303926 279038 304246 279039
rect -5974 277800 -3762 278120
rect -2007 277922 -1805 277923
rect -2674 277722 -2006 277922
rect -1806 277722 -1805 277922
rect -2007 277721 -1805 277722
rect -5203 277052 -1206 277076
rect -5203 276780 -1502 277052
rect -1230 276780 -1206 277052
rect -5203 276760 -1206 276780
rect -5203 276756 -1526 276760
rect 303926 276357 304246 276358
rect 303926 276039 303927 276357
rect 304245 276039 304246 276357
rect 303926 276038 304246 276039
rect -5974 274800 -3762 275120
rect -2007 274922 -1805 274923
rect -2674 274722 -2006 274922
rect -1806 274722 -1805 274922
rect -2007 274721 -1805 274722
rect -5203 274052 -1206 274076
rect -5203 273780 -1502 274052
rect -1230 273780 -1206 274052
rect -5203 273760 -1206 273780
rect -5203 273756 -1526 273760
rect 303926 273357 304246 273358
rect 303926 273039 303927 273357
rect 304245 273039 304246 273357
rect 303926 273038 304246 273039
rect -5974 271800 -3762 272120
rect -2007 271922 -1805 271923
rect -2674 271722 -2006 271922
rect -1806 271722 -1805 271922
rect -2007 271721 -1805 271722
rect -5203 271052 -1206 271076
rect -5203 270780 -1502 271052
rect -1230 270780 -1206 271052
rect -5203 270760 -1206 270780
rect -5203 270756 -1526 270760
rect 303926 270357 304246 270358
rect 303926 270039 303927 270357
rect 304245 270039 304246 270357
rect 303926 270038 304246 270039
rect -5974 268800 -3762 269120
rect -2007 268922 -1805 268923
rect -2674 268722 -2006 268922
rect -1806 268722 -1805 268922
rect -2007 268721 -1805 268722
rect -5203 268052 -1206 268076
rect -5203 267780 -1502 268052
rect -1230 267780 -1206 268052
rect -5203 267760 -1206 267780
rect -5203 267756 -1526 267760
rect 303926 267357 304246 267358
rect 303926 267039 303927 267357
rect 304245 267039 304246 267357
rect 303926 267038 304246 267039
rect -5974 265800 -3762 266120
rect -2007 265922 -1805 265923
rect -2674 265722 -2006 265922
rect -1806 265722 -1805 265922
rect -2007 265721 -1805 265722
rect -5203 265052 -1206 265076
rect -5203 264780 -1502 265052
rect -1230 264780 -1206 265052
rect -5203 264760 -1206 264780
rect -5203 264756 -1526 264760
rect 303926 264357 304246 264358
rect 303926 264039 303927 264357
rect 304245 264039 304246 264357
rect 303926 264038 304246 264039
rect -5974 262800 -3762 263120
rect -2007 262922 -1805 262923
rect -2674 262722 -2006 262922
rect -1806 262722 -1805 262922
rect -2007 262721 -1805 262722
rect -5203 262052 -1206 262076
rect -5203 261780 -1502 262052
rect -1230 261780 -1206 262052
rect -5203 261760 -1206 261780
rect -5203 261756 -1526 261760
rect 303926 261357 304246 261358
rect 303926 261039 303927 261357
rect 304245 261039 304246 261357
rect 303926 261038 304246 261039
rect -5974 259800 -3762 260120
rect -2007 259922 -1805 259923
rect -2674 259722 -2006 259922
rect -1806 259722 -1805 259922
rect -2007 259721 -1805 259722
rect -5203 259052 -1206 259076
rect -5203 258780 -1502 259052
rect -1230 258780 -1206 259052
rect -5203 258760 -1206 258780
rect -5203 258756 -1526 258760
rect 303926 258357 304246 258358
rect 303926 258039 303927 258357
rect 304245 258039 304246 258357
rect 303926 258038 304246 258039
rect -5974 256800 -3762 257120
rect -2007 256922 -1805 256923
rect -2674 256722 -2006 256922
rect -1806 256722 -1805 256922
rect -2007 256721 -1805 256722
rect -5203 256052 -1206 256076
rect -5203 255780 -1502 256052
rect -1230 255780 -1206 256052
rect -5203 255760 -1206 255780
rect -5203 255756 -1526 255760
rect 303926 255357 304246 255358
rect 303926 255039 303927 255357
rect 304245 255039 304246 255357
rect 303926 255038 304246 255039
rect -5974 253800 -3762 254120
rect -2007 253922 -1805 253923
rect -2674 253722 -2006 253922
rect -1806 253722 -1805 253922
rect -2007 253721 -1805 253722
rect -5203 253052 -1206 253076
rect -5203 252780 -1502 253052
rect -1230 252780 -1206 253052
rect -5203 252760 -1206 252780
rect -5203 252756 -1526 252760
rect 303926 252357 304246 252358
rect 303926 252039 303927 252357
rect 304245 252039 304246 252357
rect 303926 252038 304246 252039
rect -5974 250800 -3762 251120
rect -2007 250922 -1805 250923
rect -2674 250722 -2006 250922
rect -1806 250722 -1805 250922
rect -2007 250721 -1805 250722
rect -5203 250052 -1206 250076
rect -5203 249780 -1502 250052
rect -1230 249780 -1206 250052
rect -5203 249760 -1206 249780
rect -5203 249756 -1526 249760
rect 303926 249357 304246 249358
rect 303926 249039 303927 249357
rect 304245 249039 304246 249357
rect 303926 249038 304246 249039
rect -5974 247800 -3762 248120
rect -2007 247922 -1805 247923
rect -2674 247722 -2006 247922
rect -1806 247722 -1805 247922
rect -2007 247721 -1805 247722
rect 303926 246357 304246 246358
rect 303926 246039 303927 246357
rect 304245 246039 304246 246357
rect 303926 246038 304246 246039
rect -5974 244800 -3762 245120
rect -2007 244922 -1805 244923
rect -2674 244722 -2006 244922
rect -1806 244722 -1805 244922
rect -2007 244721 -1805 244722
rect -5203 244052 -1206 244076
rect -5203 243780 -1502 244052
rect -1230 243780 -1206 244052
rect -5203 243760 -1206 243780
rect -5203 243756 -1526 243760
rect 303926 243357 304246 243358
rect 303926 243039 303927 243357
rect 304245 243039 304246 243357
rect 303926 243038 304246 243039
rect -5974 241800 -3762 242120
rect -2007 241922 -1805 241923
rect -2674 241722 -2006 241922
rect -1806 241722 -1805 241922
rect -2007 241721 -1805 241722
rect -5203 241052 -1206 241076
rect -5203 240780 -1502 241052
rect -1230 240780 -1206 241052
rect -5203 240760 -1206 240780
rect -5203 240756 -1526 240760
rect 303926 240357 304246 240358
rect 303926 240039 303927 240357
rect 304245 240039 304246 240357
rect 303926 240038 304246 240039
rect -5974 238800 -3762 239120
rect -2007 238922 -1805 238923
rect -2674 238722 -2006 238922
rect -1806 238722 -1805 238922
rect -2007 238721 -1805 238722
rect -5203 238052 -1206 238076
rect -5203 237780 -1502 238052
rect -1230 237780 -1206 238052
rect -5203 237760 -1206 237780
rect -5203 237756 -1526 237760
rect 303926 237357 304246 237358
rect 303926 237039 303927 237357
rect 304245 237039 304246 237357
rect 303926 237038 304246 237039
rect -5974 235800 -3762 236120
rect -2007 235922 -1805 235923
rect -2674 235722 -2006 235922
rect -1806 235722 -1805 235922
rect -2007 235721 -1805 235722
rect -5203 235052 -1206 235076
rect -5203 234780 -1502 235052
rect -1230 234780 -1206 235052
rect -5203 234760 -1206 234780
rect -5203 234756 -1526 234760
rect 303926 234357 304246 234358
rect 303926 234039 303927 234357
rect 304245 234039 304246 234357
rect 303926 234038 304246 234039
rect -5974 232800 -3762 233120
rect -2007 232922 -1805 232923
rect -2674 232722 -2006 232922
rect -1806 232722 -1805 232922
rect -2007 232721 -1805 232722
rect -5203 232052 -1206 232076
rect -5203 231780 -1502 232052
rect -1230 231780 -1206 232052
rect -5203 231760 -1206 231780
rect -5203 231756 -1526 231760
rect 303926 231357 304246 231358
rect 303926 231039 303927 231357
rect 304245 231039 304246 231357
rect 303926 231038 304246 231039
rect -5974 229800 -3762 230120
rect -2007 229922 -1805 229923
rect -2674 229722 -2006 229922
rect -1806 229722 -1805 229922
rect -2007 229721 -1805 229722
rect -5203 229052 -1206 229076
rect -5203 228780 -1502 229052
rect -1230 228780 -1206 229052
rect -5203 228760 -1206 228780
rect -5203 228756 -1526 228760
rect 303926 228357 304246 228358
rect 303926 228039 303927 228357
rect 304245 228039 304246 228357
rect 303926 228038 304246 228039
rect -5974 226800 -3762 227120
rect -2007 226922 -1805 226923
rect -2674 226722 -2006 226922
rect -1806 226722 -1805 226922
rect -2007 226721 -1805 226722
rect -5203 226052 -1206 226076
rect -5203 225780 -1502 226052
rect -1230 225780 -1206 226052
rect -5203 225760 -1206 225780
rect -5203 225756 -1526 225760
rect 303926 225357 304246 225358
rect 303926 225039 303927 225357
rect 304245 225039 304246 225357
rect 303926 225038 304246 225039
rect -5974 223800 -3762 224120
rect -2007 223922 -1805 223923
rect -2674 223722 -2006 223922
rect -1806 223722 -1805 223922
rect -2007 223721 -1805 223722
rect -5203 223052 -1206 223076
rect -5203 222780 -1502 223052
rect -1230 222780 -1206 223052
rect -5203 222760 -1206 222780
rect -5203 222756 -1526 222760
rect 303926 222357 304246 222358
rect 303926 222039 303927 222357
rect 304245 222039 304246 222357
rect 303926 222038 304246 222039
rect -5974 220800 -3762 221120
rect -2007 220922 -1805 220923
rect -2674 220722 -2006 220922
rect -1806 220722 -1805 220922
rect -2007 220721 -1805 220722
rect -5203 220052 -1206 220076
rect -5203 219780 -1502 220052
rect -1230 219780 -1206 220052
rect -5203 219760 -1206 219780
rect -5203 219756 -1526 219760
rect 303926 219357 304246 219358
rect 303926 219039 303927 219357
rect 304245 219039 304246 219357
rect 303926 219038 304246 219039
rect -5974 217800 -3762 218120
rect -2007 217922 -1805 217923
rect -2674 217722 -2006 217922
rect -1806 217722 -1805 217922
rect -2007 217721 -1805 217722
rect -5203 217052 -1206 217076
rect -5203 216780 -1502 217052
rect -1230 216780 -1206 217052
rect -5203 216760 -1206 216780
rect -5203 216756 -1526 216760
rect 303926 216357 304246 216358
rect 303926 216039 303927 216357
rect 304245 216039 304246 216357
rect 303926 216038 304246 216039
rect -5974 214800 -3762 215120
rect -2007 214922 -1805 214923
rect -2674 214722 -2006 214922
rect -1806 214722 -1805 214922
rect -2007 214721 -1805 214722
rect -5203 214052 -1206 214076
rect -5203 213780 -1502 214052
rect -1230 213780 -1206 214052
rect -5203 213760 -1206 213780
rect -5203 213756 -1526 213760
rect 303926 213357 304246 213358
rect 303926 213039 303927 213357
rect 304245 213039 304246 213357
rect 303926 213038 304246 213039
rect -5974 211800 -3762 212120
rect -2007 211922 -1805 211923
rect -2674 211722 -2006 211922
rect -1806 211722 -1805 211922
rect -2007 211721 -1805 211722
rect -5203 211052 -1206 211076
rect -5203 210780 -1502 211052
rect -1230 210780 -1206 211052
rect -5203 210760 -1206 210780
rect -5203 210756 -1526 210760
rect 303926 210357 304246 210358
rect 303926 210039 303927 210357
rect 304245 210039 304246 210357
rect 303926 210038 304246 210039
rect -2007 208922 -1805 208923
rect -2674 208722 -2006 208922
rect -1806 208722 -1805 208922
rect -2007 208721 -1805 208722
rect -5203 208052 -1206 208076
rect -5203 207780 -1502 208052
rect -1230 207780 -1206 208052
rect -5203 207760 -1206 207780
rect -5203 207756 -1526 207760
rect 303926 207357 304246 207358
rect 303926 207039 303927 207357
rect 304245 207039 304246 207357
rect 303926 207038 304246 207039
rect -5974 205800 -3762 206120
rect -2007 205922 -1805 205923
rect -2674 205722 -2006 205922
rect -1806 205722 -1805 205922
rect -2007 205721 -1805 205722
rect -5203 205052 -1206 205076
rect -5203 204780 -1502 205052
rect -1230 204780 -1206 205052
rect -5203 204760 -1206 204780
rect -5203 204756 -1526 204760
rect 303926 204357 304246 204358
rect 303926 204039 303927 204357
rect 304245 204039 304246 204357
rect 303926 204038 304246 204039
rect -5974 202800 -3762 203120
rect -2007 202922 -1805 202923
rect -2674 202722 -2006 202922
rect -1806 202722 -1805 202922
rect -2007 202721 -1805 202722
rect -5203 202052 -1206 202076
rect -5203 201780 -1502 202052
rect -1230 201780 -1206 202052
rect -5203 201760 -1206 201780
rect -5203 201756 -1526 201760
rect 303926 201357 304246 201358
rect 303926 201039 303927 201357
rect 304245 201039 304246 201357
rect 303926 201038 304246 201039
rect -5974 199800 -3762 200120
rect -2007 199922 -1805 199923
rect -2674 199722 -2006 199922
rect -1806 199722 -1805 199922
rect -2007 199721 -1805 199722
rect -5203 199052 -1206 199076
rect -5203 198780 -1502 199052
rect -1230 198780 -1206 199052
rect -5203 198760 -1206 198780
rect -5203 198756 -1526 198760
rect 303926 198357 304246 198358
rect 303926 198039 303927 198357
rect 304245 198039 304246 198357
rect 303926 198038 304246 198039
rect -5974 196800 -3762 197120
rect -2007 196922 -1805 196923
rect -2674 196722 -2006 196922
rect -1806 196722 -1805 196922
rect -2007 196721 -1805 196722
rect -5203 196052 -1206 196076
rect -5203 195780 -1502 196052
rect -1230 195780 -1206 196052
rect -5203 195760 -1206 195780
rect -5203 195756 -1526 195760
rect 303926 195357 304246 195358
rect 303926 195039 303927 195357
rect 304245 195039 304246 195357
rect 303926 195038 304246 195039
rect -5974 193800 -3762 194120
rect -2007 193922 -1805 193923
rect -2674 193722 -2006 193922
rect -1806 193722 -1805 193922
rect -2007 193721 -1805 193722
rect -5203 193052 -1206 193076
rect -5203 192780 -1502 193052
rect -1230 192780 -1206 193052
rect -5203 192760 -1206 192780
rect -5203 192756 -1526 192760
rect 303926 192357 304246 192358
rect 303926 192039 303927 192357
rect 304245 192039 304246 192357
rect 303926 192038 304246 192039
rect -5974 190800 -3762 191120
rect -2007 190922 -1805 190923
rect -2674 190722 -2006 190922
rect -1806 190722 -1805 190922
rect -2007 190721 -1805 190722
rect -5203 190052 -1206 190076
rect -5203 189780 -1502 190052
rect -1230 189780 -1206 190052
rect -5203 189760 -1206 189780
rect -5203 189756 -1526 189760
rect 303926 189357 304246 189358
rect 303926 189039 303927 189357
rect 304245 189039 304246 189357
rect 303926 189038 304246 189039
rect -5974 187800 -3762 188120
rect -2007 187922 -1805 187923
rect -2674 187722 -2006 187922
rect -1806 187722 -1805 187922
rect -2007 187721 -1805 187722
rect -5203 187052 -1206 187076
rect -5203 186780 -1502 187052
rect -1230 186780 -1206 187052
rect -5203 186760 -1206 186780
rect -5203 186756 -1526 186760
rect 303926 186357 304246 186358
rect 303926 186039 303927 186357
rect 304245 186039 304246 186357
rect 303926 186038 304246 186039
rect -5974 184800 -3762 185120
rect -2007 184922 -1805 184923
rect -2674 184722 -2006 184922
rect -1806 184722 -1805 184922
rect -2007 184721 -1805 184722
rect -5203 184052 -1206 184076
rect -5203 183780 -1502 184052
rect -1230 183780 -1206 184052
rect -5203 183760 -1206 183780
rect -5203 183756 -1526 183760
rect 303926 183357 304246 183358
rect 303926 183039 303927 183357
rect 304245 183039 304246 183357
rect 303926 183038 304246 183039
rect -5974 181800 -3762 182120
rect -2007 181922 -1805 181923
rect -2674 181722 -2006 181922
rect -1806 181722 -1805 181922
rect -2007 181721 -1805 181722
rect -5203 181052 -1206 181076
rect -5203 180780 -1502 181052
rect -1230 180780 -1206 181052
rect -5203 180760 -1206 180780
rect -5203 180756 -1526 180760
rect 303926 180357 304246 180358
rect 303926 180039 303927 180357
rect 304245 180039 304246 180357
rect 303926 180038 304246 180039
rect -5974 178800 -3762 179120
rect -2007 178922 -1805 178923
rect -2674 178722 -2006 178922
rect -1806 178722 -1805 178922
rect -2007 178721 -1805 178722
rect -5203 178052 -1206 178076
rect -5203 177780 -1502 178052
rect -1230 177780 -1206 178052
rect -5203 177760 -1206 177780
rect -5203 177756 -1526 177760
rect 303926 177357 304246 177358
rect 303926 177039 303927 177357
rect 304245 177039 304246 177357
rect 303926 177038 304246 177039
rect -5974 175800 -3762 176120
rect -2007 175922 -1805 175923
rect -2674 175722 -2006 175922
rect -1806 175722 -1805 175922
rect -2007 175721 -1805 175722
rect -5203 175052 -1206 175076
rect -5203 174780 -1502 175052
rect -1230 174780 -1206 175052
rect -5203 174760 -1206 174780
rect -5203 174756 -1526 174760
rect 303926 174357 304246 174358
rect 303926 174039 303927 174357
rect 304245 174039 304246 174357
rect 303926 174038 304246 174039
rect -5974 172800 -3762 173120
rect -2007 172922 -1805 172923
rect -2674 172722 -2006 172922
rect -1806 172722 -1805 172922
rect -2007 172721 -1805 172722
rect -5203 172052 -1206 172076
rect -5203 171780 -1502 172052
rect -1230 171780 -1206 172052
rect -5203 171760 -1206 171780
rect -5203 171756 -1526 171760
rect 303926 171357 304246 171358
rect 303926 171039 303927 171357
rect 304245 171039 304246 171357
rect 303926 171038 304246 171039
rect -5974 169800 -3762 170120
rect -2007 169922 -1805 169923
rect -2674 169722 -2006 169922
rect -1806 169722 -1805 169922
rect -2007 169721 -1805 169722
rect -5203 169052 -1206 169076
rect -5203 168780 -1502 169052
rect -1230 168780 -1206 169052
rect -5203 168760 -1206 168780
rect -5203 168756 -1526 168760
rect 303926 168357 304246 168358
rect 303926 168039 303927 168357
rect 304245 168039 304246 168357
rect 303926 168038 304246 168039
rect -5974 166800 -3762 167120
rect -2007 166922 -1805 166923
rect -2674 166722 -2006 166922
rect -1806 166722 -1805 166922
rect -2007 166721 -1805 166722
rect -5203 166052 -1206 166076
rect -5203 165780 -1502 166052
rect -1230 165780 -1206 166052
rect -5203 165760 -1206 165780
rect -5203 165756 -1526 165760
rect 303926 165357 304246 165358
rect 303926 165039 303927 165357
rect 304245 165039 304246 165357
rect 303926 165038 304246 165039
rect -5974 163800 -3762 164120
rect -2007 163922 -1805 163923
rect -2674 163722 -2006 163922
rect -1806 163722 -1805 163922
rect -2007 163721 -1805 163722
rect -5203 163052 -1206 163076
rect -5203 162780 -1502 163052
rect -1230 162780 -1206 163052
rect -5203 162760 -1206 162780
rect -5203 162756 -1526 162760
rect 303926 162357 304246 162358
rect 303926 162039 303927 162357
rect 304245 162039 304246 162357
rect 303926 162038 304246 162039
rect -5974 160800 -3762 161120
rect -2007 160922 -1805 160923
rect -2674 160722 -2006 160922
rect -1806 160722 -1805 160922
rect -2007 160721 -1805 160722
rect -5203 160052 -1206 160076
rect -5203 159780 -1502 160052
rect -1230 159780 -1206 160052
rect -5203 159760 -1206 159780
rect -5203 159756 -1526 159760
rect 303926 159357 304246 159358
rect 303926 159039 303927 159357
rect 304245 159039 304246 159357
rect 303926 159038 304246 159039
rect -5974 157800 -3762 158120
rect -2007 157922 -1805 157923
rect -2674 157722 -2006 157922
rect -1806 157722 -1805 157922
rect -2007 157721 -1805 157722
rect -5203 157052 -1206 157076
rect -5203 156780 -1502 157052
rect -1230 156780 -1206 157052
rect -5203 156760 -1206 156780
rect -5203 156756 -1526 156760
rect 303926 156357 304246 156358
rect 303926 156039 303927 156357
rect 304245 156039 304246 156357
rect 303926 156038 304246 156039
rect -5974 154800 -3762 155120
rect -2007 154922 -1805 154923
rect -2674 154722 -2006 154922
rect -1806 154722 -1805 154922
rect -2007 154721 -1805 154722
rect -5203 154052 -1206 154076
rect -5203 153780 -1502 154052
rect -1230 153780 -1206 154052
rect -5203 153760 -1206 153780
rect -5203 153756 -1526 153760
rect 303926 153357 304246 153358
rect 303926 153039 303927 153357
rect 304245 153039 304246 153357
rect 303926 153038 304246 153039
rect -5974 151800 -3762 152120
rect -2007 151922 -1805 151923
rect -2674 151722 -2006 151922
rect -1806 151722 -1805 151922
rect -2007 151721 -1805 151722
rect -5203 151052 -1206 151076
rect -5203 150780 -1502 151052
rect -1230 150780 -1206 151052
rect -5203 150760 -1206 150780
rect -5203 150756 -1526 150760
rect 303926 150357 304246 150358
rect 303926 150039 303927 150357
rect 304245 150039 304246 150357
rect 303926 150038 304246 150039
rect -5974 148800 -3762 149120
rect -2007 148922 -1805 148923
rect -2674 148722 -2006 148922
rect -1806 148722 -1805 148922
rect -2007 148721 -1805 148722
rect -5203 148052 -1206 148076
rect -5203 147780 -1502 148052
rect -1230 147780 -1206 148052
rect -5203 147760 -1206 147780
rect -5203 147756 -1526 147760
rect 303926 147357 304246 147358
rect 303926 147039 303927 147357
rect 304245 147039 304246 147357
rect 303926 147038 304246 147039
rect -5974 145800 -3762 146120
rect -2007 145922 -1805 145923
rect -2674 145722 -2006 145922
rect -1806 145722 -1805 145922
rect -2007 145721 -1805 145722
rect -5203 145052 -1206 145076
rect -5203 144780 -1502 145052
rect -1230 144780 -1206 145052
rect -5203 144760 -1206 144780
rect -5203 144756 -1526 144760
rect 303926 144357 304246 144358
rect 303926 144039 303927 144357
rect 304245 144039 304246 144357
rect 303926 144038 304246 144039
rect -5974 142800 -3762 143120
rect -2007 142922 -1805 142923
rect -2674 142722 -2006 142922
rect -1806 142722 -1805 142922
rect -2007 142721 -1805 142722
rect -5203 142052 -1206 142076
rect -5203 141780 -1502 142052
rect -1230 141780 -1206 142052
rect -5203 141760 -1206 141780
rect -5203 141756 -1526 141760
rect 303926 141357 304246 141358
rect 303926 141039 303927 141357
rect 304245 141039 304246 141357
rect 303926 141038 304246 141039
rect -5974 139800 -3762 140120
rect -2007 139922 -1805 139923
rect -2674 139722 -2006 139922
rect -1806 139722 -1805 139922
rect -2007 139721 -1805 139722
rect -5203 139052 -1206 139076
rect -5203 138780 -1502 139052
rect -1230 138780 -1206 139052
rect -5203 138760 -1206 138780
rect -5203 138756 -1526 138760
rect 303926 138357 304246 138358
rect 303926 138039 303927 138357
rect 304245 138039 304246 138357
rect 303926 138038 304246 138039
rect -5974 136800 -3762 137120
rect -2007 136922 -1805 136923
rect -2674 136722 -2006 136922
rect -1806 136722 -1805 136922
rect -2007 136721 -1805 136722
rect -5203 136052 -1206 136076
rect -5203 135780 -1502 136052
rect -1230 135780 -1206 136052
rect -5203 135760 -1206 135780
rect -5203 135756 -1526 135760
rect 303926 135357 304246 135358
rect 303926 135039 303927 135357
rect 304245 135039 304246 135357
rect 303926 135038 304246 135039
rect -5974 133800 -3762 134120
rect -2007 133922 -1805 133923
rect -2674 133722 -2006 133922
rect -1806 133722 -1805 133922
rect -2007 133721 -1805 133722
rect -5203 133052 -1206 133076
rect -5203 132780 -1502 133052
rect -1230 132780 -1206 133052
rect -5203 132760 -1206 132780
rect -5203 132756 -1526 132760
rect 303926 132357 304246 132358
rect 303926 132039 303927 132357
rect 304245 132039 304246 132357
rect 303926 132038 304246 132039
rect -5974 130800 -3762 131120
rect -2007 130922 -1805 130923
rect -2674 130722 -2006 130922
rect -1806 130722 -1805 130922
rect -2007 130721 -1805 130722
rect -5203 130052 -1206 130076
rect -5203 129780 -1502 130052
rect -1230 129780 -1206 130052
rect -5203 129760 -1206 129780
rect -5203 129756 -1526 129760
rect 303926 129357 304246 129358
rect 303926 129039 303927 129357
rect 304245 129039 304246 129357
rect 303926 129038 304246 129039
rect -5974 127800 -3762 128120
rect -2007 127922 -1805 127923
rect -2674 127722 -2006 127922
rect -1806 127722 -1805 127922
rect -2007 127721 -1805 127722
rect -5203 127052 -1206 127076
rect -5203 126780 -1502 127052
rect -1230 126780 -1206 127052
rect -5203 126760 -1206 126780
rect -5203 126756 -1526 126760
rect 303926 126357 304246 126358
rect 303926 126039 303927 126357
rect 304245 126039 304246 126357
rect 303926 126038 304246 126039
rect -5974 124800 -3762 125120
rect -2007 124922 -1805 124923
rect -2674 124722 -2006 124922
rect -1806 124722 -1805 124922
rect -2007 124721 -1805 124722
rect -5203 124052 -1206 124076
rect -5203 123780 -1502 124052
rect -1230 123780 -1206 124052
rect -5203 123760 -1206 123780
rect -5203 123756 -1526 123760
rect 303926 123357 304246 123358
rect 303926 123039 303927 123357
rect 304245 123039 304246 123357
rect 303926 123038 304246 123039
rect -5974 121800 -3762 122120
rect -2007 121922 -1805 121923
rect -2674 121722 -2006 121922
rect -1806 121722 -1805 121922
rect -2007 121721 -1805 121722
rect -5203 121052 -1206 121076
rect -5203 120780 -1502 121052
rect -1230 120780 -1206 121052
rect -5203 120760 -1206 120780
rect -5203 120756 -1526 120760
rect 303926 120357 304246 120358
rect 303926 120039 303927 120357
rect 304245 120039 304246 120357
rect 303926 120038 304246 120039
rect -5974 118800 -3762 119120
rect -2007 118922 -1805 118923
rect -2674 118722 -2006 118922
rect -1806 118722 -1805 118922
rect -2007 118721 -1805 118722
rect -5203 118052 -1206 118076
rect -5203 117780 -1502 118052
rect -1230 117780 -1206 118052
rect -5203 117760 -1206 117780
rect -5203 117756 -1526 117760
rect 303926 117357 304246 117358
rect 303926 117039 303927 117357
rect 304245 117039 304246 117357
rect 303926 117038 304246 117039
rect -5974 115800 -3762 116120
rect -2007 115922 -1805 115923
rect -2674 115722 -2006 115922
rect -1806 115722 -1805 115922
rect -2007 115721 -1805 115722
rect -5203 115052 -1206 115076
rect -5203 114780 -1502 115052
rect -1230 114780 -1206 115052
rect -5203 114760 -1206 114780
rect -5203 114756 -1526 114760
rect 303926 114357 304246 114358
rect 303926 114039 303927 114357
rect 304245 114039 304246 114357
rect 303926 114038 304246 114039
rect -5974 112800 -3762 113120
rect -2007 112922 -1805 112923
rect -2674 112722 -2006 112922
rect -1806 112722 -1805 112922
rect -2007 112721 -1805 112722
rect -5203 112052 -1206 112076
rect -5203 111780 -1502 112052
rect -1230 111780 -1206 112052
rect -5203 111760 -1206 111780
rect -5203 111756 -1526 111760
rect 303926 111357 304246 111358
rect 303926 111039 303927 111357
rect 304245 111039 304246 111357
rect 303926 111038 304246 111039
rect -5974 109800 -3762 110120
rect -2007 109922 -1805 109923
rect -2674 109722 -2006 109922
rect -1806 109722 -1805 109922
rect -2007 109721 -1805 109722
rect -5203 109052 -1206 109076
rect -5203 108780 -1502 109052
rect -1230 108780 -1206 109052
rect -5203 108760 -1206 108780
rect -5203 108756 -1526 108760
rect 303926 108357 304246 108358
rect 303926 108039 303927 108357
rect 304245 108039 304246 108357
rect 303926 108038 304246 108039
rect -5974 106800 -3762 107120
rect -2007 106922 -1805 106923
rect -2674 106722 -2006 106922
rect -1806 106722 -1805 106922
rect -2007 106721 -1805 106722
rect -5203 106052 -1206 106076
rect -5203 105780 -1502 106052
rect -1230 105780 -1206 106052
rect -5203 105760 -1206 105780
rect -5203 105756 -1526 105760
rect 303926 105357 304246 105358
rect 303926 105039 303927 105357
rect 304245 105039 304246 105357
rect 303926 105038 304246 105039
rect -5974 103800 -3762 104120
rect -2007 103922 -1805 103923
rect -2674 103722 -2006 103922
rect -1806 103722 -1805 103922
rect -2007 103721 -1805 103722
rect -5203 103052 -1206 103076
rect -5203 102780 -1502 103052
rect -1230 102780 -1206 103052
rect -5203 102760 -1206 102780
rect -5203 102756 -1526 102760
rect 303926 102357 304246 102358
rect 303926 102039 303927 102357
rect 304245 102039 304246 102357
rect 303926 102038 304246 102039
rect -5974 100800 -3762 101120
rect -2007 100922 -1805 100923
rect -2674 100722 -2006 100922
rect -1806 100722 -1805 100922
rect -2007 100721 -1805 100722
rect -5203 100052 -1206 100076
rect -5203 99780 -1502 100052
rect -1230 99780 -1206 100052
rect -5203 99760 -1206 99780
rect -5203 99756 -1526 99760
rect 303926 99357 304246 99358
rect 303926 99039 303927 99357
rect 304245 99039 304246 99357
rect 303926 99038 304246 99039
rect -5974 97800 -3762 98120
rect -2007 97922 -1805 97923
rect -2674 97722 -2006 97922
rect -1806 97722 -1805 97922
rect -2007 97721 -1805 97722
rect -5203 97052 -1206 97076
rect -5203 96780 -1502 97052
rect -1230 96780 -1206 97052
rect -5203 96760 -1206 96780
rect -5203 96756 -1526 96760
rect 303926 96357 304246 96358
rect 303926 96039 303927 96357
rect 304245 96039 304246 96357
rect 303926 96038 304246 96039
rect -5974 94800 -3762 95120
rect -2007 94922 -1805 94923
rect -2674 94722 -2006 94922
rect -1806 94722 -1805 94922
rect -2007 94721 -1805 94722
rect 303926 93357 304246 93358
rect 303926 93039 303927 93357
rect 304245 93039 304246 93357
rect 303926 93038 304246 93039
rect -5974 91800 -3762 92120
rect -2007 91922 -1805 91923
rect -2674 91722 -2006 91922
rect -1806 91722 -1805 91922
rect -2007 91721 -1805 91722
rect -5203 91052 -1206 91076
rect -5203 90780 -1502 91052
rect -1230 90780 -1206 91052
rect -5203 90760 -1206 90780
rect -5203 90756 -1526 90760
rect 303926 90357 304246 90358
rect 303926 90039 303927 90357
rect 304245 90039 304246 90357
rect 303926 90038 304246 90039
rect -5974 88800 -3762 89120
rect -2007 88922 -1805 88923
rect -2674 88722 -2006 88922
rect -1806 88722 -1805 88922
rect -2007 88721 -1805 88722
rect -5203 88052 -1206 88076
rect -5203 87780 -1502 88052
rect -1230 87780 -1206 88052
rect -5203 87760 -1206 87780
rect -5203 87756 -1526 87760
rect 303926 87357 304246 87358
rect 303926 87039 303927 87357
rect 304245 87039 304246 87357
rect 303926 87038 304246 87039
rect -5974 85800 -3762 86120
rect -2007 85922 -1805 85923
rect -2674 85722 -2006 85922
rect -1806 85722 -1805 85922
rect -2007 85721 -1805 85722
rect -5203 85052 -1206 85076
rect -5203 84780 -1502 85052
rect -1230 84780 -1206 85052
rect -5203 84760 -1206 84780
rect -5203 84756 -1526 84760
rect 303926 84357 304246 84358
rect 303926 84039 303927 84357
rect 304245 84039 304246 84357
rect 303926 84038 304246 84039
rect -5974 82800 -3762 83120
rect -2007 82922 -1805 82923
rect -2674 82722 -2006 82922
rect -1806 82722 -1805 82922
rect -2007 82721 -1805 82722
rect -5203 82052 -1206 82076
rect -5203 81780 -1502 82052
rect -1230 81780 -1206 82052
rect -5203 81760 -1206 81780
rect -5203 81756 -1526 81760
rect 303926 81357 304246 81358
rect 303926 81039 303927 81357
rect 304245 81039 304246 81357
rect 303926 81038 304246 81039
rect -5974 79800 -3762 80120
rect -2007 79922 -1805 79923
rect -2674 79722 -2006 79922
rect -1806 79722 -1805 79922
rect -2007 79721 -1805 79722
rect -5203 79052 -1206 79076
rect -5203 78780 -1502 79052
rect -1230 78780 -1206 79052
rect -5203 78760 -1206 78780
rect -5203 78756 -1526 78760
rect 303926 78357 304246 78358
rect 303926 78039 303927 78357
rect 304245 78039 304246 78357
rect 303926 78038 304246 78039
rect -5974 76800 -3762 77120
rect -2007 76922 -1805 76923
rect -2674 76722 -2006 76922
rect -1806 76722 -1805 76922
rect -2007 76721 -1805 76722
rect -5203 76052 -1206 76076
rect -5203 75780 -1502 76052
rect -1230 75780 -1206 76052
rect -5203 75760 -1206 75780
rect -5203 75756 -1526 75760
rect 303926 75357 304246 75358
rect 303926 75039 303927 75357
rect 304245 75039 304246 75357
rect 303926 75038 304246 75039
rect -5974 73800 -3762 74120
rect -2007 73922 -1805 73923
rect -2674 73722 -2006 73922
rect -1806 73722 -1805 73922
rect -2007 73721 -1805 73722
rect -5203 73052 -1206 73076
rect -5203 72780 -1502 73052
rect -1230 72780 -1206 73052
rect -5203 72760 -1206 72780
rect -5203 72756 -1526 72760
rect 303926 72357 304246 72358
rect 303926 72039 303927 72357
rect 304245 72039 304246 72357
rect 303926 72038 304246 72039
rect -5974 70800 -3762 71120
rect -2007 70922 -1805 70923
rect -2674 70722 -2006 70922
rect -1806 70722 -1805 70922
rect -2007 70721 -1805 70722
rect -5203 70052 -1206 70076
rect -5203 69780 -1502 70052
rect -1230 69780 -1206 70052
rect -5203 69760 -1206 69780
rect -5203 69756 -1526 69760
rect 303926 69357 304246 69358
rect 303926 69039 303927 69357
rect 304245 69039 304246 69357
rect 303926 69038 304246 69039
rect -5974 67800 -3762 68120
rect -2007 67922 -1805 67923
rect -2674 67722 -2006 67922
rect -1806 67722 -1805 67922
rect -2007 67721 -1805 67722
rect -5203 67052 -1206 67076
rect -5203 66780 -1502 67052
rect -1230 66780 -1206 67052
rect -5203 66760 -1206 66780
rect -5203 66756 -1526 66760
rect 303926 66357 304246 66358
rect 303926 66039 303927 66357
rect 304245 66039 304246 66357
rect 303926 66038 304246 66039
rect -5974 64800 -3762 65120
rect -2007 64922 -1805 64923
rect -2674 64722 -2006 64922
rect -1806 64722 -1805 64922
rect -2007 64721 -1805 64722
rect -5203 64052 -1206 64076
rect -5203 63780 -1502 64052
rect -1230 63780 -1206 64052
rect -5203 63760 -1206 63780
rect -5203 63756 -1526 63760
rect 303926 63357 304246 63358
rect 303926 63039 303927 63357
rect 304245 63039 304246 63357
rect 303926 63038 304246 63039
rect -5974 61800 -3762 62120
rect -2007 61922 -1805 61923
rect -2674 61722 -2006 61922
rect -1806 61722 -1805 61922
rect -2007 61721 -1805 61722
rect -5203 61052 -1206 61076
rect -5203 60780 -1502 61052
rect -1230 60780 -1206 61052
rect -5203 60760 -1206 60780
rect -5203 60756 -1526 60760
rect 303926 60357 304246 60358
rect 303926 60039 303927 60357
rect 304245 60039 304246 60357
rect 303926 60038 304246 60039
rect -5974 58800 -3762 59120
rect -2007 58922 -1805 58923
rect -2674 58722 -2006 58922
rect -1806 58722 -1805 58922
rect -2007 58721 -1805 58722
rect -5203 58052 -1206 58076
rect -5203 57780 -1502 58052
rect -1230 57780 -1206 58052
rect -5203 57760 -1206 57780
rect -5203 57756 -1526 57760
rect 303926 57357 304246 57358
rect 303926 57039 303927 57357
rect 304245 57039 304246 57357
rect 303926 57038 304246 57039
rect -2007 55922 -1805 55923
rect -2674 55722 -2006 55922
rect -1806 55722 -1805 55922
rect -2007 55721 -1805 55722
rect -5203 55052 -1206 55076
rect -5203 54780 -1502 55052
rect -1230 54780 -1206 55052
rect -5203 54760 -1206 54780
rect -5203 54756 -1526 54760
rect 303926 54357 304246 54358
rect 303926 54039 303927 54357
rect 304245 54039 304246 54357
rect 303926 54038 304246 54039
rect -5974 52800 -3762 53120
rect -2007 52922 -1805 52923
rect -2674 52722 -2006 52922
rect -1806 52722 -1805 52922
rect -2007 52721 -1805 52722
rect -5203 52052 -1206 52076
rect -5203 51780 -1502 52052
rect -1230 51780 -1206 52052
rect -5203 51760 -1206 51780
rect -5203 51756 -1526 51760
rect 303926 51357 304246 51358
rect 303926 51039 303927 51357
rect 304245 51039 304246 51357
rect 303926 51038 304246 51039
rect -5974 49800 -3762 50120
rect -2007 49922 -1805 49923
rect -2674 49722 -2006 49922
rect -1806 49722 -1805 49922
rect -2007 49721 -1805 49722
rect -5203 49052 -1206 49076
rect -5203 48780 -1502 49052
rect -1230 48780 -1206 49052
rect -5203 48760 -1206 48780
rect -5203 48756 -1526 48760
rect 303926 48357 304246 48358
rect 303926 48039 303927 48357
rect 304245 48039 304246 48357
rect 303926 48038 304246 48039
rect -5974 46800 -3762 47120
rect -2007 46922 -1805 46923
rect -2674 46722 -2006 46922
rect -1806 46722 -1805 46922
rect -2007 46721 -1805 46722
rect -5203 46052 -1206 46076
rect -5203 45780 -1502 46052
rect -1230 45780 -1206 46052
rect -5203 45760 -1206 45780
rect -5203 45756 -1526 45760
rect 303926 45357 304246 45358
rect 303926 45039 303927 45357
rect 304245 45039 304246 45357
rect 303926 45038 304246 45039
rect -5974 43800 -3762 44120
rect -2007 43922 -1805 43923
rect -2674 43722 -2006 43922
rect -1806 43722 -1805 43922
rect -2007 43721 -1805 43722
rect -5203 43052 -1206 43076
rect -5203 42780 -1502 43052
rect -1230 42780 -1206 43052
rect -5203 42760 -1206 42780
rect -5203 42756 -1526 42760
rect 303926 42357 304246 42358
rect 303926 42039 303927 42357
rect 304245 42039 304246 42357
rect 303926 42038 304246 42039
rect -5974 40800 -3762 41120
rect -2007 40922 -1805 40923
rect -2674 40722 -2006 40922
rect -1806 40722 -1805 40922
rect -2007 40721 -1805 40722
rect -5203 40052 -1206 40076
rect -5203 39780 -1502 40052
rect -1230 39780 -1206 40052
rect -5203 39760 -1206 39780
rect -5203 39756 -1526 39760
rect 303926 39357 304246 39358
rect 303926 39039 303927 39357
rect 304245 39039 304246 39357
rect 303926 39038 304246 39039
rect -5974 37800 -3762 38120
rect -2007 37922 -1805 37923
rect -2674 37722 -2006 37922
rect -1806 37722 -1805 37922
rect -2007 37721 -1805 37722
rect -5203 37052 -1206 37076
rect -5203 36780 -1502 37052
rect -1230 36780 -1206 37052
rect -5203 36760 -1206 36780
rect -5203 36756 -1526 36760
rect 303926 36357 304246 36358
rect 303926 36039 303927 36357
rect 304245 36039 304246 36357
rect 303926 36038 304246 36039
rect -5974 34800 -3762 35120
rect -2007 34922 -1805 34923
rect -2674 34722 -2006 34922
rect -1806 34722 -1805 34922
rect -2007 34721 -1805 34722
rect -5203 34052 -1206 34076
rect -5203 33780 -1502 34052
rect -1230 33780 -1206 34052
rect -5203 33760 -1206 33780
rect -5203 33756 -1526 33760
rect 303926 33357 304246 33358
rect 303926 33039 303927 33357
rect 304245 33039 304246 33357
rect 303926 33038 304246 33039
rect -5974 31800 -3762 32120
rect -2007 31922 -1805 31923
rect -2674 31722 -2006 31922
rect -1806 31722 -1805 31922
rect -2007 31721 -1805 31722
rect -5203 31052 -1206 31076
rect -5203 30780 -1502 31052
rect -1230 30780 -1206 31052
rect -5203 30760 -1206 30780
rect -5203 30756 -1526 30760
rect 303926 30357 304246 30358
rect 303926 30039 303927 30357
rect 304245 30039 304246 30357
rect 303926 30038 304246 30039
rect -5974 28800 -3762 29120
rect -2007 28922 -1805 28923
rect -2674 28722 -2006 28922
rect -1806 28722 -1805 28922
rect -2007 28721 -1805 28722
rect -5203 28052 -1206 28076
rect -5203 27780 -1502 28052
rect -1230 27780 -1206 28052
rect -5203 27760 -1206 27780
rect -5203 27756 -1526 27760
rect 303926 27357 304246 27358
rect 303926 27039 303927 27357
rect 304245 27039 304246 27357
rect 303926 27038 304246 27039
rect -5974 25800 -3762 26120
rect -2007 25922 -1805 25923
rect -2674 25722 -2006 25922
rect -1806 25722 -1805 25922
rect -2007 25721 -1805 25722
rect -5203 25052 -1206 25076
rect -5203 24780 -1502 25052
rect -1230 24780 -1206 25052
rect -5203 24760 -1206 24780
rect -5203 24756 -1526 24760
rect 303926 24357 304246 24358
rect 303926 24039 303927 24357
rect 304245 24039 304246 24357
rect 303926 24038 304246 24039
rect -5974 22800 -3762 23120
rect -2007 22922 -1805 22923
rect -2674 22722 -2006 22922
rect -1806 22722 -1805 22922
rect -2007 22721 -1805 22722
rect -5203 22052 -1206 22076
rect -5203 21780 -1502 22052
rect -1230 21780 -1206 22052
rect -5203 21760 -1206 21780
rect -5203 21756 -1526 21760
rect 303926 21357 304246 21358
rect 303926 21039 303927 21357
rect 304245 21039 304246 21357
rect 303926 21038 304246 21039
rect -5974 19800 -3762 20120
rect -5203 19052 -1206 19076
rect -5203 18780 -1502 19052
rect -1230 18780 -1206 19052
rect -5203 18760 -1206 18780
rect -781 18795 1738 18905
rect -5203 18756 -1526 18760
rect -6095 17942 -5993 17943
rect -5994 17742 -5993 17942
rect -6095 17741 -5993 17742
rect -781 16797 -671 18795
rect 2328 18467 2548 19498
rect 5328 18810 5548 19607
rect 7470 18892 7720 18911
rect 8328 18892 8548 19654
rect 7470 18891 8548 18892
rect 5317 18784 5567 18810
rect 3664 18759 3984 18760
rect 2316 18439 2566 18467
rect 3664 18441 3665 18759
rect 3983 18441 3984 18759
rect 5317 18566 5329 18784
rect 5547 18566 5567 18784
rect 7470 18673 7483 18891
rect 7701 18673 8548 18891
rect 7470 18672 8548 18673
rect 10692 18836 10942 18858
rect 11328 18836 11548 19678
rect 10692 18835 11548 18836
rect 7470 18653 7720 18672
rect 10692 18617 10712 18835
rect 10930 18617 11548 18835
rect 13790 18930 14040 18950
rect 14328 18930 14548 19678
rect 13790 18929 14548 18930
rect 13790 18711 13802 18929
rect 14020 18711 14548 18929
rect 13790 18710 14548 18711
rect 16900 18817 17150 18825
rect 17328 18817 17548 19673
rect 19851 19194 20101 19202
rect 20328 19194 20548 19678
rect 19851 19193 20548 19194
rect 19851 18975 19870 19193
rect 20088 18975 20548 19193
rect 19851 18974 20548 18975
rect 19851 18944 20101 18974
rect 16900 18816 17548 18817
rect 13790 18692 14040 18710
rect 10692 18616 11548 18617
rect 10692 18600 10942 18616
rect 16900 18598 16912 18816
rect 17130 18598 17548 18816
rect 16900 18597 17548 18598
rect 18088 18759 18408 18760
rect 16900 18567 17150 18597
rect 5317 18552 5567 18566
rect 3664 18440 3984 18441
rect 18088 18441 18089 18759
rect 18407 18441 18408 18759
rect 18088 18440 18408 18441
rect 22872 18659 23189 18673
rect 23328 18659 23548 19678
rect 25909 19012 26226 19029
rect 26328 19012 26548 19678
rect 29328 19062 29548 19678
rect 25909 19011 26548 19012
rect 25909 18793 25944 19011
rect 26162 18793 26548 19011
rect 29084 19061 29548 19062
rect 29084 18843 29085 19061
rect 29303 18843 29548 19061
rect 29084 18842 29548 18843
rect 32328 18986 32548 19678
rect 35328 19066 35548 19597
rect 38328 19226 38548 19635
rect 38313 19218 38563 19226
rect 25909 18792 26548 18793
rect 25909 18763 26226 18792
rect 32328 18768 32329 18986
rect 32547 18768 32548 18986
rect 35298 19055 35585 19066
rect 35298 18837 35329 19055
rect 35547 18837 35585 19055
rect 38313 19000 38329 19218
rect 38547 19000 38563 19218
rect 38313 18968 38563 19000
rect 41328 18892 41548 19678
rect 44328 18936 44548 19673
rect 47328 19145 47548 19678
rect 47318 19130 47568 19145
rect 44320 18923 44570 18936
rect 35298 18828 35585 18837
rect 41318 18872 41568 18892
rect 32328 18767 32548 18768
rect 22872 18658 23548 18659
rect 22872 18440 22898 18658
rect 23116 18440 23548 18658
rect 32914 18759 33234 18760
rect 35328 18759 35548 18828
rect 32914 18441 32915 18759
rect 33233 18441 33234 18759
rect 41318 18654 41329 18872
rect 41547 18654 41568 18872
rect 44320 18705 44329 18923
rect 44547 18705 44570 18923
rect 47318 18912 47329 19130
rect 47547 18912 47568 19130
rect 47318 18887 47568 18912
rect 50328 19023 50548 19654
rect 53328 19065 53548 19678
rect 56328 19163 56548 19666
rect 56328 19162 56835 19163
rect 53328 19042 53770 19065
rect 50328 19011 50750 19023
rect 50328 18793 50517 19011
rect 50735 18793 50750 19011
rect 53328 18824 53538 19042
rect 53756 18824 53770 19042
rect 56328 18944 56616 19162
rect 56834 18944 56835 19162
rect 56328 18943 56835 18944
rect 53328 18823 53770 18824
rect 53520 18807 53770 18823
rect 59328 18867 59548 19678
rect 59328 18866 59850 18867
rect 50328 18792 50750 18793
rect 50500 18765 50750 18792
rect 44320 18678 44570 18705
rect 41318 18634 41568 18654
rect 59328 18648 59631 18866
rect 59849 18648 59850 18866
rect 59328 18647 59850 18648
rect 62328 18791 62548 19678
rect 65328 18882 65548 19645
rect 68328 18952 68548 19638
rect 65328 18881 65962 18882
rect 62328 18790 62852 18791
rect 62328 18572 62633 18790
rect 62851 18572 62852 18790
rect 62328 18571 62852 18572
rect 64256 18759 64576 18760
rect 32914 18440 33234 18441
rect 64256 18441 64257 18759
rect 64575 18441 64576 18759
rect 65328 18663 65743 18881
rect 65961 18663 65962 18881
rect 68328 18734 68329 18952
rect 68547 18734 68548 18952
rect 71328 19061 71548 19631
rect 71328 19060 72148 19061
rect 71328 18842 71929 19060
rect 72147 18842 72148 19060
rect 71328 18841 72148 18842
rect 74328 19031 74548 19676
rect 74328 19030 75298 19031
rect 74328 18812 75079 19030
rect 75297 18812 75298 19030
rect 74328 18811 75298 18812
rect 68328 18733 68548 18734
rect 65328 18662 65962 18663
rect 64256 18440 64576 18441
rect 2316 18221 2329 18439
rect 2547 18221 2566 18439
rect 22872 18439 23548 18440
rect 22872 18407 23189 18439
rect 2316 18209 2566 18221
rect 77328 18307 77548 19678
rect 80328 18906 80548 19677
rect 80328 18905 81410 18906
rect 80328 18687 81191 18905
rect 81409 18687 81410 18905
rect 80328 18686 81410 18687
rect 83328 18404 83548 19662
rect 83328 18403 84494 18404
rect 77328 18306 78318 18307
rect 77328 18088 78099 18306
rect 78317 18088 78318 18306
rect 83328 18185 84275 18403
rect 84493 18185 84494 18403
rect 83328 18184 84494 18185
rect 86328 18315 86548 19678
rect 89328 18838 89548 19632
rect 89328 18837 90632 18838
rect 89328 18619 90413 18837
rect 90631 18619 90632 18837
rect 89328 18618 90632 18619
rect 92328 18794 92548 19624
rect 95328 18876 95548 19632
rect 95328 18875 96673 18876
rect 92328 18793 93776 18794
rect 92328 18575 93557 18793
rect 93775 18575 93776 18793
rect 95328 18657 96454 18875
rect 96672 18657 96673 18875
rect 95328 18656 96673 18657
rect 92328 18574 93776 18575
rect 98328 18502 98548 19639
rect 101328 18741 101548 19610
rect 104328 18756 104548 19632
rect 107328 19033 107548 19624
rect 107328 19032 109121 19033
rect 107328 18814 108902 19032
rect 109120 18814 109121 19032
rect 107328 18813 109121 18814
rect 110328 18936 110548 19647
rect 113328 18985 113548 19658
rect 113328 18984 115173 18985
rect 110328 18935 112168 18936
rect 104328 18755 105895 18756
rect 101328 18740 102931 18741
rect 101328 18522 102712 18740
rect 102930 18522 102931 18740
rect 104328 18537 105676 18755
rect 105894 18537 105895 18755
rect 110328 18717 111949 18935
rect 112167 18717 112168 18935
rect 113328 18766 114954 18984
rect 115172 18766 115173 18984
rect 113328 18765 115173 18766
rect 116328 18978 116548 19613
rect 116328 18977 118188 18978
rect 116328 18759 117969 18977
rect 118187 18759 118188 18977
rect 116328 18758 118188 18759
rect 119328 18865 119548 19678
rect 119328 18864 121370 18865
rect 110328 18716 112168 18717
rect 119328 18646 121151 18864
rect 121369 18646 121370 18864
rect 122328 18852 122548 19659
rect 125328 18943 125548 19678
rect 125328 18942 127461 18943
rect 122328 18851 124338 18852
rect 119328 18645 121370 18646
rect 121678 18759 121998 18760
rect 104328 18536 105895 18537
rect 101328 18521 102931 18522
rect 98328 18501 99817 18502
rect 86328 18314 87555 18315
rect 86328 18096 87336 18314
rect 87554 18096 87555 18314
rect 98328 18283 99598 18501
rect 99816 18283 99817 18501
rect 121678 18441 121679 18759
rect 121997 18441 121998 18759
rect 122328 18633 124119 18851
rect 124337 18633 124338 18851
rect 125328 18724 127242 18942
rect 127460 18724 127461 18942
rect 125328 18723 127461 18724
rect 128328 18814 128548 19644
rect 131328 18867 131548 19675
rect 131328 18866 133632 18867
rect 128328 18813 130470 18814
rect 122328 18632 124338 18633
rect 128328 18595 130251 18813
rect 130469 18595 130470 18813
rect 131328 18648 133413 18866
rect 133631 18648 133632 18866
rect 131328 18647 133632 18648
rect 128328 18594 130470 18595
rect 121678 18440 121998 18441
rect 98328 18282 99817 18283
rect 86328 18095 87555 18096
rect 134328 18242 134548 19659
rect 137328 18601 137548 19614
rect 140328 18669 140548 19678
rect 143328 18844 143548 19675
rect 146328 18844 146548 19667
rect 143328 18843 145798 18844
rect 140328 18668 142819 18669
rect 137328 18600 139772 18601
rect 137328 18382 139553 18600
rect 139771 18382 139772 18600
rect 140328 18450 142600 18668
rect 142818 18450 142819 18668
rect 143328 18625 145579 18843
rect 145797 18625 145798 18843
rect 143328 18624 145798 18625
rect 146328 18843 148974 18844
rect 146328 18625 148755 18843
rect 148973 18625 148974 18843
rect 146328 18624 148974 18625
rect 149328 18775 149548 19658
rect 152328 18859 152548 19658
rect 155328 18998 155548 19658
rect 155328 18997 158063 18998
rect 152328 18858 155012 18859
rect 149328 18774 151992 18775
rect 149328 18556 151773 18774
rect 151991 18556 151992 18774
rect 152328 18640 154793 18858
rect 155011 18640 155012 18858
rect 155328 18779 157844 18997
rect 158062 18779 158063 18997
rect 155328 18778 158063 18779
rect 152328 18639 155012 18640
rect 158328 18759 158548 19678
rect 161328 18890 161548 19666
rect 164328 19028 164548 19666
rect 167328 19136 167548 19658
rect 158328 18758 161153 18759
rect 149328 18555 151992 18556
rect 158328 18540 160887 18758
rect 161105 18540 161153 18758
rect 161328 18670 163556 18890
rect 164328 18808 166148 19028
rect 167328 18916 169083 19136
rect 158328 18539 161153 18540
rect 140328 18449 142819 18450
rect 163238 18459 163458 18670
rect 137328 18381 139772 18382
rect 134328 18241 136687 18242
rect 77328 18087 78318 18088
rect 134328 18023 136468 18241
rect 136686 18023 136687 18241
rect 163238 18241 163239 18459
rect 163457 18241 163458 18459
rect 163238 18240 163458 18241
rect 134328 18022 136687 18023
rect 165928 18174 166148 18808
rect 167548 18759 167868 18760
rect 167548 18441 167549 18759
rect 167867 18441 167868 18759
rect 167548 18440 167868 18441
rect 165928 17956 165929 18174
rect 166147 17956 166148 18174
rect 165928 17955 166148 17956
rect 168863 17421 169083 18916
rect 170328 18490 170548 19643
rect 173328 19136 173548 19678
rect 173328 19135 174586 19136
rect 173328 18917 174367 19135
rect 174585 18917 174586 19135
rect 173328 18916 174586 18917
rect 176328 18812 176548 19628
rect 176328 18594 176329 18812
rect 176547 18594 176548 18812
rect 176328 18593 176548 18594
rect 170328 18489 173302 18490
rect 170328 18271 173083 18489
rect 173301 18271 173302 18489
rect 170328 18270 173302 18271
rect 179328 17860 179548 19678
rect 182328 18782 182548 19658
rect 180548 18759 180868 18760
rect 180548 18441 180549 18759
rect 180867 18441 180868 18759
rect 182328 18562 184230 18782
rect 180548 18440 180868 18441
rect 179328 17859 182693 17860
rect 179328 17641 182474 17859
rect 182692 17641 182693 17859
rect 179328 17640 182693 17641
rect 168863 17203 168864 17421
rect 169082 17203 169083 17421
rect 168863 17202 169083 17203
rect 184010 17152 184230 18562
rect 185328 18036 185548 19678
rect 185328 17818 185329 18036
rect 185547 17818 185548 18036
rect 185328 17817 185548 17818
rect 188328 17659 188548 19658
rect 189548 18759 189868 18760
rect 189548 18441 189549 18759
rect 189867 18441 189868 18759
rect 189548 18440 189868 18441
rect 191328 18626 191548 19634
rect 191328 18406 193685 18626
rect 188328 17441 188329 17659
rect 188547 17441 188548 17659
rect 188328 17440 188548 17441
rect 184010 16934 184011 17152
rect 184229 16934 184230 17152
rect 184010 16933 184230 16934
rect 193465 17019 193685 18406
rect 194328 17930 194548 19625
rect 197328 17957 197548 19661
rect 200328 18804 200548 19625
rect 198548 18759 198868 18760
rect 198548 18441 198549 18759
rect 198867 18441 198868 18759
rect 200328 18584 202223 18804
rect 198548 18440 198868 18441
rect 197328 17956 201135 17957
rect 194328 17929 197013 17930
rect 194328 17711 196794 17929
rect 197012 17711 197013 17929
rect 197328 17738 200916 17956
rect 201134 17738 201135 17956
rect 197328 17737 201135 17738
rect 194328 17710 197013 17711
rect 193465 16801 193466 17019
rect 193684 16801 193685 17019
rect 193465 16800 193685 16801
rect 202003 16894 202223 18584
rect 203328 17752 203548 19670
rect 204548 18759 204868 18760
rect 204548 18441 204549 18759
rect 204867 18441 204868 18759
rect 204548 18440 204868 18441
rect 206328 18455 206548 19678
rect 206328 18237 206329 18455
rect 206547 18237 206548 18455
rect 206328 18236 206548 18237
rect 209328 18099 209548 19652
rect 212328 18885 212548 19634
rect 211548 18759 211868 18760
rect 211548 18441 211549 18759
rect 211867 18441 211868 18759
rect 212328 18665 214124 18885
rect 211548 18440 211868 18441
rect 209328 18098 213375 18099
rect 209328 17880 213156 18098
rect 213374 17880 213375 18098
rect 209328 17879 213375 17880
rect 203328 17751 207219 17752
rect 203328 17533 207000 17751
rect 207218 17533 207219 17751
rect 203328 17532 207219 17533
rect 213904 17269 214124 18665
rect 215328 18563 215548 19666
rect 218328 18895 218548 19678
rect 218328 18675 220908 18895
rect 215328 18345 215329 18563
rect 215547 18345 215548 18563
rect 215328 18344 215548 18345
rect 213904 17051 213905 17269
rect 214123 17051 214124 17269
rect 213904 17050 214124 17051
rect 220688 17228 220908 18675
rect 221328 17711 221548 19666
rect 223548 18759 223868 18760
rect 223548 18441 223549 18759
rect 223867 18441 223868 18759
rect 223548 18440 223868 18441
rect 224328 18429 224548 19657
rect 227328 18940 227548 19675
rect 227328 18939 229878 18940
rect 227328 18721 229659 18939
rect 229877 18721 229878 18939
rect 227328 18720 229878 18721
rect 224328 18428 227414 18429
rect 224328 18210 227195 18428
rect 227413 18210 227414 18428
rect 224328 18209 227414 18210
rect 230328 18304 230548 19648
rect 232548 18759 232868 18760
rect 232548 18441 232549 18759
rect 232867 18441 232868 18759
rect 233328 18689 233548 19678
rect 233328 18471 233329 18689
rect 233547 18471 233548 18689
rect 233328 18470 233548 18471
rect 232548 18440 232868 18441
rect 230328 18303 234870 18304
rect 230328 18085 234651 18303
rect 234869 18085 234870 18303
rect 230328 18084 234870 18085
rect 236328 18016 236548 19498
rect 238548 18759 238868 18760
rect 238548 18441 238549 18759
rect 238867 18441 238868 18759
rect 238548 18440 238868 18441
rect 239328 18535 239548 19610
rect 242328 18570 242548 19678
rect 239328 18534 241892 18535
rect 239328 18316 241673 18534
rect 241891 18316 241892 18534
rect 242328 18352 242329 18570
rect 242547 18352 242548 18570
rect 245328 18599 245548 19678
rect 248328 19091 248548 19655
rect 248328 18871 249887 19091
rect 245328 18379 248931 18599
rect 242328 18351 242548 18352
rect 239328 18315 241892 18316
rect 236328 18015 241136 18016
rect 236328 17797 240917 18015
rect 241135 17797 241136 18015
rect 236328 17796 241136 17797
rect 221328 17493 221329 17711
rect 221547 17493 221548 17711
rect 221328 17492 221548 17493
rect 220688 17010 220689 17228
rect 220907 17010 220908 17228
rect 220688 17009 220908 17010
rect 248711 17077 248931 18379
rect 249667 17860 249887 18871
rect 250548 18759 250868 18760
rect 250548 18441 250549 18759
rect 250867 18441 250868 18759
rect 250548 18440 250868 18441
rect 251328 18510 251548 19678
rect 254328 18700 254548 19678
rect 251328 18509 254145 18510
rect 251328 18291 253926 18509
rect 254144 18291 254145 18509
rect 254328 18482 254329 18700
rect 254547 18482 254548 18700
rect 254328 18481 254548 18482
rect 257328 18577 257548 19671
rect 260328 19117 260548 19678
rect 260328 18897 261264 19117
rect 257328 18357 260273 18577
rect 251328 18290 254145 18291
rect 249667 17642 249668 17860
rect 249886 17642 249887 17860
rect 249667 17641 249887 17642
rect -4335 16687 -671 16797
rect -4335 13977 -4225 16687
rect 202003 16676 202004 16894
rect 202222 16676 202223 16894
rect 248711 16859 248712 17077
rect 248930 16859 248931 17077
rect 260053 17246 260273 18357
rect 261044 18125 261264 18897
rect 261044 17907 261045 18125
rect 261263 17907 261264 18125
rect 261044 17906 261264 17907
rect 263328 17964 263548 19678
rect 263948 18759 264268 18760
rect 263948 18441 263949 18759
rect 264267 18441 264268 18759
rect 263948 18440 264268 18441
rect 266328 18561 266548 19621
rect 266328 18560 269252 18561
rect 266328 18342 269033 18560
rect 269251 18342 269252 18560
rect 266328 18341 269252 18342
rect 269328 18268 269548 19594
rect 269948 18759 270268 18760
rect 269948 18441 269949 18759
rect 270267 18441 270268 18759
rect 269948 18440 270268 18441
rect 269328 18050 269329 18268
rect 269547 18050 269548 18268
rect 269328 18049 269548 18050
rect 263328 17963 266146 17964
rect 263328 17745 265871 17963
rect 266089 17745 266146 17963
rect 263328 17744 266146 17745
rect 272328 17583 272548 19649
rect 272948 18759 273268 18760
rect 272948 18441 272949 18759
rect 273267 18441 273268 18759
rect 272948 18440 273268 18441
rect 275328 18207 275548 19649
rect 275948 18759 276268 18760
rect 275948 18441 275949 18759
rect 276267 18441 276268 18759
rect 278328 18699 278548 19670
rect 278328 18698 279896 18699
rect 278328 18480 279677 18698
rect 279895 18480 279896 18698
rect 278328 18479 279896 18480
rect 275948 18440 276268 18441
rect 275328 18206 279098 18207
rect 275328 17988 278879 18206
rect 279097 17988 279098 18206
rect 275328 17987 279098 17988
rect 272328 17582 277913 17583
rect 272328 17364 277694 17582
rect 277912 17364 277913 17582
rect 272328 17363 277913 17364
rect 281328 17513 281548 19678
rect 281948 18759 282268 18760
rect 281948 18441 281949 18759
rect 282267 18441 282268 18759
rect 281948 18440 282268 18441
rect 284328 18137 284548 19678
rect 285948 18759 286268 18760
rect 285948 18441 285949 18759
rect 286267 18441 286268 18759
rect 285948 18440 286268 18441
rect 284328 17919 284329 18137
rect 284547 17919 284548 18137
rect 287328 18228 287548 19670
rect 290328 18955 290548 19678
rect 290328 18737 290329 18955
rect 290547 18737 290548 18955
rect 290328 18736 290548 18737
rect 287328 18227 292627 18228
rect 287328 18009 292408 18227
rect 292626 18009 292627 18227
rect 287328 18008 292627 18009
rect 284328 17918 284548 17919
rect 293328 17724 293548 19642
rect 293948 18759 294268 18760
rect 293948 18441 293949 18759
rect 294267 18441 294268 18759
rect 293948 18440 294268 18441
rect 296328 18328 296548 19655
rect 299328 19100 299548 19678
rect 299328 19099 305605 19100
rect 299328 18881 305386 19099
rect 305604 18881 305605 19099
rect 299328 18880 305605 18881
rect 296948 18759 297268 18760
rect 296948 18441 296949 18759
rect 297267 18441 297268 18759
rect 296948 18440 297268 18441
rect 299948 18759 300268 18760
rect 299948 18441 299949 18759
rect 300267 18441 300268 18759
rect 299948 18440 300268 18441
rect 302948 18759 303268 18760
rect 302948 18441 302949 18759
rect 303267 18441 303268 18759
rect 302948 18440 303268 18441
rect 296328 18108 300471 18328
rect 293328 17723 299478 17724
rect 281328 17512 287149 17513
rect 281328 17294 286930 17512
rect 287148 17294 287149 17512
rect 293328 17505 299259 17723
rect 299477 17505 299478 17723
rect 293328 17504 299478 17505
rect 281328 17293 287149 17294
rect 260053 17028 260054 17246
rect 260272 17028 260273 17246
rect 260053 17027 260273 17028
rect 300251 17105 300471 18108
rect 300251 16887 300252 17105
rect 300470 16887 300471 17105
rect 300251 16886 300471 16887
rect 303866 17265 304186 17289
rect 303866 16993 303890 17265
rect 304162 16993 304186 17265
rect 248711 16858 248931 16859
rect 202003 16675 202223 16676
rect 302941 16411 303275 16412
rect 302941 16410 302942 16411
rect 303274 16410 303275 16411
rect 18082 15707 18414 15708
rect 18082 15706 18083 15707
rect 18413 15706 18414 15707
rect 167542 15707 167874 15708
rect 167542 15706 167543 15707
rect 167873 15706 167874 15707
rect 3658 15689 3990 15690
rect 3658 15688 3659 15689
rect 3989 15688 3990 15689
rect 121672 15705 122004 15706
rect 121672 15704 121673 15705
rect 122003 15704 122004 15705
rect 64250 15691 64582 15692
rect 64250 15690 64251 15691
rect 64581 15690 64582 15691
rect 32908 15683 33240 15684
rect 32908 15682 32909 15683
rect 33239 15682 33240 15683
rect 180542 15707 180874 15708
rect 180542 15706 180543 15707
rect 180873 15706 180874 15707
rect 189542 15707 189874 15708
rect 189542 15706 189543 15707
rect 189873 15706 189874 15707
rect 198542 15707 198874 15708
rect 198542 15706 198543 15707
rect 198873 15706 198874 15707
rect 204542 15707 204874 15708
rect 204542 15706 204543 15707
rect 204873 15706 204874 15707
rect 211542 15707 211874 15708
rect 211542 15706 211543 15707
rect 211873 15706 211874 15707
rect 223542 15707 223874 15708
rect 223542 15706 223543 15707
rect 223873 15706 223874 15707
rect 232542 15707 232874 15708
rect 232542 15706 232543 15707
rect 232873 15706 232874 15707
rect 238542 15707 238874 15708
rect 238542 15706 238543 15707
rect 238873 15706 238874 15707
rect 250542 15707 250874 15708
rect 250542 15706 250543 15707
rect 250873 15706 250874 15707
rect 263942 15707 264274 15708
rect 263942 15706 263943 15707
rect 264273 15706 264274 15707
rect 269942 15707 270274 15708
rect 269942 15706 269943 15707
rect 270273 15706 270274 15707
rect 272942 15707 273274 15708
rect 272942 15706 272943 15707
rect 273273 15706 273274 15707
rect 275942 15707 276274 15708
rect 275942 15706 275943 15707
rect 276273 15706 276274 15707
rect 281942 15707 282274 15708
rect 281942 15706 281943 15707
rect 282273 15706 282274 15707
rect 285942 15707 286274 15708
rect 285942 15706 285943 15707
rect 286273 15706 286274 15707
rect 293942 15707 294274 15708
rect 293942 15706 293943 15707
rect 294273 15706 294274 15707
rect 296942 15707 297274 15708
rect 296942 15706 296943 15707
rect 297273 15706 297274 15707
rect 299942 15707 300274 15708
rect 299942 15706 299943 15707
rect 300273 15706 300274 15707
rect 302942 15707 303274 15708
rect 302942 15706 302943 15707
rect 303273 15706 303274 15707
rect 303866 15692 304186 16993
rect 303683 15396 303866 15668
<< via4 >>
rect -5523 321756 -5203 322076
rect -1502 321780 -1230 322052
rect 302448 324538 302768 324598
rect 302448 324338 302503 324538
rect 302503 324338 302713 324538
rect 302713 324338 302768 324538
rect 302448 324278 302768 324338
rect 303950 321062 304222 321334
rect -6294 319800 -5974 320120
rect -3762 319800 -3442 320120
rect -2994 319662 -2674 319982
rect -5523 318756 -5203 319076
rect -1502 318780 -1230 319052
rect 303950 318062 304222 318334
rect -6294 316800 -5974 317120
rect -3762 316800 -3442 317120
rect -2994 316662 -2674 316982
rect -5523 315756 -5203 316076
rect -1502 315780 -1230 316052
rect 303950 315062 304222 315334
rect -6294 313800 -5974 314120
rect -3762 313800 -3442 314120
rect -2994 313662 -2674 313982
rect -5523 312756 -5203 313076
rect -1502 312780 -1230 313052
rect 303950 312062 304222 312334
rect -6294 310800 -5974 311120
rect -3762 310800 -3442 311120
rect -2994 310662 -2674 310982
rect -5523 309756 -5203 310076
rect -1502 309780 -1230 310052
rect 303950 309062 304222 309334
rect -6294 307800 -5974 308120
rect -3762 307800 -3442 308120
rect -2994 307662 -2674 307982
rect -5523 306756 -5203 307076
rect -1502 306780 -1230 307052
rect 303950 306062 304222 306334
rect -6294 304800 -5974 305120
rect -3762 304800 -3442 305120
rect -2994 304662 -2674 304982
rect -5523 303756 -5203 304076
rect -1502 303780 -1230 304052
rect 303950 303062 304222 303334
rect -6294 301800 -5974 302120
rect -3762 301800 -3442 302120
rect -2994 301662 -2674 301982
rect -5523 300756 -5203 301076
rect -1502 300780 -1230 301052
rect 303950 300062 304222 300334
rect -6294 298800 -5974 299120
rect -3762 298800 -3442 299120
rect -2994 298662 -2674 298982
rect -5523 297756 -5203 298076
rect -1502 297780 -1230 298052
rect 303950 297062 304222 297334
rect -6294 295800 -5974 296120
rect -3762 295800 -3442 296120
rect -2994 295662 -2674 295982
rect -5523 294756 -5203 295076
rect -1502 294780 -1230 295052
rect 303950 294062 304222 294334
rect -6294 292800 -5974 293120
rect -3762 292800 -3442 293120
rect -2994 292662 -2674 292982
rect -5523 291756 -5203 292076
rect -1502 291780 -1230 292052
rect 303950 291062 304222 291334
rect -6294 289800 -5974 290120
rect -3762 289800 -3442 290120
rect -2994 289662 -2674 289982
rect -5523 288756 -5203 289076
rect -1502 288780 -1230 289052
rect 303950 288062 304222 288334
rect -6294 286800 -5974 287120
rect -3762 286800 -3442 287120
rect -2994 286662 -2674 286982
rect -5523 285756 -5203 286076
rect -1502 285780 -1230 286052
rect 303950 285062 304222 285334
rect -6294 283800 -5974 284120
rect -3762 283800 -3442 284120
rect -2994 283662 -2674 283982
rect -5523 282756 -5203 283076
rect -1502 282780 -1230 283052
rect 303950 282062 304222 282334
rect -6294 280800 -5974 281120
rect -3762 280800 -3442 281120
rect -2994 280662 -2674 280982
rect -5523 279756 -5203 280076
rect -1502 279780 -1230 280052
rect 303950 279062 304222 279334
rect -6294 277800 -5974 278120
rect -3762 277800 -3442 278120
rect -2994 277662 -2674 277982
rect -5523 276756 -5203 277076
rect -1502 276780 -1230 277052
rect 303950 276062 304222 276334
rect -6294 274800 -5974 275120
rect -3762 274800 -3442 275120
rect -2994 274662 -2674 274982
rect -5523 273756 -5203 274076
rect -1502 273780 -1230 274052
rect 303950 273062 304222 273334
rect -6294 271800 -5974 272120
rect -3762 271800 -3442 272120
rect -2994 271662 -2674 271982
rect -5523 270756 -5203 271076
rect -1502 270780 -1230 271052
rect 303950 270062 304222 270334
rect -6294 268800 -5974 269120
rect -3762 268800 -3442 269120
rect -2994 268662 -2674 268982
rect -5523 267756 -5203 268076
rect -1502 267780 -1230 268052
rect 303950 267062 304222 267334
rect -6294 265800 -5974 266120
rect -3762 265800 -3442 266120
rect -2994 265662 -2674 265982
rect -5523 264756 -5203 265076
rect -1502 264780 -1230 265052
rect 303950 264062 304222 264334
rect -6294 262800 -5974 263120
rect -3762 262800 -3442 263120
rect -2994 262662 -2674 262982
rect -5523 261756 -5203 262076
rect -1502 261780 -1230 262052
rect 303950 261062 304222 261334
rect -6294 259800 -5974 260120
rect -3762 259800 -3442 260120
rect -2994 259662 -2674 259982
rect -5523 258756 -5203 259076
rect -1502 258780 -1230 259052
rect 303950 258062 304222 258334
rect -6294 256800 -5974 257120
rect -3762 256800 -3442 257120
rect -2994 256662 -2674 256982
rect -5523 255756 -5203 256076
rect -1502 255780 -1230 256052
rect 303950 255062 304222 255334
rect -6294 253800 -5974 254120
rect -3762 253800 -3442 254120
rect -2994 253662 -2674 253982
rect -5523 252756 -5203 253076
rect -1502 252780 -1230 253052
rect 303950 252062 304222 252334
rect -6294 250800 -5974 251120
rect -3762 250800 -3442 251120
rect -2994 250662 -2674 250982
rect -5523 249756 -5203 250076
rect -1502 249780 -1230 250052
rect 303950 249062 304222 249334
rect -6294 247800 -5974 248120
rect -3762 247800 -3442 248120
rect -2994 247662 -2674 247982
rect 303950 246062 304222 246334
rect -6294 244800 -5974 245120
rect -3762 244800 -3442 245120
rect -2994 244662 -2674 244982
rect -5523 243756 -5203 244076
rect -1502 243780 -1230 244052
rect 303950 243062 304222 243334
rect -6294 241800 -5974 242120
rect -3762 241800 -3442 242120
rect -2994 241662 -2674 241982
rect -5523 240756 -5203 241076
rect -1502 240780 -1230 241052
rect 303950 240062 304222 240334
rect -6294 238800 -5974 239120
rect -3762 238800 -3442 239120
rect -2994 238662 -2674 238982
rect -5523 237756 -5203 238076
rect -1502 237780 -1230 238052
rect 303950 237062 304222 237334
rect -6294 235800 -5974 236120
rect -3762 235800 -3442 236120
rect -2994 235662 -2674 235982
rect -5523 234756 -5203 235076
rect -1502 234780 -1230 235052
rect 303950 234062 304222 234334
rect -6294 232800 -5974 233120
rect -3762 232800 -3442 233120
rect -2994 232662 -2674 232982
rect -5523 231756 -5203 232076
rect -1502 231780 -1230 232052
rect 303950 231062 304222 231334
rect -6294 229800 -5974 230120
rect -3762 229800 -3442 230120
rect -2994 229662 -2674 229982
rect -5523 228756 -5203 229076
rect -1502 228780 -1230 229052
rect 303950 228062 304222 228334
rect -6294 226800 -5974 227120
rect -3762 226800 -3442 227120
rect -2994 226662 -2674 226982
rect -5523 225756 -5203 226076
rect -1502 225780 -1230 226052
rect 303950 225062 304222 225334
rect -6294 223800 -5974 224120
rect -3762 223800 -3442 224120
rect -2994 223662 -2674 223982
rect -5523 222756 -5203 223076
rect -1502 222780 -1230 223052
rect 303950 222062 304222 222334
rect -6294 220800 -5974 221120
rect -3762 220800 -3442 221120
rect -2994 220662 -2674 220982
rect -5523 219756 -5203 220076
rect -1502 219780 -1230 220052
rect 303950 219062 304222 219334
rect -6294 217800 -5974 218120
rect -3762 217800 -3442 218120
rect -2994 217662 -2674 217982
rect -5523 216756 -5203 217076
rect -1502 216780 -1230 217052
rect 303950 216062 304222 216334
rect -6294 214800 -5974 215120
rect -3762 214800 -3442 215120
rect -2994 214662 -2674 214982
rect -5523 213756 -5203 214076
rect -1502 213780 -1230 214052
rect 303950 213062 304222 213334
rect -6294 211800 -5974 212120
rect -3762 211800 -3442 212120
rect -2994 211662 -2674 211982
rect -5523 210756 -5203 211076
rect -1502 210780 -1230 211052
rect 303950 210062 304222 210334
rect -2994 208662 -2674 208982
rect -5523 207756 -5203 208076
rect -1502 207780 -1230 208052
rect 303950 207062 304222 207334
rect -6294 205800 -5974 206120
rect -3762 205800 -3442 206120
rect -2994 205662 -2674 205982
rect -5523 204756 -5203 205076
rect -1502 204780 -1230 205052
rect 303950 204062 304222 204334
rect -6294 202800 -5974 203120
rect -3762 202800 -3442 203120
rect -2994 202662 -2674 202982
rect -5523 201756 -5203 202076
rect -1502 201780 -1230 202052
rect 303950 201062 304222 201334
rect -6294 199800 -5974 200120
rect -3762 199800 -3442 200120
rect -2994 199662 -2674 199982
rect -5523 198756 -5203 199076
rect -1502 198780 -1230 199052
rect 303950 198062 304222 198334
rect -6294 196800 -5974 197120
rect -3762 196800 -3442 197120
rect -2994 196662 -2674 196982
rect -5523 195756 -5203 196076
rect -1502 195780 -1230 196052
rect 303950 195062 304222 195334
rect -6294 193800 -5974 194120
rect -3762 193800 -3442 194120
rect -2994 193662 -2674 193982
rect -5523 192756 -5203 193076
rect -1502 192780 -1230 193052
rect 303950 192062 304222 192334
rect -6294 190800 -5974 191120
rect -3762 190800 -3442 191120
rect -2994 190662 -2674 190982
rect -5523 189756 -5203 190076
rect -1502 189780 -1230 190052
rect 303950 189062 304222 189334
rect -6294 187800 -5974 188120
rect -3762 187800 -3442 188120
rect -2994 187662 -2674 187982
rect -5523 186756 -5203 187076
rect -1502 186780 -1230 187052
rect 303950 186062 304222 186334
rect -6294 184800 -5974 185120
rect -3762 184800 -3442 185120
rect -2994 184662 -2674 184982
rect -5523 183756 -5203 184076
rect -1502 183780 -1230 184052
rect 303950 183062 304222 183334
rect -6294 181800 -5974 182120
rect -3762 181800 -3442 182120
rect -2994 181662 -2674 181982
rect -5523 180756 -5203 181076
rect -1502 180780 -1230 181052
rect 303950 180062 304222 180334
rect -6294 178800 -5974 179120
rect -3762 178800 -3442 179120
rect -2994 178662 -2674 178982
rect -5523 177756 -5203 178076
rect -1502 177780 -1230 178052
rect 303950 177062 304222 177334
rect -6294 175800 -5974 176120
rect -3762 175800 -3442 176120
rect -2994 175662 -2674 175982
rect -5523 174756 -5203 175076
rect -1502 174780 -1230 175052
rect 303950 174062 304222 174334
rect -6294 172800 -5974 173120
rect -3762 172800 -3442 173120
rect -2994 172662 -2674 172982
rect -5523 171756 -5203 172076
rect -1502 171780 -1230 172052
rect 303950 171062 304222 171334
rect -6294 169800 -5974 170120
rect -3762 169800 -3442 170120
rect -2994 169662 -2674 169982
rect -5523 168756 -5203 169076
rect -1502 168780 -1230 169052
rect 303950 168062 304222 168334
rect -6294 166800 -5974 167120
rect -3762 166800 -3442 167120
rect -2994 166662 -2674 166982
rect -5523 165756 -5203 166076
rect -1502 165780 -1230 166052
rect 303950 165062 304222 165334
rect -6294 163800 -5974 164120
rect -3762 163800 -3442 164120
rect -2994 163662 -2674 163982
rect -5523 162756 -5203 163076
rect -1502 162780 -1230 163052
rect 303950 162062 304222 162334
rect -6294 160800 -5974 161120
rect -3762 160800 -3442 161120
rect -2994 160662 -2674 160982
rect -5523 159756 -5203 160076
rect -1502 159780 -1230 160052
rect 303950 159062 304222 159334
rect -6294 157800 -5974 158120
rect -3762 157800 -3442 158120
rect -2994 157662 -2674 157982
rect -5523 156756 -5203 157076
rect -1502 156780 -1230 157052
rect 303950 156062 304222 156334
rect -6294 154800 -5974 155120
rect -3762 154800 -3442 155120
rect -2994 154662 -2674 154982
rect -5523 153756 -5203 154076
rect -1502 153780 -1230 154052
rect 303950 153062 304222 153334
rect -6294 151800 -5974 152120
rect -3762 151800 -3442 152120
rect -2994 151662 -2674 151982
rect -5523 150756 -5203 151076
rect -1502 150780 -1230 151052
rect 303950 150062 304222 150334
rect -6294 148800 -5974 149120
rect -3762 148800 -3442 149120
rect -2994 148662 -2674 148982
rect -5523 147756 -5203 148076
rect -1502 147780 -1230 148052
rect 303950 147062 304222 147334
rect -6294 145800 -5974 146120
rect -3762 145800 -3442 146120
rect -2994 145662 -2674 145982
rect -5523 144756 -5203 145076
rect -1502 144780 -1230 145052
rect 303950 144062 304222 144334
rect -6294 142800 -5974 143120
rect -3762 142800 -3442 143120
rect -2994 142662 -2674 142982
rect -5523 141756 -5203 142076
rect -1502 141780 -1230 142052
rect 303950 141062 304222 141334
rect -6294 139800 -5974 140120
rect -3762 139800 -3442 140120
rect -2994 139662 -2674 139982
rect -5523 138756 -5203 139076
rect -1502 138780 -1230 139052
rect 303950 138062 304222 138334
rect -6294 136800 -5974 137120
rect -3762 136800 -3442 137120
rect -2994 136662 -2674 136982
rect -5523 135756 -5203 136076
rect -1502 135780 -1230 136052
rect 303950 135062 304222 135334
rect -6294 133800 -5974 134120
rect -3762 133800 -3442 134120
rect -2994 133662 -2674 133982
rect -5523 132756 -5203 133076
rect -1502 132780 -1230 133052
rect 303950 132062 304222 132334
rect -6294 130800 -5974 131120
rect -3762 130800 -3442 131120
rect -2994 130662 -2674 130982
rect -5523 129756 -5203 130076
rect -1502 129780 -1230 130052
rect 303950 129062 304222 129334
rect -6294 127800 -5974 128120
rect -3762 127800 -3442 128120
rect -2994 127662 -2674 127982
rect -5523 126756 -5203 127076
rect -1502 126780 -1230 127052
rect 303950 126062 304222 126334
rect -6294 124800 -5974 125120
rect -3762 124800 -3442 125120
rect -2994 124662 -2674 124982
rect -5523 123756 -5203 124076
rect -1502 123780 -1230 124052
rect 303950 123062 304222 123334
rect -6294 121800 -5974 122120
rect -3762 121800 -3442 122120
rect -2994 121662 -2674 121982
rect -5523 120756 -5203 121076
rect -1502 120780 -1230 121052
rect 303950 120062 304222 120334
rect -6294 118800 -5974 119120
rect -3762 118800 -3442 119120
rect -2994 118662 -2674 118982
rect -5523 117756 -5203 118076
rect -1502 117780 -1230 118052
rect 303950 117062 304222 117334
rect -6294 115800 -5974 116120
rect -3762 115800 -3442 116120
rect -2994 115662 -2674 115982
rect -5523 114756 -5203 115076
rect -1502 114780 -1230 115052
rect 303950 114062 304222 114334
rect -6294 112800 -5974 113120
rect -3762 112800 -3442 113120
rect -2994 112662 -2674 112982
rect -5523 111756 -5203 112076
rect -1502 111780 -1230 112052
rect 303950 111062 304222 111334
rect -6294 109800 -5974 110120
rect -3762 109800 -3442 110120
rect -2994 109662 -2674 109982
rect -5523 108756 -5203 109076
rect -1502 108780 -1230 109052
rect 303950 108062 304222 108334
rect -6294 106800 -5974 107120
rect -3762 106800 -3442 107120
rect -2994 106662 -2674 106982
rect -5523 105756 -5203 106076
rect -1502 105780 -1230 106052
rect 303950 105062 304222 105334
rect -6294 103800 -5974 104120
rect -3762 103800 -3442 104120
rect -2994 103662 -2674 103982
rect -5523 102756 -5203 103076
rect -1502 102780 -1230 103052
rect 303950 102062 304222 102334
rect -6294 100800 -5974 101120
rect -3762 100800 -3442 101120
rect -2994 100662 -2674 100982
rect -5523 99756 -5203 100076
rect -1502 99780 -1230 100052
rect 303950 99062 304222 99334
rect -6294 97800 -5974 98120
rect -3762 97800 -3442 98120
rect -2994 97662 -2674 97982
rect -5523 96756 -5203 97076
rect -1502 96780 -1230 97052
rect 303950 96062 304222 96334
rect -6294 94800 -5974 95120
rect -3762 94800 -3442 95120
rect -2994 94662 -2674 94982
rect 303950 93062 304222 93334
rect -6294 91800 -5974 92120
rect -3762 91800 -3442 92120
rect -2994 91662 -2674 91982
rect -5523 90756 -5203 91076
rect -1502 90780 -1230 91052
rect 303950 90062 304222 90334
rect -6294 88800 -5974 89120
rect -3762 88800 -3442 89120
rect -2994 88662 -2674 88982
rect -5523 87756 -5203 88076
rect -1502 87780 -1230 88052
rect 303950 87062 304222 87334
rect -6294 85800 -5974 86120
rect -3762 85800 -3442 86120
rect -2994 85662 -2674 85982
rect -5523 84756 -5203 85076
rect -1502 84780 -1230 85052
rect 303950 84062 304222 84334
rect -6294 82800 -5974 83120
rect -3762 82800 -3442 83120
rect -2994 82662 -2674 82982
rect -5523 81756 -5203 82076
rect -1502 81780 -1230 82052
rect 303950 81062 304222 81334
rect -6294 79800 -5974 80120
rect -3762 79800 -3442 80120
rect -2994 79662 -2674 79982
rect -5523 78756 -5203 79076
rect -1502 78780 -1230 79052
rect 303950 78062 304222 78334
rect -6294 76800 -5974 77120
rect -3762 76800 -3442 77120
rect -2994 76662 -2674 76982
rect -5523 75756 -5203 76076
rect -1502 75780 -1230 76052
rect 303950 75062 304222 75334
rect -6294 73800 -5974 74120
rect -3762 73800 -3442 74120
rect -2994 73662 -2674 73982
rect -5523 72756 -5203 73076
rect -1502 72780 -1230 73052
rect 303950 72062 304222 72334
rect -6294 70800 -5974 71120
rect -3762 70800 -3442 71120
rect -2994 70662 -2674 70982
rect -5523 69756 -5203 70076
rect -1502 69780 -1230 70052
rect 303950 69062 304222 69334
rect -6294 67800 -5974 68120
rect -3762 67800 -3442 68120
rect -2994 67662 -2674 67982
rect -5523 66756 -5203 67076
rect -1502 66780 -1230 67052
rect 303950 66062 304222 66334
rect -6294 64800 -5974 65120
rect -3762 64800 -3442 65120
rect -2994 64662 -2674 64982
rect -5523 63756 -5203 64076
rect -1502 63780 -1230 64052
rect 303950 63062 304222 63334
rect -6294 61800 -5974 62120
rect -3762 61800 -3442 62120
rect -2994 61662 -2674 61982
rect -5523 60756 -5203 61076
rect -1502 60780 -1230 61052
rect 303950 60062 304222 60334
rect -6294 58800 -5974 59120
rect -3762 58800 -3442 59120
rect -2994 58662 -2674 58982
rect -5523 57756 -5203 58076
rect -1502 57780 -1230 58052
rect 303950 57062 304222 57334
rect -2994 55662 -2674 55982
rect -5523 54756 -5203 55076
rect -1502 54780 -1230 55052
rect 303950 54062 304222 54334
rect -6294 52800 -5974 53120
rect -3762 52800 -3442 53120
rect -2994 52662 -2674 52982
rect -5523 51756 -5203 52076
rect -1502 51780 -1230 52052
rect 303950 51062 304222 51334
rect -6294 49800 -5974 50120
rect -3762 49800 -3442 50120
rect -2994 49662 -2674 49982
rect -5523 48756 -5203 49076
rect -1502 48780 -1230 49052
rect 303950 48062 304222 48334
rect -6294 46800 -5974 47120
rect -3762 46800 -3442 47120
rect -2994 46662 -2674 46982
rect -5523 45756 -5203 46076
rect -1502 45780 -1230 46052
rect 303950 45062 304222 45334
rect -6294 43800 -5974 44120
rect -3762 43800 -3442 44120
rect -2994 43662 -2674 43982
rect -5523 42756 -5203 43076
rect -1502 42780 -1230 43052
rect 303950 42062 304222 42334
rect -6294 40800 -5974 41120
rect -3762 40800 -3442 41120
rect -2994 40662 -2674 40982
rect -5523 39756 -5203 40076
rect -1502 39780 -1230 40052
rect 303950 39062 304222 39334
rect -6294 37800 -5974 38120
rect -3762 37800 -3442 38120
rect -2994 37662 -2674 37982
rect -5523 36756 -5203 37076
rect -1502 36780 -1230 37052
rect 303950 36062 304222 36334
rect -6294 34800 -5974 35120
rect -3762 34800 -3442 35120
rect -2994 34662 -2674 34982
rect -5523 33756 -5203 34076
rect -1502 33780 -1230 34052
rect 303950 33062 304222 33334
rect -6294 31800 -5974 32120
rect -3762 31800 -3442 32120
rect -2994 31662 -2674 31982
rect -5523 30756 -5203 31076
rect -1502 30780 -1230 31052
rect 303950 30062 304222 30334
rect -6294 28800 -5974 29120
rect -3762 28800 -3442 29120
rect -2994 28662 -2674 28982
rect -5523 27756 -5203 28076
rect -1502 27780 -1230 28052
rect 303950 27062 304222 27334
rect -6294 25800 -5974 26120
rect -3762 25800 -3442 26120
rect -2994 25662 -2674 25982
rect -5523 24756 -5203 25076
rect -1502 24780 -1230 25052
rect 303950 24062 304222 24334
rect -6294 22800 -5974 23120
rect -3762 22800 -3442 23120
rect -2994 22662 -2674 22982
rect -5523 21756 -5203 22076
rect -1502 21780 -1230 22052
rect 303950 21062 304222 21334
rect -6294 19800 -5974 20120
rect -3762 19800 -3442 20120
rect -5523 18756 -5203 19076
rect -1502 18780 -1230 19052
rect -6415 17942 -6095 18002
rect -6415 17742 -6204 17942
rect -6204 17742 -6095 17942
rect -6415 17682 -6095 17742
rect 3688 18464 3960 18736
rect 18112 18464 18384 18736
rect 32938 18464 33210 18736
rect 64280 18464 64552 18736
rect 121702 18464 121974 18736
rect 167572 18464 167844 18736
rect 180572 18464 180844 18736
rect 189572 18464 189844 18736
rect 198572 18464 198844 18736
rect 204572 18464 204844 18736
rect 211572 18464 211844 18736
rect 223572 18464 223844 18736
rect 232572 18464 232844 18736
rect 238572 18464 238844 18736
rect 250572 18464 250844 18736
rect 263972 18464 264244 18736
rect 269972 18464 270244 18736
rect 272972 18464 273244 18736
rect 275972 18464 276244 18736
rect 281972 18464 282244 18736
rect 285972 18464 286244 18736
rect 293972 18464 294244 18736
rect 296972 18464 297244 18736
rect 299972 18464 300244 18736
rect 302972 18464 303244 18736
rect 303890 16993 304162 17265
rect 302941 16089 302942 16410
rect 302942 16089 303274 16410
rect 303274 16089 303275 16410
rect 302941 16088 303275 16089
rect 48 15583 368 15643
rect 48 15383 103 15583
rect 103 15383 313 15583
rect 313 15383 368 15583
rect 48 15323 368 15383
rect 3658 15369 3659 15688
rect 3659 15369 3989 15688
rect 3989 15369 3990 15688
rect 18082 15387 18083 15706
rect 18083 15387 18413 15706
rect 18413 15387 18414 15706
rect 18082 15386 18414 15387
rect 3658 15368 3990 15369
rect 32908 15363 32909 15682
rect 32909 15363 33239 15682
rect 33239 15363 33240 15682
rect 64250 15371 64251 15690
rect 64251 15371 64581 15690
rect 64581 15371 64582 15690
rect 121672 15385 121673 15704
rect 121673 15385 122003 15704
rect 122003 15385 122004 15704
rect 167542 15387 167543 15706
rect 167543 15387 167873 15706
rect 167873 15387 167874 15706
rect 167542 15386 167874 15387
rect 180542 15387 180543 15706
rect 180543 15387 180873 15706
rect 180873 15387 180874 15706
rect 180542 15386 180874 15387
rect 189542 15387 189543 15706
rect 189543 15387 189873 15706
rect 189873 15387 189874 15706
rect 189542 15386 189874 15387
rect 198542 15387 198543 15706
rect 198543 15387 198873 15706
rect 198873 15387 198874 15706
rect 198542 15386 198874 15387
rect 204542 15387 204543 15706
rect 204543 15387 204873 15706
rect 204873 15387 204874 15706
rect 204542 15386 204874 15387
rect 211542 15387 211543 15706
rect 211543 15387 211873 15706
rect 211873 15387 211874 15706
rect 211542 15386 211874 15387
rect 223542 15387 223543 15706
rect 223543 15387 223873 15706
rect 223873 15387 223874 15706
rect 223542 15386 223874 15387
rect 232542 15387 232543 15706
rect 232543 15387 232873 15706
rect 232873 15387 232874 15706
rect 232542 15386 232874 15387
rect 238542 15387 238543 15706
rect 238543 15387 238873 15706
rect 238873 15387 238874 15706
rect 238542 15386 238874 15387
rect 250542 15387 250543 15706
rect 250543 15387 250873 15706
rect 250873 15387 250874 15706
rect 250542 15386 250874 15387
rect 263942 15387 263943 15706
rect 263943 15387 264273 15706
rect 264273 15387 264274 15706
rect 263942 15386 264274 15387
rect 269942 15387 269943 15706
rect 269943 15387 270273 15706
rect 270273 15387 270274 15706
rect 269942 15386 270274 15387
rect 272942 15387 272943 15706
rect 272943 15387 273273 15706
rect 273273 15387 273274 15706
rect 272942 15386 273274 15387
rect 275942 15387 275943 15706
rect 275943 15387 276273 15706
rect 276273 15387 276274 15706
rect 275942 15386 276274 15387
rect 281942 15387 281943 15706
rect 281943 15387 282273 15706
rect 282273 15387 282274 15706
rect 281942 15386 282274 15387
rect 285942 15387 285943 15706
rect 285943 15387 286273 15706
rect 286273 15387 286274 15706
rect 285942 15386 286274 15387
rect 293942 15387 293943 15706
rect 293943 15387 294273 15706
rect 294273 15387 294274 15706
rect 293942 15386 294274 15387
rect 296942 15387 296943 15706
rect 296943 15387 297273 15706
rect 297273 15387 297274 15706
rect 296942 15386 297274 15387
rect 299942 15387 299943 15706
rect 299943 15387 300273 15706
rect 300273 15387 300274 15706
rect 299942 15386 300274 15387
rect 302942 15387 302943 15706
rect 302943 15387 303273 15706
rect 303273 15387 303274 15706
rect 302942 15386 303274 15387
rect 121672 15384 122004 15385
rect 303866 15372 304186 15692
rect 64250 15370 64582 15371
rect 32908 15362 33240 15363
<< metal5 >>
rect -2946 326542 -2626 326564
rect -1526 326542 -1206 326564
rect -2946 326222 305854 326542
rect -5547 322076 -5179 322100
rect -5547 321756 -5523 322076
rect -5203 321756 -5179 322076
rect -5547 321732 -5179 321756
rect -6318 320120 -5950 320144
rect -6318 319800 -6294 320120
rect -5974 319800 -5950 320120
rect -6318 319776 -5950 319800
rect -3786 320120 -3418 320144
rect -2946 320120 -2626 326222
rect -1526 326069 -1206 326222
rect -1526 324637 -1206 324684
rect 302448 324637 302768 324994
rect -1928 324598 304435 324637
rect -1928 324317 302448 324598
rect -3786 319800 -3762 320120
rect -3442 319982 -2626 320120
rect -3442 319800 -2994 319982
rect -3786 319776 -3418 319800
rect -3018 319662 -2994 319800
rect -2674 319662 -2626 319982
rect -3018 319638 -2626 319662
rect -5547 319076 -5179 319100
rect -5547 318756 -5523 319076
rect -5203 318756 -5179 319076
rect -5547 318732 -5179 318756
rect -6318 317120 -5950 317144
rect -6318 316800 -6294 317120
rect -5974 316800 -5950 317120
rect -6318 316776 -5950 316800
rect -3786 317120 -3418 317144
rect -2946 317120 -2626 319638
rect -3786 316800 -3762 317120
rect -3442 316982 -2626 317120
rect -3442 316800 -2994 316982
rect -3786 316776 -3418 316800
rect -3018 316662 -2994 316800
rect -2674 316662 -2626 316982
rect -1526 322052 -1206 324317
rect 302424 324278 302448 324317
rect 302768 324317 304435 324598
rect 302768 324278 302792 324317
rect 302424 324254 302792 324278
rect -1526 321780 -1502 322052
rect -1230 321780 -1206 322052
rect -1526 319052 -1206 321780
rect -1526 318780 -1502 319052
rect -1230 318780 -1206 319052
rect -1526 316960 -1206 318780
rect -3018 316638 -2626 316662
rect -1529 316640 -1206 316960
rect -5547 316076 -5179 316100
rect -5547 315756 -5523 316076
rect -5203 315756 -5179 316076
rect -5547 315732 -5179 315756
rect -6318 314120 -5950 314144
rect -6318 313800 -6294 314120
rect -5974 313800 -5950 314120
rect -6318 313776 -5950 313800
rect -3786 314120 -3418 314144
rect -2946 314120 -2626 316638
rect -3786 313800 -3762 314120
rect -3442 313982 -2626 314120
rect -3442 313800 -2994 313982
rect -3786 313776 -3418 313800
rect -3018 313662 -2994 313800
rect -2674 313662 -2626 313982
rect -1526 316052 -1206 316640
rect -1526 315780 -1502 316052
rect -1230 315780 -1206 316052
rect -1526 313960 -1206 315780
rect -3018 313638 -2626 313662
rect -1529 313640 -1206 313960
rect -5547 313076 -5179 313100
rect -5547 312756 -5523 313076
rect -5203 312756 -5179 313076
rect -5547 312732 -5179 312756
rect -6318 311120 -5950 311144
rect -6318 310800 -6294 311120
rect -5974 310800 -5950 311120
rect -6318 310776 -5950 310800
rect -3786 311120 -3418 311144
rect -2946 311120 -2626 313638
rect -3786 310800 -3762 311120
rect -3442 310982 -2626 311120
rect -3442 310800 -2994 310982
rect -3786 310776 -3418 310800
rect -3018 310662 -2994 310800
rect -2674 310662 -2626 310982
rect -1526 313052 -1206 313640
rect -1526 312780 -1502 313052
rect -1230 312780 -1206 313052
rect -1526 310960 -1206 312780
rect -3018 310638 -2626 310662
rect -1529 310640 -1206 310960
rect -5547 310076 -5179 310100
rect -5547 309756 -5523 310076
rect -5203 309756 -5179 310076
rect -5547 309732 -5179 309756
rect -6318 308120 -5950 308144
rect -6318 307800 -6294 308120
rect -5974 307800 -5950 308120
rect -6318 307776 -5950 307800
rect -3786 308120 -3418 308144
rect -2946 308120 -2626 310638
rect -3786 307800 -3762 308120
rect -3442 307982 -2626 308120
rect -3442 307800 -2994 307982
rect -3786 307776 -3418 307800
rect -3018 307662 -2994 307800
rect -2674 307662 -2626 307982
rect -1526 310052 -1206 310640
rect -1526 309780 -1502 310052
rect -1230 309780 -1206 310052
rect -1526 307960 -1206 309780
rect -3018 307638 -2626 307662
rect -1529 307640 -1206 307960
rect -5547 307076 -5179 307100
rect -5547 306756 -5523 307076
rect -5203 306756 -5179 307076
rect -5547 306732 -5179 306756
rect -6318 305120 -5950 305144
rect -6318 304800 -6294 305120
rect -5974 304800 -5950 305120
rect -6318 304776 -5950 304800
rect -3786 305120 -3418 305144
rect -2946 305120 -2626 307638
rect -3786 304800 -3762 305120
rect -3442 304982 -2626 305120
rect -3442 304800 -2994 304982
rect -3786 304776 -3418 304800
rect -3018 304662 -2994 304800
rect -2674 304662 -2626 304982
rect -1526 307052 -1206 307640
rect -1526 306780 -1502 307052
rect -1230 306780 -1206 307052
rect -1526 304960 -1206 306780
rect -3018 304638 -2626 304662
rect -1529 304640 -1206 304960
rect -5547 304076 -5179 304100
rect -5547 303756 -5523 304076
rect -5203 303756 -5179 304076
rect -5547 303732 -5179 303756
rect -6318 302120 -5950 302144
rect -6318 301800 -6294 302120
rect -5974 301800 -5950 302120
rect -6318 301776 -5950 301800
rect -3786 302120 -3418 302144
rect -2946 302120 -2626 304638
rect -3786 301800 -3762 302120
rect -3442 301982 -2626 302120
rect -3442 301800 -2994 301982
rect -3786 301776 -3418 301800
rect -3018 301662 -2994 301800
rect -2674 301662 -2626 301982
rect -1526 304052 -1206 304640
rect -1526 303780 -1502 304052
rect -1230 303780 -1206 304052
rect -1526 301960 -1206 303780
rect -3018 301638 -2626 301662
rect -1529 301640 -1206 301960
rect -5547 301076 -5179 301100
rect -5547 300756 -5523 301076
rect -5203 300756 -5179 301076
rect -5547 300732 -5179 300756
rect -6318 299120 -5950 299144
rect -6318 298800 -6294 299120
rect -5974 298800 -5950 299120
rect -6318 298776 -5950 298800
rect -3786 299120 -3418 299144
rect -2946 299120 -2626 301638
rect -3786 298800 -3762 299120
rect -3442 298982 -2626 299120
rect -3442 298800 -2994 298982
rect -3786 298776 -3418 298800
rect -3018 298662 -2994 298800
rect -2674 298662 -2626 298982
rect -1526 301052 -1206 301640
rect -1526 300780 -1502 301052
rect -1230 300780 -1206 301052
rect -1526 298960 -1206 300780
rect -3018 298638 -2626 298662
rect -1529 298640 -1206 298960
rect -5547 298076 -5179 298100
rect -5547 297756 -5523 298076
rect -5203 297756 -5179 298076
rect -5547 297732 -5179 297756
rect -6318 296120 -5950 296144
rect -6318 295800 -6294 296120
rect -5974 295800 -5950 296120
rect -6318 295776 -5950 295800
rect -3786 296120 -3418 296144
rect -2946 296120 -2626 298638
rect -3786 295800 -3762 296120
rect -3442 295982 -2626 296120
rect -3442 295800 -2994 295982
rect -3786 295776 -3418 295800
rect -3018 295662 -2994 295800
rect -2674 295662 -2626 295982
rect -1526 298052 -1206 298640
rect -1526 297780 -1502 298052
rect -1230 297780 -1206 298052
rect -1526 295960 -1206 297780
rect -3018 295638 -2626 295662
rect -1529 295640 -1206 295960
rect -5547 295076 -5179 295100
rect -5547 294756 -5523 295076
rect -5203 294756 -5179 295076
rect -5547 294732 -5179 294756
rect -6318 293120 -5950 293144
rect -6318 292800 -6294 293120
rect -5974 292800 -5950 293120
rect -6318 292776 -5950 292800
rect -3786 293120 -3418 293144
rect -2946 293120 -2626 295638
rect -3786 292800 -3762 293120
rect -3442 292982 -2626 293120
rect -3442 292800 -2994 292982
rect -3786 292776 -3418 292800
rect -3018 292662 -2994 292800
rect -2674 292662 -2626 292982
rect -1526 295052 -1206 295640
rect -1526 294780 -1502 295052
rect -1230 294780 -1206 295052
rect -1526 292960 -1206 294780
rect -3018 292638 -2626 292662
rect -1529 292640 -1206 292960
rect -5547 292076 -5179 292100
rect -5547 291756 -5523 292076
rect -5203 291756 -5179 292076
rect -5547 291732 -5179 291756
rect -6318 290120 -5950 290144
rect -6318 289800 -6294 290120
rect -5974 289800 -5950 290120
rect -6318 289776 -5950 289800
rect -3786 290120 -3418 290144
rect -2946 290120 -2626 292638
rect -3786 289800 -3762 290120
rect -3442 289982 -2626 290120
rect -3442 289800 -2994 289982
rect -3786 289776 -3418 289800
rect -3018 289662 -2994 289800
rect -2674 289662 -2626 289982
rect -1526 292052 -1206 292640
rect -1526 291780 -1502 292052
rect -1230 291780 -1206 292052
rect -1526 289960 -1206 291780
rect -3018 289638 -2626 289662
rect -1529 289640 -1206 289960
rect -5547 289076 -5179 289100
rect -5547 288756 -5523 289076
rect -5203 288756 -5179 289076
rect -5547 288732 -5179 288756
rect -6318 287120 -5950 287144
rect -6318 286800 -6294 287120
rect -5974 286800 -5950 287120
rect -6318 286776 -5950 286800
rect -3786 287120 -3418 287144
rect -2946 287120 -2626 289638
rect -3786 286800 -3762 287120
rect -3442 286982 -2626 287120
rect -3442 286800 -2994 286982
rect -3786 286776 -3418 286800
rect -3018 286662 -2994 286800
rect -2674 286662 -2626 286982
rect -1526 289052 -1206 289640
rect -1526 288780 -1502 289052
rect -1230 288780 -1206 289052
rect -1526 286960 -1206 288780
rect -3018 286638 -2626 286662
rect -1529 286640 -1206 286960
rect -5547 286076 -5179 286100
rect -5547 285756 -5523 286076
rect -5203 285756 -5179 286076
rect -5547 285732 -5179 285756
rect -6318 284120 -5950 284144
rect -6318 283800 -6294 284120
rect -5974 283800 -5950 284120
rect -6318 283776 -5950 283800
rect -3786 284120 -3418 284144
rect -2946 284120 -2626 286638
rect -3786 283800 -3762 284120
rect -3442 283982 -2626 284120
rect -3442 283800 -2994 283982
rect -3786 283776 -3418 283800
rect -3018 283662 -2994 283800
rect -2674 283662 -2626 283982
rect -1526 286052 -1206 286640
rect -1526 285780 -1502 286052
rect -1230 285780 -1206 286052
rect -1526 283960 -1206 285780
rect -3018 283638 -2626 283662
rect -1529 283640 -1206 283960
rect -5547 283076 -5179 283100
rect -5547 282756 -5523 283076
rect -5203 282756 -5179 283076
rect -5547 282732 -5179 282756
rect -6318 281120 -5950 281144
rect -6318 280800 -6294 281120
rect -5974 280800 -5950 281120
rect -6318 280776 -5950 280800
rect -3786 281120 -3418 281144
rect -2946 281120 -2626 283638
rect -3786 280800 -3762 281120
rect -3442 280982 -2626 281120
rect -3442 280800 -2994 280982
rect -3786 280776 -3418 280800
rect -3018 280662 -2994 280800
rect -2674 280662 -2626 280982
rect -1526 283052 -1206 283640
rect -1526 282780 -1502 283052
rect -1230 282780 -1206 283052
rect -1526 280960 -1206 282780
rect -3018 280638 -2626 280662
rect -1529 280640 -1206 280960
rect -5547 280076 -5179 280100
rect -5547 279756 -5523 280076
rect -5203 279756 -5179 280076
rect -5547 279732 -5179 279756
rect -6318 278120 -5950 278144
rect -6318 277800 -6294 278120
rect -5974 277800 -5950 278120
rect -6318 277776 -5950 277800
rect -3786 278120 -3418 278144
rect -2946 278120 -2626 280638
rect -3786 277800 -3762 278120
rect -3442 277982 -2626 278120
rect -3442 277800 -2994 277982
rect -3786 277776 -3418 277800
rect -3018 277662 -2994 277800
rect -2674 277662 -2626 277982
rect -1526 280052 -1206 280640
rect -1526 279780 -1502 280052
rect -1230 279780 -1206 280052
rect -1526 277960 -1206 279780
rect -3018 277638 -2626 277662
rect -1529 277640 -1206 277960
rect -5547 277076 -5179 277100
rect -5547 276756 -5523 277076
rect -5203 276756 -5179 277076
rect -5547 276732 -5179 276756
rect -6318 275120 -5950 275144
rect -6318 274800 -6294 275120
rect -5974 274800 -5950 275120
rect -6318 274776 -5950 274800
rect -3786 275120 -3418 275144
rect -2946 275120 -2626 277638
rect -3786 274800 -3762 275120
rect -3442 274982 -2626 275120
rect -3442 274800 -2994 274982
rect -3786 274776 -3418 274800
rect -3018 274662 -2994 274800
rect -2674 274662 -2626 274982
rect -1526 277052 -1206 277640
rect -1526 276780 -1502 277052
rect -1230 276780 -1206 277052
rect -1526 274960 -1206 276780
rect -3018 274638 -2626 274662
rect -1529 274640 -1206 274960
rect -5547 274076 -5179 274100
rect -5547 273756 -5523 274076
rect -5203 273756 -5179 274076
rect -5547 273732 -5179 273756
rect -6318 272120 -5950 272144
rect -6318 271800 -6294 272120
rect -5974 271800 -5950 272120
rect -6318 271776 -5950 271800
rect -3786 272120 -3418 272144
rect -2946 272120 -2626 274638
rect -3786 271800 -3762 272120
rect -3442 271982 -2626 272120
rect -3442 271800 -2994 271982
rect -3786 271776 -3418 271800
rect -3018 271662 -2994 271800
rect -2674 271662 -2626 271982
rect -1526 274052 -1206 274640
rect -1526 273780 -1502 274052
rect -1230 273780 -1206 274052
rect -1526 271960 -1206 273780
rect -3018 271638 -2626 271662
rect -1529 271640 -1206 271960
rect -5547 271076 -5179 271100
rect -5547 270756 -5523 271076
rect -5203 270756 -5179 271076
rect -5547 270732 -5179 270756
rect -6318 269120 -5950 269144
rect -6318 268800 -6294 269120
rect -5974 268800 -5950 269120
rect -6318 268776 -5950 268800
rect -3786 269120 -3418 269144
rect -2946 269120 -2626 271638
rect -3786 268800 -3762 269120
rect -3442 268982 -2626 269120
rect -3442 268800 -2994 268982
rect -3786 268776 -3418 268800
rect -3018 268662 -2994 268800
rect -2674 268662 -2626 268982
rect -1526 271052 -1206 271640
rect -1526 270780 -1502 271052
rect -1230 270780 -1206 271052
rect -1526 268960 -1206 270780
rect -3018 268638 -2626 268662
rect -1529 268640 -1206 268960
rect -5547 268076 -5179 268100
rect -5547 267756 -5523 268076
rect -5203 267756 -5179 268076
rect -5547 267732 -5179 267756
rect -6318 266120 -5950 266144
rect -6318 265800 -6294 266120
rect -5974 265800 -5950 266120
rect -6318 265776 -5950 265800
rect -3786 266120 -3418 266144
rect -2946 266120 -2626 268638
rect -3786 265800 -3762 266120
rect -3442 265982 -2626 266120
rect -3442 265800 -2994 265982
rect -3786 265776 -3418 265800
rect -3018 265662 -2994 265800
rect -2674 265662 -2626 265982
rect -1526 268052 -1206 268640
rect -1526 267780 -1502 268052
rect -1230 267780 -1206 268052
rect -1526 265960 -1206 267780
rect -3018 265638 -2626 265662
rect -1529 265640 -1206 265960
rect -5547 265076 -5179 265100
rect -5547 264756 -5523 265076
rect -5203 264756 -5179 265076
rect -5547 264732 -5179 264756
rect -6318 263120 -5950 263144
rect -6318 262800 -6294 263120
rect -5974 262800 -5950 263120
rect -6318 262776 -5950 262800
rect -3786 263120 -3418 263144
rect -2946 263120 -2626 265638
rect -3786 262800 -3762 263120
rect -3442 262982 -2626 263120
rect -3442 262800 -2994 262982
rect -3786 262776 -3418 262800
rect -3018 262662 -2994 262800
rect -2674 262662 -2626 262982
rect -1526 265052 -1206 265640
rect -1526 264780 -1502 265052
rect -1230 264780 -1206 265052
rect -1526 262960 -1206 264780
rect -3018 262638 -2626 262662
rect -1529 262640 -1206 262960
rect -5547 262076 -5179 262100
rect -5547 261756 -5523 262076
rect -5203 261756 -5179 262076
rect -5547 261732 -5179 261756
rect -6318 260120 -5950 260144
rect -6318 259800 -6294 260120
rect -5974 259800 -5950 260120
rect -6318 259776 -5950 259800
rect -3786 260120 -3418 260144
rect -2946 260120 -2626 262638
rect -3786 259800 -3762 260120
rect -3442 259982 -2626 260120
rect -3442 259800 -2994 259982
rect -3786 259776 -3418 259800
rect -3018 259662 -2994 259800
rect -2674 259662 -2626 259982
rect -1526 262052 -1206 262640
rect -1526 261780 -1502 262052
rect -1230 261780 -1206 262052
rect -1526 259960 -1206 261780
rect -3018 259638 -2626 259662
rect -1529 259640 -1206 259960
rect -5547 259076 -5179 259100
rect -5547 258756 -5523 259076
rect -5203 258756 -5179 259076
rect -5547 258732 -5179 258756
rect -6318 257120 -5950 257144
rect -6318 256800 -6294 257120
rect -5974 256800 -5950 257120
rect -6318 256776 -5950 256800
rect -3786 257120 -3418 257144
rect -2946 257120 -2626 259638
rect -3786 256800 -3762 257120
rect -3442 256982 -2626 257120
rect -3442 256800 -2994 256982
rect -3786 256776 -3418 256800
rect -3018 256662 -2994 256800
rect -2674 256662 -2626 256982
rect -1526 259052 -1206 259640
rect -1526 258780 -1502 259052
rect -1230 258780 -1206 259052
rect -1526 256960 -1206 258780
rect -3018 256638 -2626 256662
rect -1529 256640 -1206 256960
rect -5547 256076 -5179 256100
rect -5547 255756 -5523 256076
rect -5203 255756 -5179 256076
rect -5547 255732 -5179 255756
rect -6318 254120 -5950 254144
rect -6318 253800 -6294 254120
rect -5974 253800 -5950 254120
rect -6318 253776 -5950 253800
rect -3786 254120 -3418 254144
rect -2946 254120 -2626 256638
rect -3786 253800 -3762 254120
rect -3442 253982 -2626 254120
rect -3442 253800 -2994 253982
rect -3786 253776 -3418 253800
rect -3018 253662 -2994 253800
rect -2674 253662 -2626 253982
rect -1526 256052 -1206 256640
rect -1526 255780 -1502 256052
rect -1230 255780 -1206 256052
rect -1526 253960 -1206 255780
rect -3018 253638 -2626 253662
rect -1529 253640 -1206 253960
rect -5547 253076 -5179 253100
rect -5547 252756 -5523 253076
rect -5203 252756 -5179 253076
rect -5547 252732 -5179 252756
rect -6318 251120 -5950 251144
rect -6318 250800 -6294 251120
rect -5974 250800 -5950 251120
rect -6318 250776 -5950 250800
rect -3786 251120 -3418 251144
rect -2946 251120 -2626 253638
rect -3786 250800 -3762 251120
rect -3442 250982 -2626 251120
rect -3442 250800 -2994 250982
rect -3786 250776 -3418 250800
rect -3018 250662 -2994 250800
rect -2674 250662 -2626 250982
rect -1526 253052 -1206 253640
rect -1526 252780 -1502 253052
rect -1230 252780 -1206 253052
rect -1526 250960 -1206 252780
rect -3018 250638 -2626 250662
rect -1529 250640 -1206 250960
rect -5547 250076 -5179 250100
rect -5547 249756 -5523 250076
rect -5203 249756 -5179 250076
rect -5547 249732 -5179 249756
rect -6318 248120 -5950 248144
rect -6318 247800 -6294 248120
rect -5974 247800 -5950 248120
rect -6318 247776 -5950 247800
rect -3786 248120 -3418 248144
rect -2946 248120 -2626 250638
rect -3786 247800 -3762 248120
rect -3442 247982 -2626 248120
rect -3442 247800 -2994 247982
rect -3786 247776 -3418 247800
rect -3018 247662 -2994 247800
rect -2674 247662 -2626 247982
rect -1526 250052 -1206 250640
rect -1526 249780 -1502 250052
rect -1230 249780 -1206 250052
rect -1526 247960 -1206 249780
rect -3018 247638 -2626 247662
rect -1529 247640 -1206 247960
rect -6318 245120 -5950 245144
rect -6318 244800 -6294 245120
rect -5974 244800 -5950 245120
rect -6318 244776 -5950 244800
rect -3786 245120 -3418 245144
rect -2946 245120 -2626 247638
rect -3786 244800 -3762 245120
rect -3442 244982 -2626 245120
rect -3442 244800 -2994 244982
rect -3786 244776 -3418 244800
rect -3018 244662 -2994 244800
rect -2674 244662 -2626 244982
rect -1526 244960 -1206 247640
rect -3018 244638 -2626 244662
rect -1529 244640 -1206 244960
rect -5547 244076 -5179 244100
rect -5547 243756 -5523 244076
rect -5203 243756 -5179 244076
rect -5547 243732 -5179 243756
rect -6318 242120 -5950 242144
rect -6318 241800 -6294 242120
rect -5974 241800 -5950 242120
rect -6318 241776 -5950 241800
rect -3786 242120 -3418 242144
rect -2946 242120 -2626 244638
rect -3786 241800 -3762 242120
rect -3442 241982 -2626 242120
rect -3442 241800 -2994 241982
rect -3786 241776 -3418 241800
rect -3018 241662 -2994 241800
rect -2674 241662 -2626 241982
rect -1526 244052 -1206 244640
rect -1526 243780 -1502 244052
rect -1230 243780 -1206 244052
rect -1526 241960 -1206 243780
rect -3018 241638 -2626 241662
rect -1529 241640 -1206 241960
rect -5547 241076 -5179 241100
rect -5547 240756 -5523 241076
rect -5203 240756 -5179 241076
rect -5547 240732 -5179 240756
rect -6318 239120 -5950 239144
rect -6318 238800 -6294 239120
rect -5974 238800 -5950 239120
rect -6318 238776 -5950 238800
rect -3786 239120 -3418 239144
rect -2946 239120 -2626 241638
rect -3786 238800 -3762 239120
rect -3442 238982 -2626 239120
rect -3442 238800 -2994 238982
rect -3786 238776 -3418 238800
rect -3018 238662 -2994 238800
rect -2674 238662 -2626 238982
rect -1526 241052 -1206 241640
rect -1526 240780 -1502 241052
rect -1230 240780 -1206 241052
rect -1526 238960 -1206 240780
rect -3018 238638 -2626 238662
rect -1529 238640 -1206 238960
rect -5547 238076 -5179 238100
rect -5547 237756 -5523 238076
rect -5203 237756 -5179 238076
rect -5547 237732 -5179 237756
rect -6318 236120 -5950 236144
rect -6318 235800 -6294 236120
rect -5974 235800 -5950 236120
rect -6318 235776 -5950 235800
rect -3786 236120 -3418 236144
rect -2946 236120 -2626 238638
rect -3786 235800 -3762 236120
rect -3442 235982 -2626 236120
rect -3442 235800 -2994 235982
rect -3786 235776 -3418 235800
rect -3018 235662 -2994 235800
rect -2674 235662 -2626 235982
rect -1526 238052 -1206 238640
rect -1526 237780 -1502 238052
rect -1230 237780 -1206 238052
rect -1526 235960 -1206 237780
rect -3018 235638 -2626 235662
rect -1529 235640 -1206 235960
rect -5547 235076 -5179 235100
rect -5547 234756 -5523 235076
rect -5203 234756 -5179 235076
rect -5547 234732 -5179 234756
rect -6318 233120 -5950 233144
rect -6318 232800 -6294 233120
rect -5974 232800 -5950 233120
rect -6318 232776 -5950 232800
rect -3786 233120 -3418 233144
rect -2946 233120 -2626 235638
rect -3786 232800 -3762 233120
rect -3442 232982 -2626 233120
rect -3442 232800 -2994 232982
rect -3786 232776 -3418 232800
rect -3018 232662 -2994 232800
rect -2674 232662 -2626 232982
rect -1526 235052 -1206 235640
rect -1526 234780 -1502 235052
rect -1230 234780 -1206 235052
rect -1526 232960 -1206 234780
rect -3018 232638 -2626 232662
rect -1529 232640 -1206 232960
rect -5547 232076 -5179 232100
rect -5547 231756 -5523 232076
rect -5203 231756 -5179 232076
rect -5547 231732 -5179 231756
rect -6318 230120 -5950 230144
rect -6318 229800 -6294 230120
rect -5974 229800 -5950 230120
rect -6318 229776 -5950 229800
rect -3786 230120 -3418 230144
rect -2946 230120 -2626 232638
rect -3786 229800 -3762 230120
rect -3442 229982 -2626 230120
rect -3442 229800 -2994 229982
rect -3786 229776 -3418 229800
rect -3018 229662 -2994 229800
rect -2674 229662 -2626 229982
rect -1526 232052 -1206 232640
rect -1526 231780 -1502 232052
rect -1230 231780 -1206 232052
rect -1526 229960 -1206 231780
rect -3018 229638 -2626 229662
rect -1529 229640 -1206 229960
rect -5547 229076 -5179 229100
rect -5547 228756 -5523 229076
rect -5203 228756 -5179 229076
rect -5547 228732 -5179 228756
rect -6318 227120 -5950 227144
rect -6318 226800 -6294 227120
rect -5974 226800 -5950 227120
rect -6318 226776 -5950 226800
rect -3786 227120 -3418 227144
rect -2946 227120 -2626 229638
rect -3786 226800 -3762 227120
rect -3442 226982 -2626 227120
rect -3442 226800 -2994 226982
rect -3786 226776 -3418 226800
rect -3018 226662 -2994 226800
rect -2674 226662 -2626 226982
rect -1526 229052 -1206 229640
rect -1526 228780 -1502 229052
rect -1230 228780 -1206 229052
rect -1526 226960 -1206 228780
rect -3018 226638 -2626 226662
rect -1529 226640 -1206 226960
rect -5547 226076 -5179 226100
rect -5547 225756 -5523 226076
rect -5203 225756 -5179 226076
rect -5547 225732 -5179 225756
rect -6318 224120 -5950 224144
rect -6318 223800 -6294 224120
rect -5974 223800 -5950 224120
rect -6318 223776 -5950 223800
rect -3786 224120 -3418 224144
rect -2946 224120 -2626 226638
rect -3786 223800 -3762 224120
rect -3442 223982 -2626 224120
rect -3442 223800 -2994 223982
rect -3786 223776 -3418 223800
rect -3018 223662 -2994 223800
rect -2674 223662 -2626 223982
rect -1526 226052 -1206 226640
rect -1526 225780 -1502 226052
rect -1230 225780 -1206 226052
rect -1526 223960 -1206 225780
rect -3018 223638 -2626 223662
rect -1529 223640 -1206 223960
rect -5547 223076 -5179 223100
rect -5547 222756 -5523 223076
rect -5203 222756 -5179 223076
rect -5547 222732 -5179 222756
rect -6318 221120 -5950 221144
rect -6318 220800 -6294 221120
rect -5974 220800 -5950 221120
rect -6318 220776 -5950 220800
rect -3786 221120 -3418 221144
rect -2946 221120 -2626 223638
rect -3786 220800 -3762 221120
rect -3442 220982 -2626 221120
rect -3442 220800 -2994 220982
rect -3786 220776 -3418 220800
rect -3018 220662 -2994 220800
rect -2674 220662 -2626 220982
rect -1526 223052 -1206 223640
rect -1526 222780 -1502 223052
rect -1230 222780 -1206 223052
rect -1526 220960 -1206 222780
rect -3018 220638 -2626 220662
rect -1529 220640 -1206 220960
rect -5547 220076 -5179 220100
rect -5547 219756 -5523 220076
rect -5203 219756 -5179 220076
rect -5547 219732 -5179 219756
rect -6318 218120 -5950 218144
rect -6318 217800 -6294 218120
rect -5974 217800 -5950 218120
rect -6318 217776 -5950 217800
rect -3786 218120 -3418 218144
rect -2946 218120 -2626 220638
rect -3786 217800 -3762 218120
rect -3442 217982 -2626 218120
rect -3442 217800 -2994 217982
rect -3786 217776 -3418 217800
rect -3018 217662 -2994 217800
rect -2674 217662 -2626 217982
rect -1526 220052 -1206 220640
rect -1526 219780 -1502 220052
rect -1230 219780 -1206 220052
rect -1526 217960 -1206 219780
rect -3018 217638 -2626 217662
rect -1529 217640 -1206 217960
rect -5547 217076 -5179 217100
rect -5547 216756 -5523 217076
rect -5203 216756 -5179 217076
rect -5547 216732 -5179 216756
rect -6318 215120 -5950 215144
rect -6318 214800 -6294 215120
rect -5974 214800 -5950 215120
rect -6318 214776 -5950 214800
rect -3786 215120 -3418 215144
rect -2946 215120 -2626 217638
rect -3786 214800 -3762 215120
rect -3442 214982 -2626 215120
rect -3442 214800 -2994 214982
rect -3786 214776 -3418 214800
rect -3018 214662 -2994 214800
rect -2674 214662 -2626 214982
rect -1526 217052 -1206 217640
rect -1526 216780 -1502 217052
rect -1230 216780 -1206 217052
rect -1526 214960 -1206 216780
rect -3018 214638 -2626 214662
rect -1529 214640 -1206 214960
rect -5547 214076 -5179 214100
rect -5547 213756 -5523 214076
rect -5203 213756 -5179 214076
rect -5547 213732 -5179 213756
rect -6318 212120 -5950 212144
rect -6318 211800 -6294 212120
rect -5974 211800 -5950 212120
rect -6318 211776 -5950 211800
rect -3786 212120 -3418 212144
rect -2946 212120 -2626 214638
rect -3786 211800 -3762 212120
rect -3442 211982 -2626 212120
rect -3442 211800 -2994 211982
rect -3786 211776 -3418 211800
rect -3018 211662 -2994 211800
rect -2674 211662 -2626 211982
rect -1526 214052 -1206 214640
rect -1526 213780 -1502 214052
rect -1230 213780 -1206 214052
rect -1526 211960 -1206 213780
rect -3018 211638 -2626 211662
rect -1529 211640 -1206 211960
rect -5547 211076 -5179 211100
rect -5547 210756 -5523 211076
rect -5203 210756 -5179 211076
rect -5547 210732 -5179 210756
rect -2946 209120 -2626 211638
rect -3120 208982 -2626 209120
rect -3120 208800 -2994 208982
rect -3018 208662 -2994 208800
rect -2674 208662 -2626 208982
rect -1526 211052 -1206 211640
rect -1526 210780 -1502 211052
rect -1230 210780 -1206 211052
rect -1526 208960 -1206 210780
rect -3018 208638 -2626 208662
rect -1529 208640 -1206 208960
rect -5547 208076 -5179 208100
rect -5547 207756 -5523 208076
rect -5203 207756 -5179 208076
rect -5547 207732 -5179 207756
rect -6318 206120 -5950 206144
rect -6318 205800 -6294 206120
rect -5974 205800 -5950 206120
rect -6318 205776 -5950 205800
rect -3786 206120 -3418 206144
rect -2946 206120 -2626 208638
rect -3786 205800 -3762 206120
rect -3442 205982 -2626 206120
rect -3442 205800 -2994 205982
rect -3786 205776 -3418 205800
rect -3018 205662 -2994 205800
rect -2674 205662 -2626 205982
rect -1526 208052 -1206 208640
rect -1526 207780 -1502 208052
rect -1230 207780 -1206 208052
rect -1526 205960 -1206 207780
rect -3018 205638 -2626 205662
rect -1529 205640 -1206 205960
rect -5547 205076 -5179 205100
rect -5547 204756 -5523 205076
rect -5203 204756 -5179 205076
rect -5547 204732 -5179 204756
rect -6318 203120 -5950 203144
rect -6318 202800 -6294 203120
rect -5974 202800 -5950 203120
rect -6318 202776 -5950 202800
rect -3786 203120 -3418 203144
rect -2946 203120 -2626 205638
rect -3786 202800 -3762 203120
rect -3442 202982 -2626 203120
rect -3442 202800 -2994 202982
rect -3786 202776 -3418 202800
rect -3018 202662 -2994 202800
rect -2674 202662 -2626 202982
rect -1526 205052 -1206 205640
rect -1526 204780 -1502 205052
rect -1230 204780 -1206 205052
rect -1526 202960 -1206 204780
rect -3018 202638 -2626 202662
rect -1529 202640 -1206 202960
rect -5547 202076 -5179 202100
rect -5547 201756 -5523 202076
rect -5203 201756 -5179 202076
rect -5547 201732 -5179 201756
rect -6318 200120 -5950 200144
rect -6318 199800 -6294 200120
rect -5974 199800 -5950 200120
rect -6318 199776 -5950 199800
rect -3786 200120 -3418 200144
rect -2946 200120 -2626 202638
rect -3786 199800 -3762 200120
rect -3442 199982 -2626 200120
rect -3442 199800 -2994 199982
rect -3786 199776 -3418 199800
rect -3018 199662 -2994 199800
rect -2674 199662 -2626 199982
rect -1526 202052 -1206 202640
rect -1526 201780 -1502 202052
rect -1230 201780 -1206 202052
rect -1526 199960 -1206 201780
rect -3018 199638 -2626 199662
rect -1529 199640 -1206 199960
rect -5547 199076 -5179 199100
rect -5547 198756 -5523 199076
rect -5203 198756 -5179 199076
rect -5547 198732 -5179 198756
rect -6318 197120 -5950 197144
rect -6318 196800 -6294 197120
rect -5974 196800 -5950 197120
rect -6318 196776 -5950 196800
rect -3786 197120 -3418 197144
rect -2946 197120 -2626 199638
rect -3786 196800 -3762 197120
rect -3442 196982 -2626 197120
rect -3442 196800 -2994 196982
rect -3786 196776 -3418 196800
rect -3018 196662 -2994 196800
rect -2674 196662 -2626 196982
rect -1526 199052 -1206 199640
rect -1526 198780 -1502 199052
rect -1230 198780 -1206 199052
rect -1526 196960 -1206 198780
rect -3018 196638 -2626 196662
rect -1529 196640 -1206 196960
rect -5547 196076 -5179 196100
rect -5547 195756 -5523 196076
rect -5203 195756 -5179 196076
rect -5547 195732 -5179 195756
rect -6318 194120 -5950 194144
rect -6318 193800 -6294 194120
rect -5974 193800 -5950 194120
rect -6318 193776 -5950 193800
rect -3786 194120 -3418 194144
rect -2946 194120 -2626 196638
rect -3786 193800 -3762 194120
rect -3442 193982 -2626 194120
rect -3442 193800 -2994 193982
rect -3786 193776 -3418 193800
rect -3018 193662 -2994 193800
rect -2674 193662 -2626 193982
rect -1526 196052 -1206 196640
rect -1526 195780 -1502 196052
rect -1230 195780 -1206 196052
rect -1526 193960 -1206 195780
rect -3018 193638 -2626 193662
rect -1529 193640 -1206 193960
rect -5547 193076 -5179 193100
rect -5547 192756 -5523 193076
rect -5203 192756 -5179 193076
rect -5547 192732 -5179 192756
rect -6318 191120 -5950 191144
rect -6318 190800 -6294 191120
rect -5974 190800 -5950 191120
rect -6318 190776 -5950 190800
rect -3786 191120 -3418 191144
rect -2946 191120 -2626 193638
rect -3786 190800 -3762 191120
rect -3442 190982 -2626 191120
rect -3442 190800 -2994 190982
rect -3786 190776 -3418 190800
rect -3018 190662 -2994 190800
rect -2674 190662 -2626 190982
rect -1526 193052 -1206 193640
rect -1526 192780 -1502 193052
rect -1230 192780 -1206 193052
rect -1526 190960 -1206 192780
rect -3018 190638 -2626 190662
rect -1529 190640 -1206 190960
rect -5547 190076 -5179 190100
rect -5547 189756 -5523 190076
rect -5203 189756 -5179 190076
rect -5547 189732 -5179 189756
rect -6318 188120 -5950 188144
rect -6318 187800 -6294 188120
rect -5974 187800 -5950 188120
rect -6318 187776 -5950 187800
rect -3786 188120 -3418 188144
rect -2946 188120 -2626 190638
rect -3786 187800 -3762 188120
rect -3442 187982 -2626 188120
rect -3442 187800 -2994 187982
rect -3786 187776 -3418 187800
rect -3018 187662 -2994 187800
rect -2674 187662 -2626 187982
rect -1526 190052 -1206 190640
rect -1526 189780 -1502 190052
rect -1230 189780 -1206 190052
rect -1526 187960 -1206 189780
rect -3018 187638 -2626 187662
rect -1529 187640 -1206 187960
rect -5547 187076 -5179 187100
rect -5547 186756 -5523 187076
rect -5203 186756 -5179 187076
rect -5547 186732 -5179 186756
rect -6318 185120 -5950 185144
rect -6318 184800 -6294 185120
rect -5974 184800 -5950 185120
rect -6318 184776 -5950 184800
rect -3786 185120 -3418 185144
rect -2946 185120 -2626 187638
rect -3786 184800 -3762 185120
rect -3442 184982 -2626 185120
rect -3442 184800 -2994 184982
rect -3786 184776 -3418 184800
rect -3018 184662 -2994 184800
rect -2674 184662 -2626 184982
rect -1526 187052 -1206 187640
rect -1526 186780 -1502 187052
rect -1230 186780 -1206 187052
rect -1526 184960 -1206 186780
rect -3018 184638 -2626 184662
rect -1529 184640 -1206 184960
rect -5547 184076 -5179 184100
rect -5547 183756 -5523 184076
rect -5203 183756 -5179 184076
rect -5547 183732 -5179 183756
rect -6318 182120 -5950 182144
rect -6318 181800 -6294 182120
rect -5974 181800 -5950 182120
rect -6318 181776 -5950 181800
rect -3786 182120 -3418 182144
rect -2946 182120 -2626 184638
rect -3786 181800 -3762 182120
rect -3442 181982 -2626 182120
rect -3442 181800 -2994 181982
rect -3786 181776 -3418 181800
rect -3018 181662 -2994 181800
rect -2674 181662 -2626 181982
rect -1526 184052 -1206 184640
rect -1526 183780 -1502 184052
rect -1230 183780 -1206 184052
rect -1526 181960 -1206 183780
rect -3018 181638 -2626 181662
rect -1529 181640 -1206 181960
rect -5547 181076 -5179 181100
rect -5547 180756 -5523 181076
rect -5203 180756 -5179 181076
rect -5547 180732 -5179 180756
rect -6318 179120 -5950 179144
rect -6318 178800 -6294 179120
rect -5974 178800 -5950 179120
rect -6318 178776 -5950 178800
rect -3786 179120 -3418 179144
rect -2946 179120 -2626 181638
rect -3786 178800 -3762 179120
rect -3442 178982 -2626 179120
rect -3442 178800 -2994 178982
rect -3786 178776 -3418 178800
rect -3018 178662 -2994 178800
rect -2674 178662 -2626 178982
rect -1526 181052 -1206 181640
rect -1526 180780 -1502 181052
rect -1230 180780 -1206 181052
rect -1526 178960 -1206 180780
rect -3018 178638 -2626 178662
rect -1529 178640 -1206 178960
rect -5547 178076 -5179 178100
rect -5547 177756 -5523 178076
rect -5203 177756 -5179 178076
rect -5547 177732 -5179 177756
rect -6318 176120 -5950 176144
rect -6318 175800 -6294 176120
rect -5974 175800 -5950 176120
rect -6318 175776 -5950 175800
rect -3786 176120 -3418 176144
rect -2946 176120 -2626 178638
rect -3786 175800 -3762 176120
rect -3442 175982 -2626 176120
rect -3442 175800 -2994 175982
rect -3786 175776 -3418 175800
rect -3018 175662 -2994 175800
rect -2674 175662 -2626 175982
rect -1526 178052 -1206 178640
rect -1526 177780 -1502 178052
rect -1230 177780 -1206 178052
rect -1526 175960 -1206 177780
rect -3018 175638 -2626 175662
rect -1529 175640 -1206 175960
rect -5547 175076 -5179 175100
rect -5547 174756 -5523 175076
rect -5203 174756 -5179 175076
rect -5547 174732 -5179 174756
rect -6318 173120 -5950 173144
rect -6318 172800 -6294 173120
rect -5974 172800 -5950 173120
rect -6318 172776 -5950 172800
rect -3786 173120 -3418 173144
rect -2946 173120 -2626 175638
rect -3786 172800 -3762 173120
rect -3442 172982 -2626 173120
rect -3442 172800 -2994 172982
rect -3786 172776 -3418 172800
rect -3018 172662 -2994 172800
rect -2674 172662 -2626 172982
rect -1526 175052 -1206 175640
rect -1526 174780 -1502 175052
rect -1230 174780 -1206 175052
rect -1526 172960 -1206 174780
rect -3018 172638 -2626 172662
rect -1529 172640 -1206 172960
rect -5547 172076 -5179 172100
rect -5547 171756 -5523 172076
rect -5203 171756 -5179 172076
rect -5547 171732 -5179 171756
rect -6318 170120 -5950 170144
rect -6318 169800 -6294 170120
rect -5974 169800 -5950 170120
rect -6318 169776 -5950 169800
rect -3786 170120 -3418 170144
rect -2946 170120 -2626 172638
rect -3786 169800 -3762 170120
rect -3442 169982 -2626 170120
rect -3442 169800 -2994 169982
rect -3786 169776 -3418 169800
rect -3018 169662 -2994 169800
rect -2674 169662 -2626 169982
rect -1526 172052 -1206 172640
rect -1526 171780 -1502 172052
rect -1230 171780 -1206 172052
rect -1526 169960 -1206 171780
rect -3018 169638 -2626 169662
rect -1529 169640 -1206 169960
rect -5547 169076 -5179 169100
rect -5547 168756 -5523 169076
rect -5203 168756 -5179 169076
rect -5547 168732 -5179 168756
rect -6318 167120 -5950 167144
rect -6318 166800 -6294 167120
rect -5974 166800 -5950 167120
rect -6318 166776 -5950 166800
rect -3786 167120 -3418 167144
rect -2946 167120 -2626 169638
rect -3786 166800 -3762 167120
rect -3442 166982 -2626 167120
rect -3442 166800 -2994 166982
rect -3786 166776 -3418 166800
rect -3018 166662 -2994 166800
rect -2674 166662 -2626 166982
rect -1526 169052 -1206 169640
rect -1526 168780 -1502 169052
rect -1230 168780 -1206 169052
rect -1526 166960 -1206 168780
rect -3018 166638 -2626 166662
rect -1529 166640 -1206 166960
rect -5547 166076 -5179 166100
rect -5547 165756 -5523 166076
rect -5203 165756 -5179 166076
rect -5547 165732 -5179 165756
rect -6318 164120 -5950 164144
rect -6318 163800 -6294 164120
rect -5974 163800 -5950 164120
rect -6318 163776 -5950 163800
rect -3786 164120 -3418 164144
rect -2946 164120 -2626 166638
rect -3786 163800 -3762 164120
rect -3442 163982 -2626 164120
rect -3442 163800 -2994 163982
rect -3786 163776 -3418 163800
rect -3018 163662 -2994 163800
rect -2674 163662 -2626 163982
rect -1526 166052 -1206 166640
rect -1526 165780 -1502 166052
rect -1230 165780 -1206 166052
rect -1526 163960 -1206 165780
rect -3018 163638 -2626 163662
rect -1529 163640 -1206 163960
rect -5547 163076 -5179 163100
rect -5547 162756 -5523 163076
rect -5203 162756 -5179 163076
rect -5547 162732 -5179 162756
rect -6318 161120 -5950 161144
rect -6318 160800 -6294 161120
rect -5974 160800 -5950 161120
rect -6318 160776 -5950 160800
rect -3786 161120 -3418 161144
rect -2946 161120 -2626 163638
rect -3786 160800 -3762 161120
rect -3442 160982 -2626 161120
rect -3442 160800 -2994 160982
rect -3786 160776 -3418 160800
rect -3018 160662 -2994 160800
rect -2674 160662 -2626 160982
rect -1526 163052 -1206 163640
rect -1526 162780 -1502 163052
rect -1230 162780 -1206 163052
rect -1526 160960 -1206 162780
rect -3018 160638 -2626 160662
rect -1529 160640 -1206 160960
rect -5547 160076 -5179 160100
rect -5547 159756 -5523 160076
rect -5203 159756 -5179 160076
rect -5547 159732 -5179 159756
rect -6318 158120 -5950 158144
rect -6318 157800 -6294 158120
rect -5974 157800 -5950 158120
rect -6318 157776 -5950 157800
rect -3786 158120 -3418 158144
rect -2946 158120 -2626 160638
rect -3786 157800 -3762 158120
rect -3442 157982 -2626 158120
rect -3442 157800 -2994 157982
rect -3786 157776 -3418 157800
rect -3018 157662 -2994 157800
rect -2674 157662 -2626 157982
rect -1526 160052 -1206 160640
rect -1526 159780 -1502 160052
rect -1230 159780 -1206 160052
rect -1526 157960 -1206 159780
rect -3018 157638 -2626 157662
rect -1529 157640 -1206 157960
rect -5547 157076 -5179 157100
rect -5547 156756 -5523 157076
rect -5203 156756 -5179 157076
rect -5547 156732 -5179 156756
rect -6318 155120 -5950 155144
rect -6318 154800 -6294 155120
rect -5974 154800 -5950 155120
rect -6318 154776 -5950 154800
rect -3786 155120 -3418 155144
rect -2946 155120 -2626 157638
rect -3786 154800 -3762 155120
rect -3442 154982 -2626 155120
rect -3442 154800 -2994 154982
rect -3786 154776 -3418 154800
rect -3018 154662 -2994 154800
rect -2674 154662 -2626 154982
rect -1526 157052 -1206 157640
rect -1526 156780 -1502 157052
rect -1230 156780 -1206 157052
rect -1526 154960 -1206 156780
rect -3018 154638 -2626 154662
rect -1529 154640 -1206 154960
rect -5547 154076 -5179 154100
rect -5547 153756 -5523 154076
rect -5203 153756 -5179 154076
rect -5547 153732 -5179 153756
rect -6318 152120 -5950 152144
rect -6318 151800 -6294 152120
rect -5974 151800 -5950 152120
rect -6318 151776 -5950 151800
rect -3786 152120 -3418 152144
rect -2946 152120 -2626 154638
rect -3786 151800 -3762 152120
rect -3442 151982 -2626 152120
rect -3442 151800 -2994 151982
rect -3786 151776 -3418 151800
rect -3018 151662 -2994 151800
rect -2674 151662 -2626 151982
rect -1526 154052 -1206 154640
rect -1526 153780 -1502 154052
rect -1230 153780 -1206 154052
rect -1526 151960 -1206 153780
rect -3018 151638 -2626 151662
rect -1529 151640 -1206 151960
rect -5547 151076 -5179 151100
rect -5547 150756 -5523 151076
rect -5203 150756 -5179 151076
rect -5547 150732 -5179 150756
rect -6318 149120 -5950 149144
rect -6318 148800 -6294 149120
rect -5974 148800 -5950 149120
rect -6318 148776 -5950 148800
rect -3786 149120 -3418 149144
rect -2946 149120 -2626 151638
rect -3786 148800 -3762 149120
rect -3442 148982 -2626 149120
rect -3442 148800 -2994 148982
rect -3786 148776 -3418 148800
rect -3018 148662 -2994 148800
rect -2674 148662 -2626 148982
rect -1526 151052 -1206 151640
rect -1526 150780 -1502 151052
rect -1230 150780 -1206 151052
rect -1526 148960 -1206 150780
rect -3018 148638 -2626 148662
rect -1529 148640 -1206 148960
rect -5547 148076 -5179 148100
rect -5547 147756 -5523 148076
rect -5203 147756 -5179 148076
rect -5547 147732 -5179 147756
rect -6318 146120 -5950 146144
rect -6318 145800 -6294 146120
rect -5974 145800 -5950 146120
rect -6318 145776 -5950 145800
rect -3786 146120 -3418 146144
rect -2946 146120 -2626 148638
rect -3786 145800 -3762 146120
rect -3442 145982 -2626 146120
rect -3442 145800 -2994 145982
rect -3786 145776 -3418 145800
rect -3018 145662 -2994 145800
rect -2674 145662 -2626 145982
rect -1526 148052 -1206 148640
rect -1526 147780 -1502 148052
rect -1230 147780 -1206 148052
rect -1526 145960 -1206 147780
rect -3018 145638 -2626 145662
rect -1529 145640 -1206 145960
rect -5547 145076 -5179 145100
rect -5547 144756 -5523 145076
rect -5203 144756 -5179 145076
rect -5547 144732 -5179 144756
rect -6318 143120 -5950 143144
rect -6318 142800 -6294 143120
rect -5974 142800 -5950 143120
rect -6318 142776 -5950 142800
rect -3786 143120 -3418 143144
rect -2946 143120 -2626 145638
rect -3786 142800 -3762 143120
rect -3442 142982 -2626 143120
rect -3442 142800 -2994 142982
rect -3786 142776 -3418 142800
rect -3018 142662 -2994 142800
rect -2674 142662 -2626 142982
rect -1526 145052 -1206 145640
rect -1526 144780 -1502 145052
rect -1230 144780 -1206 145052
rect -1526 142960 -1206 144780
rect -3018 142638 -2626 142662
rect -1529 142640 -1206 142960
rect -5547 142076 -5179 142100
rect -5547 141756 -5523 142076
rect -5203 141756 -5179 142076
rect -5547 141732 -5179 141756
rect -6318 140120 -5950 140144
rect -6318 139800 -6294 140120
rect -5974 139800 -5950 140120
rect -6318 139776 -5950 139800
rect -3786 140120 -3418 140144
rect -2946 140120 -2626 142638
rect -3786 139800 -3762 140120
rect -3442 139982 -2626 140120
rect -3442 139800 -2994 139982
rect -3786 139776 -3418 139800
rect -3018 139662 -2994 139800
rect -2674 139662 -2626 139982
rect -1526 142052 -1206 142640
rect -1526 141780 -1502 142052
rect -1230 141780 -1206 142052
rect -1526 139960 -1206 141780
rect -3018 139638 -2626 139662
rect -1529 139640 -1206 139960
rect -5547 139076 -5179 139100
rect -5547 138756 -5523 139076
rect -5203 138756 -5179 139076
rect -5547 138732 -5179 138756
rect -6318 137120 -5950 137144
rect -6318 136800 -6294 137120
rect -5974 136800 -5950 137120
rect -6318 136776 -5950 136800
rect -3786 137120 -3418 137144
rect -2946 137120 -2626 139638
rect -3786 136800 -3762 137120
rect -3442 136982 -2626 137120
rect -3442 136800 -2994 136982
rect -3786 136776 -3418 136800
rect -3018 136662 -2994 136800
rect -2674 136662 -2626 136982
rect -1526 139052 -1206 139640
rect -1526 138780 -1502 139052
rect -1230 138780 -1206 139052
rect -1526 136960 -1206 138780
rect -3018 136638 -2626 136662
rect -1529 136640 -1206 136960
rect -5547 136076 -5179 136100
rect -5547 135756 -5523 136076
rect -5203 135756 -5179 136076
rect -5547 135732 -5179 135756
rect -6318 134120 -5950 134144
rect -6318 133800 -6294 134120
rect -5974 133800 -5950 134120
rect -6318 133776 -5950 133800
rect -3786 134120 -3418 134144
rect -2946 134120 -2626 136638
rect -3786 133800 -3762 134120
rect -3442 133982 -2626 134120
rect -3442 133800 -2994 133982
rect -3786 133776 -3418 133800
rect -3018 133662 -2994 133800
rect -2674 133662 -2626 133982
rect -1526 136052 -1206 136640
rect -1526 135780 -1502 136052
rect -1230 135780 -1206 136052
rect -1526 133960 -1206 135780
rect -3018 133638 -2626 133662
rect -1529 133640 -1206 133960
rect -5547 133076 -5179 133100
rect -5547 132756 -5523 133076
rect -5203 132756 -5179 133076
rect -5547 132732 -5179 132756
rect -6318 131120 -5950 131144
rect -6318 130800 -6294 131120
rect -5974 130800 -5950 131120
rect -6318 130776 -5950 130800
rect -3786 131120 -3418 131144
rect -2946 131120 -2626 133638
rect -3786 130800 -3762 131120
rect -3442 130982 -2626 131120
rect -3442 130800 -2994 130982
rect -3786 130776 -3418 130800
rect -3018 130662 -2994 130800
rect -2674 130662 -2626 130982
rect -1526 133052 -1206 133640
rect -1526 132780 -1502 133052
rect -1230 132780 -1206 133052
rect -1526 130960 -1206 132780
rect -3018 130638 -2626 130662
rect -1529 130640 -1206 130960
rect -5547 130076 -5179 130100
rect -5547 129756 -5523 130076
rect -5203 129756 -5179 130076
rect -5547 129732 -5179 129756
rect -6318 128120 -5950 128144
rect -6318 127800 -6294 128120
rect -5974 127800 -5950 128120
rect -6318 127776 -5950 127800
rect -3786 128120 -3418 128144
rect -2946 128120 -2626 130638
rect -3786 127800 -3762 128120
rect -3442 127982 -2626 128120
rect -3442 127800 -2994 127982
rect -3786 127776 -3418 127800
rect -3018 127662 -2994 127800
rect -2674 127662 -2626 127982
rect -1526 130052 -1206 130640
rect -1526 129780 -1502 130052
rect -1230 129780 -1206 130052
rect -1526 127960 -1206 129780
rect -3018 127638 -2626 127662
rect -1529 127640 -1206 127960
rect -5547 127076 -5179 127100
rect -5547 126756 -5523 127076
rect -5203 126756 -5179 127076
rect -5547 126732 -5179 126756
rect -6318 125120 -5950 125144
rect -6318 124800 -6294 125120
rect -5974 124800 -5950 125120
rect -6318 124776 -5950 124800
rect -3786 125120 -3418 125144
rect -2946 125120 -2626 127638
rect -3786 124800 -3762 125120
rect -3442 124982 -2626 125120
rect -3442 124800 -2994 124982
rect -3786 124776 -3418 124800
rect -3018 124662 -2994 124800
rect -2674 124662 -2626 124982
rect -1526 127052 -1206 127640
rect -1526 126780 -1502 127052
rect -1230 126780 -1206 127052
rect -1526 124960 -1206 126780
rect -3018 124638 -2626 124662
rect -1529 124640 -1206 124960
rect -5547 124076 -5179 124100
rect -5547 123756 -5523 124076
rect -5203 123756 -5179 124076
rect -5547 123732 -5179 123756
rect -6318 122120 -5950 122144
rect -6318 121800 -6294 122120
rect -5974 121800 -5950 122120
rect -6318 121776 -5950 121800
rect -3786 122120 -3418 122144
rect -2946 122120 -2626 124638
rect -3786 121800 -3762 122120
rect -3442 121982 -2626 122120
rect -3442 121800 -2994 121982
rect -3786 121776 -3418 121800
rect -3018 121662 -2994 121800
rect -2674 121662 -2626 121982
rect -1526 124052 -1206 124640
rect -1526 123780 -1502 124052
rect -1230 123780 -1206 124052
rect -1526 121960 -1206 123780
rect -3018 121638 -2626 121662
rect -1529 121640 -1206 121960
rect -5547 121076 -5179 121100
rect -5547 120756 -5523 121076
rect -5203 120756 -5179 121076
rect -5547 120732 -5179 120756
rect -6318 119120 -5950 119144
rect -6318 118800 -6294 119120
rect -5974 118800 -5950 119120
rect -6318 118776 -5950 118800
rect -3786 119120 -3418 119144
rect -2946 119120 -2626 121638
rect -3786 118800 -3762 119120
rect -3442 118982 -2626 119120
rect -3442 118800 -2994 118982
rect -3786 118776 -3418 118800
rect -3018 118662 -2994 118800
rect -2674 118662 -2626 118982
rect -1526 121052 -1206 121640
rect -1526 120780 -1502 121052
rect -1230 120780 -1206 121052
rect -1526 118960 -1206 120780
rect -3018 118638 -2626 118662
rect -1529 118640 -1206 118960
rect -5547 118076 -5179 118100
rect -5547 117756 -5523 118076
rect -5203 117756 -5179 118076
rect -5547 117732 -5179 117756
rect -6318 116120 -5950 116144
rect -6318 115800 -6294 116120
rect -5974 115800 -5950 116120
rect -6318 115776 -5950 115800
rect -3786 116120 -3418 116144
rect -2946 116120 -2626 118638
rect -3786 115800 -3762 116120
rect -3442 115982 -2626 116120
rect -3442 115800 -2994 115982
rect -3786 115776 -3418 115800
rect -3018 115662 -2994 115800
rect -2674 115662 -2626 115982
rect -1526 118052 -1206 118640
rect -1526 117780 -1502 118052
rect -1230 117780 -1206 118052
rect -1526 115960 -1206 117780
rect -3018 115638 -2626 115662
rect -1529 115640 -1206 115960
rect -5547 115076 -5179 115100
rect -5547 114756 -5523 115076
rect -5203 114756 -5179 115076
rect -5547 114732 -5179 114756
rect -6318 113120 -5950 113144
rect -6318 112800 -6294 113120
rect -5974 112800 -5950 113120
rect -6318 112776 -5950 112800
rect -3786 113120 -3418 113144
rect -2946 113120 -2626 115638
rect -3786 112800 -3762 113120
rect -3442 112982 -2626 113120
rect -3442 112800 -2994 112982
rect -3786 112776 -3418 112800
rect -3018 112662 -2994 112800
rect -2674 112662 -2626 112982
rect -1526 115052 -1206 115640
rect -1526 114780 -1502 115052
rect -1230 114780 -1206 115052
rect -1526 112960 -1206 114780
rect -3018 112638 -2626 112662
rect -1529 112640 -1206 112960
rect -5547 112076 -5179 112100
rect -5547 111756 -5523 112076
rect -5203 111756 -5179 112076
rect -5547 111732 -5179 111756
rect -6318 110120 -5950 110144
rect -6318 109800 -6294 110120
rect -5974 109800 -5950 110120
rect -6318 109776 -5950 109800
rect -3786 110120 -3418 110144
rect -2946 110120 -2626 112638
rect -3786 109800 -3762 110120
rect -3442 109982 -2626 110120
rect -3442 109800 -2994 109982
rect -3786 109776 -3418 109800
rect -3018 109662 -2994 109800
rect -2674 109662 -2626 109982
rect -1526 112052 -1206 112640
rect -1526 111780 -1502 112052
rect -1230 111780 -1206 112052
rect -1526 109960 -1206 111780
rect -3018 109638 -2626 109662
rect -1529 109640 -1206 109960
rect -5547 109076 -5179 109100
rect -5547 108756 -5523 109076
rect -5203 108756 -5179 109076
rect -5547 108732 -5179 108756
rect -6318 107120 -5950 107144
rect -6318 106800 -6294 107120
rect -5974 106800 -5950 107120
rect -6318 106776 -5950 106800
rect -3786 107120 -3418 107144
rect -2946 107120 -2626 109638
rect -3786 106800 -3762 107120
rect -3442 106982 -2626 107120
rect -3442 106800 -2994 106982
rect -3786 106776 -3418 106800
rect -3018 106662 -2994 106800
rect -2674 106662 -2626 106982
rect -1526 109052 -1206 109640
rect -1526 108780 -1502 109052
rect -1230 108780 -1206 109052
rect -1526 106960 -1206 108780
rect -3018 106638 -2626 106662
rect -1529 106640 -1206 106960
rect -5547 106076 -5179 106100
rect -5547 105756 -5523 106076
rect -5203 105756 -5179 106076
rect -5547 105732 -5179 105756
rect -6318 104120 -5950 104144
rect -6318 103800 -6294 104120
rect -5974 103800 -5950 104120
rect -6318 103776 -5950 103800
rect -3786 104120 -3418 104144
rect -2946 104120 -2626 106638
rect -3786 103800 -3762 104120
rect -3442 103982 -2626 104120
rect -3442 103800 -2994 103982
rect -3786 103776 -3418 103800
rect -3018 103662 -2994 103800
rect -2674 103662 -2626 103982
rect -1526 106052 -1206 106640
rect -1526 105780 -1502 106052
rect -1230 105780 -1206 106052
rect -1526 103960 -1206 105780
rect -3018 103638 -2626 103662
rect -1529 103640 -1206 103960
rect -5547 103076 -5179 103100
rect -5547 102756 -5523 103076
rect -5203 102756 -5179 103076
rect -5547 102732 -5179 102756
rect -6318 101120 -5950 101144
rect -6318 100800 -6294 101120
rect -5974 100800 -5950 101120
rect -6318 100776 -5950 100800
rect -3786 101120 -3418 101144
rect -2946 101120 -2626 103638
rect -3786 100800 -3762 101120
rect -3442 100982 -2626 101120
rect -3442 100800 -2994 100982
rect -3786 100776 -3418 100800
rect -3018 100662 -2994 100800
rect -2674 100662 -2626 100982
rect -1526 103052 -1206 103640
rect -1526 102780 -1502 103052
rect -1230 102780 -1206 103052
rect -1526 100960 -1206 102780
rect -3018 100638 -2626 100662
rect -1529 100640 -1206 100960
rect -5547 100076 -5179 100100
rect -5547 99756 -5523 100076
rect -5203 99756 -5179 100076
rect -5547 99732 -5179 99756
rect -6318 98120 -5950 98144
rect -6318 97800 -6294 98120
rect -5974 97800 -5950 98120
rect -6318 97776 -5950 97800
rect -3786 98120 -3418 98144
rect -2946 98120 -2626 100638
rect -3786 97800 -3762 98120
rect -3442 97982 -2626 98120
rect -3442 97800 -2994 97982
rect -3786 97776 -3418 97800
rect -3018 97662 -2994 97800
rect -2674 97662 -2626 97982
rect -1526 100052 -1206 100640
rect -1526 99780 -1502 100052
rect -1230 99780 -1206 100052
rect -1526 97960 -1206 99780
rect -3018 97638 -2626 97662
rect -1529 97640 -1206 97960
rect -5547 97076 -5179 97100
rect -5547 96756 -5523 97076
rect -5203 96756 -5179 97076
rect -5547 96732 -5179 96756
rect -6318 95120 -5950 95144
rect -6318 94800 -6294 95120
rect -5974 94800 -5950 95120
rect -6318 94776 -5950 94800
rect -3786 95120 -3418 95144
rect -2946 95120 -2626 97638
rect -3786 94800 -3762 95120
rect -3442 94982 -2626 95120
rect -3442 94800 -2994 94982
rect -3786 94776 -3418 94800
rect -3018 94662 -2994 94800
rect -2674 94662 -2626 94982
rect -1526 97052 -1206 97640
rect -1526 96780 -1502 97052
rect -1230 96780 -1206 97052
rect -1526 94960 -1206 96780
rect -3018 94638 -2626 94662
rect -1529 94640 -1206 94960
rect -6318 92120 -5950 92144
rect -6318 91800 -6294 92120
rect -5974 91800 -5950 92120
rect -6318 91776 -5950 91800
rect -3786 92120 -3418 92144
rect -2946 92120 -2626 94638
rect -3786 91800 -3762 92120
rect -3442 91982 -2626 92120
rect -3442 91800 -2994 91982
rect -3786 91776 -3418 91800
rect -3018 91662 -2994 91800
rect -2674 91662 -2626 91982
rect -1526 91960 -1206 94640
rect -3018 91638 -2626 91662
rect -1529 91640 -1206 91960
rect -5547 91076 -5179 91100
rect -5547 90756 -5523 91076
rect -5203 90756 -5179 91076
rect -5547 90732 -5179 90756
rect -6318 89120 -5950 89144
rect -6318 88800 -6294 89120
rect -5974 88800 -5950 89120
rect -6318 88776 -5950 88800
rect -3786 89120 -3418 89144
rect -2946 89120 -2626 91638
rect -3786 88800 -3762 89120
rect -3442 88982 -2626 89120
rect -3442 88800 -2994 88982
rect -3786 88776 -3418 88800
rect -3018 88662 -2994 88800
rect -2674 88662 -2626 88982
rect -1526 91052 -1206 91640
rect -1526 90780 -1502 91052
rect -1230 90780 -1206 91052
rect -1526 88960 -1206 90780
rect -3018 88638 -2626 88662
rect -1529 88640 -1206 88960
rect -5547 88076 -5179 88100
rect -5547 87756 -5523 88076
rect -5203 87756 -5179 88076
rect -5547 87732 -5179 87756
rect -6318 86120 -5950 86144
rect -6318 85800 -6294 86120
rect -5974 85800 -5950 86120
rect -6318 85776 -5950 85800
rect -3786 86120 -3418 86144
rect -2946 86120 -2626 88638
rect -3786 85800 -3762 86120
rect -3442 85982 -2626 86120
rect -3442 85800 -2994 85982
rect -3786 85776 -3418 85800
rect -3018 85662 -2994 85800
rect -2674 85662 -2626 85982
rect -1526 88052 -1206 88640
rect -1526 87780 -1502 88052
rect -1230 87780 -1206 88052
rect -1526 85960 -1206 87780
rect -3018 85638 -2626 85662
rect -1529 85640 -1206 85960
rect -5547 85076 -5179 85100
rect -5547 84756 -5523 85076
rect -5203 84756 -5179 85076
rect -5547 84732 -5179 84756
rect -6318 83120 -5950 83144
rect -6318 82800 -6294 83120
rect -5974 82800 -5950 83120
rect -6318 82776 -5950 82800
rect -3786 83120 -3418 83144
rect -2946 83120 -2626 85638
rect -3786 82800 -3762 83120
rect -3442 82982 -2626 83120
rect -3442 82800 -2994 82982
rect -3786 82776 -3418 82800
rect -3018 82662 -2994 82800
rect -2674 82662 -2626 82982
rect -1526 85052 -1206 85640
rect -1526 84780 -1502 85052
rect -1230 84780 -1206 85052
rect -1526 82960 -1206 84780
rect -3018 82638 -2626 82662
rect -1529 82640 -1206 82960
rect -5547 82076 -5179 82100
rect -5547 81756 -5523 82076
rect -5203 81756 -5179 82076
rect -5547 81732 -5179 81756
rect -6318 80120 -5950 80144
rect -6318 79800 -6294 80120
rect -5974 79800 -5950 80120
rect -6318 79776 -5950 79800
rect -3786 80120 -3418 80144
rect -2946 80120 -2626 82638
rect -3786 79800 -3762 80120
rect -3442 79982 -2626 80120
rect -3442 79800 -2994 79982
rect -3786 79776 -3418 79800
rect -3018 79662 -2994 79800
rect -2674 79662 -2626 79982
rect -1526 82052 -1206 82640
rect -1526 81780 -1502 82052
rect -1230 81780 -1206 82052
rect -1526 79960 -1206 81780
rect -3018 79638 -2626 79662
rect -1529 79640 -1206 79960
rect -5547 79076 -5179 79100
rect -5547 78756 -5523 79076
rect -5203 78756 -5179 79076
rect -5547 78732 -5179 78756
rect -6318 77120 -5950 77144
rect -6318 76800 -6294 77120
rect -5974 76800 -5950 77120
rect -6318 76776 -5950 76800
rect -3786 77120 -3418 77144
rect -2946 77120 -2626 79638
rect -3786 76800 -3762 77120
rect -3442 76982 -2626 77120
rect -3442 76800 -2994 76982
rect -3786 76776 -3418 76800
rect -3018 76662 -2994 76800
rect -2674 76662 -2626 76982
rect -1526 79052 -1206 79640
rect -1526 78780 -1502 79052
rect -1230 78780 -1206 79052
rect -1526 76960 -1206 78780
rect -3018 76638 -2626 76662
rect -1529 76640 -1206 76960
rect -5547 76076 -5179 76100
rect -5547 75756 -5523 76076
rect -5203 75756 -5179 76076
rect -5547 75732 -5179 75756
rect -6318 74120 -5950 74144
rect -6318 73800 -6294 74120
rect -5974 73800 -5950 74120
rect -6318 73776 -5950 73800
rect -3786 74120 -3418 74144
rect -2946 74120 -2626 76638
rect -3786 73800 -3762 74120
rect -3442 73982 -2626 74120
rect -3442 73800 -2994 73982
rect -3786 73776 -3418 73800
rect -3018 73662 -2994 73800
rect -2674 73662 -2626 73982
rect -1526 76052 -1206 76640
rect -1526 75780 -1502 76052
rect -1230 75780 -1206 76052
rect -1526 73960 -1206 75780
rect -3018 73638 -2626 73662
rect -1529 73640 -1206 73960
rect -5547 73076 -5179 73100
rect -5547 72756 -5523 73076
rect -5203 72756 -5179 73076
rect -5547 72732 -5179 72756
rect -6318 71120 -5950 71144
rect -6318 70800 -6294 71120
rect -5974 70800 -5950 71120
rect -6318 70776 -5950 70800
rect -3786 71120 -3418 71144
rect -2946 71120 -2626 73638
rect -3786 70800 -3762 71120
rect -3442 70982 -2626 71120
rect -3442 70800 -2994 70982
rect -3786 70776 -3418 70800
rect -3018 70662 -2994 70800
rect -2674 70662 -2626 70982
rect -1526 73052 -1206 73640
rect -1526 72780 -1502 73052
rect -1230 72780 -1206 73052
rect -1526 70960 -1206 72780
rect -3018 70638 -2626 70662
rect -1529 70640 -1206 70960
rect -5547 70076 -5179 70100
rect -5547 69756 -5523 70076
rect -5203 69756 -5179 70076
rect -5547 69732 -5179 69756
rect -6318 68120 -5950 68144
rect -6318 67800 -6294 68120
rect -5974 67800 -5950 68120
rect -6318 67776 -5950 67800
rect -3786 68120 -3418 68144
rect -2946 68120 -2626 70638
rect -3786 67800 -3762 68120
rect -3442 67982 -2626 68120
rect -3442 67800 -2994 67982
rect -3786 67776 -3418 67800
rect -3018 67662 -2994 67800
rect -2674 67662 -2626 67982
rect -1526 70052 -1206 70640
rect -1526 69780 -1502 70052
rect -1230 69780 -1206 70052
rect -1526 67960 -1206 69780
rect -3018 67638 -2626 67662
rect -1529 67640 -1206 67960
rect -5547 67076 -5179 67100
rect -5547 66756 -5523 67076
rect -5203 66756 -5179 67076
rect -5547 66732 -5179 66756
rect -6318 65120 -5950 65144
rect -6318 64800 -6294 65120
rect -5974 64800 -5950 65120
rect -6318 64776 -5950 64800
rect -3786 65120 -3418 65144
rect -2946 65120 -2626 67638
rect -3786 64800 -3762 65120
rect -3442 64982 -2626 65120
rect -3442 64800 -2994 64982
rect -3786 64776 -3418 64800
rect -3018 64662 -2994 64800
rect -2674 64662 -2626 64982
rect -1526 67052 -1206 67640
rect -1526 66780 -1502 67052
rect -1230 66780 -1206 67052
rect -1526 64960 -1206 66780
rect -3018 64638 -2626 64662
rect -1529 64640 -1206 64960
rect -5547 64076 -5179 64100
rect -5547 63756 -5523 64076
rect -5203 63756 -5179 64076
rect -5547 63732 -5179 63756
rect -6318 62120 -5950 62144
rect -6318 61800 -6294 62120
rect -5974 61800 -5950 62120
rect -6318 61776 -5950 61800
rect -3786 62120 -3418 62144
rect -2946 62120 -2626 64638
rect -3786 61800 -3762 62120
rect -3442 61982 -2626 62120
rect -3442 61800 -2994 61982
rect -3786 61776 -3418 61800
rect -3018 61662 -2994 61800
rect -2674 61662 -2626 61982
rect -1526 64052 -1206 64640
rect -1526 63780 -1502 64052
rect -1230 63780 -1206 64052
rect -1526 61960 -1206 63780
rect -3018 61638 -2626 61662
rect -1529 61640 -1206 61960
rect -5547 61076 -5179 61100
rect -5547 60756 -5523 61076
rect -5203 60756 -5179 61076
rect -5547 60732 -5179 60756
rect -6318 59120 -5950 59144
rect -6318 58800 -6294 59120
rect -5974 58800 -5950 59120
rect -6318 58776 -5950 58800
rect -3786 59120 -3418 59144
rect -2946 59120 -2626 61638
rect -3786 58800 -3762 59120
rect -3442 58982 -2626 59120
rect -3442 58800 -2994 58982
rect -3786 58776 -3418 58800
rect -3018 58662 -2994 58800
rect -2674 58662 -2626 58982
rect -1526 61052 -1206 61640
rect -1526 60780 -1502 61052
rect -1230 60780 -1206 61052
rect -1526 58960 -1206 60780
rect -3018 58638 -2626 58662
rect -1529 58640 -1206 58960
rect -5547 58076 -5179 58100
rect -5547 57756 -5523 58076
rect -5203 57756 -5179 58076
rect -5547 57732 -5179 57756
rect -2946 56120 -2626 58638
rect -3120 55982 -2626 56120
rect -3120 55800 -2994 55982
rect -3018 55662 -2994 55800
rect -2674 55662 -2626 55982
rect -1526 58052 -1206 58640
rect -1526 57780 -1502 58052
rect -1230 57780 -1206 58052
rect -1526 55960 -1206 57780
rect -3018 55638 -2626 55662
rect -1529 55640 -1206 55960
rect -5547 55076 -5179 55100
rect -5547 54756 -5523 55076
rect -5203 54756 -5179 55076
rect -5547 54732 -5179 54756
rect -6318 53120 -5950 53144
rect -6318 52800 -6294 53120
rect -5974 52800 -5950 53120
rect -6318 52776 -5950 52800
rect -3786 53120 -3418 53144
rect -2946 53120 -2626 55638
rect -3786 52800 -3762 53120
rect -3442 52982 -2626 53120
rect -3442 52800 -2994 52982
rect -3786 52776 -3418 52800
rect -3018 52662 -2994 52800
rect -2674 52662 -2626 52982
rect -1526 55052 -1206 55640
rect -1526 54780 -1502 55052
rect -1230 54780 -1206 55052
rect -1526 52960 -1206 54780
rect -3018 52638 -2626 52662
rect -1529 52640 -1206 52960
rect -5547 52076 -5179 52100
rect -5547 51756 -5523 52076
rect -5203 51756 -5179 52076
rect -5547 51732 -5179 51756
rect -6318 50120 -5950 50144
rect -6318 49800 -6294 50120
rect -5974 49800 -5950 50120
rect -6318 49776 -5950 49800
rect -3786 50120 -3418 50144
rect -2946 50120 -2626 52638
rect -3786 49800 -3762 50120
rect -3442 49982 -2626 50120
rect -3442 49800 -2994 49982
rect -3786 49776 -3418 49800
rect -3018 49662 -2994 49800
rect -2674 49662 -2626 49982
rect -1526 52052 -1206 52640
rect -1526 51780 -1502 52052
rect -1230 51780 -1206 52052
rect -1526 49960 -1206 51780
rect -3018 49638 -2626 49662
rect -1529 49640 -1206 49960
rect -5547 49076 -5179 49100
rect -5547 48756 -5523 49076
rect -5203 48756 -5179 49076
rect -5547 48732 -5179 48756
rect -6318 47120 -5950 47144
rect -6318 46800 -6294 47120
rect -5974 46800 -5950 47120
rect -6318 46776 -5950 46800
rect -3786 47120 -3418 47144
rect -2946 47120 -2626 49638
rect -3786 46800 -3762 47120
rect -3442 46982 -2626 47120
rect -3442 46800 -2994 46982
rect -3786 46776 -3418 46800
rect -3018 46662 -2994 46800
rect -2674 46662 -2626 46982
rect -1526 49052 -1206 49640
rect -1526 48780 -1502 49052
rect -1230 48780 -1206 49052
rect -1526 46960 -1206 48780
rect -3018 46638 -2626 46662
rect -1529 46640 -1206 46960
rect -5547 46076 -5179 46100
rect -5547 45756 -5523 46076
rect -5203 45756 -5179 46076
rect -5547 45732 -5179 45756
rect -6318 44120 -5950 44144
rect -6318 43800 -6294 44120
rect -5974 43800 -5950 44120
rect -6318 43776 -5950 43800
rect -3786 44120 -3418 44144
rect -2946 44120 -2626 46638
rect -3786 43800 -3762 44120
rect -3442 43982 -2626 44120
rect -3442 43800 -2994 43982
rect -3786 43776 -3418 43800
rect -3018 43662 -2994 43800
rect -2674 43662 -2626 43982
rect -1526 46052 -1206 46640
rect -1526 45780 -1502 46052
rect -1230 45780 -1206 46052
rect -1526 43960 -1206 45780
rect -3018 43638 -2626 43662
rect -1529 43640 -1206 43960
rect -5547 43076 -5179 43100
rect -5547 42756 -5523 43076
rect -5203 42756 -5179 43076
rect -5547 42732 -5179 42756
rect -6318 41120 -5950 41144
rect -6318 40800 -6294 41120
rect -5974 40800 -5950 41120
rect -6318 40776 -5950 40800
rect -3786 41120 -3418 41144
rect -2946 41120 -2626 43638
rect -3786 40800 -3762 41120
rect -3442 40982 -2626 41120
rect -3442 40800 -2994 40982
rect -3786 40776 -3418 40800
rect -3018 40662 -2994 40800
rect -2674 40662 -2626 40982
rect -1526 43052 -1206 43640
rect -1526 42780 -1502 43052
rect -1230 42780 -1206 43052
rect -1526 40960 -1206 42780
rect -3018 40638 -2626 40662
rect -1529 40640 -1206 40960
rect -5547 40076 -5179 40100
rect -5547 39756 -5523 40076
rect -5203 39756 -5179 40076
rect -5547 39732 -5179 39756
rect -6318 38120 -5950 38144
rect -6318 37800 -6294 38120
rect -5974 37800 -5950 38120
rect -6318 37776 -5950 37800
rect -3786 38120 -3418 38144
rect -2946 38120 -2626 40638
rect -3786 37800 -3762 38120
rect -3442 37982 -2626 38120
rect -3442 37800 -2994 37982
rect -3786 37776 -3418 37800
rect -3018 37662 -2994 37800
rect -2674 37662 -2626 37982
rect -1526 40052 -1206 40640
rect -1526 39780 -1502 40052
rect -1230 39780 -1206 40052
rect -1526 37960 -1206 39780
rect -3018 37638 -2626 37662
rect -1529 37640 -1206 37960
rect -5547 37076 -5179 37100
rect -5547 36756 -5523 37076
rect -5203 36756 -5179 37076
rect -5547 36732 -5179 36756
rect -6318 35120 -5950 35144
rect -6318 34800 -6294 35120
rect -5974 34800 -5950 35120
rect -6318 34776 -5950 34800
rect -3786 35120 -3418 35144
rect -2946 35120 -2626 37638
rect -3786 34800 -3762 35120
rect -3442 34982 -2626 35120
rect -3442 34800 -2994 34982
rect -3786 34776 -3418 34800
rect -3018 34662 -2994 34800
rect -2674 34662 -2626 34982
rect -1526 37052 -1206 37640
rect -1526 36780 -1502 37052
rect -1230 36780 -1206 37052
rect -1526 34960 -1206 36780
rect -3018 34638 -2626 34662
rect -1529 34640 -1206 34960
rect -5547 34076 -5179 34100
rect -5547 33756 -5523 34076
rect -5203 33756 -5179 34076
rect -5547 33732 -5179 33756
rect -6318 32120 -5950 32144
rect -6318 31800 -6294 32120
rect -5974 31800 -5950 32120
rect -6318 31776 -5950 31800
rect -3786 32120 -3418 32144
rect -2946 32120 -2626 34638
rect -3786 31800 -3762 32120
rect -3442 31982 -2626 32120
rect -3442 31800 -2994 31982
rect -3786 31776 -3418 31800
rect -3018 31662 -2994 31800
rect -2674 31662 -2626 31982
rect -1526 34052 -1206 34640
rect -1526 33780 -1502 34052
rect -1230 33780 -1206 34052
rect -1526 31960 -1206 33780
rect -3018 31638 -2626 31662
rect -1529 31640 -1206 31960
rect -5547 31076 -5179 31100
rect -5547 30756 -5523 31076
rect -5203 30756 -5179 31076
rect -5547 30732 -5179 30756
rect -6318 29120 -5950 29144
rect -6318 28800 -6294 29120
rect -5974 28800 -5950 29120
rect -6318 28776 -5950 28800
rect -3786 29120 -3418 29144
rect -2946 29120 -2626 31638
rect -3786 28800 -3762 29120
rect -3442 28982 -2626 29120
rect -3442 28800 -2994 28982
rect -3786 28776 -3418 28800
rect -3018 28662 -2994 28800
rect -2674 28662 -2626 28982
rect -1526 31052 -1206 31640
rect -1526 30780 -1502 31052
rect -1230 30780 -1206 31052
rect -1526 28960 -1206 30780
rect -3018 28638 -2626 28662
rect -1529 28640 -1206 28960
rect -5547 28076 -5179 28100
rect -5547 27756 -5523 28076
rect -5203 27756 -5179 28076
rect -5547 27732 -5179 27756
rect -6318 26120 -5950 26144
rect -6318 25800 -6294 26120
rect -5974 25800 -5950 26120
rect -6318 25776 -5950 25800
rect -3786 26120 -3418 26144
rect -2946 26120 -2626 28638
rect -3786 25800 -3762 26120
rect -3442 25982 -2626 26120
rect -3442 25800 -2994 25982
rect -3786 25776 -3418 25800
rect -3018 25662 -2994 25800
rect -2674 25662 -2626 25982
rect -1526 28052 -1206 28640
rect -1526 27780 -1502 28052
rect -1230 27780 -1206 28052
rect -1526 25960 -1206 27780
rect -3018 25638 -2626 25662
rect -1529 25640 -1206 25960
rect -5547 25076 -5179 25100
rect -5547 24756 -5523 25076
rect -5203 24756 -5179 25076
rect -5547 24732 -5179 24756
rect -6318 23120 -5950 23144
rect -6318 22800 -6294 23120
rect -5974 22800 -5950 23120
rect -6318 22776 -5950 22800
rect -3786 23120 -3418 23144
rect -2946 23120 -2626 25638
rect -3786 22800 -3762 23120
rect -3442 22982 -2626 23120
rect -3442 22800 -2994 22982
rect -3786 22776 -3418 22800
rect -3018 22662 -2994 22800
rect -2674 22662 -2626 22982
rect -1526 25052 -1206 25640
rect -1526 24780 -1502 25052
rect -1230 24780 -1206 25052
rect -1526 22960 -1206 24780
rect -3018 22638 -2626 22662
rect -1529 22640 -1206 22960
rect -5547 22076 -5179 22100
rect -5547 21756 -5523 22076
rect -5203 21756 -5179 22076
rect -5547 21732 -5179 21756
rect -6318 20120 -5950 20144
rect -6318 19800 -6294 20120
rect -5974 19800 -5950 20120
rect -6318 19776 -5950 19800
rect -3786 20120 -3418 20144
rect -2946 20120 -2626 22638
rect -3786 19800 -3762 20120
rect -3442 19800 -2626 20120
rect -1526 22052 -1206 22640
rect -1526 21780 -1502 22052
rect -1230 21780 -1206 22052
rect -1526 19960 -1206 21780
rect -3786 19776 -3418 19800
rect -5547 19076 -5179 19100
rect -5547 18756 -5523 19076
rect -5203 18756 -5179 19076
rect -5547 18732 -5179 18756
rect -6415 18026 -6095 18186
rect -6439 18002 -6071 18026
rect -6439 17682 -6415 18002
rect -6095 17682 -6071 18002
rect -6439 17658 -6071 17682
rect -6415 17375 -6095 17658
rect -2946 17289 -2626 19800
rect -1529 19640 -1206 19960
rect -1526 19052 -1206 19640
rect -1526 18780 -1502 19052
rect -1230 18780 -1206 19052
rect 303926 321334 304246 324317
rect 303926 321062 303950 321334
rect 304222 321062 304246 321334
rect 303926 318334 304246 321062
rect 303926 318062 303950 318334
rect 304222 318062 304246 318334
rect 303926 315334 304246 318062
rect 303926 315062 303950 315334
rect 304222 315062 304246 315334
rect 303926 312334 304246 315062
rect 303926 312062 303950 312334
rect 304222 312062 304246 312334
rect 303926 309334 304246 312062
rect 303926 309062 303950 309334
rect 304222 309062 304246 309334
rect 303926 306334 304246 309062
rect 303926 306062 303950 306334
rect 304222 306062 304246 306334
rect 303926 303334 304246 306062
rect 303926 303062 303950 303334
rect 304222 303062 304246 303334
rect 303926 300334 304246 303062
rect 303926 300062 303950 300334
rect 304222 300062 304246 300334
rect 303926 297334 304246 300062
rect 303926 297062 303950 297334
rect 304222 297062 304246 297334
rect 303926 294334 304246 297062
rect 303926 294062 303950 294334
rect 304222 294062 304246 294334
rect 303926 291334 304246 294062
rect 303926 291062 303950 291334
rect 304222 291062 304246 291334
rect 303926 288334 304246 291062
rect 303926 288062 303950 288334
rect 304222 288062 304246 288334
rect 303926 285334 304246 288062
rect 303926 285062 303950 285334
rect 304222 285062 304246 285334
rect 303926 282334 304246 285062
rect 303926 282062 303950 282334
rect 304222 282062 304246 282334
rect 303926 279334 304246 282062
rect 303926 279062 303950 279334
rect 304222 279062 304246 279334
rect 303926 276334 304246 279062
rect 303926 276062 303950 276334
rect 304222 276062 304246 276334
rect 303926 273334 304246 276062
rect 303926 273062 303950 273334
rect 304222 273062 304246 273334
rect 303926 270334 304246 273062
rect 303926 270062 303950 270334
rect 304222 270062 304246 270334
rect 303926 267334 304246 270062
rect 303926 267062 303950 267334
rect 304222 267062 304246 267334
rect 303926 264334 304246 267062
rect 303926 264062 303950 264334
rect 304222 264062 304246 264334
rect 303926 261334 304246 264062
rect 303926 261062 303950 261334
rect 304222 261062 304246 261334
rect 303926 258334 304246 261062
rect 303926 258062 303950 258334
rect 304222 258062 304246 258334
rect 303926 255334 304246 258062
rect 303926 255062 303950 255334
rect 304222 255062 304246 255334
rect 303926 252334 304246 255062
rect 303926 252062 303950 252334
rect 304222 252062 304246 252334
rect 303926 249334 304246 252062
rect 303926 249062 303950 249334
rect 304222 249062 304246 249334
rect 303926 246334 304246 249062
rect 303926 246062 303950 246334
rect 304222 246062 304246 246334
rect 303926 243334 304246 246062
rect 303926 243062 303950 243334
rect 304222 243062 304246 243334
rect 303926 240334 304246 243062
rect 303926 240062 303950 240334
rect 304222 240062 304246 240334
rect 303926 237334 304246 240062
rect 303926 237062 303950 237334
rect 304222 237062 304246 237334
rect 303926 234334 304246 237062
rect 303926 234062 303950 234334
rect 304222 234062 304246 234334
rect 303926 231334 304246 234062
rect 303926 231062 303950 231334
rect 304222 231062 304246 231334
rect 303926 228334 304246 231062
rect 303926 228062 303950 228334
rect 304222 228062 304246 228334
rect 303926 225334 304246 228062
rect 303926 225062 303950 225334
rect 304222 225062 304246 225334
rect 303926 222334 304246 225062
rect 303926 222062 303950 222334
rect 304222 222062 304246 222334
rect 303926 219334 304246 222062
rect 303926 219062 303950 219334
rect 304222 219062 304246 219334
rect 303926 216334 304246 219062
rect 303926 216062 303950 216334
rect 304222 216062 304246 216334
rect 303926 213334 304246 216062
rect 303926 213062 303950 213334
rect 304222 213062 304246 213334
rect 303926 210334 304246 213062
rect 303926 210062 303950 210334
rect 304222 210062 304246 210334
rect 303926 207334 304246 210062
rect 303926 207062 303950 207334
rect 304222 207062 304246 207334
rect 303926 204334 304246 207062
rect 303926 204062 303950 204334
rect 304222 204062 304246 204334
rect 303926 201334 304246 204062
rect 303926 201062 303950 201334
rect 304222 201062 304246 201334
rect 303926 198334 304246 201062
rect 303926 198062 303950 198334
rect 304222 198062 304246 198334
rect 303926 195334 304246 198062
rect 303926 195062 303950 195334
rect 304222 195062 304246 195334
rect 303926 192334 304246 195062
rect 303926 192062 303950 192334
rect 304222 192062 304246 192334
rect 303926 189334 304246 192062
rect 303926 189062 303950 189334
rect 304222 189062 304246 189334
rect 303926 186334 304246 189062
rect 303926 186062 303950 186334
rect 304222 186062 304246 186334
rect 303926 183334 304246 186062
rect 303926 183062 303950 183334
rect 304222 183062 304246 183334
rect 303926 180334 304246 183062
rect 303926 180062 303950 180334
rect 304222 180062 304246 180334
rect 303926 177334 304246 180062
rect 303926 177062 303950 177334
rect 304222 177062 304246 177334
rect 303926 174334 304246 177062
rect 303926 174062 303950 174334
rect 304222 174062 304246 174334
rect 303926 171334 304246 174062
rect 303926 171062 303950 171334
rect 304222 171062 304246 171334
rect 303926 168334 304246 171062
rect 303926 168062 303950 168334
rect 304222 168062 304246 168334
rect 303926 165334 304246 168062
rect 303926 165062 303950 165334
rect 304222 165062 304246 165334
rect 303926 162334 304246 165062
rect 303926 162062 303950 162334
rect 304222 162062 304246 162334
rect 303926 159334 304246 162062
rect 303926 159062 303950 159334
rect 304222 159062 304246 159334
rect 303926 156334 304246 159062
rect 303926 156062 303950 156334
rect 304222 156062 304246 156334
rect 303926 153334 304246 156062
rect 303926 153062 303950 153334
rect 304222 153062 304246 153334
rect 303926 150334 304246 153062
rect 303926 150062 303950 150334
rect 304222 150062 304246 150334
rect 303926 147334 304246 150062
rect 303926 147062 303950 147334
rect 304222 147062 304246 147334
rect 303926 144334 304246 147062
rect 303926 144062 303950 144334
rect 304222 144062 304246 144334
rect 303926 141334 304246 144062
rect 303926 141062 303950 141334
rect 304222 141062 304246 141334
rect 303926 138334 304246 141062
rect 303926 138062 303950 138334
rect 304222 138062 304246 138334
rect 303926 135334 304246 138062
rect 303926 135062 303950 135334
rect 304222 135062 304246 135334
rect 303926 132334 304246 135062
rect 303926 132062 303950 132334
rect 304222 132062 304246 132334
rect 303926 129334 304246 132062
rect 303926 129062 303950 129334
rect 304222 129062 304246 129334
rect 303926 126334 304246 129062
rect 303926 126062 303950 126334
rect 304222 126062 304246 126334
rect 303926 123334 304246 126062
rect 303926 123062 303950 123334
rect 304222 123062 304246 123334
rect 303926 120334 304246 123062
rect 303926 120062 303950 120334
rect 304222 120062 304246 120334
rect 303926 117334 304246 120062
rect 303926 117062 303950 117334
rect 304222 117062 304246 117334
rect 303926 114334 304246 117062
rect 303926 114062 303950 114334
rect 304222 114062 304246 114334
rect 303926 111334 304246 114062
rect 303926 111062 303950 111334
rect 304222 111062 304246 111334
rect 303926 108334 304246 111062
rect 303926 108062 303950 108334
rect 304222 108062 304246 108334
rect 303926 105334 304246 108062
rect 303926 105062 303950 105334
rect 304222 105062 304246 105334
rect 303926 102334 304246 105062
rect 303926 102062 303950 102334
rect 304222 102062 304246 102334
rect 303926 99334 304246 102062
rect 303926 99062 303950 99334
rect 304222 99062 304246 99334
rect 303926 96334 304246 99062
rect 303926 96062 303950 96334
rect 304222 96062 304246 96334
rect 303926 93334 304246 96062
rect 303926 93062 303950 93334
rect 304222 93062 304246 93334
rect 303926 90334 304246 93062
rect 303926 90062 303950 90334
rect 304222 90062 304246 90334
rect 303926 87334 304246 90062
rect 303926 87062 303950 87334
rect 304222 87062 304246 87334
rect 303926 84334 304246 87062
rect 303926 84062 303950 84334
rect 304222 84062 304246 84334
rect 303926 81334 304246 84062
rect 303926 81062 303950 81334
rect 304222 81062 304246 81334
rect 303926 78334 304246 81062
rect 303926 78062 303950 78334
rect 304222 78062 304246 78334
rect 303926 75334 304246 78062
rect 303926 75062 303950 75334
rect 304222 75062 304246 75334
rect 303926 72334 304246 75062
rect 303926 72062 303950 72334
rect 304222 72062 304246 72334
rect 303926 69334 304246 72062
rect 303926 69062 303950 69334
rect 304222 69062 304246 69334
rect 303926 66334 304246 69062
rect 303926 66062 303950 66334
rect 304222 66062 304246 66334
rect 303926 63334 304246 66062
rect 303926 63062 303950 63334
rect 304222 63062 304246 63334
rect 303926 60334 304246 63062
rect 303926 60062 303950 60334
rect 304222 60062 304246 60334
rect 303926 57334 304246 60062
rect 303926 57062 303950 57334
rect 304222 57062 304246 57334
rect 303926 54334 304246 57062
rect 303926 54062 303950 54334
rect 304222 54062 304246 54334
rect 303926 51334 304246 54062
rect 303926 51062 303950 51334
rect 304222 51062 304246 51334
rect 303926 48334 304246 51062
rect 303926 48062 303950 48334
rect 304222 48062 304246 48334
rect 303926 45334 304246 48062
rect 303926 45062 303950 45334
rect 304222 45062 304246 45334
rect 303926 42334 304246 45062
rect 303926 42062 303950 42334
rect 304222 42062 304246 42334
rect 303926 39334 304246 42062
rect 303926 39062 303950 39334
rect 304222 39062 304246 39334
rect 303926 36334 304246 39062
rect 303926 36062 303950 36334
rect 304222 36062 304246 36334
rect 303926 33334 304246 36062
rect 303926 33062 303950 33334
rect 304222 33062 304246 33334
rect 303926 30334 304246 33062
rect 303926 30062 303950 30334
rect 304222 30062 304246 30334
rect 303926 27334 304246 30062
rect 303926 27062 303950 27334
rect 304222 27062 304246 27334
rect 303926 24334 304246 27062
rect 303926 24062 303950 24334
rect 304222 24062 304246 24334
rect 303926 21334 304246 24062
rect 303926 21062 303950 21334
rect 304222 21062 304246 21334
rect -1526 18760 -1206 18780
rect 289572 18760 289952 18790
rect 303926 18760 304246 21062
rect -1579 18736 304262 18760
rect -1579 18464 3688 18736
rect 3960 18464 18112 18736
rect 18384 18464 32938 18736
rect 33210 18464 64280 18736
rect 64552 18464 121702 18736
rect 121974 18464 167572 18736
rect 167844 18464 180572 18736
rect 180844 18464 189572 18736
rect 189844 18464 198572 18736
rect 198844 18464 204572 18736
rect 204844 18464 211572 18736
rect 211844 18464 223572 18736
rect 223844 18464 232572 18736
rect 232844 18464 238572 18736
rect 238844 18464 250572 18736
rect 250844 18464 263972 18736
rect 264244 18464 269972 18736
rect 270244 18464 272972 18736
rect 273244 18464 275972 18736
rect 276244 18464 281972 18736
rect 282244 18464 285972 18736
rect 286244 18464 293972 18736
rect 294244 18464 296972 18736
rect 297244 18464 299972 18736
rect 300244 18464 302972 18736
rect 303244 18464 304262 18736
rect -1579 18440 304262 18464
rect 289572 18422 289952 18440
rect 303926 18104 304246 18440
rect 305437 17289 305757 326222
rect -2982 17265 305757 17289
rect -2982 16993 303890 17265
rect 304162 16993 305757 17265
rect -2982 16969 305757 16993
rect -2946 16904 -2626 16969
rect 644 16875 964 16969
rect 3644 16875 3964 16969
rect 6644 16875 6964 16969
rect 9644 16875 9964 16969
rect 12644 16875 12964 16969
rect 15644 16875 15964 16969
rect 18644 16875 18964 16969
rect 21644 16875 21964 16969
rect 24644 16875 24964 16969
rect 27644 16875 27964 16969
rect 30644 16875 30964 16969
rect 33644 16875 33964 16969
rect 36644 16875 36964 16969
rect 39644 16875 39964 16969
rect 42644 16875 42964 16969
rect 45644 16875 45964 16969
rect 48644 16875 48964 16969
rect 51644 16875 51964 16969
rect 54644 16875 54964 16969
rect 57644 16875 57964 16969
rect 60644 16875 60964 16969
rect 63644 16875 63964 16969
rect 66644 16875 66964 16969
rect 69644 16875 69964 16969
rect 72644 16875 72964 16969
rect 75644 16875 75964 16969
rect 78644 16875 78964 16969
rect 81644 16875 81964 16969
rect 84644 16875 84964 16969
rect 87644 16875 87964 16969
rect 90644 16875 90964 16969
rect 93644 16875 93964 16969
rect 96644 16875 96964 16969
rect 99644 16875 99964 16969
rect 102644 16875 102964 16969
rect 105644 16875 105964 16969
rect 108644 16875 108964 16969
rect 111644 16875 111964 16969
rect 114644 16875 114964 16969
rect 117644 16875 117964 16969
rect 120644 16875 120964 16969
rect 123644 16875 123964 16969
rect 126644 16875 126964 16969
rect 129644 16875 129964 16969
rect 132644 16875 132964 16969
rect 135644 16875 135964 16969
rect 138644 16875 138964 16969
rect 141644 16875 141964 16969
rect 144644 16875 144964 16969
rect 147644 16875 147964 16969
rect 150644 16875 150964 16969
rect 153644 16875 153964 16969
rect 156644 16875 156964 16969
rect 159644 16875 159964 16969
rect 162644 16875 162964 16969
rect 165644 16875 165964 16969
rect 168644 16875 168964 16969
rect 171644 16875 171964 16969
rect 174644 16875 174964 16969
rect 177644 16875 177964 16969
rect 180644 16875 180964 16969
rect 183644 16875 183964 16969
rect 186644 16875 186964 16969
rect 189644 16875 189964 16969
rect 192644 16875 192964 16969
rect 195644 16875 195964 16969
rect 198644 16875 198964 16969
rect 201644 16875 201964 16969
rect 204644 16875 204964 16969
rect 207644 16875 207964 16969
rect 210644 16875 210964 16969
rect 213644 16875 213964 16969
rect 216644 16875 216964 16969
rect 219644 16875 219964 16969
rect 222644 16875 222964 16969
rect 225644 16875 225964 16969
rect 228644 16875 228964 16969
rect 231644 16875 231964 16969
rect 234644 16875 234964 16969
rect 237644 16875 237964 16969
rect 240644 16875 240964 16969
rect 243644 16875 243964 16969
rect 246644 16875 246964 16969
rect 249644 16875 249964 16969
rect 252644 16875 252964 16969
rect 255644 16875 255964 16969
rect 258644 16875 258964 16969
rect 261644 16875 261964 16969
rect 264644 16875 264964 16969
rect 270644 16875 270964 16969
rect 273644 16875 273964 16969
rect 276644 16875 276964 16969
rect 279644 16875 279964 16969
rect 282644 16875 282964 16969
rect 285644 16875 285964 16969
rect 288644 16875 288964 16969
rect 291644 16875 291964 16969
rect 294644 16875 294964 16969
rect 297644 16875 297964 16969
rect 300644 16875 300964 16969
rect 302917 16410 303299 16434
rect 302917 16088 302941 16410
rect 303275 16088 303299 16410
rect 302917 16064 303299 16088
rect 306874 16049 307194 16842
rect 3634 15688 4014 15712
rect 24 15643 392 15667
rect 24 15323 48 15643
rect 368 15323 837 15643
rect 3634 15368 3658 15688
rect 3990 15368 4014 15688
rect 3634 15344 4014 15368
rect 18058 15706 18438 15730
rect 18058 15386 18082 15706
rect 18414 15386 18438 15706
rect 18058 15362 18438 15386
rect 32884 15682 33264 15706
rect 32884 15362 32908 15682
rect 33240 15362 33264 15682
rect 32884 15338 33264 15362
rect 64226 15690 64606 15714
rect 64226 15370 64250 15690
rect 64582 15370 64606 15690
rect 64226 15346 64606 15370
rect 121648 15704 122028 15728
rect 121648 15384 121672 15704
rect 122004 15384 122028 15704
rect 121648 15360 122028 15384
rect 167518 15706 167898 15730
rect 167518 15386 167542 15706
rect 167874 15386 167898 15706
rect 167518 15362 167898 15386
rect 180518 15706 180898 15730
rect 180518 15386 180542 15706
rect 180874 15386 180898 15706
rect 180518 15362 180898 15386
rect 189518 15706 189898 15730
rect 189518 15386 189542 15706
rect 189874 15386 189898 15706
rect 189518 15362 189898 15386
rect 198518 15706 198898 15730
rect 198518 15386 198542 15706
rect 198874 15386 198898 15706
rect 198518 15362 198898 15386
rect 204518 15706 204898 15730
rect 204518 15386 204542 15706
rect 204874 15386 204898 15706
rect 204518 15362 204898 15386
rect 211518 15706 211898 15730
rect 211518 15386 211542 15706
rect 211874 15386 211898 15706
rect 211518 15362 211898 15386
rect 223518 15706 223898 15730
rect 223518 15386 223542 15706
rect 223874 15386 223898 15706
rect 223518 15362 223898 15386
rect 232518 15706 232898 15730
rect 232518 15386 232542 15706
rect 232874 15386 232898 15706
rect 232518 15362 232898 15386
rect 238518 15706 238898 15730
rect 238518 15386 238542 15706
rect 238874 15386 238898 15706
rect 238518 15362 238898 15386
rect 250518 15706 250898 15730
rect 250518 15386 250542 15706
rect 250874 15386 250898 15706
rect 250518 15362 250898 15386
rect 263918 15706 264298 15730
rect 263918 15386 263942 15706
rect 264274 15386 264298 15706
rect 263918 15362 264298 15386
rect 269918 15706 270298 15730
rect 269918 15386 269942 15706
rect 270274 15386 270298 15706
rect 269918 15362 270298 15386
rect 272918 15706 273298 15730
rect 272918 15386 272942 15706
rect 273274 15386 273298 15706
rect 272918 15362 273298 15386
rect 275918 15706 276298 15730
rect 275918 15386 275942 15706
rect 276274 15386 276298 15706
rect 275918 15362 276298 15386
rect 281918 15706 282298 15730
rect 281918 15386 281942 15706
rect 282274 15386 282298 15706
rect 281918 15362 282298 15386
rect 285918 15706 286298 15730
rect 285918 15386 285942 15706
rect 286274 15386 286298 15706
rect 285918 15362 286298 15386
rect 293918 15706 294298 15730
rect 293918 15386 293942 15706
rect 294274 15386 294298 15706
rect 293918 15362 294298 15386
rect 296918 15706 297298 15730
rect 296918 15386 296942 15706
rect 297274 15386 297298 15706
rect 296918 15362 297298 15386
rect 299918 15706 300298 15730
rect 299918 15386 299942 15706
rect 300274 15386 300298 15706
rect 299918 15362 300298 15386
rect 302918 15706 303298 15730
rect 302918 15386 302942 15706
rect 303274 15386 303298 15706
rect 302918 15362 303298 15386
rect 303842 15692 304210 15716
rect 303842 15372 303866 15692
rect 304186 15372 304210 15692
rect 303842 15348 304210 15372
rect 24 15299 392 15323
use pixel_array100x100  pixel_array100x100_0
timestamp 1654904798
transform 1 0 2108 0 1 317378
box -3000 -298600 300740 5750
use shift_registerC  shift_registerC_0
timestamp 1654744971
transform 1 0 58 0 1 590
box -1076 -4 307988 16000
use shift_register  shift_register_0
timestamp 1654744971
transform 0 1 -21072 -1 0 323984
box -1076 -4 307988 16000
<< labels >>
rlabel metal5 -2842 18751 -2834 18760 1 VDD
<< end >>
