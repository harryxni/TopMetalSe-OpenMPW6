magic
tech sky130A
magscale 1 2
timestamp 1654709783
<< error_p >>
rect 452877 671886 452911 672462
rect 452995 671886 453029 672462
rect 453113 671886 453147 672462
rect 453231 671886 453265 672462
rect 453349 671886 453383 672462
rect 453467 671886 453501 672462
rect 453585 671886 453619 672462
rect 453703 671886 453737 672462
rect 453821 671886 453855 672462
rect 453939 671886 453973 672462
rect 454057 671886 454091 672462
rect 454175 671886 454209 672462
rect 454293 671886 454327 672462
rect 454411 671886 454445 672462
rect 454529 671886 454563 672462
rect 454647 671886 454681 672462
rect 454765 671886 454799 672462
rect 454883 671886 454917 672462
rect 455001 671886 455035 672462
rect 455119 671886 455153 672462
rect 455237 671886 455271 672462
rect 455355 671886 455389 672462
rect 455473 671886 455507 672462
rect 455591 671886 455625 672462
rect 457000 671886 457034 672462
rect 457118 671886 457152 672462
rect 457236 671886 457270 672462
rect 457354 671886 457388 672462
rect 457472 671886 457506 672462
rect 457590 671886 457624 672462
rect 457708 671886 457742 672462
rect 457826 671886 457860 672462
rect 457944 671886 457978 672462
rect 458062 671886 458096 672462
rect 458180 671886 458214 672462
rect 458298 671886 458332 672462
rect 458416 671886 458450 672462
rect 458534 671886 458568 672462
rect 458652 671886 458686 672462
rect 458770 671886 458804 672462
rect 458888 671886 458922 672462
rect 459006 671886 459040 672462
rect 459124 671886 459158 672462
rect 459242 671886 459276 672462
rect 459360 671886 459394 672462
rect 459478 671886 459512 672462
rect 459596 671886 459630 672462
rect 459714 671886 459748 672462
rect 461123 671886 461157 672462
rect 461241 671886 461275 672462
rect 461359 671886 461393 672462
rect 461477 671886 461511 672462
rect 461595 671886 461629 672462
rect 461713 671886 461747 672462
rect 461831 671886 461865 672462
rect 461949 671886 461983 672462
rect 462067 671886 462101 672462
rect 462185 671886 462219 672462
rect 462303 671886 462337 672462
rect 462421 671886 462455 672462
rect 462539 671886 462573 672462
rect 462657 671886 462691 672462
rect 462775 671886 462809 672462
rect 462893 671886 462927 672462
rect 463011 671886 463045 672462
rect 463129 671886 463163 672462
rect 463247 671886 463281 672462
rect 463365 671886 463399 672462
rect 463483 671886 463517 672462
rect 463601 671886 463635 672462
rect 463719 671886 463753 672462
rect 463837 671886 463871 672462
rect 448064 671127 450903 671161
rect 448137 670390 448171 670966
rect 448255 670390 448289 670966
rect 448373 670390 448407 670966
rect 448491 670390 448525 670966
rect 448609 670390 448643 670966
rect 448727 670390 448761 670966
rect 448845 670390 448879 670966
rect 448963 670390 448997 670966
rect 449081 670390 449115 670966
rect 449199 670390 449233 670966
rect 449317 670390 449351 670966
rect 449435 670390 449469 670966
rect 449553 670390 449587 670966
rect 449671 670390 449705 670966
rect 449789 670390 449823 670966
rect 449907 670390 449941 670966
rect 450025 670390 450059 670966
rect 450143 670390 450177 670966
rect 450261 670390 450295 670966
rect 450379 670390 450413 670966
rect 450497 670390 450531 670966
rect 450615 670390 450649 670966
rect 450733 670390 450767 670966
rect 450851 670390 450885 670966
rect 448137 669554 448171 670130
rect 448255 669554 448289 670130
rect 448373 669554 448407 670130
rect 448491 669554 448525 670130
rect 448609 669554 448643 670130
rect 448727 669554 448761 670130
rect 448845 669554 448879 670130
rect 448963 669554 448997 670130
rect 449081 669554 449115 670130
rect 449199 669554 449233 670130
rect 449317 669554 449351 670130
rect 449435 669554 449469 670130
rect 449553 669554 449587 670130
rect 449671 669554 449705 670130
rect 449789 669554 449823 670130
rect 449907 669554 449941 670130
rect 450025 669554 450059 670130
rect 450143 669554 450177 670130
rect 450261 669554 450295 670130
rect 450379 669554 450413 670130
rect 450497 669554 450531 670130
rect 450615 669554 450649 670130
rect 450733 669554 450767 670130
rect 450851 669554 450885 670130
rect 450965 669455 450999 671065
rect 452641 671050 452675 671626
rect 452759 671050 452793 671626
rect 452877 671050 452911 671626
rect 452995 671050 453029 671626
rect 453113 671050 453147 671626
rect 453231 671050 453265 671626
rect 453349 671050 453383 671626
rect 453467 671050 453501 671626
rect 453585 671050 453619 671626
rect 453703 671050 453737 671626
rect 453821 671050 453855 671626
rect 453939 671050 453973 671626
rect 454057 671050 454091 671626
rect 454175 671050 454209 671626
rect 454293 671050 454327 671626
rect 454411 671050 454445 671626
rect 454529 671050 454563 671626
rect 454647 671050 454681 671626
rect 454765 671050 454799 671626
rect 454883 671050 454917 671626
rect 455001 671050 455035 671626
rect 455119 671050 455153 671626
rect 455237 671050 455271 671626
rect 455355 671050 455389 671626
rect 455473 671050 455507 671626
rect 455591 671050 455625 671626
rect 456764 671050 456798 671626
rect 456882 671050 456916 671626
rect 457000 671050 457034 671626
rect 457118 671050 457152 671626
rect 457236 671050 457270 671626
rect 457354 671050 457388 671626
rect 457472 671050 457506 671626
rect 457590 671050 457624 671626
rect 457708 671050 457742 671626
rect 457826 671050 457860 671626
rect 457944 671050 457978 671626
rect 458062 671050 458096 671626
rect 458180 671050 458214 671626
rect 458298 671050 458332 671626
rect 458416 671050 458450 671626
rect 458534 671050 458568 671626
rect 458652 671050 458686 671626
rect 458770 671050 458804 671626
rect 458888 671050 458922 671626
rect 459006 671050 459040 671626
rect 459124 671050 459158 671626
rect 459242 671050 459276 671626
rect 459360 671050 459394 671626
rect 459478 671050 459512 671626
rect 459596 671050 459630 671626
rect 459714 671050 459748 671626
rect 460887 671050 460921 671626
rect 461005 671050 461039 671626
rect 461123 671050 461157 671626
rect 461241 671050 461275 671626
rect 461359 671050 461393 671626
rect 461477 671050 461511 671626
rect 461595 671050 461629 671626
rect 461713 671050 461747 671626
rect 461831 671050 461865 671626
rect 461949 671050 461983 671626
rect 462067 671050 462101 671626
rect 462185 671050 462219 671626
rect 462303 671050 462337 671626
rect 462421 671050 462455 671626
rect 462539 671050 462573 671626
rect 462657 671050 462691 671626
rect 462775 671050 462809 671626
rect 462893 671050 462927 671626
rect 463011 671050 463045 671626
rect 463129 671050 463163 671626
rect 463247 671050 463281 671626
rect 463365 671050 463399 671626
rect 463483 671050 463517 671626
rect 463601 671050 463635 671626
rect 463719 671050 463753 671626
rect 463837 671050 463871 671626
rect 448064 669359 450903 669393
rect 448064 669077 450903 669111
rect 448727 668340 448761 668916
rect 448845 668340 448879 668916
rect 448963 668340 448997 668916
rect 449081 668340 449115 668916
rect 449199 668340 449233 668916
rect 449317 668340 449351 668916
rect 449435 668340 449469 668916
rect 449553 668340 449587 668916
rect 449671 668340 449705 668916
rect 449789 668340 449823 668916
rect 449907 668340 449941 668916
rect 450025 668340 450059 668916
rect 450143 668340 450177 668916
rect 450261 668340 450295 668916
rect 450379 668340 450413 668916
rect 450497 668340 450531 668916
rect 450615 668340 450649 668916
rect 450733 668340 450767 668916
rect 450851 668340 450885 668916
rect 448727 667504 448761 668080
rect 448845 667504 448879 668080
rect 448963 667504 448997 668080
rect 449081 667504 449115 668080
rect 449199 667504 449233 668080
rect 449317 667504 449351 668080
rect 449435 667504 449469 668080
rect 449553 667504 449587 668080
rect 449671 667504 449705 668080
rect 449789 667504 449823 668080
rect 449907 667504 449941 668080
rect 450025 667504 450059 668080
rect 450143 667504 450177 668080
rect 450261 667504 450295 668080
rect 450379 667504 450413 668080
rect 450497 667504 450531 668080
rect 450615 667504 450649 668080
rect 450733 667504 450767 668080
rect 450851 667504 450885 668080
rect 450965 667405 450999 669015
rect 448704 667309 450903 667343
rect 448704 667027 450903 667061
rect 448727 666290 448761 666866
rect 448845 666290 448879 666866
rect 448963 666290 448997 666866
rect 449081 666290 449115 666866
rect 449199 666290 449233 666866
rect 449317 666290 449351 666866
rect 449435 666290 449469 666866
rect 449553 666290 449587 666866
rect 449671 666290 449705 666866
rect 449789 666290 449823 666866
rect 449907 666290 449941 666866
rect 450025 666290 450059 666866
rect 450143 666290 450177 666866
rect 450261 666290 450295 666866
rect 450379 666290 450413 666866
rect 450497 666290 450531 666866
rect 450615 666290 450649 666866
rect 450733 666290 450767 666866
rect 450851 666290 450885 666866
rect 448727 665454 448761 666030
rect 448845 665454 448879 666030
rect 448963 665454 448997 666030
rect 449081 665454 449115 666030
rect 449199 665454 449233 666030
rect 449317 665454 449351 666030
rect 449435 665454 449469 666030
rect 449553 665454 449587 666030
rect 449671 665454 449705 666030
rect 449789 665454 449823 666030
rect 449907 665454 449941 666030
rect 450025 665454 450059 666030
rect 450143 665454 450177 666030
rect 450261 665454 450295 666030
rect 450379 665454 450413 666030
rect 450497 665454 450531 666030
rect 450615 665454 450649 666030
rect 450733 665454 450767 666030
rect 450851 665454 450885 666030
rect 450965 665355 450999 666965
rect 448704 665259 450903 665293
rect 448727 664240 448761 664816
rect 448845 664240 448879 664816
rect 448963 664240 448997 664816
rect 449081 664240 449115 664816
rect 449199 664240 449233 664816
rect 449317 664240 449351 664816
rect 449435 664240 449469 664816
rect 449553 664240 449587 664816
rect 449671 664240 449705 664816
rect 449789 664240 449823 664816
rect 449907 664240 449941 664816
rect 450025 664240 450059 664816
rect 450143 664240 450177 664816
rect 450261 664240 450295 664816
rect 450379 664240 450413 664816
rect 450497 664240 450531 664816
rect 450615 664240 450649 664816
rect 450733 664240 450767 664816
rect 450851 664240 450885 664816
rect 448727 663404 448761 663980
rect 448845 663404 448879 663980
rect 448963 663404 448997 663980
rect 449081 663404 449115 663980
rect 449199 663404 449233 663980
rect 449317 663404 449351 663980
rect 449435 663404 449469 663980
rect 449553 663404 449587 663980
rect 449671 663404 449705 663980
rect 449789 663404 449823 663980
rect 449907 663404 449941 663980
rect 450025 663404 450059 663980
rect 450143 663404 450177 663980
rect 450261 663404 450295 663980
rect 450379 663404 450413 663980
rect 450497 663404 450531 663980
rect 450615 663404 450649 663980
rect 450733 663404 450767 663980
rect 450851 663404 450885 663980
rect 448723 661997 448757 662573
rect 448841 661997 448875 662573
rect 448959 661997 448993 662573
rect 449077 661997 449111 662573
rect 449195 661997 449229 662573
rect 449313 661997 449347 662573
rect 449431 661997 449465 662573
rect 449549 661997 449583 662573
rect 449667 661997 449701 662573
rect 449785 661997 449819 662573
rect 450878 662195 450912 662501
rect 450992 662285 451026 662411
rect 451080 662285 451114 662411
rect 451194 662195 451228 662501
rect 451308 662285 451342 662411
rect 451396 662285 451430 662411
rect 451510 662195 451544 662501
rect 451624 662285 451658 662411
rect 451712 662285 451746 662411
rect 451826 662195 451860 662501
rect 451940 662285 451974 662411
rect 452028 662285 452062 662411
rect 452142 662195 452176 662501
rect 452256 662285 452290 662411
rect 452344 662285 452378 662411
rect 452458 662195 452492 662501
rect 448723 661179 448757 661755
rect 448841 661179 448875 661755
rect 448959 661179 448993 661755
rect 449077 661179 449111 661755
rect 449195 661179 449229 661755
rect 449313 661179 449347 661755
rect 449431 661179 449465 661755
rect 449549 661179 449583 661755
rect 449667 661179 449701 661755
rect 449785 661179 449819 661755
rect 452675 661697 452709 662573
rect 452823 661697 452857 662573
rect 452971 661697 453005 662573
rect 453119 661697 453153 662573
rect 453267 661697 453301 662573
rect 453415 661697 453449 662573
rect 453563 661697 453597 662573
rect 453711 661697 453745 662573
rect 453859 661697 453893 662573
rect 454007 661697 454041 662573
rect 454155 661697 454189 662573
rect 454303 661697 454337 662573
rect 454451 661697 454485 662573
rect 454599 661697 454633 662573
rect 454747 661697 454781 662573
rect 454895 661697 454929 662573
rect 455043 661697 455077 662573
rect 455191 661697 455225 662573
rect 455339 661697 455373 662573
rect 455487 661697 455521 662573
rect 455635 661697 455669 662573
rect 455783 661697 455817 662573
rect 455931 661697 455965 662573
rect 456079 661697 456113 662573
rect 456227 661697 456261 662573
rect 456375 661697 456409 662573
rect 456523 661697 456557 662573
rect 456671 661697 456705 662573
rect 456819 661697 456853 662573
rect 456967 661697 457001 662573
rect 457115 661697 457149 662573
rect 457263 661697 457297 662573
rect 457411 661697 457445 662573
rect 457559 661697 457593 662573
rect 457707 661697 457741 662573
rect 457855 661697 457889 662573
rect 458003 661697 458037 662573
rect 458151 661697 458185 662573
rect 458299 661697 458333 662573
rect 458447 661697 458481 662573
rect 458595 661697 458629 662573
rect 458743 661697 458777 662573
rect 458891 661697 458925 662573
rect 459039 661697 459073 662573
rect 459187 661697 459221 662573
rect 459335 661697 459369 662573
rect 459483 661697 459517 662573
rect 459631 661697 459665 662573
rect 459779 661697 459813 662573
rect 459927 661697 459961 662573
rect 460075 661697 460109 662573
rect 460223 661697 460257 662573
rect 460371 661697 460405 662573
rect 460519 661697 460553 662573
rect 460667 661697 460701 662573
rect 460815 661697 460849 662573
rect 460963 661697 460997 662573
rect 461111 661697 461145 662573
rect 461259 661697 461293 662573
rect 461407 661697 461441 662573
rect 461555 661697 461589 662573
rect 461703 661697 461737 662573
rect 461851 661697 461885 662573
rect 461999 661697 462033 662573
rect 462147 661697 462181 662573
rect 462295 661697 462329 662573
rect 462443 661697 462477 662573
rect 462591 661697 462625 662573
rect 462739 661697 462773 662573
rect 462887 661697 462921 662573
rect 463035 661697 463069 662573
rect 463183 661697 463217 662573
rect 463331 661697 463365 662573
rect 463479 661697 463513 662573
rect 463775 661697 463809 662573
rect 452885 661613 452943 661647
rect 453033 661613 453091 661647
rect 453181 661613 453239 661647
rect 453329 661613 453387 661647
rect 453477 661613 453535 661647
rect 453625 661613 453683 661647
rect 453773 661613 453831 661647
rect 453921 661613 453979 661647
rect 454069 661613 454127 661647
rect 454217 661613 454275 661647
rect 454365 661613 454423 661647
rect 454513 661613 454571 661647
rect 454661 661613 454719 661647
rect 454809 661613 454867 661647
rect 454957 661613 455015 661647
rect 455105 661613 455163 661647
rect 455253 661613 455311 661647
rect 455401 661613 455459 661647
rect 455549 661613 455607 661647
rect 455697 661613 455755 661647
rect 455845 661613 455903 661647
rect 455993 661613 456051 661647
rect 456141 661613 456199 661647
rect 456289 661613 456347 661647
rect 456437 661613 456495 661647
rect 456585 661613 456643 661647
rect 456733 661613 456791 661647
rect 456881 661613 456939 661647
rect 457029 661613 457087 661647
rect 457177 661613 457235 661647
rect 457325 661613 457383 661647
rect 457473 661613 457531 661647
rect 457621 661613 457679 661647
rect 457769 661613 457827 661647
rect 457917 661613 457975 661647
rect 458065 661613 458123 661647
rect 458213 661613 458271 661647
rect 458361 661613 458419 661647
rect 458509 661613 458567 661647
rect 458657 661613 458715 661647
rect 458805 661613 458863 661647
rect 458953 661613 459011 661647
rect 459101 661613 459159 661647
rect 459249 661613 459307 661647
rect 459397 661613 459455 661647
rect 459545 661613 459603 661647
rect 459693 661613 459751 661647
rect 459841 661613 459899 661647
rect 459989 661613 460047 661647
rect 460137 661613 460195 661647
rect 460285 661613 460343 661647
rect 460433 661613 460491 661647
rect 460581 661613 460639 661647
rect 460729 661613 460787 661647
rect 460877 661613 460935 661647
rect 461025 661613 461083 661647
rect 461173 661613 461231 661647
rect 461321 661613 461379 661647
rect 461469 661613 461527 661647
rect 461617 661613 461675 661647
rect 461765 661613 461823 661647
rect 461913 661613 461971 661647
rect 462061 661613 462119 661647
rect 462209 661613 462267 661647
rect 462357 661613 462415 661647
rect 462505 661613 462563 661647
rect 462653 661613 462711 661647
rect 462801 661613 462859 661647
rect 462949 661613 463007 661647
rect 463097 661613 463155 661647
rect 463245 661613 463303 661647
rect 463393 661613 463451 661647
rect 463541 661613 463599 661647
rect 463689 661613 463747 661647
rect 452885 661505 452943 661539
rect 453033 661505 453091 661539
rect 453181 661505 453239 661539
rect 453329 661505 453387 661539
rect 453477 661505 453535 661539
rect 453625 661505 453683 661539
rect 453773 661505 453831 661539
rect 453921 661505 453979 661539
rect 454069 661505 454127 661539
rect 454217 661505 454275 661539
rect 454365 661505 454423 661539
rect 454513 661505 454571 661539
rect 454661 661505 454719 661539
rect 454809 661505 454867 661539
rect 454957 661505 455015 661539
rect 455105 661505 455163 661539
rect 455253 661505 455311 661539
rect 455401 661505 455459 661539
rect 455549 661505 455607 661539
rect 455697 661505 455755 661539
rect 455845 661505 455903 661539
rect 455993 661505 456051 661539
rect 456141 661505 456199 661539
rect 456289 661505 456347 661539
rect 456437 661505 456495 661539
rect 456585 661505 456643 661539
rect 456733 661505 456791 661539
rect 456881 661505 456939 661539
rect 457029 661505 457087 661539
rect 457177 661505 457235 661539
rect 457325 661505 457383 661539
rect 457473 661505 457531 661539
rect 457621 661505 457679 661539
rect 457769 661505 457827 661539
rect 457917 661505 457975 661539
rect 458065 661505 458123 661539
rect 458213 661505 458271 661539
rect 458361 661505 458419 661539
rect 458509 661505 458567 661539
rect 458657 661505 458715 661539
rect 458805 661505 458863 661539
rect 458953 661505 459011 661539
rect 459101 661505 459159 661539
rect 459249 661505 459307 661539
rect 459397 661505 459455 661539
rect 459545 661505 459603 661539
rect 459693 661505 459751 661539
rect 459841 661505 459899 661539
rect 459989 661505 460047 661539
rect 460137 661505 460195 661539
rect 460285 661505 460343 661539
rect 460433 661505 460491 661539
rect 460581 661505 460639 661539
rect 460729 661505 460787 661539
rect 460877 661505 460935 661539
rect 461025 661505 461083 661539
rect 461173 661505 461231 661539
rect 461321 661505 461379 661539
rect 461469 661505 461527 661539
rect 461617 661505 461675 661539
rect 461765 661505 461823 661539
rect 461913 661505 461971 661539
rect 462061 661505 462119 661539
rect 462209 661505 462267 661539
rect 462357 661505 462415 661539
rect 462505 661505 462563 661539
rect 462653 661505 462711 661539
rect 462801 661505 462859 661539
rect 462949 661505 463007 661539
rect 463097 661505 463155 661539
rect 463245 661505 463303 661539
rect 463393 661505 463451 661539
rect 463541 661505 463599 661539
rect 463689 661505 463747 661539
rect 452675 660579 452709 661455
rect 452823 660579 452857 661455
rect 452971 660579 453005 661455
rect 453119 660579 453153 661455
rect 453267 660579 453301 661455
rect 453415 660579 453449 661455
rect 453563 660579 453597 661455
rect 453711 660579 453745 661455
rect 453859 660579 453893 661455
rect 454007 660579 454041 661455
rect 454155 660579 454189 661455
rect 454303 660579 454337 661455
rect 454451 660579 454485 661455
rect 454599 660579 454633 661455
rect 454747 660579 454781 661455
rect 454895 660579 454929 661455
rect 455043 660579 455077 661455
rect 455191 660579 455225 661455
rect 455339 660579 455373 661455
rect 455487 660579 455521 661455
rect 455635 660579 455669 661455
rect 455783 660579 455817 661455
rect 455931 660579 455965 661455
rect 456079 660579 456113 661455
rect 456227 660579 456261 661455
rect 456375 660579 456409 661455
rect 456523 660579 456557 661455
rect 456671 660579 456705 661455
rect 456819 660579 456853 661455
rect 456967 660579 457001 661455
rect 457115 660579 457149 661455
rect 457263 660579 457297 661455
rect 457411 660579 457445 661455
rect 457559 660579 457593 661455
rect 457707 660579 457741 661455
rect 457855 660579 457889 661455
rect 458003 660579 458037 661455
rect 458151 660579 458185 661455
rect 458299 660579 458333 661455
rect 458447 660579 458481 661455
rect 458595 660579 458629 661455
rect 458743 660579 458777 661455
rect 458891 660579 458925 661455
rect 459039 660579 459073 661455
rect 459187 660579 459221 661455
rect 459335 660579 459369 661455
rect 459483 660579 459517 661455
rect 459631 660579 459665 661455
rect 459779 660579 459813 661455
rect 459927 660579 459961 661455
rect 460075 660579 460109 661455
rect 460223 660579 460257 661455
rect 460371 660579 460405 661455
rect 460519 660579 460553 661455
rect 460667 660579 460701 661455
rect 460815 660579 460849 661455
rect 460963 660579 460997 661455
rect 461111 660579 461145 661455
rect 461259 660579 461293 661455
rect 461407 660579 461441 661455
rect 461555 660579 461589 661455
rect 461703 660579 461737 661455
rect 461851 660579 461885 661455
rect 461999 660579 462033 661455
rect 462147 660579 462181 661455
rect 462295 660579 462329 661455
rect 462443 660579 462477 661455
rect 462591 660579 462625 661455
rect 462739 660579 462773 661455
rect 462887 660579 462921 661455
rect 463035 660579 463069 661455
rect 463183 660579 463217 661455
rect 463331 660579 463365 661455
rect 463479 660579 463513 661455
<< error_ps >>
rect 447539 671887 447573 672463
rect 444933 671127 448064 671161
rect 444837 669455 444871 671065
rect 444951 670390 444985 670966
rect 445069 670390 445103 670966
rect 445187 670390 445221 670966
rect 445305 670390 445339 670966
rect 445423 670390 445457 670966
rect 445541 670390 445575 670966
rect 445659 670390 445693 670966
rect 445777 670390 445811 670966
rect 445895 670390 445929 670966
rect 446013 670390 446047 670966
rect 446131 670390 446165 670966
rect 446249 670390 446283 670966
rect 446367 670390 446401 670966
rect 446485 670390 446519 670966
rect 446603 670390 446637 670966
rect 446721 670390 446755 670966
rect 446839 670390 446873 670966
rect 446957 670390 446991 670966
rect 447075 670390 447109 670966
rect 447193 670390 447227 670966
rect 447311 670390 447345 670966
rect 447429 670390 447463 670966
rect 447547 670390 447581 670966
rect 447665 670390 447699 670966
rect 447783 670390 447817 670966
rect 447901 670390 447935 670966
rect 448019 670390 448053 670966
rect 444951 669554 444985 670130
rect 445069 669554 445103 670130
rect 445187 669554 445221 670130
rect 445305 669554 445339 670130
rect 445423 669554 445457 670130
rect 445541 669554 445575 670130
rect 445659 669554 445693 670130
rect 445777 669554 445811 670130
rect 445895 669554 445929 670130
rect 446013 669554 446047 670130
rect 446131 669554 446165 670130
rect 446249 669554 446283 670130
rect 446367 669554 446401 670130
rect 446485 669554 446519 670130
rect 446603 669554 446637 670130
rect 446721 669554 446755 670130
rect 446839 669554 446873 670130
rect 446957 669554 446991 670130
rect 447075 669554 447109 670130
rect 447193 669554 447227 670130
rect 447311 669554 447345 670130
rect 447429 669554 447463 670130
rect 447547 669554 447581 670130
rect 447665 669554 447699 670130
rect 447783 669554 447817 670130
rect 447901 669554 447935 670130
rect 448019 669554 448053 670130
rect 444933 669359 448064 669393
rect 444933 669077 448064 669111
rect 444837 667405 444871 669015
rect 444951 668340 444985 668916
rect 445069 668340 445103 668916
rect 445187 668340 445221 668916
rect 445305 668340 445339 668916
rect 445423 668340 445457 668916
rect 445541 668340 445575 668916
rect 445659 668340 445693 668916
rect 445777 668340 445811 668916
rect 445895 668340 445929 668916
rect 446013 668340 446047 668916
rect 446131 668340 446165 668916
rect 446249 668340 446283 668916
rect 446367 668340 446401 668916
rect 446485 668340 446519 668916
rect 446603 668340 446637 668916
rect 446721 668340 446755 668916
rect 446839 668340 446873 668916
rect 446957 668340 446991 668916
rect 447075 668340 447109 668916
rect 447193 668340 447227 668916
rect 447311 668340 447345 668916
rect 447429 668340 447463 668916
rect 447547 668340 447581 668916
rect 447665 668340 447699 668916
rect 447783 668340 447817 668916
rect 447901 668340 447935 668916
rect 448019 668340 448053 668916
rect 448137 668340 448171 668916
rect 448255 668340 448289 668916
rect 448373 668340 448407 668916
rect 448491 668340 448525 668916
rect 448609 668340 448643 668916
rect 444951 667504 444985 668080
rect 445069 667504 445103 668080
rect 445187 667504 445221 668080
rect 445305 667504 445339 668080
rect 445423 667504 445457 668080
rect 445541 667504 445575 668080
rect 445659 667504 445693 668080
rect 445777 667504 445811 668080
rect 445895 667504 445929 668080
rect 446013 667504 446047 668080
rect 446131 667504 446165 668080
rect 446249 667504 446283 668080
rect 446367 667504 446401 668080
rect 446485 667504 446519 668080
rect 446603 667504 446637 668080
rect 446721 667504 446755 668080
rect 446839 667504 446873 668080
rect 446957 667504 446991 668080
rect 447075 667504 447109 668080
rect 447193 667504 447227 668080
rect 447311 667504 447345 668080
rect 447429 667504 447463 668080
rect 447547 667504 447581 668080
rect 447665 667504 447699 668080
rect 447783 667504 447817 668080
rect 447901 667504 447935 668080
rect 448019 667504 448053 668080
rect 448137 667504 448171 668080
rect 448255 667504 448289 668080
rect 448373 667504 448407 668080
rect 448491 667504 448525 668080
rect 448609 667504 448643 668080
rect 444933 667309 448704 667343
rect 444933 667027 448704 667061
rect 444837 665355 444871 666965
rect 444951 666290 444985 666866
rect 445069 666290 445103 666866
rect 445187 666290 445221 666866
rect 445305 666290 445339 666866
rect 445423 666290 445457 666866
rect 445541 666290 445575 666866
rect 445659 666290 445693 666866
rect 445777 666290 445811 666866
rect 445895 666290 445929 666866
rect 446013 666290 446047 666866
rect 446131 666290 446165 666866
rect 446249 666290 446283 666866
rect 446367 666290 446401 666866
rect 446485 666290 446519 666866
rect 446603 666290 446637 666866
rect 446721 666290 446755 666866
rect 446839 666290 446873 666866
rect 446957 666290 446991 666866
rect 447075 666290 447109 666866
rect 447193 666290 447227 666866
rect 447311 666290 447345 666866
rect 447429 666290 447463 666866
rect 447547 666290 447581 666866
rect 447665 666290 447699 666866
rect 447783 666290 447817 666866
rect 447901 666290 447935 666866
rect 448019 666290 448053 666866
rect 448137 666290 448171 666866
rect 448255 666290 448289 666866
rect 448373 666290 448407 666866
rect 448491 666290 448525 666866
rect 448609 666290 448643 666866
rect 444951 665454 444985 666030
rect 445069 665454 445103 666030
rect 445187 665454 445221 666030
rect 445305 665454 445339 666030
rect 445423 665454 445457 666030
rect 445541 665454 445575 666030
rect 445659 665454 445693 666030
rect 445777 665454 445811 666030
rect 445895 665454 445929 666030
rect 446013 665454 446047 666030
rect 446131 665454 446165 666030
rect 446249 665454 446283 666030
rect 446367 665454 446401 666030
rect 446485 665454 446519 666030
rect 446603 665454 446637 666030
rect 446721 665454 446755 666030
rect 446839 665454 446873 666030
rect 446957 665454 446991 666030
rect 447075 665454 447109 666030
rect 447193 665454 447227 666030
rect 447311 665454 447345 666030
rect 447429 665454 447463 666030
rect 447547 665454 447581 666030
rect 447665 665454 447699 666030
rect 447783 665454 447817 666030
rect 447901 665454 447935 666030
rect 448019 665454 448053 666030
rect 448137 665454 448171 666030
rect 448255 665454 448289 666030
rect 448373 665454 448407 666030
rect 448491 665454 448525 666030
rect 448609 665454 448643 666030
rect 444933 665259 448704 665293
rect 445187 664240 445221 664816
rect 445305 664240 445339 664816
rect 445423 664240 445457 664816
rect 445541 664240 445575 664816
rect 445659 664240 445693 664816
rect 445777 664240 445811 664816
rect 445895 664240 445929 664816
rect 446013 664240 446047 664816
rect 446131 664240 446165 664816
rect 446249 664240 446283 664816
rect 446367 664240 446401 664816
rect 446485 664240 446519 664816
rect 446603 664240 446637 664816
rect 446721 664240 446755 664816
rect 446839 664240 446873 664816
rect 446957 664240 446991 664816
rect 447075 664240 447109 664816
rect 447193 664240 447227 664816
rect 447311 664240 447345 664816
rect 447429 664240 447463 664816
rect 447547 664240 447581 664816
rect 447665 664240 447699 664816
rect 447783 664240 447817 664816
rect 447901 664240 447935 664816
rect 448019 664240 448053 664816
rect 448137 664240 448171 664816
rect 448255 664240 448289 664816
rect 448373 664240 448407 664816
rect 448491 664240 448525 664816
rect 448609 664240 448643 664816
rect 444951 663404 444985 663980
rect 445069 663404 445103 663980
rect 445187 663404 445221 663980
rect 445305 663404 445339 663980
rect 445423 663404 445457 663980
rect 445541 663404 445575 663980
rect 445659 663404 445693 663980
rect 445777 663404 445811 663980
rect 445895 663404 445929 663980
rect 446013 663404 446047 663980
rect 446131 663404 446165 663980
rect 446249 663404 446283 663980
rect 446367 663404 446401 663980
rect 446485 663404 446519 663980
rect 446603 663404 446637 663980
rect 446721 663404 446755 663980
rect 446839 663404 446873 663980
rect 446957 663404 446991 663980
rect 447075 663404 447109 663980
rect 447193 663404 447227 663980
rect 447311 663404 447345 663980
rect 447429 663404 447463 663980
rect 447547 663404 447581 663980
rect 447665 663404 447699 663980
rect 447783 663404 447817 663980
rect 447901 663404 447935 663980
rect 448019 663404 448053 663980
rect 448137 663404 448171 663980
rect 448255 663404 448289 663980
rect 448373 663404 448407 663980
rect 448491 663404 448525 663980
rect 448609 663404 448643 663980
rect 446253 661997 446287 662573
rect 446371 661997 446405 662573
rect 446489 661997 446523 662573
rect 446607 661997 446641 662573
rect 446725 661997 446759 662573
rect 446843 661997 446877 662573
rect 446961 661997 446995 662573
rect 447079 661997 447113 662573
rect 447197 661997 447231 662573
rect 447315 661997 447349 662573
rect 447433 661997 447467 662573
rect 447551 661997 447585 662573
rect 447669 661997 447703 662573
rect 447787 661997 447821 662573
rect 448015 661997 448049 662573
rect 448133 661997 448167 662573
rect 448251 661997 448285 662573
rect 448369 661997 448403 662573
rect 448487 661997 448521 662573
rect 448605 661997 448639 662573
rect 446017 661179 446051 661755
rect 446135 661179 446169 661755
rect 446253 661179 446287 661755
rect 446371 661179 446405 661755
rect 446489 661179 446523 661755
rect 446607 661179 446641 661755
rect 446725 661179 446759 661755
rect 446843 661179 446877 661755
rect 446961 661179 446995 661755
rect 447079 661179 447113 661755
rect 447197 661179 447231 661755
rect 447315 661179 447349 661755
rect 447433 661179 447467 661755
rect 447551 661179 447585 661755
rect 447669 661179 447703 661755
rect 447787 661179 447821 661755
rect 448015 661179 448049 661755
rect 448133 661179 448167 661755
rect 448251 661179 448285 661755
rect 448369 661179 448403 661755
rect 448487 661179 448521 661755
rect 448605 661179 448639 661755
<< metal1 >>
rect 418200 691950 481296 691952
rect 416234 690440 481296 691950
rect 416234 675250 417746 690440
rect 475450 686940 477450 687220
rect 420280 686830 444000 686940
rect 416234 674110 416380 675250
rect 417490 674110 417746 675250
rect 416234 651066 417746 674110
rect 420230 685320 444000 686830
rect 473700 685320 477450 686940
rect 420230 676726 422230 685320
rect 420230 676336 428895 676726
rect 420230 670410 422230 676336
rect 428600 675416 428900 675430
rect 427204 674776 427210 675416
rect 428770 674776 429790 675416
rect 428600 674760 428900 674776
rect 475450 672970 477450 685320
rect 465755 672680 477450 672970
rect 420230 670210 426010 670410
rect 420230 667590 422230 670210
rect 420230 667390 426010 667590
rect 420230 664600 422230 667390
rect 420230 664400 426010 664600
rect 420230 661860 422230 664400
rect 420230 661660 426010 661860
rect 420230 655560 422230 661660
rect 469740 659830 469900 660130
rect 475450 655560 477450 672680
rect 420230 653560 477450 655560
rect 479784 660320 481296 690440
rect 479784 659910 479970 660320
rect 479784 659060 479960 659910
rect 481070 659470 481296 660320
rect 481060 659060 481296 659470
rect 479784 651066 481296 659060
rect 416234 649554 436784 651066
rect 438296 651030 481296 651066
rect 438296 650980 462600 651030
rect 438296 649580 452970 650980
rect 455460 649690 462600 650980
rect 464980 651020 481296 651030
rect 464980 649710 470790 651020
rect 473190 650930 481296 651020
rect 473190 649710 478570 650930
rect 464980 649690 478570 649710
rect 455460 649580 478570 649690
rect 438296 649570 478570 649580
rect 481250 649570 481296 650930
rect 438296 649554 481296 649570
<< via1 >>
rect 416380 674110 417490 675250
rect 444000 685320 473700 686940
rect 427210 674776 428770 675416
rect 437230 661710 437390 670670
rect 467660 659830 469740 660130
rect 479970 659910 481070 660320
rect 479960 659470 481070 659910
rect 479960 659060 481060 659470
rect 436784 649554 438296 651066
rect 452970 649580 455460 650980
rect 462600 649690 464980 651030
rect 470790 649710 473190 651020
rect 478570 649570 481250 650930
<< metal2 >>
rect 329590 703898 334190 703950
rect 329590 701295 329727 703898
rect 329385 700562 329727 701295
rect 334023 701295 334190 703898
rect 334023 700562 431530 701295
rect 329385 700405 431530 700562
rect 329590 700390 334190 700405
rect 430640 691190 431530 700405
rect 429890 690283 431530 691190
rect 429890 688627 430087 690283
rect 431423 688627 431530 690283
rect 429890 688420 431530 688627
rect 443980 686940 474650 687220
rect 443980 685320 444000 686940
rect 473700 685320 474650 686940
rect 443980 684550 474650 685320
rect 428371 675905 428445 675914
rect 428371 675806 428445 675815
rect 427180 675416 427880 675440
rect 428600 675416 428900 675430
rect 416340 675270 417560 675410
rect 416340 675250 416410 675270
rect 416340 674110 416380 675250
rect 417490 674110 417560 675270
rect 427180 674776 427210 675416
rect 428770 674776 428900 675416
rect 427180 674750 427880 674776
rect 428600 674760 428900 674776
rect 416340 673900 417560 674110
rect 423285 671010 424775 671120
rect 18660 668210 21180 668340
rect 18660 666130 18750 668210
rect 20950 666825 21180 668210
rect 423285 666825 423395 671010
rect 437210 670670 437410 670690
rect 424356 669140 424365 669230
rect 424455 669140 424645 669230
rect 20950 666715 423395 666825
rect 20950 666130 21180 666715
rect 424226 666140 424235 666230
rect 424325 666140 424565 666230
rect 18660 666030 21180 666130
rect 424585 663015 424675 663230
rect 424585 662916 424675 662925
rect 437210 661710 437230 670670
rect 437390 661710 437410 670670
rect 437210 661690 437410 661710
rect 479880 660330 481170 660450
rect 467633 660320 481170 660330
rect 467633 660155 479970 660320
rect 467535 660130 479970 660155
rect 467535 659830 467660 660130
rect 469740 659910 479970 660130
rect 469740 659830 479960 659910
rect 467535 659805 479960 659830
rect 467633 659060 479960 659805
rect 481070 659725 481170 660320
rect 481070 659470 481195 659725
rect 481060 659060 481195 659470
rect 467633 658935 481195 659060
rect 436590 651066 438530 651300
rect 436590 649554 436784 651066
rect 438296 649554 438530 651066
rect 452910 650980 455590 651380
rect 452910 649580 452970 650980
rect 455460 649580 455590 650980
rect 452910 649560 455590 649580
rect 462490 651030 465070 651320
rect 462490 649690 462600 651030
rect 464980 649690 465070 651030
rect 436590 649320 438530 649554
rect 462490 649550 465070 649690
rect 470650 651020 473280 651240
rect 470650 649710 470790 651020
rect 473190 649710 473280 651020
rect 470650 649630 473280 649710
rect 478470 650930 481370 651020
rect 478470 649570 478570 650930
rect 481250 649570 481370 650930
rect 478470 649490 481370 649570
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 329727 700562 334023 703898
rect 430087 688627 431423 690283
rect 444000 685320 473700 686940
rect 428371 675815 428445 675905
rect 416410 675250 417490 675270
rect 416410 674120 417490 675250
rect 427210 674776 427850 675416
rect 18750 666130 20950 668210
rect 424365 669140 424455 669230
rect 424235 666140 424325 666230
rect 424585 662925 424675 663015
rect 437230 661710 437390 670670
rect 436784 649554 438296 651066
rect 452970 649580 455460 650980
rect 462600 649690 464980 651030
rect 470790 649710 473190 651020
rect 478570 649570 481250 650930
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 703898 334294 704800
rect 329294 703862 329727 703898
rect 334023 703862 334294 703898
rect 329294 702300 329723 703862
rect -800 682742 1700 685242
rect -800 680242 8830 682742
rect 6330 658270 8830 680242
rect 18694 668340 21194 702300
rect 68940 680457 71440 702300
rect 68940 677513 69183 680457
rect 71087 677513 71440 680457
rect 68940 677160 71440 677513
rect 122330 673460 124830 702300
rect 177230 690870 179730 702300
rect 329590 700598 329723 702300
rect 334027 702300 334294 703862
rect 413394 703390 418394 704800
rect 413394 703190 427730 703390
rect 413394 702300 418394 703190
rect 334027 700598 334190 702300
rect 329590 700562 329727 700598
rect 334023 700562 334190 700598
rect 329590 700390 334190 700562
rect 177230 690670 420840 690870
rect 177230 690420 179730 690670
rect 420590 677600 420790 690670
rect 427530 679000 427730 703190
rect 465394 702720 470394 704800
rect 465394 702300 466100 702720
rect 465730 695550 466100 702300
rect 469420 702300 470394 702720
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 469420 695550 469710 702300
rect 465730 695030 469710 695550
rect 430080 690283 431430 690300
rect 428070 690142 429420 690170
rect 428070 688398 428073 690142
rect 429417 689404 429420 690142
rect 429417 688398 429424 689404
rect 430080 688627 430087 690283
rect 431423 689290 431430 690283
rect 431423 689170 433700 689290
rect 431423 688627 431430 689170
rect 430080 688610 431430 688627
rect 428070 688370 429424 688398
rect 428080 687660 429424 688370
rect 428360 687430 428480 687660
rect 428360 687310 431630 687430
rect 430490 679000 430690 679020
rect 427530 678800 430860 679000
rect 420590 677400 430230 677600
rect 429980 676650 430180 677400
rect 430490 676640 430690 678800
rect 431510 676350 431630 687310
rect 433580 676440 433700 689170
rect 442150 687830 476150 688490
rect 510594 687830 513054 702340
rect 566594 702300 571594 704800
rect 442150 686940 513054 687830
rect 442150 685320 444000 686940
rect 473700 685370 513054 686940
rect 473700 685320 476150 685370
rect 442150 684090 476150 685320
rect 574600 682984 582176 683000
rect 574600 682800 584800 682984
rect 574440 682402 584800 682800
rect 574440 678818 575238 682402
rect 582000 678818 584800 682402
rect 574440 678370 584800 678818
rect 582300 677984 584800 678370
rect 424900 675905 428470 675910
rect 424900 675815 428371 675905
rect 428445 675815 428470 675905
rect 424900 675810 428470 675815
rect 424900 675765 425140 675810
rect 413295 675675 425140 675765
rect 122330 671020 134005 673460
rect 413295 671020 413385 675675
rect 424900 675670 425140 675675
rect 427180 675416 427880 675440
rect 416340 675270 427210 675416
rect 416340 674120 416410 675270
rect 417490 674776 427210 675270
rect 427850 674776 428540 675416
rect 417490 674120 417550 674776
rect 427180 674750 427880 674776
rect 416340 673900 417550 674120
rect 122330 670960 413415 671020
rect 122330 670490 124830 670960
rect 125145 670930 413415 670960
rect 437210 670670 437410 670690
rect 424360 669230 424460 669235
rect 424360 669140 424365 669230
rect 424455 669140 424460 669230
rect 424360 669135 424460 669140
rect 424365 668465 424455 669135
rect 18660 668210 21194 668340
rect 18660 666130 18750 668210
rect 20950 667230 21194 668210
rect 423635 668375 424455 668465
rect 20950 666130 21180 667230
rect 423635 666465 423725 668375
rect 18660 666030 21180 666130
rect 412735 666375 423725 666465
rect 279474 665526 283616 665616
rect 412735 665526 412825 666375
rect 424230 666230 424330 666235
rect 424230 666140 424235 666230
rect 424325 666140 424330 666230
rect 424230 666135 424330 666140
rect 279474 665444 413031 665526
rect 279474 665440 279760 665444
rect 6330 655770 53060 658270
rect 47050 649732 53060 655770
rect -800 643842 1660 648642
rect 47050 644468 47678 649732
rect 51662 644468 53060 649732
rect 47050 643640 53060 644468
rect 47050 643620 52370 643640
rect -800 633842 1660 638642
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 279474 269342 279586 665440
rect 424235 665325 424325 666135
rect 422835 665235 424325 665325
rect 292684 662530 292796 662596
rect 422835 662530 422925 665235
rect 424580 663015 424680 663020
rect 424580 662925 424585 663015
rect 424675 662925 424680 663015
rect 424580 662920 424680 662925
rect 291330 662440 422925 662530
rect 292684 313764 292796 662440
rect 422835 662415 422925 662440
rect 384641 659530 384720 659540
rect 412770 659530 413900 659890
rect 384640 659450 413900 659530
rect 384640 358986 384720 659450
rect 412770 659425 413900 659450
rect 424585 659425 424675 662920
rect 412770 659335 424675 659425
rect 437210 661710 437230 670670
rect 437390 661760 437410 670670
rect 437390 661710 437900 661760
rect 412770 659220 413900 659335
rect 437210 651300 437900 661710
rect 436590 651066 438530 651300
rect 436590 649554 436784 651066
rect 438296 649554 438530 651066
rect 452910 650980 455590 651380
rect 452910 649580 452970 650980
rect 455460 649580 455590 650980
rect 452910 649560 455590 649580
rect 462480 651030 465120 651390
rect 462480 649690 462600 651030
rect 464980 649690 465120 651030
rect 462480 649560 465120 649690
rect 470650 651020 473280 651240
rect 470650 649710 470790 651020
rect 473190 649710 473280 651020
rect 470650 649630 473280 649710
rect 478470 650930 481370 651020
rect 436590 649320 438530 649554
rect 453010 642244 455470 649560
rect 462600 642244 465060 649560
rect 470690 642244 473150 649630
rect 478470 649570 478570 650930
rect 481250 649570 481370 650930
rect 478470 649490 481370 649570
rect 478710 642244 481170 649490
rect 582340 642244 584800 644584
rect 453010 639784 584800 642244
rect 431430 632842 431660 632910
rect 431430 632698 431478 632842
rect 431622 632746 431660 632842
rect 431622 632698 434196 632746
rect 431430 632640 434196 632698
rect 431434 632634 434196 632640
rect 424960 629437 425750 629530
rect 417534 629116 417646 629126
rect 424960 629116 425058 629437
rect 417534 629004 425058 629116
rect 417534 449830 417646 629004
rect 424960 628653 425058 629004
rect 425682 628653 425750 629437
rect 424960 628570 425750 628653
rect 425010 618052 425650 618150
rect 425010 617428 425063 618052
rect 425607 617428 425650 618052
rect 425010 617320 425650 617428
rect 425244 494252 425356 617320
rect 434084 583674 434196 632634
rect 582340 629784 584800 634584
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 434084 583562 584800 583674
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 425244 494140 584800 494252
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 416110 449718 584800 449830
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 382590 358874 584800 358986
rect 384640 347160 384720 358874
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 292684 313652 584800 313764
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 279474 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 69183 677513 71087 680457
rect 329723 700598 329727 703862
rect 329727 700598 334023 703862
rect 334023 700598 334027 703862
rect 466100 695550 469420 702720
rect 428073 688398 429417 690142
rect 575238 678818 582000 682402
rect 47678 644468 51662 649732
rect 431478 632698 431622 632842
rect 425058 628653 425682 629437
rect 425063 617428 425607 618052
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 703862 334294 704800
rect 329294 702300 329723 703862
rect 329590 700598 329723 702300
rect 334027 702300 334294 703862
rect 465730 702720 469710 702920
rect 334027 700598 334190 702300
rect 329590 700390 334190 700598
rect 229190 699708 231690 699960
rect 229190 698530 229597 699708
rect 228350 697552 229597 698530
rect 231433 698530 231690 699708
rect 231433 697552 429260 698530
rect 228350 697490 429260 697552
rect 229190 697460 231690 697490
rect 428220 691210 429260 697490
rect 465730 695550 466100 702720
rect 469420 695550 469710 702720
rect 465730 695030 469710 695550
rect 427960 690142 429520 691210
rect 427960 688398 428073 690142
rect 429417 688398 429520 690142
rect 427960 688310 429520 688398
rect 574553 682650 577887 682687
rect 574553 682402 582200 682650
rect 69000 680457 71280 680620
rect 69000 677513 69183 680457
rect 71087 677513 71280 680457
rect 69000 677445 71280 677513
rect 574553 678818 575238 682402
rect 582000 678818 582200 682402
rect 574553 678570 582200 678818
rect 68975 668080 71305 677445
rect 414355 671210 424765 671320
rect 412730 668125 413270 668290
rect 414355 668125 414465 671210
rect 469630 668230 472820 669090
rect 412730 668080 414465 668125
rect 51105 668015 414465 668080
rect 51105 667990 413270 668015
rect 291955 666770 292045 667715
rect 471960 665164 472820 668230
rect 574553 665164 577887 678570
rect 471883 661830 577887 665164
rect 427330 652525 427440 660015
rect 423975 652415 427440 652525
rect 47040 649732 52410 650020
rect 47040 644468 47678 649732
rect 51662 644468 52410 649732
rect 47040 643860 52410 644468
rect 291955 643860 292045 644510
rect 423975 643860 424085 652415
rect 428030 648860 428250 660290
rect 425300 648640 428250 648860
rect 46850 643760 424530 643860
rect 47040 643620 52410 643760
rect 291955 643670 292045 643760
rect 423975 643735 424085 643760
rect 425300 643110 425660 648640
rect 431030 647240 431250 660390
rect 428460 647020 431250 647240
rect 428460 644040 428680 647020
rect 425440 629530 425660 643110
rect 428440 642840 428680 644040
rect 431440 643660 431660 644250
rect 434030 643660 434250 660140
rect 431440 643440 434250 643660
rect 424960 629437 425750 629530
rect 424960 628653 425058 629437
rect 425682 628653 425750 629437
rect 424960 628570 425750 628653
rect 425440 628500 425660 628570
rect 425010 618052 425650 618150
rect 425010 617428 425063 618052
rect 425607 617910 425650 618052
rect 428440 617910 428660 642840
rect 431440 632842 431660 643440
rect 431440 632698 431478 632842
rect 431622 632698 431660 632842
rect 431440 632650 431660 632698
rect 425607 617690 428660 617910
rect 425607 617428 425650 617690
rect 425010 617320 425650 617428
<< via4 >>
rect 329837 700672 333913 703788
rect 229597 697552 231433 699708
rect 466100 695550 469420 702720
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 703788 334294 704800
rect 329294 702300 329837 703788
rect 229160 699708 231660 702300
rect 329590 700672 329837 702300
rect 333913 702300 334294 703788
rect 465730 702960 468080 702970
rect 465730 702720 469630 702960
rect 333913 700672 334230 702300
rect 329590 700360 334230 700672
rect 229160 697552 229597 699708
rect 231433 697552 231660 699708
rect 229160 697490 231660 697552
rect 465730 695550 466100 702720
rect 469420 695550 469630 702720
rect 465730 695350 469630 695550
rect 424660 695030 469730 695350
rect 424660 670500 424980 695030
use test  test_0
timestamp 1654648307
transform 1 0 431360 0 1 656230
box -6885 3561 39290 20620
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1400 0 0 0 gpio_analog[0]
port 1 nsew
flabel metal3 s -800 381864 480 381976 0 FreeSans 1400 0 0 0 gpio_analog[10]
port 2 nsew
flabel metal3 s -800 338642 480 338754 0 FreeSans 1400 0 0 0 gpio_analog[11]
port 3 nsew
flabel metal3 s -800 295420 480 295532 0 FreeSans 1400 0 0 0 gpio_analog[12]
port 4 nsew
flabel metal3 s -800 252398 480 252510 0 FreeSans 1400 0 0 0 gpio_analog[13]
port 5 nsew
flabel metal3 s -800 124776 480 124888 0 FreeSans 1400 0 0 0 gpio_analog[14]
port 6 nsew
flabel metal3 s -800 81554 480 81666 0 FreeSans 1400 0 0 0 gpio_analog[15]
port 7 nsew
flabel metal3 s -800 38332 480 38444 0 FreeSans 1400 0 0 0 gpio_analog[16]
port 8 nsew
flabel metal3 s -800 16910 480 17022 0 FreeSans 1400 0 0 0 gpio_analog[17]
port 9 nsew
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1400 0 0 0 gpio_analog[1]
port 10 nsew
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1400 0 0 0 gpio_analog[2]
port 11 nsew
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1400 0 0 0 gpio_analog[3]
port 12 nsew
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1400 0 0 0 gpio_analog[4]
port 13 nsew
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1400 0 0 0 gpio_analog[5]
port 14 nsew
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1400 0 0 0 gpio_analog[6]
port 15 nsew
flabel metal3 s -800 511530 480 511642 0 FreeSans 1400 0 0 0 gpio_analog[7]
port 16 nsew
flabel metal3 s -800 468308 480 468420 0 FreeSans 1400 0 0 0 gpio_analog[8]
port 17 nsew
flabel metal3 s -800 425086 480 425198 0 FreeSans 1400 0 0 0 gpio_analog[9]
port 18 nsew
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1400 0 0 0 gpio_noesd[0]
port 19 nsew
flabel metal3 s -800 380682 480 380794 0 FreeSans 1400 0 0 0 gpio_noesd[10]
port 20 nsew
flabel metal3 s -800 337460 480 337572 0 FreeSans 1400 0 0 0 gpio_noesd[11]
port 21 nsew
flabel metal3 s -800 294238 480 294350 0 FreeSans 1400 0 0 0 gpio_noesd[12]
port 22 nsew
flabel metal3 s -800 251216 480 251328 0 FreeSans 1400 0 0 0 gpio_noesd[13]
port 23 nsew
flabel metal3 s -800 123594 480 123706 0 FreeSans 1400 0 0 0 gpio_noesd[14]
port 24 nsew
flabel metal3 s -800 80372 480 80484 0 FreeSans 1400 0 0 0 gpio_noesd[15]
port 25 nsew
flabel metal3 s -800 37150 480 37262 0 FreeSans 1400 0 0 0 gpio_noesd[16]
port 26 nsew
flabel metal3 s -800 15728 480 15840 0 FreeSans 1400 0 0 0 gpio_noesd[17]
port 27 nsew
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1400 0 0 0 gpio_noesd[1]
port 28 nsew
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1400 0 0 0 gpio_noesd[2]
port 29 nsew
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1400 0 0 0 gpio_noesd[3]
port 30 nsew
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1400 0 0 0 gpio_noesd[4]
port 31 nsew
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1400 0 0 0 gpio_noesd[5]
port 32 nsew
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1400 0 0 0 gpio_noesd[6]
port 33 nsew
flabel metal3 s -800 510348 480 510460 0 FreeSans 1400 0 0 0 gpio_noesd[7]
port 34 nsew
flabel metal3 s -800 467126 480 467238 0 FreeSans 1400 0 0 0 gpio_noesd[8]
port 35 nsew
flabel metal3 s -800 423904 480 424016 0 FreeSans 1400 0 0 0 gpio_noesd[9]
port 36 nsew
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1400 0 0 0 io_analog[0]
port 37 nsew
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1400 0 0 0 io_analog[10]
port 38 nsew
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 2400 180 0 0 io_analog[1]
port 39 nsew
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 2400 180 0 0 io_analog[2]
port 40 nsew
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 2400 180 0 0 io_analog[3]
port 41 nsew
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 2400 180 0 0 io_analog[7]
port 45 nsew
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 2400 180 0 0 io_analog[8]
port 46 nsew
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 2400 180 0 0 io_analog[9]
port 47 nsew
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 2400 180 0 0 io_clamp_high[0]
port 48 nsew
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 2400 180 0 0 io_clamp_high[1]
port 49 nsew
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 2400 180 0 0 io_clamp_high[2]
port 50 nsew
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 2400 180 0 0 io_clamp_low[0]
port 51 nsew
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 2400 180 0 0 io_clamp_low[1]
port 52 nsew
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 2400 180 0 0 io_clamp_low[2]
port 53 nsew
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1400 0 0 0 io_in[0]
port 54 nsew
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1400 0 0 0 io_in[10]
port 55 nsew
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1400 0 0 0 io_in[11]
port 56 nsew
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1400 0 0 0 io_in[12]
port 57 nsew
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1400 0 0 0 io_in[13]
port 58 nsew
flabel metal3 s -800 507984 480 508096 0 FreeSans 1400 0 0 0 io_in[14]
port 59 nsew
flabel metal3 s -800 464762 480 464874 0 FreeSans 1400 0 0 0 io_in[15]
port 60 nsew
flabel metal3 s -800 421540 480 421652 0 FreeSans 1400 0 0 0 io_in[16]
port 61 nsew
flabel metal3 s -800 378318 480 378430 0 FreeSans 1400 0 0 0 io_in[17]
port 62 nsew
flabel metal3 s -800 335096 480 335208 0 FreeSans 1400 0 0 0 io_in[18]
port 63 nsew
flabel metal3 s -800 291874 480 291986 0 FreeSans 1400 0 0 0 io_in[19]
port 64 nsew
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1400 0 0 0 io_in[1]
port 65 nsew
flabel metal3 s -800 248852 480 248964 0 FreeSans 1400 0 0 0 io_in[20]
port 66 nsew
flabel metal3 s -800 121230 480 121342 0 FreeSans 1400 0 0 0 io_in[21]
port 67 nsew
flabel metal3 s -800 78008 480 78120 0 FreeSans 1400 0 0 0 io_in[22]
port 68 nsew
flabel metal3 s -800 34786 480 34898 0 FreeSans 1400 0 0 0 io_in[23]
port 69 nsew
flabel metal3 s -800 13364 480 13476 0 FreeSans 1400 0 0 0 io_in[24]
port 70 nsew
flabel metal3 s -800 8636 480 8748 0 FreeSans 1400 0 0 0 io_in[25]
port 71 nsew
flabel metal3 s -800 3908 480 4020 0 FreeSans 1400 0 0 0 io_in[26]
port 72 nsew
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1400 0 0 0 io_in[2]
port 73 nsew
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1400 0 0 0 io_in[3]
port 74 nsew
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1400 0 0 0 io_in[4]
port 75 nsew
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1400 0 0 0 io_in[5]
port 76 nsew
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1400 0 0 0 io_in[6]
port 77 nsew
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1400 0 0 0 io_in[7]
port 78 nsew
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1400 0 0 0 io_in[8]
port 79 nsew
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1400 0 0 0 io_in[9]
port 80 nsew
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1400 0 0 0 io_in_3v3[0]
port 81 nsew
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1400 0 0 0 io_in_3v3[10]
port 82 nsew
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1400 0 0 0 io_in_3v3[11]
port 83 nsew
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1400 0 0 0 io_in_3v3[12]
port 84 nsew
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1400 0 0 0 io_in_3v3[13]
port 85 nsew
flabel metal3 s -800 509166 480 509278 0 FreeSans 1400 0 0 0 io_in_3v3[14]
port 86 nsew
flabel metal3 s -800 465944 480 466056 0 FreeSans 1400 0 0 0 io_in_3v3[15]
port 87 nsew
flabel metal3 s -800 422722 480 422834 0 FreeSans 1400 0 0 0 io_in_3v3[16]
port 88 nsew
flabel metal3 s -800 379500 480 379612 0 FreeSans 1400 0 0 0 io_in_3v3[17]
port 89 nsew
flabel metal3 s -800 336278 480 336390 0 FreeSans 1400 0 0 0 io_in_3v3[18]
port 90 nsew
flabel metal3 s -800 293056 480 293168 0 FreeSans 1400 0 0 0 io_in_3v3[19]
port 91 nsew
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1400 0 0 0 io_in_3v3[1]
port 92 nsew
flabel metal3 s -800 250034 480 250146 0 FreeSans 1400 0 0 0 io_in_3v3[20]
port 93 nsew
flabel metal3 s -800 122412 480 122524 0 FreeSans 1400 0 0 0 io_in_3v3[21]
port 94 nsew
flabel metal3 s -800 79190 480 79302 0 FreeSans 1400 0 0 0 io_in_3v3[22]
port 95 nsew
flabel metal3 s -800 35968 480 36080 0 FreeSans 1400 0 0 0 io_in_3v3[23]
port 96 nsew
flabel metal3 s -800 14546 480 14658 0 FreeSans 1400 0 0 0 io_in_3v3[24]
port 97 nsew
flabel metal3 s -800 9818 480 9930 0 FreeSans 1400 0 0 0 io_in_3v3[25]
port 98 nsew
flabel metal3 s -800 5090 480 5202 0 FreeSans 1400 0 0 0 io_in_3v3[26]
port 99 nsew
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1400 0 0 0 io_in_3v3[2]
port 100 nsew
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1400 0 0 0 io_in_3v3[3]
port 101 nsew
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1400 0 0 0 io_in_3v3[4]
port 102 nsew
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1400 0 0 0 io_in_3v3[5]
port 103 nsew
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1400 0 0 0 io_in_3v3[6]
port 104 nsew
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1400 0 0 0 io_in_3v3[7]
port 105 nsew
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1400 0 0 0 io_in_3v3[8]
port 106 nsew
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1400 0 0 0 io_in_3v3[9]
port 107 nsew
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1400 0 0 0 io_oeb[0]
port 108 nsew
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1400 0 0 0 io_oeb[10]
port 109 nsew
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1400 0 0 0 io_oeb[11]
port 110 nsew
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1400 0 0 0 io_oeb[12]
port 111 nsew
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1400 0 0 0 io_oeb[13]
port 112 nsew
flabel metal3 s -800 505620 480 505732 0 FreeSans 1400 0 0 0 io_oeb[14]
port 113 nsew
flabel metal3 s -800 462398 480 462510 0 FreeSans 1400 0 0 0 io_oeb[15]
port 114 nsew
flabel metal3 s -800 419176 480 419288 0 FreeSans 1400 0 0 0 io_oeb[16]
port 115 nsew
flabel metal3 s -800 375954 480 376066 0 FreeSans 1400 0 0 0 io_oeb[17]
port 116 nsew
flabel metal3 s -800 332732 480 332844 0 FreeSans 1400 0 0 0 io_oeb[18]
port 117 nsew
flabel metal3 s -800 289510 480 289622 0 FreeSans 1400 0 0 0 io_oeb[19]
port 118 nsew
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1400 0 0 0 io_oeb[1]
port 119 nsew
flabel metal3 s -800 246488 480 246600 0 FreeSans 1400 0 0 0 io_oeb[20]
port 120 nsew
flabel metal3 s -800 118866 480 118978 0 FreeSans 1400 0 0 0 io_oeb[21]
port 121 nsew
flabel metal3 s -800 75644 480 75756 0 FreeSans 1400 0 0 0 io_oeb[22]
port 122 nsew
flabel metal3 s -800 32422 480 32534 0 FreeSans 1400 0 0 0 io_oeb[23]
port 123 nsew
flabel metal3 s -800 11000 480 11112 0 FreeSans 1400 0 0 0 io_oeb[24]
port 124 nsew
flabel metal3 s -800 6272 480 6384 0 FreeSans 1400 0 0 0 io_oeb[25]
port 125 nsew
flabel metal3 s -800 1544 480 1656 0 FreeSans 1400 0 0 0 io_oeb[26]
port 126 nsew
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1400 0 0 0 io_oeb[2]
port 127 nsew
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1400 0 0 0 io_oeb[3]
port 128 nsew
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1400 0 0 0 io_oeb[4]
port 129 nsew
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1400 0 0 0 io_oeb[5]
port 130 nsew
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1400 0 0 0 io_oeb[6]
port 131 nsew
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1400 0 0 0 io_oeb[7]
port 132 nsew
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1400 0 0 0 io_oeb[8]
port 133 nsew
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1400 0 0 0 io_oeb[9]
port 134 nsew
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1400 0 0 0 io_out[0]
port 135 nsew
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1400 0 0 0 io_out[10]
port 136 nsew
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1400 0 0 0 io_out[11]
port 137 nsew
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1400 0 0 0 io_out[12]
port 138 nsew
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1400 0 0 0 io_out[13]
port 139 nsew
flabel metal3 s -800 506802 480 506914 0 FreeSans 1400 0 0 0 io_out[14]
port 140 nsew
flabel metal3 s -800 463580 480 463692 0 FreeSans 1400 0 0 0 io_out[15]
port 141 nsew
flabel metal3 s -800 420358 480 420470 0 FreeSans 1400 0 0 0 io_out[16]
port 142 nsew
flabel metal3 s -800 377136 480 377248 0 FreeSans 1400 0 0 0 io_out[17]
port 143 nsew
flabel metal3 s -800 333914 480 334026 0 FreeSans 1400 0 0 0 io_out[18]
port 144 nsew
flabel metal3 s -800 290692 480 290804 0 FreeSans 1400 0 0 0 io_out[19]
port 145 nsew
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1400 0 0 0 io_out[1]
port 146 nsew
flabel metal3 s -800 247670 480 247782 0 FreeSans 1400 0 0 0 io_out[20]
port 147 nsew
flabel metal3 s -800 120048 480 120160 0 FreeSans 1400 0 0 0 io_out[21]
port 148 nsew
flabel metal3 s -800 76826 480 76938 0 FreeSans 1400 0 0 0 io_out[22]
port 149 nsew
flabel metal3 s -800 33604 480 33716 0 FreeSans 1400 0 0 0 io_out[23]
port 150 nsew
flabel metal3 s -800 12182 480 12294 0 FreeSans 1400 0 0 0 io_out[24]
port 151 nsew
flabel metal3 s -800 7454 480 7566 0 FreeSans 1400 0 0 0 io_out[25]
port 152 nsew
flabel metal3 s -800 2726 480 2838 0 FreeSans 1400 0 0 0 io_out[26]
port 153 nsew
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1400 0 0 0 io_out[2]
port 154 nsew
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1400 0 0 0 io_out[3]
port 155 nsew
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1400 0 0 0 io_out[4]
port 156 nsew
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1400 0 0 0 io_out[5]
port 157 nsew
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1400 0 0 0 io_out[6]
port 158 nsew
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1400 0 0 0 io_out[7]
port 159 nsew
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1400 0 0 0 io_out[8]
port 160 nsew
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1400 0 0 0 io_out[9]
port 161 nsew
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1400 90 0 0 la_data_in[0]
port 162 nsew
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1400 90 0 0 la_data_in[100]
port 163 nsew
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1400 90 0 0 la_data_in[101]
port 164 nsew
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1400 90 0 0 la_data_in[102]
port 165 nsew
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1400 90 0 0 la_data_in[103]
port 166 nsew
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1400 90 0 0 la_data_in[104]
port 167 nsew
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1400 90 0 0 la_data_in[105]
port 168 nsew
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1400 90 0 0 la_data_in[106]
port 169 nsew
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1400 90 0 0 la_data_in[107]
port 170 nsew
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1400 90 0 0 la_data_in[108]
port 171 nsew
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1400 90 0 0 la_data_in[109]
port 172 nsew
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1400 90 0 0 la_data_in[10]
port 173 nsew
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1400 90 0 0 la_data_in[110]
port 174 nsew
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1400 90 0 0 la_data_in[111]
port 175 nsew
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1400 90 0 0 la_data_in[112]
port 176 nsew
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1400 90 0 0 la_data_in[113]
port 177 nsew
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1400 90 0 0 la_data_in[114]
port 178 nsew
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1400 90 0 0 la_data_in[115]
port 179 nsew
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1400 90 0 0 la_data_in[116]
port 180 nsew
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1400 90 0 0 la_data_in[117]
port 181 nsew
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1400 90 0 0 la_data_in[118]
port 182 nsew
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1400 90 0 0 la_data_in[119]
port 183 nsew
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1400 90 0 0 la_data_in[11]
port 184 nsew
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1400 90 0 0 la_data_in[120]
port 185 nsew
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1400 90 0 0 la_data_in[121]
port 186 nsew
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1400 90 0 0 la_data_in[122]
port 187 nsew
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1400 90 0 0 la_data_in[123]
port 188 nsew
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1400 90 0 0 la_data_in[124]
port 189 nsew
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1400 90 0 0 la_data_in[125]
port 190 nsew
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1400 90 0 0 la_data_in[126]
port 191 nsew
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1400 90 0 0 la_data_in[127]
port 192 nsew
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1400 90 0 0 la_data_in[12]
port 193 nsew
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1400 90 0 0 la_data_in[13]
port 194 nsew
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1400 90 0 0 la_data_in[14]
port 195 nsew
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1400 90 0 0 la_data_in[15]
port 196 nsew
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1400 90 0 0 la_data_in[16]
port 197 nsew
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1400 90 0 0 la_data_in[17]
port 198 nsew
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1400 90 0 0 la_data_in[18]
port 199 nsew
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1400 90 0 0 la_data_in[19]
port 200 nsew
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1400 90 0 0 la_data_in[1]
port 201 nsew
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1400 90 0 0 la_data_in[20]
port 202 nsew
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1400 90 0 0 la_data_in[21]
port 203 nsew
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1400 90 0 0 la_data_in[22]
port 204 nsew
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1400 90 0 0 la_data_in[23]
port 205 nsew
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1400 90 0 0 la_data_in[24]
port 206 nsew
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1400 90 0 0 la_data_in[25]
port 207 nsew
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1400 90 0 0 la_data_in[26]
port 208 nsew
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1400 90 0 0 la_data_in[27]
port 209 nsew
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1400 90 0 0 la_data_in[28]
port 210 nsew
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1400 90 0 0 la_data_in[29]
port 211 nsew
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1400 90 0 0 la_data_in[2]
port 212 nsew
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1400 90 0 0 la_data_in[30]
port 213 nsew
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1400 90 0 0 la_data_in[31]
port 214 nsew
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1400 90 0 0 la_data_in[32]
port 215 nsew
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1400 90 0 0 la_data_in[33]
port 216 nsew
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1400 90 0 0 la_data_in[34]
port 217 nsew
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1400 90 0 0 la_data_in[35]
port 218 nsew
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1400 90 0 0 la_data_in[36]
port 219 nsew
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1400 90 0 0 la_data_in[37]
port 220 nsew
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1400 90 0 0 la_data_in[38]
port 221 nsew
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1400 90 0 0 la_data_in[39]
port 222 nsew
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1400 90 0 0 la_data_in[3]
port 223 nsew
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1400 90 0 0 la_data_in[40]
port 224 nsew
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1400 90 0 0 la_data_in[41]
port 225 nsew
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1400 90 0 0 la_data_in[42]
port 226 nsew
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1400 90 0 0 la_data_in[43]
port 227 nsew
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1400 90 0 0 la_data_in[44]
port 228 nsew
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1400 90 0 0 la_data_in[45]
port 229 nsew
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1400 90 0 0 la_data_in[46]
port 230 nsew
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1400 90 0 0 la_data_in[47]
port 231 nsew
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1400 90 0 0 la_data_in[48]
port 232 nsew
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1400 90 0 0 la_data_in[49]
port 233 nsew
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1400 90 0 0 la_data_in[4]
port 234 nsew
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1400 90 0 0 la_data_in[50]
port 235 nsew
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1400 90 0 0 la_data_in[51]
port 236 nsew
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1400 90 0 0 la_data_in[52]
port 237 nsew
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1400 90 0 0 la_data_in[53]
port 238 nsew
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1400 90 0 0 la_data_in[54]
port 239 nsew
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1400 90 0 0 la_data_in[55]
port 240 nsew
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1400 90 0 0 la_data_in[56]
port 241 nsew
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1400 90 0 0 la_data_in[57]
port 242 nsew
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1400 90 0 0 la_data_in[58]
port 243 nsew
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1400 90 0 0 la_data_in[59]
port 244 nsew
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1400 90 0 0 la_data_in[5]
port 245 nsew
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1400 90 0 0 la_data_in[60]
port 246 nsew
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1400 90 0 0 la_data_in[61]
port 247 nsew
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1400 90 0 0 la_data_in[62]
port 248 nsew
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1400 90 0 0 la_data_in[63]
port 249 nsew
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1400 90 0 0 la_data_in[64]
port 250 nsew
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1400 90 0 0 la_data_in[65]
port 251 nsew
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1400 90 0 0 la_data_in[66]
port 252 nsew
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1400 90 0 0 la_data_in[67]
port 253 nsew
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1400 90 0 0 la_data_in[68]
port 254 nsew
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1400 90 0 0 la_data_in[69]
port 255 nsew
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1400 90 0 0 la_data_in[6]
port 256 nsew
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1400 90 0 0 la_data_in[70]
port 257 nsew
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1400 90 0 0 la_data_in[71]
port 258 nsew
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1400 90 0 0 la_data_in[72]
port 259 nsew
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1400 90 0 0 la_data_in[73]
port 260 nsew
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1400 90 0 0 la_data_in[74]
port 261 nsew
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1400 90 0 0 la_data_in[75]
port 262 nsew
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1400 90 0 0 la_data_in[76]
port 263 nsew
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1400 90 0 0 la_data_in[77]
port 264 nsew
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1400 90 0 0 la_data_in[78]
port 265 nsew
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1400 90 0 0 la_data_in[79]
port 266 nsew
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1400 90 0 0 la_data_in[7]
port 267 nsew
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1400 90 0 0 la_data_in[80]
port 268 nsew
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1400 90 0 0 la_data_in[81]
port 269 nsew
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1400 90 0 0 la_data_in[82]
port 270 nsew
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1400 90 0 0 la_data_in[83]
port 271 nsew
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1400 90 0 0 la_data_in[84]
port 272 nsew
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1400 90 0 0 la_data_in[85]
port 273 nsew
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1400 90 0 0 la_data_in[86]
port 274 nsew
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1400 90 0 0 la_data_in[87]
port 275 nsew
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1400 90 0 0 la_data_in[88]
port 276 nsew
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1400 90 0 0 la_data_in[89]
port 277 nsew
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1400 90 0 0 la_data_in[8]
port 278 nsew
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1400 90 0 0 la_data_in[90]
port 279 nsew
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1400 90 0 0 la_data_in[91]
port 280 nsew
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1400 90 0 0 la_data_in[92]
port 281 nsew
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1400 90 0 0 la_data_in[93]
port 282 nsew
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1400 90 0 0 la_data_in[94]
port 283 nsew
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1400 90 0 0 la_data_in[95]
port 284 nsew
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1400 90 0 0 la_data_in[96]
port 285 nsew
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1400 90 0 0 la_data_in[97]
port 286 nsew
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1400 90 0 0 la_data_in[98]
port 287 nsew
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1400 90 0 0 la_data_in[99]
port 288 nsew
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1400 90 0 0 la_data_in[9]
port 289 nsew
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1400 90 0 0 la_data_out[0]
port 290 nsew
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1400 90 0 0 la_data_out[100]
port 291 nsew
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1400 90 0 0 la_data_out[101]
port 292 nsew
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1400 90 0 0 la_data_out[102]
port 293 nsew
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1400 90 0 0 la_data_out[103]
port 294 nsew
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1400 90 0 0 la_data_out[104]
port 295 nsew
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1400 90 0 0 la_data_out[105]
port 296 nsew
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1400 90 0 0 la_data_out[106]
port 297 nsew
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1400 90 0 0 la_data_out[107]
port 298 nsew
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1400 90 0 0 la_data_out[108]
port 299 nsew
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1400 90 0 0 la_data_out[109]
port 300 nsew
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1400 90 0 0 la_data_out[10]
port 301 nsew
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1400 90 0 0 la_data_out[110]
port 302 nsew
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1400 90 0 0 la_data_out[111]
port 303 nsew
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1400 90 0 0 la_data_out[112]
port 304 nsew
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1400 90 0 0 la_data_out[113]
port 305 nsew
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1400 90 0 0 la_data_out[114]
port 306 nsew
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1400 90 0 0 la_data_out[115]
port 307 nsew
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1400 90 0 0 la_data_out[116]
port 308 nsew
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1400 90 0 0 la_data_out[117]
port 309 nsew
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1400 90 0 0 la_data_out[118]
port 310 nsew
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1400 90 0 0 la_data_out[119]
port 311 nsew
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1400 90 0 0 la_data_out[11]
port 312 nsew
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1400 90 0 0 la_data_out[120]
port 313 nsew
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1400 90 0 0 la_data_out[121]
port 314 nsew
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1400 90 0 0 la_data_out[122]
port 315 nsew
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1400 90 0 0 la_data_out[123]
port 316 nsew
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1400 90 0 0 la_data_out[124]
port 317 nsew
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1400 90 0 0 la_data_out[125]
port 318 nsew
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1400 90 0 0 la_data_out[126]
port 319 nsew
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1400 90 0 0 la_data_out[127]
port 320 nsew
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1400 90 0 0 la_data_out[12]
port 321 nsew
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1400 90 0 0 la_data_out[13]
port 322 nsew
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1400 90 0 0 la_data_out[14]
port 323 nsew
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1400 90 0 0 la_data_out[15]
port 324 nsew
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1400 90 0 0 la_data_out[16]
port 325 nsew
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1400 90 0 0 la_data_out[17]
port 326 nsew
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1400 90 0 0 la_data_out[18]
port 327 nsew
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1400 90 0 0 la_data_out[19]
port 328 nsew
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1400 90 0 0 la_data_out[1]
port 329 nsew
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1400 90 0 0 la_data_out[20]
port 330 nsew
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1400 90 0 0 la_data_out[21]
port 331 nsew
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1400 90 0 0 la_data_out[22]
port 332 nsew
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1400 90 0 0 la_data_out[23]
port 333 nsew
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1400 90 0 0 la_data_out[24]
port 334 nsew
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1400 90 0 0 la_data_out[25]
port 335 nsew
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1400 90 0 0 la_data_out[26]
port 336 nsew
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1400 90 0 0 la_data_out[27]
port 337 nsew
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1400 90 0 0 la_data_out[28]
port 338 nsew
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1400 90 0 0 la_data_out[29]
port 339 nsew
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1400 90 0 0 la_data_out[2]
port 340 nsew
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1400 90 0 0 la_data_out[30]
port 341 nsew
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1400 90 0 0 la_data_out[31]
port 342 nsew
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1400 90 0 0 la_data_out[32]
port 343 nsew
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1400 90 0 0 la_data_out[33]
port 344 nsew
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1400 90 0 0 la_data_out[34]
port 345 nsew
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1400 90 0 0 la_data_out[35]
port 346 nsew
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1400 90 0 0 la_data_out[36]
port 347 nsew
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1400 90 0 0 la_data_out[37]
port 348 nsew
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1400 90 0 0 la_data_out[38]
port 349 nsew
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1400 90 0 0 la_data_out[39]
port 350 nsew
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1400 90 0 0 la_data_out[3]
port 351 nsew
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1400 90 0 0 la_data_out[40]
port 352 nsew
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1400 90 0 0 la_data_out[41]
port 353 nsew
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1400 90 0 0 la_data_out[42]
port 354 nsew
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1400 90 0 0 la_data_out[43]
port 355 nsew
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1400 90 0 0 la_data_out[44]
port 356 nsew
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1400 90 0 0 la_data_out[45]
port 357 nsew
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1400 90 0 0 la_data_out[46]
port 358 nsew
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1400 90 0 0 la_data_out[47]
port 359 nsew
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1400 90 0 0 la_data_out[48]
port 360 nsew
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1400 90 0 0 la_data_out[49]
port 361 nsew
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1400 90 0 0 la_data_out[4]
port 362 nsew
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1400 90 0 0 la_data_out[50]
port 363 nsew
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1400 90 0 0 la_data_out[51]
port 364 nsew
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1400 90 0 0 la_data_out[52]
port 365 nsew
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1400 90 0 0 la_data_out[53]
port 366 nsew
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1400 90 0 0 la_data_out[54]
port 367 nsew
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1400 90 0 0 la_data_out[55]
port 368 nsew
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1400 90 0 0 la_data_out[56]
port 369 nsew
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1400 90 0 0 la_data_out[57]
port 370 nsew
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1400 90 0 0 la_data_out[58]
port 371 nsew
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1400 90 0 0 la_data_out[59]
port 372 nsew
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1400 90 0 0 la_data_out[5]
port 373 nsew
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1400 90 0 0 la_data_out[60]
port 374 nsew
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1400 90 0 0 la_data_out[61]
port 375 nsew
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1400 90 0 0 la_data_out[62]
port 376 nsew
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1400 90 0 0 la_data_out[63]
port 377 nsew
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1400 90 0 0 la_data_out[64]
port 378 nsew
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1400 90 0 0 la_data_out[65]
port 379 nsew
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1400 90 0 0 la_data_out[66]
port 380 nsew
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1400 90 0 0 la_data_out[67]
port 381 nsew
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1400 90 0 0 la_data_out[68]
port 382 nsew
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1400 90 0 0 la_data_out[69]
port 383 nsew
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1400 90 0 0 la_data_out[6]
port 384 nsew
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1400 90 0 0 la_data_out[70]
port 385 nsew
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1400 90 0 0 la_data_out[71]
port 386 nsew
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1400 90 0 0 la_data_out[72]
port 387 nsew
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1400 90 0 0 la_data_out[73]
port 388 nsew
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1400 90 0 0 la_data_out[74]
port 389 nsew
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1400 90 0 0 la_data_out[75]
port 390 nsew
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1400 90 0 0 la_data_out[76]
port 391 nsew
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1400 90 0 0 la_data_out[77]
port 392 nsew
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1400 90 0 0 la_data_out[78]
port 393 nsew
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1400 90 0 0 la_data_out[79]
port 394 nsew
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1400 90 0 0 la_data_out[7]
port 395 nsew
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1400 90 0 0 la_data_out[80]
port 396 nsew
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1400 90 0 0 la_data_out[81]
port 397 nsew
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1400 90 0 0 la_data_out[82]
port 398 nsew
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1400 90 0 0 la_data_out[83]
port 399 nsew
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1400 90 0 0 la_data_out[84]
port 400 nsew
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1400 90 0 0 la_data_out[85]
port 401 nsew
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1400 90 0 0 la_data_out[86]
port 402 nsew
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1400 90 0 0 la_data_out[87]
port 403 nsew
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1400 90 0 0 la_data_out[88]
port 404 nsew
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1400 90 0 0 la_data_out[89]
port 405 nsew
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1400 90 0 0 la_data_out[8]
port 406 nsew
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1400 90 0 0 la_data_out[90]
port 407 nsew
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1400 90 0 0 la_data_out[91]
port 408 nsew
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1400 90 0 0 la_data_out[92]
port 409 nsew
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1400 90 0 0 la_data_out[93]
port 410 nsew
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1400 90 0 0 la_data_out[94]
port 411 nsew
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1400 90 0 0 la_data_out[95]
port 412 nsew
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1400 90 0 0 la_data_out[96]
port 413 nsew
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1400 90 0 0 la_data_out[97]
port 414 nsew
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1400 90 0 0 la_data_out[98]
port 415 nsew
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1400 90 0 0 la_data_out[99]
port 416 nsew
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1400 90 0 0 la_data_out[9]
port 417 nsew
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1400 90 0 0 la_oenb[0]
port 418 nsew
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1400 90 0 0 la_oenb[100]
port 419 nsew
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1400 90 0 0 la_oenb[101]
port 420 nsew
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1400 90 0 0 la_oenb[102]
port 421 nsew
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1400 90 0 0 la_oenb[103]
port 422 nsew
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1400 90 0 0 la_oenb[104]
port 423 nsew
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1400 90 0 0 la_oenb[105]
port 424 nsew
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1400 90 0 0 la_oenb[106]
port 425 nsew
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1400 90 0 0 la_oenb[107]
port 426 nsew
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1400 90 0 0 la_oenb[108]
port 427 nsew
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1400 90 0 0 la_oenb[109]
port 428 nsew
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1400 90 0 0 la_oenb[10]
port 429 nsew
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1400 90 0 0 la_oenb[110]
port 430 nsew
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1400 90 0 0 la_oenb[111]
port 431 nsew
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1400 90 0 0 la_oenb[112]
port 432 nsew
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1400 90 0 0 la_oenb[113]
port 433 nsew
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1400 90 0 0 la_oenb[114]
port 434 nsew
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1400 90 0 0 la_oenb[115]
port 435 nsew
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1400 90 0 0 la_oenb[116]
port 436 nsew
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1400 90 0 0 la_oenb[117]
port 437 nsew
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1400 90 0 0 la_oenb[118]
port 438 nsew
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1400 90 0 0 la_oenb[119]
port 439 nsew
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1400 90 0 0 la_oenb[11]
port 440 nsew
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1400 90 0 0 la_oenb[120]
port 441 nsew
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1400 90 0 0 la_oenb[121]
port 442 nsew
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1400 90 0 0 la_oenb[122]
port 443 nsew
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1400 90 0 0 la_oenb[123]
port 444 nsew
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1400 90 0 0 la_oenb[124]
port 445 nsew
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1400 90 0 0 la_oenb[125]
port 446 nsew
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1400 90 0 0 la_oenb[126]
port 447 nsew
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1400 90 0 0 la_oenb[127]
port 448 nsew
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1400 90 0 0 la_oenb[12]
port 449 nsew
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1400 90 0 0 la_oenb[13]
port 450 nsew
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1400 90 0 0 la_oenb[14]
port 451 nsew
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1400 90 0 0 la_oenb[15]
port 452 nsew
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1400 90 0 0 la_oenb[16]
port 453 nsew
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1400 90 0 0 la_oenb[17]
port 454 nsew
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1400 90 0 0 la_oenb[18]
port 455 nsew
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1400 90 0 0 la_oenb[19]
port 456 nsew
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1400 90 0 0 la_oenb[1]
port 457 nsew
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1400 90 0 0 la_oenb[20]
port 458 nsew
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1400 90 0 0 la_oenb[21]
port 459 nsew
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1400 90 0 0 la_oenb[22]
port 460 nsew
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1400 90 0 0 la_oenb[23]
port 461 nsew
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1400 90 0 0 la_oenb[24]
port 462 nsew
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1400 90 0 0 la_oenb[25]
port 463 nsew
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1400 90 0 0 la_oenb[26]
port 464 nsew
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1400 90 0 0 la_oenb[27]
port 465 nsew
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1400 90 0 0 la_oenb[28]
port 466 nsew
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1400 90 0 0 la_oenb[29]
port 467 nsew
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1400 90 0 0 la_oenb[2]
port 468 nsew
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1400 90 0 0 la_oenb[30]
port 469 nsew
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1400 90 0 0 la_oenb[31]
port 470 nsew
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1400 90 0 0 la_oenb[32]
port 471 nsew
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1400 90 0 0 la_oenb[33]
port 472 nsew
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1400 90 0 0 la_oenb[34]
port 473 nsew
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1400 90 0 0 la_oenb[35]
port 474 nsew
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1400 90 0 0 la_oenb[36]
port 475 nsew
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1400 90 0 0 la_oenb[37]
port 476 nsew
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1400 90 0 0 la_oenb[38]
port 477 nsew
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1400 90 0 0 la_oenb[39]
port 478 nsew
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1400 90 0 0 la_oenb[3]
port 479 nsew
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1400 90 0 0 la_oenb[40]
port 480 nsew
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1400 90 0 0 la_oenb[41]
port 481 nsew
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1400 90 0 0 la_oenb[42]
port 482 nsew
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1400 90 0 0 la_oenb[43]
port 483 nsew
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1400 90 0 0 la_oenb[44]
port 484 nsew
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1400 90 0 0 la_oenb[45]
port 485 nsew
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1400 90 0 0 la_oenb[46]
port 486 nsew
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1400 90 0 0 la_oenb[47]
port 487 nsew
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1400 90 0 0 la_oenb[48]
port 488 nsew
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1400 90 0 0 la_oenb[49]
port 489 nsew
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1400 90 0 0 la_oenb[4]
port 490 nsew
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1400 90 0 0 la_oenb[50]
port 491 nsew
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1400 90 0 0 la_oenb[51]
port 492 nsew
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1400 90 0 0 la_oenb[52]
port 493 nsew
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1400 90 0 0 la_oenb[53]
port 494 nsew
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1400 90 0 0 la_oenb[54]
port 495 nsew
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1400 90 0 0 la_oenb[55]
port 496 nsew
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1400 90 0 0 la_oenb[56]
port 497 nsew
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1400 90 0 0 la_oenb[57]
port 498 nsew
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1400 90 0 0 la_oenb[58]
port 499 nsew
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1400 90 0 0 la_oenb[59]
port 500 nsew
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1400 90 0 0 la_oenb[5]
port 501 nsew
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1400 90 0 0 la_oenb[60]
port 502 nsew
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1400 90 0 0 la_oenb[61]
port 503 nsew
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1400 90 0 0 la_oenb[62]
port 504 nsew
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1400 90 0 0 la_oenb[63]
port 505 nsew
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1400 90 0 0 la_oenb[64]
port 506 nsew
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1400 90 0 0 la_oenb[65]
port 507 nsew
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1400 90 0 0 la_oenb[66]
port 508 nsew
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1400 90 0 0 la_oenb[67]
port 509 nsew
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1400 90 0 0 la_oenb[68]
port 510 nsew
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1400 90 0 0 la_oenb[69]
port 511 nsew
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1400 90 0 0 la_oenb[6]
port 512 nsew
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1400 90 0 0 la_oenb[70]
port 513 nsew
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1400 90 0 0 la_oenb[71]
port 514 nsew
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1400 90 0 0 la_oenb[72]
port 515 nsew
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1400 90 0 0 la_oenb[73]
port 516 nsew
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1400 90 0 0 la_oenb[74]
port 517 nsew
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1400 90 0 0 la_oenb[75]
port 518 nsew
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1400 90 0 0 la_oenb[76]
port 519 nsew
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1400 90 0 0 la_oenb[77]
port 520 nsew
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1400 90 0 0 la_oenb[78]
port 521 nsew
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1400 90 0 0 la_oenb[79]
port 522 nsew
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1400 90 0 0 la_oenb[7]
port 523 nsew
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1400 90 0 0 la_oenb[80]
port 524 nsew
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1400 90 0 0 la_oenb[81]
port 525 nsew
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1400 90 0 0 la_oenb[82]
port 526 nsew
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1400 90 0 0 la_oenb[83]
port 527 nsew
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1400 90 0 0 la_oenb[84]
port 528 nsew
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1400 90 0 0 la_oenb[85]
port 529 nsew
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1400 90 0 0 la_oenb[86]
port 530 nsew
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1400 90 0 0 la_oenb[87]
port 531 nsew
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1400 90 0 0 la_oenb[88]
port 532 nsew
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1400 90 0 0 la_oenb[89]
port 533 nsew
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1400 90 0 0 la_oenb[8]
port 534 nsew
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1400 90 0 0 la_oenb[90]
port 535 nsew
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1400 90 0 0 la_oenb[91]
port 536 nsew
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1400 90 0 0 la_oenb[92]
port 537 nsew
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1400 90 0 0 la_oenb[93]
port 538 nsew
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1400 90 0 0 la_oenb[94]
port 539 nsew
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1400 90 0 0 la_oenb[95]
port 540 nsew
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1400 90 0 0 la_oenb[96]
port 541 nsew
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1400 90 0 0 la_oenb[97]
port 542 nsew
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1400 90 0 0 la_oenb[98]
port 543 nsew
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1400 90 0 0 la_oenb[99]
port 544 nsew
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1400 90 0 0 la_oenb[9]
port 545 nsew
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1400 90 0 0 user_clock2
port 546 nsew
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1400 90 0 0 user_irq[0]
port 547 nsew
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1400 90 0 0 user_irq[1]
port 548 nsew
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1400 90 0 0 user_irq[2]
port 549 nsew
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1400 0 0 0 vccd1
port 550 nsew
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1400 0 0 0 vccd1
port 550 nsew
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1400 0 0 0 vccd2
port 551 nsew
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1400 0 0 0 vccd2
port 551 nsew
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1400 0 0 0 vdda2
port 553 nsew
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1400 0 0 0 vdda2
port 553 nsew
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 2400 180 0 0 vssa1
port 554 nsew
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 2400 180 0 0 vssa1
port 554 nsew
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1400 0 0 0 vssa1
port 554 nsew
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1400 0 0 0 vssa1
port 554 nsew
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1400 0 0 0 vssa2
port 555 nsew
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1400 0 0 0 vssa2
port 555 nsew
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1400 0 0 0 vssd1
port 556 nsew
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1400 0 0 0 vssd1
port 556 nsew
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1400 0 0 0 vssd2
port 557 nsew
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1400 0 0 0 vssd2
port 557 nsew
flabel metal2 s 524 -800 636 480 0 FreeSans 1400 90 0 0 wb_clk_i
port 558 nsew
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1400 90 0 0 wb_rst_i
port 559 nsew
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1400 90 0 0 wbs_ack_o
port 560 nsew
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1400 90 0 0 wbs_adr_i[0]
port 561 nsew
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1400 90 0 0 wbs_adr_i[10]
port 562 nsew
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1400 90 0 0 wbs_adr_i[11]
port 563 nsew
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1400 90 0 0 wbs_adr_i[12]
port 564 nsew
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1400 90 0 0 wbs_adr_i[13]
port 565 nsew
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1400 90 0 0 wbs_adr_i[14]
port 566 nsew
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1400 90 0 0 wbs_adr_i[15]
port 567 nsew
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1400 90 0 0 wbs_adr_i[16]
port 568 nsew
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1400 90 0 0 wbs_adr_i[17]
port 569 nsew
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1400 90 0 0 wbs_adr_i[18]
port 570 nsew
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1400 90 0 0 wbs_adr_i[19]
port 571 nsew
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1400 90 0 0 wbs_adr_i[1]
port 572 nsew
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1400 90 0 0 wbs_adr_i[20]
port 573 nsew
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1400 90 0 0 wbs_adr_i[21]
port 574 nsew
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1400 90 0 0 wbs_adr_i[22]
port 575 nsew
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1400 90 0 0 wbs_adr_i[23]
port 576 nsew
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1400 90 0 0 wbs_adr_i[24]
port 577 nsew
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1400 90 0 0 wbs_adr_i[25]
port 578 nsew
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1400 90 0 0 wbs_adr_i[26]
port 579 nsew
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1400 90 0 0 wbs_adr_i[27]
port 580 nsew
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1400 90 0 0 wbs_adr_i[28]
port 581 nsew
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1400 90 0 0 wbs_adr_i[29]
port 582 nsew
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1400 90 0 0 wbs_adr_i[2]
port 583 nsew
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1400 90 0 0 wbs_adr_i[30]
port 584 nsew
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1400 90 0 0 wbs_adr_i[31]
port 585 nsew
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1400 90 0 0 wbs_adr_i[3]
port 586 nsew
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1400 90 0 0 wbs_adr_i[4]
port 587 nsew
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1400 90 0 0 wbs_adr_i[5]
port 588 nsew
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1400 90 0 0 wbs_adr_i[6]
port 589 nsew
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1400 90 0 0 wbs_adr_i[7]
port 590 nsew
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1400 90 0 0 wbs_adr_i[8]
port 591 nsew
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1400 90 0 0 wbs_adr_i[9]
port 592 nsew
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1400 90 0 0 wbs_cyc_i
port 593 nsew
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1400 90 0 0 wbs_dat_i[0]
port 594 nsew
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1400 90 0 0 wbs_dat_i[10]
port 595 nsew
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1400 90 0 0 wbs_dat_i[11]
port 596 nsew
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1400 90 0 0 wbs_dat_i[12]
port 597 nsew
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1400 90 0 0 wbs_dat_i[13]
port 598 nsew
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1400 90 0 0 wbs_dat_i[14]
port 599 nsew
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1400 90 0 0 wbs_dat_i[15]
port 600 nsew
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1400 90 0 0 wbs_dat_i[16]
port 601 nsew
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1400 90 0 0 wbs_dat_i[17]
port 602 nsew
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1400 90 0 0 wbs_dat_i[18]
port 603 nsew
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1400 90 0 0 wbs_dat_i[19]
port 604 nsew
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1400 90 0 0 wbs_dat_i[1]
port 605 nsew
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1400 90 0 0 wbs_dat_i[20]
port 606 nsew
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1400 90 0 0 wbs_dat_i[21]
port 607 nsew
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1400 90 0 0 wbs_dat_i[22]
port 608 nsew
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1400 90 0 0 wbs_dat_i[23]
port 609 nsew
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1400 90 0 0 wbs_dat_i[24]
port 610 nsew
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1400 90 0 0 wbs_dat_i[25]
port 611 nsew
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1400 90 0 0 wbs_dat_i[26]
port 612 nsew
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1400 90 0 0 wbs_dat_i[27]
port 613 nsew
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1400 90 0 0 wbs_dat_i[28]
port 614 nsew
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1400 90 0 0 wbs_dat_i[29]
port 615 nsew
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1400 90 0 0 wbs_dat_i[2]
port 616 nsew
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1400 90 0 0 wbs_dat_i[30]
port 617 nsew
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1400 90 0 0 wbs_dat_i[31]
port 618 nsew
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1400 90 0 0 wbs_dat_i[3]
port 619 nsew
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1400 90 0 0 wbs_dat_i[4]
port 620 nsew
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1400 90 0 0 wbs_dat_i[5]
port 621 nsew
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1400 90 0 0 wbs_dat_i[6]
port 622 nsew
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1400 90 0 0 wbs_dat_i[7]
port 623 nsew
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1400 90 0 0 wbs_dat_i[8]
port 624 nsew
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1400 90 0 0 wbs_dat_i[9]
port 625 nsew
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1400 90 0 0 wbs_dat_o[0]
port 626 nsew
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1400 90 0 0 wbs_dat_o[10]
port 627 nsew
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1400 90 0 0 wbs_dat_o[11]
port 628 nsew
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1400 90 0 0 wbs_dat_o[12]
port 629 nsew
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1400 90 0 0 wbs_dat_o[13]
port 630 nsew
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1400 90 0 0 wbs_dat_o[14]
port 631 nsew
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1400 90 0 0 wbs_dat_o[15]
port 632 nsew
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1400 90 0 0 wbs_dat_o[16]
port 633 nsew
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1400 90 0 0 wbs_dat_o[17]
port 634 nsew
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1400 90 0 0 wbs_dat_o[18]
port 635 nsew
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1400 90 0 0 wbs_dat_o[19]
port 636 nsew
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1400 90 0 0 wbs_dat_o[1]
port 637 nsew
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1400 90 0 0 wbs_dat_o[20]
port 638 nsew
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1400 90 0 0 wbs_dat_o[21]
port 639 nsew
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1400 90 0 0 wbs_dat_o[22]
port 640 nsew
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1400 90 0 0 wbs_dat_o[23]
port 641 nsew
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1400 90 0 0 wbs_dat_o[24]
port 642 nsew
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1400 90 0 0 wbs_dat_o[25]
port 643 nsew
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1400 90 0 0 wbs_dat_o[26]
port 644 nsew
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1400 90 0 0 wbs_dat_o[27]
port 645 nsew
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1400 90 0 0 wbs_dat_o[28]
port 646 nsew
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1400 90 0 0 wbs_dat_o[29]
port 647 nsew
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1400 90 0 0 wbs_dat_o[2]
port 648 nsew
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1400 90 0 0 wbs_dat_o[30]
port 649 nsew
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1400 90 0 0 wbs_dat_o[31]
port 650 nsew
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1400 90 0 0 wbs_dat_o[3]
port 651 nsew
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1400 90 0 0 wbs_dat_o[4]
port 652 nsew
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1400 90 0 0 wbs_dat_o[5]
port 653 nsew
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1400 90 0 0 wbs_dat_o[6]
port 654 nsew
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1400 90 0 0 wbs_dat_o[7]
port 655 nsew
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1400 90 0 0 wbs_dat_o[8]
port 656 nsew
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1400 90 0 0 wbs_dat_o[9]
port 657 nsew
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1400 90 0 0 wbs_sel_i[0]
port 658 nsew
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1400 90 0 0 wbs_sel_i[1]
port 659 nsew
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1400 90 0 0 wbs_sel_i[2]
port 660 nsew
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1400 90 0 0 wbs_sel_i[3]
port 661 nsew
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1400 90 0 0 wbs_stb_i
port 662 nsew
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1400 90 0 0 wbs_we_i
port 663 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
