magic
tech sky130A
magscale 1 2
timestamp 1654711683
<< error_p >>
rect -855 -347 -797 -341
rect -737 -347 -679 -341
rect -619 -347 -561 -341
rect -501 -347 -443 -341
rect -383 -347 -325 -341
rect -265 -347 -207 -341
rect -147 -347 -89 -341
rect -29 -347 29 -341
rect 89 -347 147 -341
rect 207 -347 265 -341
rect 325 -347 383 -341
rect 443 -347 501 -341
rect 561 -347 619 -341
rect 679 -347 737 -341
rect 797 -347 855 -341
rect -855 -381 -843 -347
rect -737 -381 -725 -347
rect -619 -381 -607 -347
rect -501 -381 -489 -347
rect -383 -381 -371 -347
rect -265 -381 -253 -347
rect -147 -381 -135 -347
rect -29 -381 -17 -347
rect 89 -381 101 -347
rect 207 -381 219 -347
rect 325 -381 337 -347
rect 443 -381 455 -347
rect 561 -381 573 -347
rect 679 -381 691 -347
rect 797 -381 809 -347
rect -855 -387 -797 -381
rect -737 -387 -679 -381
rect -619 -387 -561 -381
rect -501 -387 -443 -381
rect -383 -387 -325 -381
rect -265 -387 -207 -381
rect -147 -387 -89 -381
rect -29 -387 29 -381
rect 89 -387 147 -381
rect 207 -387 265 -381
rect 325 -387 383 -381
rect 443 -387 501 -381
rect 561 -387 619 -381
rect 679 -387 737 -381
rect 797 -387 855 -381
<< nwell >>
rect -1052 -519 1052 519
<< pmos >>
rect -856 -300 -796 300
rect -738 -300 -678 300
rect -620 -300 -560 300
rect -502 -300 -442 300
rect -384 -300 -324 300
rect -266 -300 -206 300
rect -148 -300 -88 300
rect -30 -300 30 300
rect 88 -300 148 300
rect 206 -300 266 300
rect 324 -300 384 300
rect 442 -300 502 300
rect 560 -300 620 300
rect 678 -300 738 300
rect 796 -300 856 300
<< pdiff >>
rect -914 288 -856 300
rect -914 -288 -902 288
rect -868 -288 -856 288
rect -914 -300 -856 -288
rect -796 288 -738 300
rect -796 -288 -784 288
rect -750 -288 -738 288
rect -796 -300 -738 -288
rect -678 288 -620 300
rect -678 -288 -666 288
rect -632 -288 -620 288
rect -678 -300 -620 -288
rect -560 288 -502 300
rect -560 -288 -548 288
rect -514 -288 -502 288
rect -560 -300 -502 -288
rect -442 288 -384 300
rect -442 -288 -430 288
rect -396 -288 -384 288
rect -442 -300 -384 -288
rect -324 288 -266 300
rect -324 -288 -312 288
rect -278 -288 -266 288
rect -324 -300 -266 -288
rect -206 288 -148 300
rect -206 -288 -194 288
rect -160 -288 -148 288
rect -206 -300 -148 -288
rect -88 288 -30 300
rect -88 -288 -76 288
rect -42 -288 -30 288
rect -88 -300 -30 -288
rect 30 288 88 300
rect 30 -288 42 288
rect 76 -288 88 288
rect 30 -300 88 -288
rect 148 288 206 300
rect 148 -288 160 288
rect 194 -288 206 288
rect 148 -300 206 -288
rect 266 288 324 300
rect 266 -288 278 288
rect 312 -288 324 288
rect 266 -300 324 -288
rect 384 288 442 300
rect 384 -288 396 288
rect 430 -288 442 288
rect 384 -300 442 -288
rect 502 288 560 300
rect 502 -288 514 288
rect 548 -288 560 288
rect 502 -300 560 -288
rect 620 288 678 300
rect 620 -288 632 288
rect 666 -288 678 288
rect 620 -300 678 -288
rect 738 288 796 300
rect 738 -288 750 288
rect 784 -288 796 288
rect 738 -300 796 -288
rect 856 288 914 300
rect 856 -288 868 288
rect 902 -288 914 288
rect 856 -300 914 -288
<< pdiffc >>
rect -902 -288 -868 288
rect -784 -288 -750 288
rect -666 -288 -632 288
rect -548 -288 -514 288
rect -430 -288 -396 288
rect -312 -288 -278 288
rect -194 -288 -160 288
rect -76 -288 -42 288
rect 42 -288 76 288
rect 160 -288 194 288
rect 278 -288 312 288
rect 396 -288 430 288
rect 514 -288 548 288
rect 632 -288 666 288
rect 750 -288 784 288
rect 868 -288 902 288
<< nsubdiff >>
rect -1016 449 -920 483
rect 920 449 1016 483
rect -1016 387 -982 449
rect 982 387 1016 449
rect -1016 -449 -982 -387
rect 982 -449 1016 -387
rect -1016 -483 -920 -449
rect 920 -483 1016 -449
<< nsubdiffcont >>
rect -920 449 920 483
rect -1016 -387 -982 387
rect 982 -387 1016 387
rect -920 -483 920 -449
<< poly >>
rect -731 397 -682 399
rect -859 331 -793 397
rect -741 331 -675 397
rect -623 331 -557 397
rect -505 331 -439 397
rect -387 331 -321 397
rect -269 331 -203 397
rect -151 331 -85 397
rect -33 331 33 397
rect 85 331 151 397
rect 203 331 269 397
rect 321 331 387 397
rect 439 331 505 397
rect 557 331 623 397
rect 675 331 741 397
rect 793 331 859 397
rect -856 300 -796 331
rect -738 300 -678 331
rect -620 300 -560 331
rect -502 300 -442 331
rect -384 300 -324 331
rect -266 300 -206 331
rect -148 300 -88 331
rect -30 300 30 331
rect 88 300 148 331
rect 206 300 266 331
rect 324 300 384 331
rect 442 300 502 331
rect 560 300 620 331
rect 678 300 738 331
rect 796 300 856 331
rect -856 -331 -796 -300
rect -738 -331 -678 -300
rect -620 -331 -560 -300
rect -502 -331 -442 -300
rect -384 -331 -324 -300
rect -266 -331 -206 -300
rect -148 -331 -88 -300
rect -30 -331 30 -300
rect 88 -331 148 -300
rect 206 -331 266 -300
rect 324 -331 384 -300
rect 442 -331 502 -300
rect 560 -331 620 -300
rect 678 -331 738 -300
rect 796 -331 856 -300
rect -859 -347 -793 -331
rect -859 -381 -843 -347
rect -809 -381 -793 -347
rect -859 -397 -793 -381
rect -741 -347 -675 -331
rect -741 -381 -725 -347
rect -691 -381 -675 -347
rect -741 -397 -675 -381
rect -623 -347 -557 -331
rect -623 -381 -607 -347
rect -573 -381 -557 -347
rect -623 -397 -557 -381
rect -505 -347 -439 -331
rect -505 -381 -489 -347
rect -455 -381 -439 -347
rect -505 -397 -439 -381
rect -387 -347 -321 -331
rect -387 -381 -371 -347
rect -337 -381 -321 -347
rect -387 -397 -321 -381
rect -269 -347 -203 -331
rect -269 -381 -253 -347
rect -219 -381 -203 -347
rect -269 -397 -203 -381
rect -151 -347 -85 -331
rect -151 -381 -135 -347
rect -101 -381 -85 -347
rect -151 -397 -85 -381
rect -33 -347 33 -331
rect -33 -381 -17 -347
rect 17 -381 33 -347
rect -33 -397 33 -381
rect 85 -347 151 -331
rect 85 -381 101 -347
rect 135 -381 151 -347
rect 85 -397 151 -381
rect 203 -347 269 -331
rect 203 -381 219 -347
rect 253 -381 269 -347
rect 203 -397 269 -381
rect 321 -347 387 -331
rect 321 -381 337 -347
rect 371 -381 387 -347
rect 321 -397 387 -381
rect 439 -347 505 -331
rect 439 -381 455 -347
rect 489 -381 505 -347
rect 439 -397 505 -381
rect 557 -347 623 -331
rect 557 -381 573 -347
rect 607 -381 623 -347
rect 557 -397 623 -381
rect 675 -347 741 -331
rect 675 -381 691 -347
rect 725 -381 741 -347
rect 675 -397 741 -381
rect 793 -347 859 -331
rect 793 -381 809 -347
rect 843 -381 859 -347
rect 793 -397 859 -381
<< polycont >>
rect -843 -381 -809 -347
rect -725 -381 -691 -347
rect -607 -381 -573 -347
rect -489 -381 -455 -347
rect -371 -381 -337 -347
rect -253 -381 -219 -347
rect -135 -381 -101 -347
rect -17 -381 17 -347
rect 101 -381 135 -347
rect 219 -381 253 -347
rect 337 -381 371 -347
rect 455 -381 489 -347
rect 573 -381 607 -347
rect 691 -381 725 -347
rect 809 -381 843 -347
<< locali >>
rect -1016 449 -920 483
rect 920 449 1016 483
rect -1016 387 -982 449
rect 982 387 1016 449
rect -902 288 -868 304
rect -902 -304 -868 -288
rect -784 288 -750 304
rect -784 -304 -750 -288
rect -666 288 -632 304
rect -666 -304 -632 -288
rect -548 288 -514 304
rect -548 -304 -514 -288
rect -430 288 -396 304
rect -430 -304 -396 -288
rect -312 288 -278 304
rect -312 -304 -278 -288
rect -194 288 -160 304
rect -194 -304 -160 -288
rect -76 288 -42 304
rect -76 -304 -42 -288
rect 42 288 76 304
rect 42 -304 76 -288
rect 160 288 194 304
rect 160 -304 194 -288
rect 278 288 312 304
rect 278 -304 312 -288
rect 396 288 430 304
rect 396 -304 430 -288
rect 514 288 548 304
rect 514 -304 548 -288
rect 632 288 666 304
rect 632 -304 666 -288
rect 750 288 784 304
rect 750 -304 784 -288
rect 868 288 902 304
rect 868 -304 902 -288
rect -859 -381 -843 -347
rect -809 -381 -793 -347
rect -741 -381 -725 -347
rect -691 -381 -675 -347
rect -623 -381 -607 -347
rect -573 -381 -557 -347
rect -505 -381 -489 -347
rect -455 -381 -439 -347
rect -387 -381 -371 -347
rect -337 -381 -321 -347
rect -269 -381 -253 -347
rect -219 -381 -203 -347
rect -151 -381 -135 -347
rect -101 -381 -85 -347
rect -33 -381 -17 -347
rect 17 -381 33 -347
rect 85 -381 101 -347
rect 135 -381 151 -347
rect 203 -381 219 -347
rect 253 -381 269 -347
rect 321 -381 337 -347
rect 371 -381 387 -347
rect 439 -381 455 -347
rect 489 -381 505 -347
rect 557 -381 573 -347
rect 607 -381 623 -347
rect 675 -381 691 -347
rect 725 -381 741 -347
rect 793 -381 809 -347
rect 843 -381 859 -347
rect -1016 -449 -982 -387
rect 982 -449 1016 -387
rect -1016 -483 -920 -449
rect 920 -483 1016 -449
<< viali >>
rect -902 -288 -868 288
rect -784 -288 -750 288
rect -666 -288 -632 288
rect -548 -288 -514 288
rect -430 -288 -396 288
rect -312 -288 -278 288
rect -194 -288 -160 288
rect -76 -288 -42 288
rect 42 -288 76 288
rect 160 -288 194 288
rect 278 -288 312 288
rect 396 -288 430 288
rect 514 -288 548 288
rect 632 -288 666 288
rect 750 -288 784 288
rect 868 -288 902 288
rect -843 -381 -809 -347
rect -725 -381 -691 -347
rect -607 -381 -573 -347
rect -489 -381 -455 -347
rect -371 -381 -337 -347
rect -253 -381 -219 -347
rect -135 -381 -101 -347
rect -17 -381 17 -347
rect 101 -381 135 -347
rect 219 -381 253 -347
rect 337 -381 371 -347
rect 455 -381 489 -347
rect 573 -381 607 -347
rect 691 -381 725 -347
rect 809 -381 843 -347
<< metal1 >>
rect -908 288 -862 300
rect -908 -288 -902 288
rect -868 -288 -862 288
rect -908 -300 -862 -288
rect -790 288 -744 300
rect -790 -288 -784 288
rect -750 -288 -744 288
rect -790 -300 -744 -288
rect -672 288 -626 300
rect -672 -288 -666 288
rect -632 -288 -626 288
rect -672 -300 -626 -288
rect -554 288 -508 300
rect -554 -288 -548 288
rect -514 -288 -508 288
rect -554 -300 -508 -288
rect -436 288 -390 300
rect -436 -288 -430 288
rect -396 -288 -390 288
rect -436 -300 -390 -288
rect -318 288 -272 300
rect -318 -288 -312 288
rect -278 -288 -272 288
rect -318 -300 -272 -288
rect -200 288 -154 300
rect -200 -288 -194 288
rect -160 -288 -154 288
rect -200 -300 -154 -288
rect -82 288 -36 300
rect -82 -288 -76 288
rect -42 -288 -36 288
rect -82 -300 -36 -288
rect 36 288 82 300
rect 36 -288 42 288
rect 76 -288 82 288
rect 36 -300 82 -288
rect 154 288 200 300
rect 154 -288 160 288
rect 194 -288 200 288
rect 154 -300 200 -288
rect 272 288 318 300
rect 272 -288 278 288
rect 312 -288 318 288
rect 272 -300 318 -288
rect 390 288 436 300
rect 390 -288 396 288
rect 430 -288 436 288
rect 390 -300 436 -288
rect 508 288 554 300
rect 508 -288 514 288
rect 548 -288 554 288
rect 508 -300 554 -288
rect 626 288 672 300
rect 626 -288 632 288
rect 666 -288 672 288
rect 626 -300 672 -288
rect 744 288 790 300
rect 744 -288 750 288
rect 784 -288 790 288
rect 744 -300 790 -288
rect 862 288 908 300
rect 862 -288 868 288
rect 902 -288 908 288
rect 862 -300 908 -288
rect -855 -347 -797 -341
rect -855 -381 -843 -347
rect -809 -381 -797 -347
rect -855 -387 -797 -381
rect -737 -347 -679 -341
rect -737 -381 -725 -347
rect -691 -381 -679 -347
rect -737 -387 -679 -381
rect -619 -347 -561 -341
rect -619 -381 -607 -347
rect -573 -381 -561 -347
rect -619 -387 -561 -381
rect -501 -347 -443 -341
rect -501 -381 -489 -347
rect -455 -381 -443 -347
rect -501 -387 -443 -381
rect -383 -347 -325 -341
rect -383 -381 -371 -347
rect -337 -381 -325 -347
rect -383 -387 -325 -381
rect -265 -347 -207 -341
rect -265 -381 -253 -347
rect -219 -381 -207 -347
rect -265 -387 -207 -381
rect -147 -347 -89 -341
rect -147 -381 -135 -347
rect -101 -381 -89 -347
rect -147 -387 -89 -381
rect -29 -347 29 -341
rect -29 -381 -17 -347
rect 17 -381 29 -347
rect -29 -387 29 -381
rect 89 -347 147 -341
rect 89 -381 101 -347
rect 135 -381 147 -347
rect 89 -387 147 -381
rect 207 -347 265 -341
rect 207 -381 219 -347
rect 253 -381 265 -347
rect 207 -387 265 -381
rect 325 -347 383 -341
rect 325 -381 337 -347
rect 371 -381 383 -347
rect 325 -387 383 -381
rect 443 -347 501 -341
rect 443 -381 455 -347
rect 489 -381 501 -347
rect 443 -387 501 -381
rect 561 -347 619 -341
rect 561 -381 573 -347
rect 607 -381 619 -347
rect 561 -387 619 -381
rect 679 -347 737 -341
rect 679 -381 691 -347
rect 725 -381 737 -347
rect 679 -387 737 -381
rect 797 -347 855 -341
rect 797 -381 809 -347
rect 843 -381 855 -347
rect 797 -387 855 -381
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -999 -466 999 466
string parameters w 3 l 0.3 m 1 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
