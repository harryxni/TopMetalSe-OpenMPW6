magic
tech sky130A
magscale 1 2
timestamp 1654643737
<< error_p >>
rect -855 71 -797 77
rect -737 71 -679 77
rect -619 71 -561 77
rect -501 71 -443 77
rect -383 71 -325 77
rect -265 71 -207 77
rect -147 71 -89 77
rect -29 71 29 77
rect 89 71 147 77
rect 207 71 265 77
rect 325 71 383 77
rect 443 71 501 77
rect 561 71 619 77
rect 679 71 737 77
rect 797 71 855 77
rect -855 37 -843 71
rect -737 37 -725 71
rect -619 37 -607 71
rect -501 37 -489 71
rect -383 37 -371 71
rect -265 37 -253 71
rect -147 37 -135 71
rect -29 37 -17 71
rect 89 37 101 71
rect 207 37 219 71
rect 325 37 337 71
rect 443 37 455 71
rect 561 37 573 71
rect 679 37 691 71
rect 797 37 809 71
rect -855 31 -797 37
rect -737 31 -679 37
rect -619 31 -561 37
rect -501 31 -443 37
rect -383 31 -325 37
rect -265 31 -207 37
rect -147 31 -89 37
rect -29 31 29 37
rect 89 31 147 37
rect 207 31 265 37
rect 325 31 383 37
rect 443 31 501 37
rect 561 31 619 37
rect 679 31 737 37
rect 797 31 855 37
rect -855 -37 -797 -31
rect -737 -37 -679 -31
rect -619 -37 -561 -31
rect -501 -37 -443 -31
rect -383 -37 -325 -31
rect -265 -37 -207 -31
rect -147 -37 -89 -31
rect -29 -37 29 -31
rect 89 -37 147 -31
rect 207 -37 265 -31
rect 325 -37 383 -31
rect 443 -37 501 -31
rect 561 -37 619 -31
rect 679 -37 737 -31
rect 797 -37 855 -31
rect -855 -71 -843 -37
rect -737 -71 -725 -37
rect -619 -71 -607 -37
rect -501 -71 -489 -37
rect -383 -71 -371 -37
rect -265 -71 -253 -37
rect -147 -71 -135 -37
rect -29 -71 -17 -37
rect 89 -71 101 -37
rect 207 -71 219 -37
rect 325 -71 337 -37
rect 443 -71 455 -37
rect 561 -71 573 -37
rect 679 -71 691 -37
rect 797 -71 809 -37
rect -855 -77 -797 -71
rect -737 -77 -679 -71
rect -619 -77 -561 -71
rect -501 -77 -443 -71
rect -383 -77 -325 -71
rect -265 -77 -207 -71
rect -147 -77 -89 -71
rect -29 -77 29 -71
rect 89 -77 147 -71
rect 207 -77 265 -71
rect 325 -77 383 -71
rect 443 -77 501 -71
rect 561 -77 619 -71
rect 679 -77 737 -71
rect 797 -77 855 -71
<< pwell >>
rect -1042 -909 1042 909
<< nmos >>
rect -856 109 -796 709
rect -738 109 -678 709
rect -620 109 -560 709
rect -502 109 -442 709
rect -384 109 -324 709
rect -266 109 -206 709
rect -148 109 -88 709
rect -30 109 30 709
rect 88 109 148 709
rect 206 109 266 709
rect 324 109 384 709
rect 442 109 502 709
rect 560 109 620 709
rect 678 109 738 709
rect 796 109 856 709
rect -856 -709 -796 -109
rect -738 -709 -678 -109
rect -620 -709 -560 -109
rect -502 -709 -442 -109
rect -384 -709 -324 -109
rect -266 -709 -206 -109
rect -148 -709 -88 -109
rect -30 -709 30 -109
rect 88 -709 148 -109
rect 206 -709 266 -109
rect 324 -709 384 -109
rect 442 -709 502 -109
rect 560 -709 620 -109
rect 678 -709 738 -109
rect 796 -709 856 -109
<< ndiff >>
rect -914 664 -856 709
rect -914 630 -902 664
rect -868 630 -856 664
rect -914 596 -856 630
rect -914 562 -902 596
rect -868 562 -856 596
rect -914 528 -856 562
rect -914 494 -902 528
rect -868 494 -856 528
rect -914 460 -856 494
rect -914 426 -902 460
rect -868 426 -856 460
rect -914 392 -856 426
rect -914 358 -902 392
rect -868 358 -856 392
rect -914 324 -856 358
rect -914 290 -902 324
rect -868 290 -856 324
rect -914 256 -856 290
rect -914 222 -902 256
rect -868 222 -856 256
rect -914 188 -856 222
rect -914 154 -902 188
rect -868 154 -856 188
rect -914 109 -856 154
rect -796 664 -738 709
rect -796 630 -784 664
rect -750 630 -738 664
rect -796 596 -738 630
rect -796 562 -784 596
rect -750 562 -738 596
rect -796 528 -738 562
rect -796 494 -784 528
rect -750 494 -738 528
rect -796 460 -738 494
rect -796 426 -784 460
rect -750 426 -738 460
rect -796 392 -738 426
rect -796 358 -784 392
rect -750 358 -738 392
rect -796 324 -738 358
rect -796 290 -784 324
rect -750 290 -738 324
rect -796 256 -738 290
rect -796 222 -784 256
rect -750 222 -738 256
rect -796 188 -738 222
rect -796 154 -784 188
rect -750 154 -738 188
rect -796 109 -738 154
rect -678 664 -620 709
rect -678 630 -666 664
rect -632 630 -620 664
rect -678 596 -620 630
rect -678 562 -666 596
rect -632 562 -620 596
rect -678 528 -620 562
rect -678 494 -666 528
rect -632 494 -620 528
rect -678 460 -620 494
rect -678 426 -666 460
rect -632 426 -620 460
rect -678 392 -620 426
rect -678 358 -666 392
rect -632 358 -620 392
rect -678 324 -620 358
rect -678 290 -666 324
rect -632 290 -620 324
rect -678 256 -620 290
rect -678 222 -666 256
rect -632 222 -620 256
rect -678 188 -620 222
rect -678 154 -666 188
rect -632 154 -620 188
rect -678 109 -620 154
rect -560 664 -502 709
rect -560 630 -548 664
rect -514 630 -502 664
rect -560 596 -502 630
rect -560 562 -548 596
rect -514 562 -502 596
rect -560 528 -502 562
rect -560 494 -548 528
rect -514 494 -502 528
rect -560 460 -502 494
rect -560 426 -548 460
rect -514 426 -502 460
rect -560 392 -502 426
rect -560 358 -548 392
rect -514 358 -502 392
rect -560 324 -502 358
rect -560 290 -548 324
rect -514 290 -502 324
rect -560 256 -502 290
rect -560 222 -548 256
rect -514 222 -502 256
rect -560 188 -502 222
rect -560 154 -548 188
rect -514 154 -502 188
rect -560 109 -502 154
rect -442 664 -384 709
rect -442 630 -430 664
rect -396 630 -384 664
rect -442 596 -384 630
rect -442 562 -430 596
rect -396 562 -384 596
rect -442 528 -384 562
rect -442 494 -430 528
rect -396 494 -384 528
rect -442 460 -384 494
rect -442 426 -430 460
rect -396 426 -384 460
rect -442 392 -384 426
rect -442 358 -430 392
rect -396 358 -384 392
rect -442 324 -384 358
rect -442 290 -430 324
rect -396 290 -384 324
rect -442 256 -384 290
rect -442 222 -430 256
rect -396 222 -384 256
rect -442 188 -384 222
rect -442 154 -430 188
rect -396 154 -384 188
rect -442 109 -384 154
rect -324 664 -266 709
rect -324 630 -312 664
rect -278 630 -266 664
rect -324 596 -266 630
rect -324 562 -312 596
rect -278 562 -266 596
rect -324 528 -266 562
rect -324 494 -312 528
rect -278 494 -266 528
rect -324 460 -266 494
rect -324 426 -312 460
rect -278 426 -266 460
rect -324 392 -266 426
rect -324 358 -312 392
rect -278 358 -266 392
rect -324 324 -266 358
rect -324 290 -312 324
rect -278 290 -266 324
rect -324 256 -266 290
rect -324 222 -312 256
rect -278 222 -266 256
rect -324 188 -266 222
rect -324 154 -312 188
rect -278 154 -266 188
rect -324 109 -266 154
rect -206 664 -148 709
rect -206 630 -194 664
rect -160 630 -148 664
rect -206 596 -148 630
rect -206 562 -194 596
rect -160 562 -148 596
rect -206 528 -148 562
rect -206 494 -194 528
rect -160 494 -148 528
rect -206 460 -148 494
rect -206 426 -194 460
rect -160 426 -148 460
rect -206 392 -148 426
rect -206 358 -194 392
rect -160 358 -148 392
rect -206 324 -148 358
rect -206 290 -194 324
rect -160 290 -148 324
rect -206 256 -148 290
rect -206 222 -194 256
rect -160 222 -148 256
rect -206 188 -148 222
rect -206 154 -194 188
rect -160 154 -148 188
rect -206 109 -148 154
rect -88 664 -30 709
rect -88 630 -76 664
rect -42 630 -30 664
rect -88 596 -30 630
rect -88 562 -76 596
rect -42 562 -30 596
rect -88 528 -30 562
rect -88 494 -76 528
rect -42 494 -30 528
rect -88 460 -30 494
rect -88 426 -76 460
rect -42 426 -30 460
rect -88 392 -30 426
rect -88 358 -76 392
rect -42 358 -30 392
rect -88 324 -30 358
rect -88 290 -76 324
rect -42 290 -30 324
rect -88 256 -30 290
rect -88 222 -76 256
rect -42 222 -30 256
rect -88 188 -30 222
rect -88 154 -76 188
rect -42 154 -30 188
rect -88 109 -30 154
rect 30 664 88 709
rect 30 630 42 664
rect 76 630 88 664
rect 30 596 88 630
rect 30 562 42 596
rect 76 562 88 596
rect 30 528 88 562
rect 30 494 42 528
rect 76 494 88 528
rect 30 460 88 494
rect 30 426 42 460
rect 76 426 88 460
rect 30 392 88 426
rect 30 358 42 392
rect 76 358 88 392
rect 30 324 88 358
rect 30 290 42 324
rect 76 290 88 324
rect 30 256 88 290
rect 30 222 42 256
rect 76 222 88 256
rect 30 188 88 222
rect 30 154 42 188
rect 76 154 88 188
rect 30 109 88 154
rect 148 664 206 709
rect 148 630 160 664
rect 194 630 206 664
rect 148 596 206 630
rect 148 562 160 596
rect 194 562 206 596
rect 148 528 206 562
rect 148 494 160 528
rect 194 494 206 528
rect 148 460 206 494
rect 148 426 160 460
rect 194 426 206 460
rect 148 392 206 426
rect 148 358 160 392
rect 194 358 206 392
rect 148 324 206 358
rect 148 290 160 324
rect 194 290 206 324
rect 148 256 206 290
rect 148 222 160 256
rect 194 222 206 256
rect 148 188 206 222
rect 148 154 160 188
rect 194 154 206 188
rect 148 109 206 154
rect 266 664 324 709
rect 266 630 278 664
rect 312 630 324 664
rect 266 596 324 630
rect 266 562 278 596
rect 312 562 324 596
rect 266 528 324 562
rect 266 494 278 528
rect 312 494 324 528
rect 266 460 324 494
rect 266 426 278 460
rect 312 426 324 460
rect 266 392 324 426
rect 266 358 278 392
rect 312 358 324 392
rect 266 324 324 358
rect 266 290 278 324
rect 312 290 324 324
rect 266 256 324 290
rect 266 222 278 256
rect 312 222 324 256
rect 266 188 324 222
rect 266 154 278 188
rect 312 154 324 188
rect 266 109 324 154
rect 384 664 442 709
rect 384 630 396 664
rect 430 630 442 664
rect 384 596 442 630
rect 384 562 396 596
rect 430 562 442 596
rect 384 528 442 562
rect 384 494 396 528
rect 430 494 442 528
rect 384 460 442 494
rect 384 426 396 460
rect 430 426 442 460
rect 384 392 442 426
rect 384 358 396 392
rect 430 358 442 392
rect 384 324 442 358
rect 384 290 396 324
rect 430 290 442 324
rect 384 256 442 290
rect 384 222 396 256
rect 430 222 442 256
rect 384 188 442 222
rect 384 154 396 188
rect 430 154 442 188
rect 384 109 442 154
rect 502 664 560 709
rect 502 630 514 664
rect 548 630 560 664
rect 502 596 560 630
rect 502 562 514 596
rect 548 562 560 596
rect 502 528 560 562
rect 502 494 514 528
rect 548 494 560 528
rect 502 460 560 494
rect 502 426 514 460
rect 548 426 560 460
rect 502 392 560 426
rect 502 358 514 392
rect 548 358 560 392
rect 502 324 560 358
rect 502 290 514 324
rect 548 290 560 324
rect 502 256 560 290
rect 502 222 514 256
rect 548 222 560 256
rect 502 188 560 222
rect 502 154 514 188
rect 548 154 560 188
rect 502 109 560 154
rect 620 664 678 709
rect 620 630 632 664
rect 666 630 678 664
rect 620 596 678 630
rect 620 562 632 596
rect 666 562 678 596
rect 620 528 678 562
rect 620 494 632 528
rect 666 494 678 528
rect 620 460 678 494
rect 620 426 632 460
rect 666 426 678 460
rect 620 392 678 426
rect 620 358 632 392
rect 666 358 678 392
rect 620 324 678 358
rect 620 290 632 324
rect 666 290 678 324
rect 620 256 678 290
rect 620 222 632 256
rect 666 222 678 256
rect 620 188 678 222
rect 620 154 632 188
rect 666 154 678 188
rect 620 109 678 154
rect 738 664 796 709
rect 738 630 750 664
rect 784 630 796 664
rect 738 596 796 630
rect 738 562 750 596
rect 784 562 796 596
rect 738 528 796 562
rect 738 494 750 528
rect 784 494 796 528
rect 738 460 796 494
rect 738 426 750 460
rect 784 426 796 460
rect 738 392 796 426
rect 738 358 750 392
rect 784 358 796 392
rect 738 324 796 358
rect 738 290 750 324
rect 784 290 796 324
rect 738 256 796 290
rect 738 222 750 256
rect 784 222 796 256
rect 738 188 796 222
rect 738 154 750 188
rect 784 154 796 188
rect 738 109 796 154
rect 856 664 914 709
rect 856 630 868 664
rect 902 630 914 664
rect 856 596 914 630
rect 856 562 868 596
rect 902 562 914 596
rect 856 528 914 562
rect 856 494 868 528
rect 902 494 914 528
rect 856 460 914 494
rect 856 426 868 460
rect 902 426 914 460
rect 856 392 914 426
rect 856 358 868 392
rect 902 358 914 392
rect 856 324 914 358
rect 856 290 868 324
rect 902 290 914 324
rect 856 256 914 290
rect 856 222 868 256
rect 902 222 914 256
rect 856 188 914 222
rect 856 154 868 188
rect 902 154 914 188
rect 856 109 914 154
rect -914 -154 -856 -109
rect -914 -188 -902 -154
rect -868 -188 -856 -154
rect -914 -222 -856 -188
rect -914 -256 -902 -222
rect -868 -256 -856 -222
rect -914 -290 -856 -256
rect -914 -324 -902 -290
rect -868 -324 -856 -290
rect -914 -358 -856 -324
rect -914 -392 -902 -358
rect -868 -392 -856 -358
rect -914 -426 -856 -392
rect -914 -460 -902 -426
rect -868 -460 -856 -426
rect -914 -494 -856 -460
rect -914 -528 -902 -494
rect -868 -528 -856 -494
rect -914 -562 -856 -528
rect -914 -596 -902 -562
rect -868 -596 -856 -562
rect -914 -630 -856 -596
rect -914 -664 -902 -630
rect -868 -664 -856 -630
rect -914 -709 -856 -664
rect -796 -154 -738 -109
rect -796 -188 -784 -154
rect -750 -188 -738 -154
rect -796 -222 -738 -188
rect -796 -256 -784 -222
rect -750 -256 -738 -222
rect -796 -290 -738 -256
rect -796 -324 -784 -290
rect -750 -324 -738 -290
rect -796 -358 -738 -324
rect -796 -392 -784 -358
rect -750 -392 -738 -358
rect -796 -426 -738 -392
rect -796 -460 -784 -426
rect -750 -460 -738 -426
rect -796 -494 -738 -460
rect -796 -528 -784 -494
rect -750 -528 -738 -494
rect -796 -562 -738 -528
rect -796 -596 -784 -562
rect -750 -596 -738 -562
rect -796 -630 -738 -596
rect -796 -664 -784 -630
rect -750 -664 -738 -630
rect -796 -709 -738 -664
rect -678 -154 -620 -109
rect -678 -188 -666 -154
rect -632 -188 -620 -154
rect -678 -222 -620 -188
rect -678 -256 -666 -222
rect -632 -256 -620 -222
rect -678 -290 -620 -256
rect -678 -324 -666 -290
rect -632 -324 -620 -290
rect -678 -358 -620 -324
rect -678 -392 -666 -358
rect -632 -392 -620 -358
rect -678 -426 -620 -392
rect -678 -460 -666 -426
rect -632 -460 -620 -426
rect -678 -494 -620 -460
rect -678 -528 -666 -494
rect -632 -528 -620 -494
rect -678 -562 -620 -528
rect -678 -596 -666 -562
rect -632 -596 -620 -562
rect -678 -630 -620 -596
rect -678 -664 -666 -630
rect -632 -664 -620 -630
rect -678 -709 -620 -664
rect -560 -154 -502 -109
rect -560 -188 -548 -154
rect -514 -188 -502 -154
rect -560 -222 -502 -188
rect -560 -256 -548 -222
rect -514 -256 -502 -222
rect -560 -290 -502 -256
rect -560 -324 -548 -290
rect -514 -324 -502 -290
rect -560 -358 -502 -324
rect -560 -392 -548 -358
rect -514 -392 -502 -358
rect -560 -426 -502 -392
rect -560 -460 -548 -426
rect -514 -460 -502 -426
rect -560 -494 -502 -460
rect -560 -528 -548 -494
rect -514 -528 -502 -494
rect -560 -562 -502 -528
rect -560 -596 -548 -562
rect -514 -596 -502 -562
rect -560 -630 -502 -596
rect -560 -664 -548 -630
rect -514 -664 -502 -630
rect -560 -709 -502 -664
rect -442 -154 -384 -109
rect -442 -188 -430 -154
rect -396 -188 -384 -154
rect -442 -222 -384 -188
rect -442 -256 -430 -222
rect -396 -256 -384 -222
rect -442 -290 -384 -256
rect -442 -324 -430 -290
rect -396 -324 -384 -290
rect -442 -358 -384 -324
rect -442 -392 -430 -358
rect -396 -392 -384 -358
rect -442 -426 -384 -392
rect -442 -460 -430 -426
rect -396 -460 -384 -426
rect -442 -494 -384 -460
rect -442 -528 -430 -494
rect -396 -528 -384 -494
rect -442 -562 -384 -528
rect -442 -596 -430 -562
rect -396 -596 -384 -562
rect -442 -630 -384 -596
rect -442 -664 -430 -630
rect -396 -664 -384 -630
rect -442 -709 -384 -664
rect -324 -154 -266 -109
rect -324 -188 -312 -154
rect -278 -188 -266 -154
rect -324 -222 -266 -188
rect -324 -256 -312 -222
rect -278 -256 -266 -222
rect -324 -290 -266 -256
rect -324 -324 -312 -290
rect -278 -324 -266 -290
rect -324 -358 -266 -324
rect -324 -392 -312 -358
rect -278 -392 -266 -358
rect -324 -426 -266 -392
rect -324 -460 -312 -426
rect -278 -460 -266 -426
rect -324 -494 -266 -460
rect -324 -528 -312 -494
rect -278 -528 -266 -494
rect -324 -562 -266 -528
rect -324 -596 -312 -562
rect -278 -596 -266 -562
rect -324 -630 -266 -596
rect -324 -664 -312 -630
rect -278 -664 -266 -630
rect -324 -709 -266 -664
rect -206 -154 -148 -109
rect -206 -188 -194 -154
rect -160 -188 -148 -154
rect -206 -222 -148 -188
rect -206 -256 -194 -222
rect -160 -256 -148 -222
rect -206 -290 -148 -256
rect -206 -324 -194 -290
rect -160 -324 -148 -290
rect -206 -358 -148 -324
rect -206 -392 -194 -358
rect -160 -392 -148 -358
rect -206 -426 -148 -392
rect -206 -460 -194 -426
rect -160 -460 -148 -426
rect -206 -494 -148 -460
rect -206 -528 -194 -494
rect -160 -528 -148 -494
rect -206 -562 -148 -528
rect -206 -596 -194 -562
rect -160 -596 -148 -562
rect -206 -630 -148 -596
rect -206 -664 -194 -630
rect -160 -664 -148 -630
rect -206 -709 -148 -664
rect -88 -154 -30 -109
rect -88 -188 -76 -154
rect -42 -188 -30 -154
rect -88 -222 -30 -188
rect -88 -256 -76 -222
rect -42 -256 -30 -222
rect -88 -290 -30 -256
rect -88 -324 -76 -290
rect -42 -324 -30 -290
rect -88 -358 -30 -324
rect -88 -392 -76 -358
rect -42 -392 -30 -358
rect -88 -426 -30 -392
rect -88 -460 -76 -426
rect -42 -460 -30 -426
rect -88 -494 -30 -460
rect -88 -528 -76 -494
rect -42 -528 -30 -494
rect -88 -562 -30 -528
rect -88 -596 -76 -562
rect -42 -596 -30 -562
rect -88 -630 -30 -596
rect -88 -664 -76 -630
rect -42 -664 -30 -630
rect -88 -709 -30 -664
rect 30 -154 88 -109
rect 30 -188 42 -154
rect 76 -188 88 -154
rect 30 -222 88 -188
rect 30 -256 42 -222
rect 76 -256 88 -222
rect 30 -290 88 -256
rect 30 -324 42 -290
rect 76 -324 88 -290
rect 30 -358 88 -324
rect 30 -392 42 -358
rect 76 -392 88 -358
rect 30 -426 88 -392
rect 30 -460 42 -426
rect 76 -460 88 -426
rect 30 -494 88 -460
rect 30 -528 42 -494
rect 76 -528 88 -494
rect 30 -562 88 -528
rect 30 -596 42 -562
rect 76 -596 88 -562
rect 30 -630 88 -596
rect 30 -664 42 -630
rect 76 -664 88 -630
rect 30 -709 88 -664
rect 148 -154 206 -109
rect 148 -188 160 -154
rect 194 -188 206 -154
rect 148 -222 206 -188
rect 148 -256 160 -222
rect 194 -256 206 -222
rect 148 -290 206 -256
rect 148 -324 160 -290
rect 194 -324 206 -290
rect 148 -358 206 -324
rect 148 -392 160 -358
rect 194 -392 206 -358
rect 148 -426 206 -392
rect 148 -460 160 -426
rect 194 -460 206 -426
rect 148 -494 206 -460
rect 148 -528 160 -494
rect 194 -528 206 -494
rect 148 -562 206 -528
rect 148 -596 160 -562
rect 194 -596 206 -562
rect 148 -630 206 -596
rect 148 -664 160 -630
rect 194 -664 206 -630
rect 148 -709 206 -664
rect 266 -154 324 -109
rect 266 -188 278 -154
rect 312 -188 324 -154
rect 266 -222 324 -188
rect 266 -256 278 -222
rect 312 -256 324 -222
rect 266 -290 324 -256
rect 266 -324 278 -290
rect 312 -324 324 -290
rect 266 -358 324 -324
rect 266 -392 278 -358
rect 312 -392 324 -358
rect 266 -426 324 -392
rect 266 -460 278 -426
rect 312 -460 324 -426
rect 266 -494 324 -460
rect 266 -528 278 -494
rect 312 -528 324 -494
rect 266 -562 324 -528
rect 266 -596 278 -562
rect 312 -596 324 -562
rect 266 -630 324 -596
rect 266 -664 278 -630
rect 312 -664 324 -630
rect 266 -709 324 -664
rect 384 -154 442 -109
rect 384 -188 396 -154
rect 430 -188 442 -154
rect 384 -222 442 -188
rect 384 -256 396 -222
rect 430 -256 442 -222
rect 384 -290 442 -256
rect 384 -324 396 -290
rect 430 -324 442 -290
rect 384 -358 442 -324
rect 384 -392 396 -358
rect 430 -392 442 -358
rect 384 -426 442 -392
rect 384 -460 396 -426
rect 430 -460 442 -426
rect 384 -494 442 -460
rect 384 -528 396 -494
rect 430 -528 442 -494
rect 384 -562 442 -528
rect 384 -596 396 -562
rect 430 -596 442 -562
rect 384 -630 442 -596
rect 384 -664 396 -630
rect 430 -664 442 -630
rect 384 -709 442 -664
rect 502 -154 560 -109
rect 502 -188 514 -154
rect 548 -188 560 -154
rect 502 -222 560 -188
rect 502 -256 514 -222
rect 548 -256 560 -222
rect 502 -290 560 -256
rect 502 -324 514 -290
rect 548 -324 560 -290
rect 502 -358 560 -324
rect 502 -392 514 -358
rect 548 -392 560 -358
rect 502 -426 560 -392
rect 502 -460 514 -426
rect 548 -460 560 -426
rect 502 -494 560 -460
rect 502 -528 514 -494
rect 548 -528 560 -494
rect 502 -562 560 -528
rect 502 -596 514 -562
rect 548 -596 560 -562
rect 502 -630 560 -596
rect 502 -664 514 -630
rect 548 -664 560 -630
rect 502 -709 560 -664
rect 620 -154 678 -109
rect 620 -188 632 -154
rect 666 -188 678 -154
rect 620 -222 678 -188
rect 620 -256 632 -222
rect 666 -256 678 -222
rect 620 -290 678 -256
rect 620 -324 632 -290
rect 666 -324 678 -290
rect 620 -358 678 -324
rect 620 -392 632 -358
rect 666 -392 678 -358
rect 620 -426 678 -392
rect 620 -460 632 -426
rect 666 -460 678 -426
rect 620 -494 678 -460
rect 620 -528 632 -494
rect 666 -528 678 -494
rect 620 -562 678 -528
rect 620 -596 632 -562
rect 666 -596 678 -562
rect 620 -630 678 -596
rect 620 -664 632 -630
rect 666 -664 678 -630
rect 620 -709 678 -664
rect 738 -154 796 -109
rect 738 -188 750 -154
rect 784 -188 796 -154
rect 738 -222 796 -188
rect 738 -256 750 -222
rect 784 -256 796 -222
rect 738 -290 796 -256
rect 738 -324 750 -290
rect 784 -324 796 -290
rect 738 -358 796 -324
rect 738 -392 750 -358
rect 784 -392 796 -358
rect 738 -426 796 -392
rect 738 -460 750 -426
rect 784 -460 796 -426
rect 738 -494 796 -460
rect 738 -528 750 -494
rect 784 -528 796 -494
rect 738 -562 796 -528
rect 738 -596 750 -562
rect 784 -596 796 -562
rect 738 -630 796 -596
rect 738 -664 750 -630
rect 784 -664 796 -630
rect 738 -709 796 -664
rect 856 -154 914 -109
rect 856 -188 868 -154
rect 902 -188 914 -154
rect 856 -222 914 -188
rect 856 -256 868 -222
rect 902 -256 914 -222
rect 856 -290 914 -256
rect 856 -324 868 -290
rect 902 -324 914 -290
rect 856 -358 914 -324
rect 856 -392 868 -358
rect 902 -392 914 -358
rect 856 -426 914 -392
rect 856 -460 868 -426
rect 902 -460 914 -426
rect 856 -494 914 -460
rect 856 -528 868 -494
rect 902 -528 914 -494
rect 856 -562 914 -528
rect 856 -596 868 -562
rect 902 -596 914 -562
rect 856 -630 914 -596
rect 856 -664 868 -630
rect 902 -664 914 -630
rect 856 -709 914 -664
<< ndiffc >>
rect -902 630 -868 664
rect -902 562 -868 596
rect -902 494 -868 528
rect -902 426 -868 460
rect -902 358 -868 392
rect -902 290 -868 324
rect -902 222 -868 256
rect -902 154 -868 188
rect -784 630 -750 664
rect -784 562 -750 596
rect -784 494 -750 528
rect -784 426 -750 460
rect -784 358 -750 392
rect -784 290 -750 324
rect -784 222 -750 256
rect -784 154 -750 188
rect -666 630 -632 664
rect -666 562 -632 596
rect -666 494 -632 528
rect -666 426 -632 460
rect -666 358 -632 392
rect -666 290 -632 324
rect -666 222 -632 256
rect -666 154 -632 188
rect -548 630 -514 664
rect -548 562 -514 596
rect -548 494 -514 528
rect -548 426 -514 460
rect -548 358 -514 392
rect -548 290 -514 324
rect -548 222 -514 256
rect -548 154 -514 188
rect -430 630 -396 664
rect -430 562 -396 596
rect -430 494 -396 528
rect -430 426 -396 460
rect -430 358 -396 392
rect -430 290 -396 324
rect -430 222 -396 256
rect -430 154 -396 188
rect -312 630 -278 664
rect -312 562 -278 596
rect -312 494 -278 528
rect -312 426 -278 460
rect -312 358 -278 392
rect -312 290 -278 324
rect -312 222 -278 256
rect -312 154 -278 188
rect -194 630 -160 664
rect -194 562 -160 596
rect -194 494 -160 528
rect -194 426 -160 460
rect -194 358 -160 392
rect -194 290 -160 324
rect -194 222 -160 256
rect -194 154 -160 188
rect -76 630 -42 664
rect -76 562 -42 596
rect -76 494 -42 528
rect -76 426 -42 460
rect -76 358 -42 392
rect -76 290 -42 324
rect -76 222 -42 256
rect -76 154 -42 188
rect 42 630 76 664
rect 42 562 76 596
rect 42 494 76 528
rect 42 426 76 460
rect 42 358 76 392
rect 42 290 76 324
rect 42 222 76 256
rect 42 154 76 188
rect 160 630 194 664
rect 160 562 194 596
rect 160 494 194 528
rect 160 426 194 460
rect 160 358 194 392
rect 160 290 194 324
rect 160 222 194 256
rect 160 154 194 188
rect 278 630 312 664
rect 278 562 312 596
rect 278 494 312 528
rect 278 426 312 460
rect 278 358 312 392
rect 278 290 312 324
rect 278 222 312 256
rect 278 154 312 188
rect 396 630 430 664
rect 396 562 430 596
rect 396 494 430 528
rect 396 426 430 460
rect 396 358 430 392
rect 396 290 430 324
rect 396 222 430 256
rect 396 154 430 188
rect 514 630 548 664
rect 514 562 548 596
rect 514 494 548 528
rect 514 426 548 460
rect 514 358 548 392
rect 514 290 548 324
rect 514 222 548 256
rect 514 154 548 188
rect 632 630 666 664
rect 632 562 666 596
rect 632 494 666 528
rect 632 426 666 460
rect 632 358 666 392
rect 632 290 666 324
rect 632 222 666 256
rect 632 154 666 188
rect 750 630 784 664
rect 750 562 784 596
rect 750 494 784 528
rect 750 426 784 460
rect 750 358 784 392
rect 750 290 784 324
rect 750 222 784 256
rect 750 154 784 188
rect 868 630 902 664
rect 868 562 902 596
rect 868 494 902 528
rect 868 426 902 460
rect 868 358 902 392
rect 868 290 902 324
rect 868 222 902 256
rect 868 154 902 188
rect -902 -188 -868 -154
rect -902 -256 -868 -222
rect -902 -324 -868 -290
rect -902 -392 -868 -358
rect -902 -460 -868 -426
rect -902 -528 -868 -494
rect -902 -596 -868 -562
rect -902 -664 -868 -630
rect -784 -188 -750 -154
rect -784 -256 -750 -222
rect -784 -324 -750 -290
rect -784 -392 -750 -358
rect -784 -460 -750 -426
rect -784 -528 -750 -494
rect -784 -596 -750 -562
rect -784 -664 -750 -630
rect -666 -188 -632 -154
rect -666 -256 -632 -222
rect -666 -324 -632 -290
rect -666 -392 -632 -358
rect -666 -460 -632 -426
rect -666 -528 -632 -494
rect -666 -596 -632 -562
rect -666 -664 -632 -630
rect -548 -188 -514 -154
rect -548 -256 -514 -222
rect -548 -324 -514 -290
rect -548 -392 -514 -358
rect -548 -460 -514 -426
rect -548 -528 -514 -494
rect -548 -596 -514 -562
rect -548 -664 -514 -630
rect -430 -188 -396 -154
rect -430 -256 -396 -222
rect -430 -324 -396 -290
rect -430 -392 -396 -358
rect -430 -460 -396 -426
rect -430 -528 -396 -494
rect -430 -596 -396 -562
rect -430 -664 -396 -630
rect -312 -188 -278 -154
rect -312 -256 -278 -222
rect -312 -324 -278 -290
rect -312 -392 -278 -358
rect -312 -460 -278 -426
rect -312 -528 -278 -494
rect -312 -596 -278 -562
rect -312 -664 -278 -630
rect -194 -188 -160 -154
rect -194 -256 -160 -222
rect -194 -324 -160 -290
rect -194 -392 -160 -358
rect -194 -460 -160 -426
rect -194 -528 -160 -494
rect -194 -596 -160 -562
rect -194 -664 -160 -630
rect -76 -188 -42 -154
rect -76 -256 -42 -222
rect -76 -324 -42 -290
rect -76 -392 -42 -358
rect -76 -460 -42 -426
rect -76 -528 -42 -494
rect -76 -596 -42 -562
rect -76 -664 -42 -630
rect 42 -188 76 -154
rect 42 -256 76 -222
rect 42 -324 76 -290
rect 42 -392 76 -358
rect 42 -460 76 -426
rect 42 -528 76 -494
rect 42 -596 76 -562
rect 42 -664 76 -630
rect 160 -188 194 -154
rect 160 -256 194 -222
rect 160 -324 194 -290
rect 160 -392 194 -358
rect 160 -460 194 -426
rect 160 -528 194 -494
rect 160 -596 194 -562
rect 160 -664 194 -630
rect 278 -188 312 -154
rect 278 -256 312 -222
rect 278 -324 312 -290
rect 278 -392 312 -358
rect 278 -460 312 -426
rect 278 -528 312 -494
rect 278 -596 312 -562
rect 278 -664 312 -630
rect 396 -188 430 -154
rect 396 -256 430 -222
rect 396 -324 430 -290
rect 396 -392 430 -358
rect 396 -460 430 -426
rect 396 -528 430 -494
rect 396 -596 430 -562
rect 396 -664 430 -630
rect 514 -188 548 -154
rect 514 -256 548 -222
rect 514 -324 548 -290
rect 514 -392 548 -358
rect 514 -460 548 -426
rect 514 -528 548 -494
rect 514 -596 548 -562
rect 514 -664 548 -630
rect 632 -188 666 -154
rect 632 -256 666 -222
rect 632 -324 666 -290
rect 632 -392 666 -358
rect 632 -460 666 -426
rect 632 -528 666 -494
rect 632 -596 666 -562
rect 632 -664 666 -630
rect 750 -188 784 -154
rect 750 -256 784 -222
rect 750 -324 784 -290
rect 750 -392 784 -358
rect 750 -460 784 -426
rect 750 -528 784 -494
rect 750 -596 784 -562
rect 750 -664 784 -630
rect 868 -188 902 -154
rect 868 -256 902 -222
rect 868 -324 902 -290
rect 868 -392 902 -358
rect 868 -460 902 -426
rect 868 -528 902 -494
rect 868 -596 902 -562
rect 868 -664 902 -630
<< psubdiff >>
rect -1016 849 -901 883
rect -867 849 -833 883
rect -799 849 -765 883
rect -731 849 -697 883
rect -663 849 -629 883
rect -595 849 -561 883
rect -527 849 -493 883
rect -459 849 -425 883
rect -391 849 -357 883
rect -323 849 -289 883
rect -255 849 -221 883
rect -187 849 -153 883
rect -119 849 -85 883
rect -51 849 -17 883
rect 17 849 51 883
rect 85 849 119 883
rect 153 849 187 883
rect 221 849 255 883
rect 289 849 323 883
rect 357 849 391 883
rect 425 849 459 883
rect 493 849 527 883
rect 561 849 595 883
rect 629 849 663 883
rect 697 849 731 883
rect 765 849 799 883
rect 833 849 867 883
rect 901 849 1016 883
rect -1016 765 -982 849
rect 982 765 1016 849
rect -1016 697 -982 731
rect -1016 629 -982 663
rect -1016 561 -982 595
rect -1016 493 -982 527
rect -1016 425 -982 459
rect -1016 357 -982 391
rect -1016 289 -982 323
rect -1016 221 -982 255
rect -1016 153 -982 187
rect -1016 85 -982 119
rect 982 697 1016 731
rect 982 629 1016 663
rect 982 561 1016 595
rect 982 493 1016 527
rect 982 425 1016 459
rect 982 357 1016 391
rect 982 289 1016 323
rect 982 221 1016 255
rect 982 153 1016 187
rect -1016 17 -982 51
rect 982 85 1016 119
rect -1016 -51 -982 -17
rect 982 17 1016 51
rect -1016 -119 -982 -85
rect 982 -51 1016 -17
rect -1016 -187 -982 -153
rect -1016 -255 -982 -221
rect -1016 -323 -982 -289
rect -1016 -391 -982 -357
rect -1016 -459 -982 -425
rect -1016 -527 -982 -493
rect -1016 -595 -982 -561
rect -1016 -663 -982 -629
rect -1016 -731 -982 -697
rect 982 -119 1016 -85
rect 982 -187 1016 -153
rect 982 -255 1016 -221
rect 982 -323 1016 -289
rect 982 -391 1016 -357
rect 982 -459 1016 -425
rect 982 -527 1016 -493
rect 982 -595 1016 -561
rect 982 -663 1016 -629
rect 982 -731 1016 -697
rect -1016 -849 -982 -765
rect 982 -849 1016 -765
rect -1016 -883 -901 -849
rect -867 -883 -833 -849
rect -799 -883 -765 -849
rect -731 -883 -697 -849
rect -663 -883 -629 -849
rect -595 -883 -561 -849
rect -527 -883 -493 -849
rect -459 -883 -425 -849
rect -391 -883 -357 -849
rect -323 -883 -289 -849
rect -255 -883 -221 -849
rect -187 -883 -153 -849
rect -119 -883 -85 -849
rect -51 -883 -17 -849
rect 17 -883 51 -849
rect 85 -883 119 -849
rect 153 -883 187 -849
rect 221 -883 255 -849
rect 289 -883 323 -849
rect 357 -883 391 -849
rect 425 -883 459 -849
rect 493 -883 527 -849
rect 561 -883 595 -849
rect 629 -883 663 -849
rect 697 -883 731 -849
rect 765 -883 799 -849
rect 833 -883 867 -849
rect 901 -883 1016 -849
<< psubdiffcont >>
rect -901 849 -867 883
rect -833 849 -799 883
rect -765 849 -731 883
rect -697 849 -663 883
rect -629 849 -595 883
rect -561 849 -527 883
rect -493 849 -459 883
rect -425 849 -391 883
rect -357 849 -323 883
rect -289 849 -255 883
rect -221 849 -187 883
rect -153 849 -119 883
rect -85 849 -51 883
rect -17 849 17 883
rect 51 849 85 883
rect 119 849 153 883
rect 187 849 221 883
rect 255 849 289 883
rect 323 849 357 883
rect 391 849 425 883
rect 459 849 493 883
rect 527 849 561 883
rect 595 849 629 883
rect 663 849 697 883
rect 731 849 765 883
rect 799 849 833 883
rect 867 849 901 883
rect -1016 731 -982 765
rect 982 731 1016 765
rect -1016 663 -982 697
rect -1016 595 -982 629
rect -1016 527 -982 561
rect -1016 459 -982 493
rect -1016 391 -982 425
rect -1016 323 -982 357
rect -1016 255 -982 289
rect -1016 187 -982 221
rect -1016 119 -982 153
rect 982 663 1016 697
rect 982 595 1016 629
rect 982 527 1016 561
rect 982 459 1016 493
rect 982 391 1016 425
rect 982 323 1016 357
rect 982 255 1016 289
rect 982 187 1016 221
rect 982 119 1016 153
rect -1016 51 -982 85
rect 982 51 1016 85
rect -1016 -17 -982 17
rect 982 -17 1016 17
rect -1016 -85 -982 -51
rect 982 -85 1016 -51
rect -1016 -153 -982 -119
rect -1016 -221 -982 -187
rect -1016 -289 -982 -255
rect -1016 -357 -982 -323
rect -1016 -425 -982 -391
rect -1016 -493 -982 -459
rect -1016 -561 -982 -527
rect -1016 -629 -982 -595
rect -1016 -697 -982 -663
rect 982 -153 1016 -119
rect 982 -221 1016 -187
rect 982 -289 1016 -255
rect 982 -357 1016 -323
rect 982 -425 1016 -391
rect 982 -493 1016 -459
rect 982 -561 1016 -527
rect 982 -629 1016 -595
rect 982 -697 1016 -663
rect -1016 -765 -982 -731
rect 982 -765 1016 -731
rect -901 -883 -867 -849
rect -833 -883 -799 -849
rect -765 -883 -731 -849
rect -697 -883 -663 -849
rect -629 -883 -595 -849
rect -561 -883 -527 -849
rect -493 -883 -459 -849
rect -425 -883 -391 -849
rect -357 -883 -323 -849
rect -289 -883 -255 -849
rect -221 -883 -187 -849
rect -153 -883 -119 -849
rect -85 -883 -51 -849
rect -17 -883 17 -849
rect 51 -883 85 -849
rect 119 -883 153 -849
rect 187 -883 221 -849
rect 255 -883 289 -849
rect 323 -883 357 -849
rect 391 -883 425 -849
rect 459 -883 493 -849
rect 527 -883 561 -849
rect 595 -883 629 -849
rect 663 -883 697 -849
rect 731 -883 765 -849
rect 799 -883 833 -849
rect 867 -883 901 -849
<< poly >>
rect -859 731 -793 797
rect -741 731 -675 797
rect -623 731 -557 797
rect -505 731 -439 797
rect -387 731 -321 797
rect -269 731 -203 797
rect -151 731 -85 797
rect -33 731 33 797
rect 85 731 151 797
rect 203 731 269 797
rect 321 731 387 797
rect 439 731 505 797
rect 557 731 623 797
rect 675 731 741 797
rect 793 731 859 797
rect -856 709 -796 731
rect -738 709 -678 731
rect -620 709 -560 731
rect -502 709 -442 731
rect -384 709 -324 731
rect -266 709 -206 731
rect -148 709 -88 731
rect -30 709 30 731
rect 88 709 148 731
rect 206 709 266 731
rect 324 709 384 731
rect 442 709 502 731
rect 560 709 620 731
rect 678 709 738 731
rect 796 709 856 731
rect -856 87 -796 109
rect -738 87 -678 109
rect -620 87 -560 109
rect -502 87 -442 109
rect -384 87 -324 109
rect -266 87 -206 109
rect -148 87 -88 109
rect -30 87 30 109
rect 88 87 148 109
rect 206 87 266 109
rect 324 87 384 109
rect 442 87 502 109
rect 560 87 620 109
rect 678 87 738 109
rect 796 87 856 109
rect -859 71 -793 87
rect -859 37 -843 71
rect -809 37 -793 71
rect -859 21 -793 37
rect -741 71 -675 87
rect -741 37 -725 71
rect -691 37 -675 71
rect -741 21 -675 37
rect -623 71 -557 87
rect -623 37 -607 71
rect -573 37 -557 71
rect -623 21 -557 37
rect -505 71 -439 87
rect -505 37 -489 71
rect -455 37 -439 71
rect -505 21 -439 37
rect -387 71 -321 87
rect -387 37 -371 71
rect -337 37 -321 71
rect -387 21 -321 37
rect -269 71 -203 87
rect -269 37 -253 71
rect -219 37 -203 71
rect -269 21 -203 37
rect -151 71 -85 87
rect -151 37 -135 71
rect -101 37 -85 71
rect -151 21 -85 37
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect 85 71 151 87
rect 85 37 101 71
rect 135 37 151 71
rect 85 21 151 37
rect 203 71 269 87
rect 203 37 219 71
rect 253 37 269 71
rect 203 21 269 37
rect 321 71 387 87
rect 321 37 337 71
rect 371 37 387 71
rect 321 21 387 37
rect 439 71 505 87
rect 439 37 455 71
rect 489 37 505 71
rect 439 21 505 37
rect 557 71 623 87
rect 557 37 573 71
rect 607 37 623 71
rect 557 21 623 37
rect 675 71 741 87
rect 675 37 691 71
rect 725 37 741 71
rect 675 21 741 37
rect 793 71 859 87
rect 793 37 809 71
rect 843 37 859 71
rect 793 21 859 37
rect -859 -37 -793 -21
rect -859 -71 -843 -37
rect -809 -71 -793 -37
rect -859 -87 -793 -71
rect -741 -37 -675 -21
rect -741 -71 -725 -37
rect -691 -71 -675 -37
rect -741 -87 -675 -71
rect -623 -37 -557 -21
rect -623 -71 -607 -37
rect -573 -71 -557 -37
rect -623 -87 -557 -71
rect -505 -37 -439 -21
rect -505 -71 -489 -37
rect -455 -71 -439 -37
rect -505 -87 -439 -71
rect -387 -37 -321 -21
rect -387 -71 -371 -37
rect -337 -71 -321 -37
rect -387 -87 -321 -71
rect -269 -37 -203 -21
rect -269 -71 -253 -37
rect -219 -71 -203 -37
rect -269 -87 -203 -71
rect -151 -37 -85 -21
rect -151 -71 -135 -37
rect -101 -71 -85 -37
rect -151 -87 -85 -71
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect 85 -37 151 -21
rect 85 -71 101 -37
rect 135 -71 151 -37
rect 85 -87 151 -71
rect 203 -37 269 -21
rect 203 -71 219 -37
rect 253 -71 269 -37
rect 203 -87 269 -71
rect 321 -37 387 -21
rect 321 -71 337 -37
rect 371 -71 387 -37
rect 321 -87 387 -71
rect 439 -37 505 -21
rect 439 -71 455 -37
rect 489 -71 505 -37
rect 439 -87 505 -71
rect 557 -37 623 -21
rect 557 -71 573 -37
rect 607 -71 623 -37
rect 557 -87 623 -71
rect 675 -37 741 -21
rect 675 -71 691 -37
rect 725 -71 741 -37
rect 675 -87 741 -71
rect 793 -37 859 -21
rect 793 -71 809 -37
rect 843 -71 859 -37
rect 793 -87 859 -71
rect -856 -109 -796 -87
rect -738 -109 -678 -87
rect -620 -109 -560 -87
rect -502 -109 -442 -87
rect -384 -109 -324 -87
rect -266 -109 -206 -87
rect -148 -109 -88 -87
rect -30 -109 30 -87
rect 88 -109 148 -87
rect 206 -109 266 -87
rect 324 -109 384 -87
rect 442 -109 502 -87
rect 560 -109 620 -87
rect 678 -109 738 -87
rect 796 -109 856 -87
rect -856 -731 -796 -709
rect -738 -731 -678 -709
rect -620 -731 -560 -709
rect -502 -731 -442 -709
rect -384 -731 -324 -709
rect -266 -731 -206 -709
rect -148 -731 -88 -709
rect -30 -731 30 -709
rect 88 -731 148 -709
rect 206 -731 266 -709
rect 324 -731 384 -709
rect 442 -731 502 -709
rect 560 -731 620 -709
rect 678 -731 738 -709
rect 796 -731 856 -709
rect -859 -797 -793 -731
rect -741 -797 -675 -731
rect -623 -797 -557 -731
rect -505 -797 -439 -731
rect -387 -797 -321 -731
rect -269 -797 -203 -731
rect -151 -797 -85 -731
rect -33 -797 33 -731
rect 85 -797 151 -731
rect 203 -797 269 -731
rect 321 -797 387 -731
rect 439 -797 505 -731
rect 557 -797 623 -731
rect 675 -797 741 -731
rect 793 -797 859 -731
<< polycont >>
rect -843 37 -809 71
rect -725 37 -691 71
rect -607 37 -573 71
rect -489 37 -455 71
rect -371 37 -337 71
rect -253 37 -219 71
rect -135 37 -101 71
rect -17 37 17 71
rect 101 37 135 71
rect 219 37 253 71
rect 337 37 371 71
rect 455 37 489 71
rect 573 37 607 71
rect 691 37 725 71
rect 809 37 843 71
rect -843 -71 -809 -37
rect -725 -71 -691 -37
rect -607 -71 -573 -37
rect -489 -71 -455 -37
rect -371 -71 -337 -37
rect -253 -71 -219 -37
rect -135 -71 -101 -37
rect -17 -71 17 -37
rect 101 -71 135 -37
rect 219 -71 253 -37
rect 337 -71 371 -37
rect 455 -71 489 -37
rect 573 -71 607 -37
rect 691 -71 725 -37
rect 809 -71 843 -37
<< locali >>
rect -1016 849 -901 883
rect -867 849 -833 883
rect -799 849 -765 883
rect -731 849 -697 883
rect -663 849 -629 883
rect -595 849 -561 883
rect -527 849 -493 883
rect -459 849 -425 883
rect -391 849 -357 883
rect -323 849 -289 883
rect -255 849 -221 883
rect -187 849 -153 883
rect -119 849 -85 883
rect -51 849 -17 883
rect 17 849 51 883
rect 85 849 119 883
rect 153 849 187 883
rect 221 849 255 883
rect 289 849 323 883
rect 357 849 391 883
rect 425 849 459 883
rect 493 849 527 883
rect 561 849 595 883
rect 629 849 663 883
rect 697 849 731 883
rect 765 849 799 883
rect 833 849 867 883
rect 901 849 1016 883
rect -1016 765 -982 849
rect -1016 697 -982 731
rect 982 765 1016 849
rect -1016 629 -982 663
rect -1016 561 -982 595
rect -1016 493 -982 527
rect -1016 425 -982 459
rect -1016 357 -982 391
rect -1016 289 -982 323
rect -1016 221 -982 255
rect -1016 153 -982 187
rect -1016 85 -982 119
rect -902 678 -868 713
rect -902 606 -868 630
rect -902 534 -868 562
rect -902 462 -868 494
rect -902 392 -868 426
rect -902 324 -868 356
rect -902 256 -868 284
rect -902 188 -868 212
rect -902 105 -868 140
rect -784 678 -750 713
rect -784 606 -750 630
rect -784 534 -750 562
rect -784 462 -750 494
rect -784 392 -750 426
rect -784 324 -750 356
rect -784 256 -750 284
rect -784 188 -750 212
rect -784 105 -750 140
rect -666 678 -632 713
rect -666 606 -632 630
rect -666 534 -632 562
rect -666 462 -632 494
rect -666 392 -632 426
rect -666 324 -632 356
rect -666 256 -632 284
rect -666 188 -632 212
rect -666 105 -632 140
rect -548 678 -514 713
rect -548 606 -514 630
rect -548 534 -514 562
rect -548 462 -514 494
rect -548 392 -514 426
rect -548 324 -514 356
rect -548 256 -514 284
rect -548 188 -514 212
rect -548 105 -514 140
rect -430 678 -396 713
rect -430 606 -396 630
rect -430 534 -396 562
rect -430 462 -396 494
rect -430 392 -396 426
rect -430 324 -396 356
rect -430 256 -396 284
rect -430 188 -396 212
rect -430 105 -396 140
rect -312 678 -278 713
rect -312 606 -278 630
rect -312 534 -278 562
rect -312 462 -278 494
rect -312 392 -278 426
rect -312 324 -278 356
rect -312 256 -278 284
rect -312 188 -278 212
rect -312 105 -278 140
rect -194 678 -160 713
rect -194 606 -160 630
rect -194 534 -160 562
rect -194 462 -160 494
rect -194 392 -160 426
rect -194 324 -160 356
rect -194 256 -160 284
rect -194 188 -160 212
rect -194 105 -160 140
rect -76 678 -42 713
rect -76 606 -42 630
rect -76 534 -42 562
rect -76 462 -42 494
rect -76 392 -42 426
rect -76 324 -42 356
rect -76 256 -42 284
rect -76 188 -42 212
rect -76 105 -42 140
rect 42 678 76 713
rect 42 606 76 630
rect 42 534 76 562
rect 42 462 76 494
rect 42 392 76 426
rect 42 324 76 356
rect 42 256 76 284
rect 42 188 76 212
rect 42 105 76 140
rect 160 678 194 713
rect 160 606 194 630
rect 160 534 194 562
rect 160 462 194 494
rect 160 392 194 426
rect 160 324 194 356
rect 160 256 194 284
rect 160 188 194 212
rect 160 105 194 140
rect 278 678 312 713
rect 278 606 312 630
rect 278 534 312 562
rect 278 462 312 494
rect 278 392 312 426
rect 278 324 312 356
rect 278 256 312 284
rect 278 188 312 212
rect 278 105 312 140
rect 396 678 430 713
rect 396 606 430 630
rect 396 534 430 562
rect 396 462 430 494
rect 396 392 430 426
rect 396 324 430 356
rect 396 256 430 284
rect 396 188 430 212
rect 396 105 430 140
rect 514 678 548 713
rect 514 606 548 630
rect 514 534 548 562
rect 514 462 548 494
rect 514 392 548 426
rect 514 324 548 356
rect 514 256 548 284
rect 514 188 548 212
rect 514 105 548 140
rect 632 678 666 713
rect 632 606 666 630
rect 632 534 666 562
rect 632 462 666 494
rect 632 392 666 426
rect 632 324 666 356
rect 632 256 666 284
rect 632 188 666 212
rect 632 105 666 140
rect 750 678 784 713
rect 750 606 784 630
rect 750 534 784 562
rect 750 462 784 494
rect 750 392 784 426
rect 750 324 784 356
rect 750 256 784 284
rect 750 188 784 212
rect 750 105 784 140
rect 868 678 902 713
rect 868 606 902 630
rect 868 534 902 562
rect 868 462 902 494
rect 868 392 902 426
rect 868 324 902 356
rect 868 256 902 284
rect 868 188 902 212
rect 868 105 902 140
rect 982 697 1016 731
rect 982 629 1016 663
rect 982 561 1016 595
rect 982 493 1016 527
rect 982 425 1016 459
rect 982 357 1016 391
rect 982 289 1016 323
rect 982 221 1016 255
rect 982 153 1016 187
rect 982 85 1016 119
rect -1016 17 -982 51
rect -859 37 -843 71
rect -809 37 -793 71
rect -741 37 -725 71
rect -691 37 -675 71
rect -623 37 -607 71
rect -573 37 -557 71
rect -505 37 -489 71
rect -455 37 -439 71
rect -387 37 -371 71
rect -337 37 -321 71
rect -269 37 -253 71
rect -219 37 -203 71
rect -151 37 -135 71
rect -101 37 -85 71
rect -33 37 -17 71
rect 17 37 33 71
rect 85 37 101 71
rect 135 37 151 71
rect 203 37 219 71
rect 253 37 269 71
rect 321 37 337 71
rect 371 37 387 71
rect 439 37 455 71
rect 489 37 505 71
rect 557 37 573 71
rect 607 37 623 71
rect 675 37 691 71
rect 725 37 741 71
rect 793 37 809 71
rect 843 37 859 71
rect -1016 -51 -982 -17
rect 982 17 1016 51
rect -859 -71 -843 -37
rect -809 -71 -793 -37
rect -741 -71 -725 -37
rect -691 -71 -675 -37
rect -623 -71 -607 -37
rect -573 -71 -557 -37
rect -505 -71 -489 -37
rect -455 -71 -439 -37
rect -387 -71 -371 -37
rect -337 -71 -321 -37
rect -269 -71 -253 -37
rect -219 -71 -203 -37
rect -151 -71 -135 -37
rect -101 -71 -85 -37
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect 85 -71 101 -37
rect 135 -71 151 -37
rect 203 -71 219 -37
rect 253 -71 269 -37
rect 321 -71 337 -37
rect 371 -71 387 -37
rect 439 -71 455 -37
rect 489 -71 505 -37
rect 557 -71 573 -37
rect 607 -71 623 -37
rect 675 -71 691 -37
rect 725 -71 741 -37
rect 793 -71 809 -37
rect 843 -71 859 -37
rect 982 -51 1016 -17
rect -1016 -119 -982 -85
rect -1016 -187 -982 -153
rect -1016 -255 -982 -221
rect -1016 -323 -982 -289
rect -1016 -391 -982 -357
rect -1016 -459 -982 -425
rect -1016 -527 -982 -493
rect -1016 -595 -982 -561
rect -1016 -663 -982 -629
rect -1016 -731 -982 -697
rect -902 -140 -868 -105
rect -902 -212 -868 -188
rect -902 -284 -868 -256
rect -902 -356 -868 -324
rect -902 -426 -868 -392
rect -902 -494 -868 -462
rect -902 -562 -868 -534
rect -902 -630 -868 -606
rect -902 -713 -868 -678
rect -784 -140 -750 -105
rect -784 -212 -750 -188
rect -784 -284 -750 -256
rect -784 -356 -750 -324
rect -784 -426 -750 -392
rect -784 -494 -750 -462
rect -784 -562 -750 -534
rect -784 -630 -750 -606
rect -784 -713 -750 -678
rect -666 -140 -632 -105
rect -666 -212 -632 -188
rect -666 -284 -632 -256
rect -666 -356 -632 -324
rect -666 -426 -632 -392
rect -666 -494 -632 -462
rect -666 -562 -632 -534
rect -666 -630 -632 -606
rect -666 -713 -632 -678
rect -548 -140 -514 -105
rect -548 -212 -514 -188
rect -548 -284 -514 -256
rect -548 -356 -514 -324
rect -548 -426 -514 -392
rect -548 -494 -514 -462
rect -548 -562 -514 -534
rect -548 -630 -514 -606
rect -548 -713 -514 -678
rect -430 -140 -396 -105
rect -430 -212 -396 -188
rect -430 -284 -396 -256
rect -430 -356 -396 -324
rect -430 -426 -396 -392
rect -430 -494 -396 -462
rect -430 -562 -396 -534
rect -430 -630 -396 -606
rect -430 -713 -396 -678
rect -312 -140 -278 -105
rect -312 -212 -278 -188
rect -312 -284 -278 -256
rect -312 -356 -278 -324
rect -312 -426 -278 -392
rect -312 -494 -278 -462
rect -312 -562 -278 -534
rect -312 -630 -278 -606
rect -312 -713 -278 -678
rect -194 -140 -160 -105
rect -194 -212 -160 -188
rect -194 -284 -160 -256
rect -194 -356 -160 -324
rect -194 -426 -160 -392
rect -194 -494 -160 -462
rect -194 -562 -160 -534
rect -194 -630 -160 -606
rect -194 -713 -160 -678
rect -76 -140 -42 -105
rect -76 -212 -42 -188
rect -76 -284 -42 -256
rect -76 -356 -42 -324
rect -76 -426 -42 -392
rect -76 -494 -42 -462
rect -76 -562 -42 -534
rect -76 -630 -42 -606
rect -76 -713 -42 -678
rect 42 -140 76 -105
rect 42 -212 76 -188
rect 42 -284 76 -256
rect 42 -356 76 -324
rect 42 -426 76 -392
rect 42 -494 76 -462
rect 42 -562 76 -534
rect 42 -630 76 -606
rect 42 -713 76 -678
rect 160 -140 194 -105
rect 160 -212 194 -188
rect 160 -284 194 -256
rect 160 -356 194 -324
rect 160 -426 194 -392
rect 160 -494 194 -462
rect 160 -562 194 -534
rect 160 -630 194 -606
rect 160 -713 194 -678
rect 278 -140 312 -105
rect 278 -212 312 -188
rect 278 -284 312 -256
rect 278 -356 312 -324
rect 278 -426 312 -392
rect 278 -494 312 -462
rect 278 -562 312 -534
rect 278 -630 312 -606
rect 278 -713 312 -678
rect 396 -140 430 -105
rect 396 -212 430 -188
rect 396 -284 430 -256
rect 396 -356 430 -324
rect 396 -426 430 -392
rect 396 -494 430 -462
rect 396 -562 430 -534
rect 396 -630 430 -606
rect 396 -713 430 -678
rect 514 -140 548 -105
rect 514 -212 548 -188
rect 514 -284 548 -256
rect 514 -356 548 -324
rect 514 -426 548 -392
rect 514 -494 548 -462
rect 514 -562 548 -534
rect 514 -630 548 -606
rect 514 -713 548 -678
rect 632 -140 666 -105
rect 632 -212 666 -188
rect 632 -284 666 -256
rect 632 -356 666 -324
rect 632 -426 666 -392
rect 632 -494 666 -462
rect 632 -562 666 -534
rect 632 -630 666 -606
rect 632 -713 666 -678
rect 750 -140 784 -105
rect 750 -212 784 -188
rect 750 -284 784 -256
rect 750 -356 784 -324
rect 750 -426 784 -392
rect 750 -494 784 -462
rect 750 -562 784 -534
rect 750 -630 784 -606
rect 750 -713 784 -678
rect 868 -140 902 -105
rect 868 -212 902 -188
rect 868 -284 902 -256
rect 868 -356 902 -324
rect 868 -426 902 -392
rect 868 -494 902 -462
rect 868 -562 902 -534
rect 868 -630 902 -606
rect 868 -713 902 -678
rect 982 -119 1016 -85
rect 982 -187 1016 -153
rect 982 -255 1016 -221
rect 982 -323 1016 -289
rect 982 -391 1016 -357
rect 982 -459 1016 -425
rect 982 -527 1016 -493
rect 982 -595 1016 -561
rect 982 -663 1016 -629
rect -1016 -849 -982 -765
rect 982 -731 1016 -697
rect 982 -849 1016 -765
rect -1016 -883 -901 -849
rect -867 -883 -833 -849
rect -799 -883 -765 -849
rect -731 -883 -697 -849
rect -663 -883 -629 -849
rect -595 -883 -561 -849
rect -527 -883 -493 -849
rect -459 -883 -425 -849
rect -391 -883 -357 -849
rect -323 -883 -289 -849
rect -255 -883 -221 -849
rect -187 -883 -153 -849
rect -119 -883 -85 -849
rect -51 -883 -17 -849
rect 17 -883 51 -849
rect 85 -883 119 -849
rect 153 -883 187 -849
rect 221 -883 255 -849
rect 289 -883 323 -849
rect 357 -883 391 -849
rect 425 -883 459 -849
rect 493 -883 527 -849
rect 561 -883 595 -849
rect 629 -883 663 -849
rect 697 -883 731 -849
rect 765 -883 799 -849
rect 833 -883 867 -849
rect 901 -883 1016 -849
<< viali >>
rect -902 664 -868 678
rect -902 644 -868 664
rect -902 596 -868 606
rect -902 572 -868 596
rect -902 528 -868 534
rect -902 500 -868 528
rect -902 460 -868 462
rect -902 428 -868 460
rect -902 358 -868 390
rect -902 356 -868 358
rect -902 290 -868 318
rect -902 284 -868 290
rect -902 222 -868 246
rect -902 212 -868 222
rect -902 154 -868 174
rect -902 140 -868 154
rect -784 664 -750 678
rect -784 644 -750 664
rect -784 596 -750 606
rect -784 572 -750 596
rect -784 528 -750 534
rect -784 500 -750 528
rect -784 460 -750 462
rect -784 428 -750 460
rect -784 358 -750 390
rect -784 356 -750 358
rect -784 290 -750 318
rect -784 284 -750 290
rect -784 222 -750 246
rect -784 212 -750 222
rect -784 154 -750 174
rect -784 140 -750 154
rect -666 664 -632 678
rect -666 644 -632 664
rect -666 596 -632 606
rect -666 572 -632 596
rect -666 528 -632 534
rect -666 500 -632 528
rect -666 460 -632 462
rect -666 428 -632 460
rect -666 358 -632 390
rect -666 356 -632 358
rect -666 290 -632 318
rect -666 284 -632 290
rect -666 222 -632 246
rect -666 212 -632 222
rect -666 154 -632 174
rect -666 140 -632 154
rect -548 664 -514 678
rect -548 644 -514 664
rect -548 596 -514 606
rect -548 572 -514 596
rect -548 528 -514 534
rect -548 500 -514 528
rect -548 460 -514 462
rect -548 428 -514 460
rect -548 358 -514 390
rect -548 356 -514 358
rect -548 290 -514 318
rect -548 284 -514 290
rect -548 222 -514 246
rect -548 212 -514 222
rect -548 154 -514 174
rect -548 140 -514 154
rect -430 664 -396 678
rect -430 644 -396 664
rect -430 596 -396 606
rect -430 572 -396 596
rect -430 528 -396 534
rect -430 500 -396 528
rect -430 460 -396 462
rect -430 428 -396 460
rect -430 358 -396 390
rect -430 356 -396 358
rect -430 290 -396 318
rect -430 284 -396 290
rect -430 222 -396 246
rect -430 212 -396 222
rect -430 154 -396 174
rect -430 140 -396 154
rect -312 664 -278 678
rect -312 644 -278 664
rect -312 596 -278 606
rect -312 572 -278 596
rect -312 528 -278 534
rect -312 500 -278 528
rect -312 460 -278 462
rect -312 428 -278 460
rect -312 358 -278 390
rect -312 356 -278 358
rect -312 290 -278 318
rect -312 284 -278 290
rect -312 222 -278 246
rect -312 212 -278 222
rect -312 154 -278 174
rect -312 140 -278 154
rect -194 664 -160 678
rect -194 644 -160 664
rect -194 596 -160 606
rect -194 572 -160 596
rect -194 528 -160 534
rect -194 500 -160 528
rect -194 460 -160 462
rect -194 428 -160 460
rect -194 358 -160 390
rect -194 356 -160 358
rect -194 290 -160 318
rect -194 284 -160 290
rect -194 222 -160 246
rect -194 212 -160 222
rect -194 154 -160 174
rect -194 140 -160 154
rect -76 664 -42 678
rect -76 644 -42 664
rect -76 596 -42 606
rect -76 572 -42 596
rect -76 528 -42 534
rect -76 500 -42 528
rect -76 460 -42 462
rect -76 428 -42 460
rect -76 358 -42 390
rect -76 356 -42 358
rect -76 290 -42 318
rect -76 284 -42 290
rect -76 222 -42 246
rect -76 212 -42 222
rect -76 154 -42 174
rect -76 140 -42 154
rect 42 664 76 678
rect 42 644 76 664
rect 42 596 76 606
rect 42 572 76 596
rect 42 528 76 534
rect 42 500 76 528
rect 42 460 76 462
rect 42 428 76 460
rect 42 358 76 390
rect 42 356 76 358
rect 42 290 76 318
rect 42 284 76 290
rect 42 222 76 246
rect 42 212 76 222
rect 42 154 76 174
rect 42 140 76 154
rect 160 664 194 678
rect 160 644 194 664
rect 160 596 194 606
rect 160 572 194 596
rect 160 528 194 534
rect 160 500 194 528
rect 160 460 194 462
rect 160 428 194 460
rect 160 358 194 390
rect 160 356 194 358
rect 160 290 194 318
rect 160 284 194 290
rect 160 222 194 246
rect 160 212 194 222
rect 160 154 194 174
rect 160 140 194 154
rect 278 664 312 678
rect 278 644 312 664
rect 278 596 312 606
rect 278 572 312 596
rect 278 528 312 534
rect 278 500 312 528
rect 278 460 312 462
rect 278 428 312 460
rect 278 358 312 390
rect 278 356 312 358
rect 278 290 312 318
rect 278 284 312 290
rect 278 222 312 246
rect 278 212 312 222
rect 278 154 312 174
rect 278 140 312 154
rect 396 664 430 678
rect 396 644 430 664
rect 396 596 430 606
rect 396 572 430 596
rect 396 528 430 534
rect 396 500 430 528
rect 396 460 430 462
rect 396 428 430 460
rect 396 358 430 390
rect 396 356 430 358
rect 396 290 430 318
rect 396 284 430 290
rect 396 222 430 246
rect 396 212 430 222
rect 396 154 430 174
rect 396 140 430 154
rect 514 664 548 678
rect 514 644 548 664
rect 514 596 548 606
rect 514 572 548 596
rect 514 528 548 534
rect 514 500 548 528
rect 514 460 548 462
rect 514 428 548 460
rect 514 358 548 390
rect 514 356 548 358
rect 514 290 548 318
rect 514 284 548 290
rect 514 222 548 246
rect 514 212 548 222
rect 514 154 548 174
rect 514 140 548 154
rect 632 664 666 678
rect 632 644 666 664
rect 632 596 666 606
rect 632 572 666 596
rect 632 528 666 534
rect 632 500 666 528
rect 632 460 666 462
rect 632 428 666 460
rect 632 358 666 390
rect 632 356 666 358
rect 632 290 666 318
rect 632 284 666 290
rect 632 222 666 246
rect 632 212 666 222
rect 632 154 666 174
rect 632 140 666 154
rect 750 664 784 678
rect 750 644 784 664
rect 750 596 784 606
rect 750 572 784 596
rect 750 528 784 534
rect 750 500 784 528
rect 750 460 784 462
rect 750 428 784 460
rect 750 358 784 390
rect 750 356 784 358
rect 750 290 784 318
rect 750 284 784 290
rect 750 222 784 246
rect 750 212 784 222
rect 750 154 784 174
rect 750 140 784 154
rect 868 664 902 678
rect 868 644 902 664
rect 868 596 902 606
rect 868 572 902 596
rect 868 528 902 534
rect 868 500 902 528
rect 868 460 902 462
rect 868 428 902 460
rect 868 358 902 390
rect 868 356 902 358
rect 868 290 902 318
rect 868 284 902 290
rect 868 222 902 246
rect 868 212 902 222
rect 868 154 902 174
rect 868 140 902 154
rect -843 37 -809 71
rect -725 37 -691 71
rect -607 37 -573 71
rect -489 37 -455 71
rect -371 37 -337 71
rect -253 37 -219 71
rect -135 37 -101 71
rect -17 37 17 71
rect 101 37 135 71
rect 219 37 253 71
rect 337 37 371 71
rect 455 37 489 71
rect 573 37 607 71
rect 691 37 725 71
rect 809 37 843 71
rect -843 -71 -809 -37
rect -725 -71 -691 -37
rect -607 -71 -573 -37
rect -489 -71 -455 -37
rect -371 -71 -337 -37
rect -253 -71 -219 -37
rect -135 -71 -101 -37
rect -17 -71 17 -37
rect 101 -71 135 -37
rect 219 -71 253 -37
rect 337 -71 371 -37
rect 455 -71 489 -37
rect 573 -71 607 -37
rect 691 -71 725 -37
rect 809 -71 843 -37
rect -902 -154 -868 -140
rect -902 -174 -868 -154
rect -902 -222 -868 -212
rect -902 -246 -868 -222
rect -902 -290 -868 -284
rect -902 -318 -868 -290
rect -902 -358 -868 -356
rect -902 -390 -868 -358
rect -902 -460 -868 -428
rect -902 -462 -868 -460
rect -902 -528 -868 -500
rect -902 -534 -868 -528
rect -902 -596 -868 -572
rect -902 -606 -868 -596
rect -902 -664 -868 -644
rect -902 -678 -868 -664
rect -784 -154 -750 -140
rect -784 -174 -750 -154
rect -784 -222 -750 -212
rect -784 -246 -750 -222
rect -784 -290 -750 -284
rect -784 -318 -750 -290
rect -784 -358 -750 -356
rect -784 -390 -750 -358
rect -784 -460 -750 -428
rect -784 -462 -750 -460
rect -784 -528 -750 -500
rect -784 -534 -750 -528
rect -784 -596 -750 -572
rect -784 -606 -750 -596
rect -784 -664 -750 -644
rect -784 -678 -750 -664
rect -666 -154 -632 -140
rect -666 -174 -632 -154
rect -666 -222 -632 -212
rect -666 -246 -632 -222
rect -666 -290 -632 -284
rect -666 -318 -632 -290
rect -666 -358 -632 -356
rect -666 -390 -632 -358
rect -666 -460 -632 -428
rect -666 -462 -632 -460
rect -666 -528 -632 -500
rect -666 -534 -632 -528
rect -666 -596 -632 -572
rect -666 -606 -632 -596
rect -666 -664 -632 -644
rect -666 -678 -632 -664
rect -548 -154 -514 -140
rect -548 -174 -514 -154
rect -548 -222 -514 -212
rect -548 -246 -514 -222
rect -548 -290 -514 -284
rect -548 -318 -514 -290
rect -548 -358 -514 -356
rect -548 -390 -514 -358
rect -548 -460 -514 -428
rect -548 -462 -514 -460
rect -548 -528 -514 -500
rect -548 -534 -514 -528
rect -548 -596 -514 -572
rect -548 -606 -514 -596
rect -548 -664 -514 -644
rect -548 -678 -514 -664
rect -430 -154 -396 -140
rect -430 -174 -396 -154
rect -430 -222 -396 -212
rect -430 -246 -396 -222
rect -430 -290 -396 -284
rect -430 -318 -396 -290
rect -430 -358 -396 -356
rect -430 -390 -396 -358
rect -430 -460 -396 -428
rect -430 -462 -396 -460
rect -430 -528 -396 -500
rect -430 -534 -396 -528
rect -430 -596 -396 -572
rect -430 -606 -396 -596
rect -430 -664 -396 -644
rect -430 -678 -396 -664
rect -312 -154 -278 -140
rect -312 -174 -278 -154
rect -312 -222 -278 -212
rect -312 -246 -278 -222
rect -312 -290 -278 -284
rect -312 -318 -278 -290
rect -312 -358 -278 -356
rect -312 -390 -278 -358
rect -312 -460 -278 -428
rect -312 -462 -278 -460
rect -312 -528 -278 -500
rect -312 -534 -278 -528
rect -312 -596 -278 -572
rect -312 -606 -278 -596
rect -312 -664 -278 -644
rect -312 -678 -278 -664
rect -194 -154 -160 -140
rect -194 -174 -160 -154
rect -194 -222 -160 -212
rect -194 -246 -160 -222
rect -194 -290 -160 -284
rect -194 -318 -160 -290
rect -194 -358 -160 -356
rect -194 -390 -160 -358
rect -194 -460 -160 -428
rect -194 -462 -160 -460
rect -194 -528 -160 -500
rect -194 -534 -160 -528
rect -194 -596 -160 -572
rect -194 -606 -160 -596
rect -194 -664 -160 -644
rect -194 -678 -160 -664
rect -76 -154 -42 -140
rect -76 -174 -42 -154
rect -76 -222 -42 -212
rect -76 -246 -42 -222
rect -76 -290 -42 -284
rect -76 -318 -42 -290
rect -76 -358 -42 -356
rect -76 -390 -42 -358
rect -76 -460 -42 -428
rect -76 -462 -42 -460
rect -76 -528 -42 -500
rect -76 -534 -42 -528
rect -76 -596 -42 -572
rect -76 -606 -42 -596
rect -76 -664 -42 -644
rect -76 -678 -42 -664
rect 42 -154 76 -140
rect 42 -174 76 -154
rect 42 -222 76 -212
rect 42 -246 76 -222
rect 42 -290 76 -284
rect 42 -318 76 -290
rect 42 -358 76 -356
rect 42 -390 76 -358
rect 42 -460 76 -428
rect 42 -462 76 -460
rect 42 -528 76 -500
rect 42 -534 76 -528
rect 42 -596 76 -572
rect 42 -606 76 -596
rect 42 -664 76 -644
rect 42 -678 76 -664
rect 160 -154 194 -140
rect 160 -174 194 -154
rect 160 -222 194 -212
rect 160 -246 194 -222
rect 160 -290 194 -284
rect 160 -318 194 -290
rect 160 -358 194 -356
rect 160 -390 194 -358
rect 160 -460 194 -428
rect 160 -462 194 -460
rect 160 -528 194 -500
rect 160 -534 194 -528
rect 160 -596 194 -572
rect 160 -606 194 -596
rect 160 -664 194 -644
rect 160 -678 194 -664
rect 278 -154 312 -140
rect 278 -174 312 -154
rect 278 -222 312 -212
rect 278 -246 312 -222
rect 278 -290 312 -284
rect 278 -318 312 -290
rect 278 -358 312 -356
rect 278 -390 312 -358
rect 278 -460 312 -428
rect 278 -462 312 -460
rect 278 -528 312 -500
rect 278 -534 312 -528
rect 278 -596 312 -572
rect 278 -606 312 -596
rect 278 -664 312 -644
rect 278 -678 312 -664
rect 396 -154 430 -140
rect 396 -174 430 -154
rect 396 -222 430 -212
rect 396 -246 430 -222
rect 396 -290 430 -284
rect 396 -318 430 -290
rect 396 -358 430 -356
rect 396 -390 430 -358
rect 396 -460 430 -428
rect 396 -462 430 -460
rect 396 -528 430 -500
rect 396 -534 430 -528
rect 396 -596 430 -572
rect 396 -606 430 -596
rect 396 -664 430 -644
rect 396 -678 430 -664
rect 514 -154 548 -140
rect 514 -174 548 -154
rect 514 -222 548 -212
rect 514 -246 548 -222
rect 514 -290 548 -284
rect 514 -318 548 -290
rect 514 -358 548 -356
rect 514 -390 548 -358
rect 514 -460 548 -428
rect 514 -462 548 -460
rect 514 -528 548 -500
rect 514 -534 548 -528
rect 514 -596 548 -572
rect 514 -606 548 -596
rect 514 -664 548 -644
rect 514 -678 548 -664
rect 632 -154 666 -140
rect 632 -174 666 -154
rect 632 -222 666 -212
rect 632 -246 666 -222
rect 632 -290 666 -284
rect 632 -318 666 -290
rect 632 -358 666 -356
rect 632 -390 666 -358
rect 632 -460 666 -428
rect 632 -462 666 -460
rect 632 -528 666 -500
rect 632 -534 666 -528
rect 632 -596 666 -572
rect 632 -606 666 -596
rect 632 -664 666 -644
rect 632 -678 666 -664
rect 750 -154 784 -140
rect 750 -174 784 -154
rect 750 -222 784 -212
rect 750 -246 784 -222
rect 750 -290 784 -284
rect 750 -318 784 -290
rect 750 -358 784 -356
rect 750 -390 784 -358
rect 750 -460 784 -428
rect 750 -462 784 -460
rect 750 -528 784 -500
rect 750 -534 784 -528
rect 750 -596 784 -572
rect 750 -606 784 -596
rect 750 -664 784 -644
rect 750 -678 784 -664
rect 868 -154 902 -140
rect 868 -174 902 -154
rect 868 -222 902 -212
rect 868 -246 902 -222
rect 868 -290 902 -284
rect 868 -318 902 -290
rect 868 -358 902 -356
rect 868 -390 902 -358
rect 868 -460 902 -428
rect 868 -462 902 -460
rect 868 -528 902 -500
rect 868 -534 902 -528
rect 868 -596 902 -572
rect 868 -606 902 -596
rect 868 -664 902 -644
rect 868 -678 902 -664
<< metal1 >>
rect -908 678 -862 709
rect -908 644 -902 678
rect -868 644 -862 678
rect -908 606 -862 644
rect -908 572 -902 606
rect -868 572 -862 606
rect -908 534 -862 572
rect -908 500 -902 534
rect -868 500 -862 534
rect -908 462 -862 500
rect -908 428 -902 462
rect -868 428 -862 462
rect -908 390 -862 428
rect -908 356 -902 390
rect -868 356 -862 390
rect -908 318 -862 356
rect -908 284 -902 318
rect -868 284 -862 318
rect -908 246 -862 284
rect -908 212 -902 246
rect -868 212 -862 246
rect -908 174 -862 212
rect -908 140 -902 174
rect -868 140 -862 174
rect -908 109 -862 140
rect -790 678 -744 709
rect -790 644 -784 678
rect -750 644 -744 678
rect -790 606 -744 644
rect -790 572 -784 606
rect -750 572 -744 606
rect -790 534 -744 572
rect -790 500 -784 534
rect -750 500 -744 534
rect -790 462 -744 500
rect -790 428 -784 462
rect -750 428 -744 462
rect -790 390 -744 428
rect -790 356 -784 390
rect -750 356 -744 390
rect -790 318 -744 356
rect -790 284 -784 318
rect -750 284 -744 318
rect -790 246 -744 284
rect -790 212 -784 246
rect -750 212 -744 246
rect -790 174 -744 212
rect -790 140 -784 174
rect -750 140 -744 174
rect -790 109 -744 140
rect -672 678 -626 709
rect -672 644 -666 678
rect -632 644 -626 678
rect -672 606 -626 644
rect -672 572 -666 606
rect -632 572 -626 606
rect -672 534 -626 572
rect -672 500 -666 534
rect -632 500 -626 534
rect -672 462 -626 500
rect -672 428 -666 462
rect -632 428 -626 462
rect -672 390 -626 428
rect -672 356 -666 390
rect -632 356 -626 390
rect -672 318 -626 356
rect -672 284 -666 318
rect -632 284 -626 318
rect -672 246 -626 284
rect -672 212 -666 246
rect -632 212 -626 246
rect -672 174 -626 212
rect -672 140 -666 174
rect -632 140 -626 174
rect -672 109 -626 140
rect -554 678 -508 709
rect -554 644 -548 678
rect -514 644 -508 678
rect -554 606 -508 644
rect -554 572 -548 606
rect -514 572 -508 606
rect -554 534 -508 572
rect -554 500 -548 534
rect -514 500 -508 534
rect -554 462 -508 500
rect -554 428 -548 462
rect -514 428 -508 462
rect -554 390 -508 428
rect -554 356 -548 390
rect -514 356 -508 390
rect -554 318 -508 356
rect -554 284 -548 318
rect -514 284 -508 318
rect -554 246 -508 284
rect -554 212 -548 246
rect -514 212 -508 246
rect -554 174 -508 212
rect -554 140 -548 174
rect -514 140 -508 174
rect -554 109 -508 140
rect -436 678 -390 709
rect -436 644 -430 678
rect -396 644 -390 678
rect -436 606 -390 644
rect -436 572 -430 606
rect -396 572 -390 606
rect -436 534 -390 572
rect -436 500 -430 534
rect -396 500 -390 534
rect -436 462 -390 500
rect -436 428 -430 462
rect -396 428 -390 462
rect -436 390 -390 428
rect -436 356 -430 390
rect -396 356 -390 390
rect -436 318 -390 356
rect -436 284 -430 318
rect -396 284 -390 318
rect -436 246 -390 284
rect -436 212 -430 246
rect -396 212 -390 246
rect -436 174 -390 212
rect -436 140 -430 174
rect -396 140 -390 174
rect -436 109 -390 140
rect -318 678 -272 709
rect -318 644 -312 678
rect -278 644 -272 678
rect -318 606 -272 644
rect -318 572 -312 606
rect -278 572 -272 606
rect -318 534 -272 572
rect -318 500 -312 534
rect -278 500 -272 534
rect -318 462 -272 500
rect -318 428 -312 462
rect -278 428 -272 462
rect -318 390 -272 428
rect -318 356 -312 390
rect -278 356 -272 390
rect -318 318 -272 356
rect -318 284 -312 318
rect -278 284 -272 318
rect -318 246 -272 284
rect -318 212 -312 246
rect -278 212 -272 246
rect -318 174 -272 212
rect -318 140 -312 174
rect -278 140 -272 174
rect -318 109 -272 140
rect -200 678 -154 709
rect -200 644 -194 678
rect -160 644 -154 678
rect -200 606 -154 644
rect -200 572 -194 606
rect -160 572 -154 606
rect -200 534 -154 572
rect -200 500 -194 534
rect -160 500 -154 534
rect -200 462 -154 500
rect -200 428 -194 462
rect -160 428 -154 462
rect -200 390 -154 428
rect -200 356 -194 390
rect -160 356 -154 390
rect -200 318 -154 356
rect -200 284 -194 318
rect -160 284 -154 318
rect -200 246 -154 284
rect -200 212 -194 246
rect -160 212 -154 246
rect -200 174 -154 212
rect -200 140 -194 174
rect -160 140 -154 174
rect -200 109 -154 140
rect -82 678 -36 709
rect -82 644 -76 678
rect -42 644 -36 678
rect -82 606 -36 644
rect -82 572 -76 606
rect -42 572 -36 606
rect -82 534 -36 572
rect -82 500 -76 534
rect -42 500 -36 534
rect -82 462 -36 500
rect -82 428 -76 462
rect -42 428 -36 462
rect -82 390 -36 428
rect -82 356 -76 390
rect -42 356 -36 390
rect -82 318 -36 356
rect -82 284 -76 318
rect -42 284 -36 318
rect -82 246 -36 284
rect -82 212 -76 246
rect -42 212 -36 246
rect -82 174 -36 212
rect -82 140 -76 174
rect -42 140 -36 174
rect -82 109 -36 140
rect 36 678 82 709
rect 36 644 42 678
rect 76 644 82 678
rect 36 606 82 644
rect 36 572 42 606
rect 76 572 82 606
rect 36 534 82 572
rect 36 500 42 534
rect 76 500 82 534
rect 36 462 82 500
rect 36 428 42 462
rect 76 428 82 462
rect 36 390 82 428
rect 36 356 42 390
rect 76 356 82 390
rect 36 318 82 356
rect 36 284 42 318
rect 76 284 82 318
rect 36 246 82 284
rect 36 212 42 246
rect 76 212 82 246
rect 36 174 82 212
rect 36 140 42 174
rect 76 140 82 174
rect 36 109 82 140
rect 154 678 200 709
rect 154 644 160 678
rect 194 644 200 678
rect 154 606 200 644
rect 154 572 160 606
rect 194 572 200 606
rect 154 534 200 572
rect 154 500 160 534
rect 194 500 200 534
rect 154 462 200 500
rect 154 428 160 462
rect 194 428 200 462
rect 154 390 200 428
rect 154 356 160 390
rect 194 356 200 390
rect 154 318 200 356
rect 154 284 160 318
rect 194 284 200 318
rect 154 246 200 284
rect 154 212 160 246
rect 194 212 200 246
rect 154 174 200 212
rect 154 140 160 174
rect 194 140 200 174
rect 154 109 200 140
rect 272 678 318 709
rect 272 644 278 678
rect 312 644 318 678
rect 272 606 318 644
rect 272 572 278 606
rect 312 572 318 606
rect 272 534 318 572
rect 272 500 278 534
rect 312 500 318 534
rect 272 462 318 500
rect 272 428 278 462
rect 312 428 318 462
rect 272 390 318 428
rect 272 356 278 390
rect 312 356 318 390
rect 272 318 318 356
rect 272 284 278 318
rect 312 284 318 318
rect 272 246 318 284
rect 272 212 278 246
rect 312 212 318 246
rect 272 174 318 212
rect 272 140 278 174
rect 312 140 318 174
rect 272 109 318 140
rect 390 678 436 709
rect 390 644 396 678
rect 430 644 436 678
rect 390 606 436 644
rect 390 572 396 606
rect 430 572 436 606
rect 390 534 436 572
rect 390 500 396 534
rect 430 500 436 534
rect 390 462 436 500
rect 390 428 396 462
rect 430 428 436 462
rect 390 390 436 428
rect 390 356 396 390
rect 430 356 436 390
rect 390 318 436 356
rect 390 284 396 318
rect 430 284 436 318
rect 390 246 436 284
rect 390 212 396 246
rect 430 212 436 246
rect 390 174 436 212
rect 390 140 396 174
rect 430 140 436 174
rect 390 109 436 140
rect 508 678 554 709
rect 508 644 514 678
rect 548 644 554 678
rect 508 606 554 644
rect 508 572 514 606
rect 548 572 554 606
rect 508 534 554 572
rect 508 500 514 534
rect 548 500 554 534
rect 508 462 554 500
rect 508 428 514 462
rect 548 428 554 462
rect 508 390 554 428
rect 508 356 514 390
rect 548 356 554 390
rect 508 318 554 356
rect 508 284 514 318
rect 548 284 554 318
rect 508 246 554 284
rect 508 212 514 246
rect 548 212 554 246
rect 508 174 554 212
rect 508 140 514 174
rect 548 140 554 174
rect 508 109 554 140
rect 626 678 672 709
rect 626 644 632 678
rect 666 644 672 678
rect 626 606 672 644
rect 626 572 632 606
rect 666 572 672 606
rect 626 534 672 572
rect 626 500 632 534
rect 666 500 672 534
rect 626 462 672 500
rect 626 428 632 462
rect 666 428 672 462
rect 626 390 672 428
rect 626 356 632 390
rect 666 356 672 390
rect 626 318 672 356
rect 626 284 632 318
rect 666 284 672 318
rect 626 246 672 284
rect 626 212 632 246
rect 666 212 672 246
rect 626 174 672 212
rect 626 140 632 174
rect 666 140 672 174
rect 626 109 672 140
rect 744 678 790 709
rect 744 644 750 678
rect 784 644 790 678
rect 744 606 790 644
rect 744 572 750 606
rect 784 572 790 606
rect 744 534 790 572
rect 744 500 750 534
rect 784 500 790 534
rect 744 462 790 500
rect 744 428 750 462
rect 784 428 790 462
rect 744 390 790 428
rect 744 356 750 390
rect 784 356 790 390
rect 744 318 790 356
rect 744 284 750 318
rect 784 284 790 318
rect 744 246 790 284
rect 744 212 750 246
rect 784 212 790 246
rect 744 174 790 212
rect 744 140 750 174
rect 784 140 790 174
rect 744 109 790 140
rect 862 678 908 709
rect 862 644 868 678
rect 902 644 908 678
rect 862 606 908 644
rect 862 572 868 606
rect 902 572 908 606
rect 862 534 908 572
rect 862 500 868 534
rect 902 500 908 534
rect 862 462 908 500
rect 862 428 868 462
rect 902 428 908 462
rect 862 390 908 428
rect 862 356 868 390
rect 902 356 908 390
rect 862 318 908 356
rect 862 284 868 318
rect 902 284 908 318
rect 862 246 908 284
rect 862 212 868 246
rect 902 212 908 246
rect 862 174 908 212
rect 862 140 868 174
rect 902 140 908 174
rect 862 109 908 140
rect -855 71 -797 77
rect -855 37 -843 71
rect -809 37 -797 71
rect -855 31 -797 37
rect -737 71 -679 77
rect -737 37 -725 71
rect -691 37 -679 71
rect -737 31 -679 37
rect -619 71 -561 77
rect -619 37 -607 71
rect -573 37 -561 71
rect -619 31 -561 37
rect -501 71 -443 77
rect -501 37 -489 71
rect -455 37 -443 71
rect -501 31 -443 37
rect -383 71 -325 77
rect -383 37 -371 71
rect -337 37 -325 71
rect -383 31 -325 37
rect -265 71 -207 77
rect -265 37 -253 71
rect -219 37 -207 71
rect -265 31 -207 37
rect -147 71 -89 77
rect -147 37 -135 71
rect -101 37 -89 71
rect -147 31 -89 37
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect 89 71 147 77
rect 89 37 101 71
rect 135 37 147 71
rect 89 31 147 37
rect 207 71 265 77
rect 207 37 219 71
rect 253 37 265 71
rect 207 31 265 37
rect 325 71 383 77
rect 325 37 337 71
rect 371 37 383 71
rect 325 31 383 37
rect 443 71 501 77
rect 443 37 455 71
rect 489 37 501 71
rect 443 31 501 37
rect 561 71 619 77
rect 561 37 573 71
rect 607 37 619 71
rect 561 31 619 37
rect 679 71 737 77
rect 679 37 691 71
rect 725 37 737 71
rect 679 31 737 37
rect 797 71 855 77
rect 797 37 809 71
rect 843 37 855 71
rect 797 31 855 37
rect -855 -37 -797 -31
rect -855 -71 -843 -37
rect -809 -71 -797 -37
rect -855 -77 -797 -71
rect -737 -37 -679 -31
rect -737 -71 -725 -37
rect -691 -71 -679 -37
rect -737 -77 -679 -71
rect -619 -37 -561 -31
rect -619 -71 -607 -37
rect -573 -71 -561 -37
rect -619 -77 -561 -71
rect -501 -37 -443 -31
rect -501 -71 -489 -37
rect -455 -71 -443 -37
rect -501 -77 -443 -71
rect -383 -37 -325 -31
rect -383 -71 -371 -37
rect -337 -71 -325 -37
rect -383 -77 -325 -71
rect -265 -37 -207 -31
rect -265 -71 -253 -37
rect -219 -71 -207 -37
rect -265 -77 -207 -71
rect -147 -37 -89 -31
rect -147 -71 -135 -37
rect -101 -71 -89 -37
rect -147 -77 -89 -71
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect 89 -37 147 -31
rect 89 -71 101 -37
rect 135 -71 147 -37
rect 89 -77 147 -71
rect 207 -37 265 -31
rect 207 -71 219 -37
rect 253 -71 265 -37
rect 207 -77 265 -71
rect 325 -37 383 -31
rect 325 -71 337 -37
rect 371 -71 383 -37
rect 325 -77 383 -71
rect 443 -37 501 -31
rect 443 -71 455 -37
rect 489 -71 501 -37
rect 443 -77 501 -71
rect 561 -37 619 -31
rect 561 -71 573 -37
rect 607 -71 619 -37
rect 561 -77 619 -71
rect 679 -37 737 -31
rect 679 -71 691 -37
rect 725 -71 737 -37
rect 679 -77 737 -71
rect 797 -37 855 -31
rect 797 -71 809 -37
rect 843 -71 855 -37
rect 797 -77 855 -71
rect -908 -140 -862 -109
rect -908 -174 -902 -140
rect -868 -174 -862 -140
rect -908 -212 -862 -174
rect -908 -246 -902 -212
rect -868 -246 -862 -212
rect -908 -284 -862 -246
rect -908 -318 -902 -284
rect -868 -318 -862 -284
rect -908 -356 -862 -318
rect -908 -390 -902 -356
rect -868 -390 -862 -356
rect -908 -428 -862 -390
rect -908 -462 -902 -428
rect -868 -462 -862 -428
rect -908 -500 -862 -462
rect -908 -534 -902 -500
rect -868 -534 -862 -500
rect -908 -572 -862 -534
rect -908 -606 -902 -572
rect -868 -606 -862 -572
rect -908 -644 -862 -606
rect -908 -678 -902 -644
rect -868 -678 -862 -644
rect -908 -709 -862 -678
rect -790 -140 -744 -109
rect -790 -174 -784 -140
rect -750 -174 -744 -140
rect -790 -212 -744 -174
rect -790 -246 -784 -212
rect -750 -246 -744 -212
rect -790 -284 -744 -246
rect -790 -318 -784 -284
rect -750 -318 -744 -284
rect -790 -356 -744 -318
rect -790 -390 -784 -356
rect -750 -390 -744 -356
rect -790 -428 -744 -390
rect -790 -462 -784 -428
rect -750 -462 -744 -428
rect -790 -500 -744 -462
rect -790 -534 -784 -500
rect -750 -534 -744 -500
rect -790 -572 -744 -534
rect -790 -606 -784 -572
rect -750 -606 -744 -572
rect -790 -644 -744 -606
rect -790 -678 -784 -644
rect -750 -678 -744 -644
rect -790 -709 -744 -678
rect -672 -140 -626 -109
rect -672 -174 -666 -140
rect -632 -174 -626 -140
rect -672 -212 -626 -174
rect -672 -246 -666 -212
rect -632 -246 -626 -212
rect -672 -284 -626 -246
rect -672 -318 -666 -284
rect -632 -318 -626 -284
rect -672 -356 -626 -318
rect -672 -390 -666 -356
rect -632 -390 -626 -356
rect -672 -428 -626 -390
rect -672 -462 -666 -428
rect -632 -462 -626 -428
rect -672 -500 -626 -462
rect -672 -534 -666 -500
rect -632 -534 -626 -500
rect -672 -572 -626 -534
rect -672 -606 -666 -572
rect -632 -606 -626 -572
rect -672 -644 -626 -606
rect -672 -678 -666 -644
rect -632 -678 -626 -644
rect -672 -709 -626 -678
rect -554 -140 -508 -109
rect -554 -174 -548 -140
rect -514 -174 -508 -140
rect -554 -212 -508 -174
rect -554 -246 -548 -212
rect -514 -246 -508 -212
rect -554 -284 -508 -246
rect -554 -318 -548 -284
rect -514 -318 -508 -284
rect -554 -356 -508 -318
rect -554 -390 -548 -356
rect -514 -390 -508 -356
rect -554 -428 -508 -390
rect -554 -462 -548 -428
rect -514 -462 -508 -428
rect -554 -500 -508 -462
rect -554 -534 -548 -500
rect -514 -534 -508 -500
rect -554 -572 -508 -534
rect -554 -606 -548 -572
rect -514 -606 -508 -572
rect -554 -644 -508 -606
rect -554 -678 -548 -644
rect -514 -678 -508 -644
rect -554 -709 -508 -678
rect -436 -140 -390 -109
rect -436 -174 -430 -140
rect -396 -174 -390 -140
rect -436 -212 -390 -174
rect -436 -246 -430 -212
rect -396 -246 -390 -212
rect -436 -284 -390 -246
rect -436 -318 -430 -284
rect -396 -318 -390 -284
rect -436 -356 -390 -318
rect -436 -390 -430 -356
rect -396 -390 -390 -356
rect -436 -428 -390 -390
rect -436 -462 -430 -428
rect -396 -462 -390 -428
rect -436 -500 -390 -462
rect -436 -534 -430 -500
rect -396 -534 -390 -500
rect -436 -572 -390 -534
rect -436 -606 -430 -572
rect -396 -606 -390 -572
rect -436 -644 -390 -606
rect -436 -678 -430 -644
rect -396 -678 -390 -644
rect -436 -709 -390 -678
rect -318 -140 -272 -109
rect -318 -174 -312 -140
rect -278 -174 -272 -140
rect -318 -212 -272 -174
rect -318 -246 -312 -212
rect -278 -246 -272 -212
rect -318 -284 -272 -246
rect -318 -318 -312 -284
rect -278 -318 -272 -284
rect -318 -356 -272 -318
rect -318 -390 -312 -356
rect -278 -390 -272 -356
rect -318 -428 -272 -390
rect -318 -462 -312 -428
rect -278 -462 -272 -428
rect -318 -500 -272 -462
rect -318 -534 -312 -500
rect -278 -534 -272 -500
rect -318 -572 -272 -534
rect -318 -606 -312 -572
rect -278 -606 -272 -572
rect -318 -644 -272 -606
rect -318 -678 -312 -644
rect -278 -678 -272 -644
rect -318 -709 -272 -678
rect -200 -140 -154 -109
rect -200 -174 -194 -140
rect -160 -174 -154 -140
rect -200 -212 -154 -174
rect -200 -246 -194 -212
rect -160 -246 -154 -212
rect -200 -284 -154 -246
rect -200 -318 -194 -284
rect -160 -318 -154 -284
rect -200 -356 -154 -318
rect -200 -390 -194 -356
rect -160 -390 -154 -356
rect -200 -428 -154 -390
rect -200 -462 -194 -428
rect -160 -462 -154 -428
rect -200 -500 -154 -462
rect -200 -534 -194 -500
rect -160 -534 -154 -500
rect -200 -572 -154 -534
rect -200 -606 -194 -572
rect -160 -606 -154 -572
rect -200 -644 -154 -606
rect -200 -678 -194 -644
rect -160 -678 -154 -644
rect -200 -709 -154 -678
rect -82 -140 -36 -109
rect -82 -174 -76 -140
rect -42 -174 -36 -140
rect -82 -212 -36 -174
rect -82 -246 -76 -212
rect -42 -246 -36 -212
rect -82 -284 -36 -246
rect -82 -318 -76 -284
rect -42 -318 -36 -284
rect -82 -356 -36 -318
rect -82 -390 -76 -356
rect -42 -390 -36 -356
rect -82 -428 -36 -390
rect -82 -462 -76 -428
rect -42 -462 -36 -428
rect -82 -500 -36 -462
rect -82 -534 -76 -500
rect -42 -534 -36 -500
rect -82 -572 -36 -534
rect -82 -606 -76 -572
rect -42 -606 -36 -572
rect -82 -644 -36 -606
rect -82 -678 -76 -644
rect -42 -678 -36 -644
rect -82 -709 -36 -678
rect 36 -140 82 -109
rect 36 -174 42 -140
rect 76 -174 82 -140
rect 36 -212 82 -174
rect 36 -246 42 -212
rect 76 -246 82 -212
rect 36 -284 82 -246
rect 36 -318 42 -284
rect 76 -318 82 -284
rect 36 -356 82 -318
rect 36 -390 42 -356
rect 76 -390 82 -356
rect 36 -428 82 -390
rect 36 -462 42 -428
rect 76 -462 82 -428
rect 36 -500 82 -462
rect 36 -534 42 -500
rect 76 -534 82 -500
rect 36 -572 82 -534
rect 36 -606 42 -572
rect 76 -606 82 -572
rect 36 -644 82 -606
rect 36 -678 42 -644
rect 76 -678 82 -644
rect 36 -709 82 -678
rect 154 -140 200 -109
rect 154 -174 160 -140
rect 194 -174 200 -140
rect 154 -212 200 -174
rect 154 -246 160 -212
rect 194 -246 200 -212
rect 154 -284 200 -246
rect 154 -318 160 -284
rect 194 -318 200 -284
rect 154 -356 200 -318
rect 154 -390 160 -356
rect 194 -390 200 -356
rect 154 -428 200 -390
rect 154 -462 160 -428
rect 194 -462 200 -428
rect 154 -500 200 -462
rect 154 -534 160 -500
rect 194 -534 200 -500
rect 154 -572 200 -534
rect 154 -606 160 -572
rect 194 -606 200 -572
rect 154 -644 200 -606
rect 154 -678 160 -644
rect 194 -678 200 -644
rect 154 -709 200 -678
rect 272 -140 318 -109
rect 272 -174 278 -140
rect 312 -174 318 -140
rect 272 -212 318 -174
rect 272 -246 278 -212
rect 312 -246 318 -212
rect 272 -284 318 -246
rect 272 -318 278 -284
rect 312 -318 318 -284
rect 272 -356 318 -318
rect 272 -390 278 -356
rect 312 -390 318 -356
rect 272 -428 318 -390
rect 272 -462 278 -428
rect 312 -462 318 -428
rect 272 -500 318 -462
rect 272 -534 278 -500
rect 312 -534 318 -500
rect 272 -572 318 -534
rect 272 -606 278 -572
rect 312 -606 318 -572
rect 272 -644 318 -606
rect 272 -678 278 -644
rect 312 -678 318 -644
rect 272 -709 318 -678
rect 390 -140 436 -109
rect 390 -174 396 -140
rect 430 -174 436 -140
rect 390 -212 436 -174
rect 390 -246 396 -212
rect 430 -246 436 -212
rect 390 -284 436 -246
rect 390 -318 396 -284
rect 430 -318 436 -284
rect 390 -356 436 -318
rect 390 -390 396 -356
rect 430 -390 436 -356
rect 390 -428 436 -390
rect 390 -462 396 -428
rect 430 -462 436 -428
rect 390 -500 436 -462
rect 390 -534 396 -500
rect 430 -534 436 -500
rect 390 -572 436 -534
rect 390 -606 396 -572
rect 430 -606 436 -572
rect 390 -644 436 -606
rect 390 -678 396 -644
rect 430 -678 436 -644
rect 390 -709 436 -678
rect 508 -140 554 -109
rect 508 -174 514 -140
rect 548 -174 554 -140
rect 508 -212 554 -174
rect 508 -246 514 -212
rect 548 -246 554 -212
rect 508 -284 554 -246
rect 508 -318 514 -284
rect 548 -318 554 -284
rect 508 -356 554 -318
rect 508 -390 514 -356
rect 548 -390 554 -356
rect 508 -428 554 -390
rect 508 -462 514 -428
rect 548 -462 554 -428
rect 508 -500 554 -462
rect 508 -534 514 -500
rect 548 -534 554 -500
rect 508 -572 554 -534
rect 508 -606 514 -572
rect 548 -606 554 -572
rect 508 -644 554 -606
rect 508 -678 514 -644
rect 548 -678 554 -644
rect 508 -709 554 -678
rect 626 -140 672 -109
rect 626 -174 632 -140
rect 666 -174 672 -140
rect 626 -212 672 -174
rect 626 -246 632 -212
rect 666 -246 672 -212
rect 626 -284 672 -246
rect 626 -318 632 -284
rect 666 -318 672 -284
rect 626 -356 672 -318
rect 626 -390 632 -356
rect 666 -390 672 -356
rect 626 -428 672 -390
rect 626 -462 632 -428
rect 666 -462 672 -428
rect 626 -500 672 -462
rect 626 -534 632 -500
rect 666 -534 672 -500
rect 626 -572 672 -534
rect 626 -606 632 -572
rect 666 -606 672 -572
rect 626 -644 672 -606
rect 626 -678 632 -644
rect 666 -678 672 -644
rect 626 -709 672 -678
rect 744 -140 790 -109
rect 744 -174 750 -140
rect 784 -174 790 -140
rect 744 -212 790 -174
rect 744 -246 750 -212
rect 784 -246 790 -212
rect 744 -284 790 -246
rect 744 -318 750 -284
rect 784 -318 790 -284
rect 744 -356 790 -318
rect 744 -390 750 -356
rect 784 -390 790 -356
rect 744 -428 790 -390
rect 744 -462 750 -428
rect 784 -462 790 -428
rect 744 -500 790 -462
rect 744 -534 750 -500
rect 784 -534 790 -500
rect 744 -572 790 -534
rect 744 -606 750 -572
rect 784 -606 790 -572
rect 744 -644 790 -606
rect 744 -678 750 -644
rect 784 -678 790 -644
rect 744 -709 790 -678
rect 862 -140 908 -109
rect 862 -174 868 -140
rect 902 -174 908 -140
rect 862 -212 908 -174
rect 862 -246 868 -212
rect 902 -246 908 -212
rect 862 -284 908 -246
rect 862 -318 868 -284
rect 902 -318 908 -284
rect 862 -356 908 -318
rect 862 -390 868 -356
rect 902 -390 908 -356
rect 862 -428 908 -390
rect 862 -462 868 -428
rect 902 -462 908 -428
rect 862 -500 908 -462
rect 862 -534 868 -500
rect 902 -534 908 -500
rect 862 -572 908 -534
rect 862 -606 868 -572
rect 902 -606 908 -572
rect 862 -644 908 -606
rect 862 -678 868 -644
rect 902 -678 908 -644
rect 862 -709 908 -678
<< properties >>
string FIXED_BBOX -999 -866 999 866
<< end >>
