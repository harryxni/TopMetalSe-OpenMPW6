magic
tech sky130A
magscale 1 2
timestamp 1608254796
<< nwell >>
rect -211 -436 211 459
<< pmos >>
rect -15 -240 15 240
<< pdiff >>
rect -73 228 -15 240
rect -73 -228 -61 228
rect -27 -228 -15 228
rect -73 -240 -15 -228
rect 15 228 73 240
rect 15 -228 27 228
rect 61 -228 73 228
rect 15 -240 73 -228
<< pdiffc >>
rect -61 -228 -27 228
rect 27 -228 61 228
<< nsubdiff >>
rect -175 389 -79 423
rect 79 389 175 423
rect -175 327 -141 389
rect 141 327 175 389
rect -175 -364 -141 -327
rect 141 -384 175 -327
<< nsubdiffcont >>
rect -79 389 79 423
rect -175 -327 -141 327
rect 141 -327 175 327
<< poly >>
rect -15 240 15 338
rect -15 -321 15 -240
<< locali >>
rect -175 389 -79 423
rect 79 389 175 423
rect -175 327 -141 389
rect 141 327 175 389
rect -61 228 -27 244
rect -61 -244 -27 -228
rect 27 228 61 244
rect 27 -244 61 -228
rect -175 -364 -141 -327
rect 141 -384 175 -327
<< viali >>
rect -61 -228 -27 228
rect 27 -228 61 228
<< metal1 >>
rect -67 228 -21 240
rect -67 -228 -61 228
rect -27 -228 -21 228
rect -67 -240 -21 -228
rect 21 228 67 240
rect 21 -228 27 228
rect 61 -228 67 228
rect 21 -240 67 -228
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -158 -406 158 406
string parameters w 2.4 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
