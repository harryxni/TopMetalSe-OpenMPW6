magic
tech sky130A
magscale 1 2
timestamp 1654749028
<< error_p >>
rect 13533 16441 13541 16463
rect 13793 16441 13895 16450
rect 14265 16441 14367 16462
rect 14973 16441 15075 16447
rect 15791 16441 15893 16462
rect 16027 16441 16129 16447
rect 16499 16441 16601 16450
rect 16971 16441 17073 16459
rect 17789 16441 17891 16462
rect 18025 16441 18127 16447
rect 18497 16441 18599 16450
rect 18969 16441 19071 16459
rect 13561 16419 13569 16441
rect 13557 16374 13569 16419
rect 13821 16413 13867 16422
rect 14293 16413 14339 16434
rect 15001 16413 15047 16419
rect 15819 16413 15865 16434
rect 16055 16413 16101 16419
rect 16527 16413 16573 16422
rect 16999 16413 17045 16431
rect 17817 16413 17863 16434
rect 18053 16413 18099 16419
rect 18525 16413 18571 16422
rect 18997 16413 19043 16431
rect 27379 16393 27413 16427
rect 32612 16401 32639 16439
rect 32640 16429 32667 16439
rect 13585 16346 13589 16391
rect 32628 16373 32639 16401
rect 14389 16245 14479 16261
rect 14389 16233 14411 16245
rect 14417 16233 14451 16245
rect 14417 16225 14439 16233
rect 14457 16225 14479 16245
rect 14625 16245 14715 16261
rect 14625 16233 14647 16245
rect 14653 16233 14687 16245
rect 14653 16225 14675 16233
rect 14693 16225 14715 16245
rect 14861 16245 14951 16261
rect 14861 16233 14883 16245
rect 14889 16233 14923 16245
rect 14889 16225 14911 16233
rect 14929 16225 14951 16245
rect 15097 16245 15187 16261
rect 15097 16233 15119 16245
rect 15125 16233 15159 16245
rect 15125 16225 15147 16233
rect 15165 16225 15187 16245
rect 15333 16245 15423 16261
rect 15333 16233 15355 16245
rect 15361 16233 15395 16245
rect 15361 16225 15383 16233
rect 15401 16225 15423 16245
rect 16623 16245 16713 16261
rect 16623 16233 16645 16245
rect 16651 16233 16685 16245
rect 16651 16225 16673 16233
rect 16691 16225 16713 16245
rect 17095 16245 17185 16261
rect 17095 16233 17117 16245
rect 17123 16233 17157 16245
rect 17123 16225 17145 16233
rect 17163 16225 17185 16245
rect 17677 16245 17767 16261
rect 17677 16233 17699 16245
rect 17705 16233 17739 16245
rect 17705 16225 17727 16233
rect 17745 16225 17767 16245
rect 18149 16245 18239 16261
rect 18149 16233 18171 16245
rect 18177 16233 18211 16245
rect 18177 16225 18199 16233
rect 18217 16225 18239 16245
rect 18621 16245 18711 16261
rect 18621 16233 18643 16245
rect 18649 16233 18683 16245
rect 18649 16225 18671 16233
rect 18689 16225 18711 16245
rect 19093 16245 19183 16261
rect 19093 16233 19115 16245
rect 19121 16233 19155 16245
rect 19121 16225 19143 16233
rect 19161 16225 19183 16245
rect 21753 16232 21769 16248
rect 21771 16232 21787 16248
rect 21871 16232 21887 16248
rect 21889 16232 21905 16248
rect 21989 16232 22005 16248
rect 22007 16232 22023 16248
rect 22107 16232 22123 16248
rect 22125 16232 22141 16248
rect 22225 16232 22241 16248
rect 22243 16232 22259 16248
rect 22343 16232 22359 16248
rect 22361 16232 22377 16248
rect 22461 16232 22477 16248
rect 22479 16232 22495 16248
rect 22579 16232 22595 16248
rect 22597 16232 22613 16248
rect 22697 16232 22713 16248
rect 22715 16232 22731 16248
rect 22815 16232 22831 16248
rect 22833 16232 22849 16248
rect 22933 16232 22949 16248
rect 22951 16232 22967 16248
rect 23051 16232 23067 16248
rect 23069 16232 23085 16248
rect 23169 16232 23185 16248
rect 23187 16232 23203 16248
rect 23287 16232 23303 16248
rect 23305 16232 23321 16248
rect 23405 16232 23421 16248
rect 23423 16232 23439 16248
rect 23523 16232 23539 16248
rect 23541 16232 23557 16248
rect 23641 16232 23657 16248
rect 23659 16232 23675 16248
rect 23759 16232 23775 16248
rect 23777 16232 23793 16248
rect 23877 16232 23893 16248
rect 23895 16232 23911 16248
rect 23995 16232 24011 16248
rect 24013 16232 24029 16248
rect 24113 16232 24129 16248
rect 24131 16232 24147 16248
rect 24231 16232 24247 16248
rect 24249 16232 24265 16248
rect 25876 16232 25892 16248
rect 25894 16232 25910 16248
rect 25994 16232 26010 16248
rect 26012 16232 26028 16248
rect 26112 16232 26128 16248
rect 26130 16232 26146 16248
rect 26230 16232 26246 16248
rect 26248 16232 26264 16248
rect 26348 16232 26364 16248
rect 26366 16232 26382 16248
rect 26466 16232 26482 16248
rect 26484 16232 26500 16248
rect 26584 16232 26600 16248
rect 26602 16232 26618 16248
rect 26702 16232 26718 16248
rect 26720 16232 26736 16248
rect 26820 16232 26836 16248
rect 26838 16232 26854 16248
rect 26938 16232 26954 16248
rect 26956 16232 26972 16248
rect 27056 16232 27072 16248
rect 27074 16232 27090 16248
rect 27174 16232 27190 16248
rect 27192 16232 27208 16248
rect 27292 16232 27308 16248
rect 27310 16232 27326 16248
rect 27410 16232 27426 16248
rect 27428 16232 27444 16248
rect 27528 16232 27544 16248
rect 27546 16232 27562 16248
rect 27646 16232 27662 16248
rect 27664 16232 27680 16248
rect 27764 16232 27780 16248
rect 27782 16232 27798 16248
rect 27882 16232 27898 16248
rect 27900 16232 27916 16248
rect 28000 16232 28016 16248
rect 28018 16232 28034 16248
rect 28118 16232 28134 16248
rect 28136 16232 28152 16248
rect 28236 16232 28252 16248
rect 28254 16232 28270 16248
rect 28354 16232 28370 16248
rect 28372 16232 28388 16248
rect 29999 16232 30015 16248
rect 30017 16232 30033 16248
rect 30117 16232 30133 16248
rect 30135 16232 30151 16248
rect 30235 16232 30251 16248
rect 30253 16232 30269 16248
rect 30353 16232 30369 16248
rect 30371 16232 30387 16248
rect 30471 16232 30487 16248
rect 30489 16232 30505 16248
rect 30589 16232 30605 16248
rect 30607 16232 30623 16248
rect 30707 16232 30723 16248
rect 30725 16232 30741 16248
rect 30825 16232 30841 16248
rect 30843 16232 30859 16248
rect 30943 16232 30959 16248
rect 30961 16232 30977 16248
rect 31061 16232 31077 16248
rect 31079 16232 31095 16248
rect 31179 16232 31195 16248
rect 31197 16232 31213 16248
rect 31297 16232 31313 16248
rect 31315 16232 31331 16248
rect 31415 16232 31431 16248
rect 31433 16232 31449 16248
rect 31533 16232 31549 16248
rect 31551 16232 31567 16248
rect 31651 16232 31667 16248
rect 31669 16232 31685 16248
rect 31769 16232 31785 16248
rect 31787 16232 31803 16248
rect 31887 16232 31903 16248
rect 31905 16232 31921 16248
rect 32005 16232 32021 16248
rect 32023 16232 32039 16248
rect 32123 16232 32139 16248
rect 32141 16232 32157 16248
rect 32241 16232 32257 16248
rect 32259 16232 32275 16248
rect 32359 16232 32375 16248
rect 32377 16232 32393 16248
rect 32477 16232 32493 16248
rect 32495 16232 32511 16248
rect 14417 16205 14451 16225
rect 14653 16205 14687 16225
rect 14889 16205 14923 16225
rect 15125 16205 15159 16225
rect 15361 16205 15395 16225
rect 16651 16205 16685 16225
rect 17123 16205 17157 16225
rect 17705 16205 17739 16225
rect 18177 16205 18211 16225
rect 18649 16205 18683 16225
rect 19121 16205 19155 16225
rect 21737 16224 21803 16232
rect 21737 16216 21761 16224
rect 14389 15665 14398 15693
rect 14417 15645 14451 15685
rect 14470 15665 14479 15693
rect 14625 15665 14634 15693
rect 14457 15657 14479 15665
rect 14653 15645 14687 15685
rect 14706 15665 14715 15693
rect 14861 15665 14870 15693
rect 14693 15657 14715 15665
rect 14889 15645 14923 15685
rect 14942 15665 14951 15693
rect 15097 15665 15106 15693
rect 14929 15657 14951 15665
rect 15125 15645 15159 15685
rect 15178 15665 15187 15693
rect 15333 15665 15342 15693
rect 15165 15657 15187 15665
rect 15361 15645 15395 15685
rect 15414 15665 15423 15693
rect 16623 15665 16632 15693
rect 15401 15657 15423 15665
rect 16651 15645 16685 15685
rect 16704 15665 16713 15693
rect 17095 15665 17104 15693
rect 16691 15657 16713 15665
rect 17123 15645 17157 15685
rect 17176 15665 17185 15693
rect 17677 15665 17686 15693
rect 17163 15657 17185 15665
rect 17705 15645 17739 15685
rect 17758 15665 17767 15693
rect 18149 15665 18158 15693
rect 17745 15657 17767 15665
rect 18177 15645 18211 15685
rect 18230 15665 18239 15693
rect 18621 15665 18630 15693
rect 18217 15657 18239 15665
rect 18649 15645 18683 15685
rect 18702 15665 18711 15693
rect 19093 15665 19102 15693
rect 18689 15657 18711 15665
rect 19121 15645 19155 15685
rect 19174 15665 19183 15693
rect 21753 15672 21761 16216
rect 19161 15657 19183 15665
rect 21737 15664 21761 15672
rect 21779 16216 21803 16224
rect 21855 16224 21921 16232
rect 21855 16216 21879 16224
rect 21779 15672 21787 16216
rect 21871 15672 21879 16216
rect 21779 15664 21803 15672
rect 21737 15656 21803 15664
rect 21855 15664 21879 15672
rect 21897 16216 21921 16224
rect 21973 16224 22039 16232
rect 21973 16216 21997 16224
rect 21897 15672 21905 16216
rect 21989 15672 21997 16216
rect 21897 15664 21921 15672
rect 21855 15656 21921 15664
rect 21973 15664 21997 15672
rect 22015 16216 22039 16224
rect 22091 16224 22157 16232
rect 22091 16216 22115 16224
rect 22015 15672 22023 16216
rect 22107 15672 22115 16216
rect 22015 15664 22039 15672
rect 21973 15656 22039 15664
rect 22091 15664 22115 15672
rect 22133 16216 22157 16224
rect 22209 16224 22275 16232
rect 22209 16216 22233 16224
rect 22133 15672 22141 16216
rect 22225 15672 22233 16216
rect 22133 15664 22157 15672
rect 22091 15656 22157 15664
rect 22209 15664 22233 15672
rect 22251 16216 22275 16224
rect 22327 16224 22393 16232
rect 22327 16216 22351 16224
rect 22251 15672 22259 16216
rect 22343 15672 22351 16216
rect 22251 15664 22275 15672
rect 22209 15656 22275 15664
rect 22327 15664 22351 15672
rect 22369 16216 22393 16224
rect 22445 16224 22511 16232
rect 22445 16216 22469 16224
rect 22369 15672 22377 16216
rect 22461 15672 22469 16216
rect 22369 15664 22393 15672
rect 22327 15656 22393 15664
rect 22445 15664 22469 15672
rect 22487 16216 22511 16224
rect 22563 16224 22629 16232
rect 22563 16216 22587 16224
rect 22487 15672 22495 16216
rect 22579 15672 22587 16216
rect 22487 15664 22511 15672
rect 22445 15656 22511 15664
rect 22563 15664 22587 15672
rect 22605 16216 22629 16224
rect 22681 16224 22747 16232
rect 22681 16216 22705 16224
rect 22605 15672 22613 16216
rect 22697 15672 22705 16216
rect 22605 15664 22629 15672
rect 22563 15656 22629 15664
rect 22681 15664 22705 15672
rect 22723 16216 22747 16224
rect 22799 16224 22865 16232
rect 22799 16216 22823 16224
rect 22723 15672 22731 16216
rect 22815 15672 22823 16216
rect 22723 15664 22747 15672
rect 22681 15656 22747 15664
rect 22799 15664 22823 15672
rect 22841 16216 22865 16224
rect 22917 16224 22983 16232
rect 22917 16216 22941 16224
rect 22841 15672 22849 16216
rect 22933 15672 22941 16216
rect 22841 15664 22865 15672
rect 22799 15656 22865 15664
rect 22917 15664 22941 15672
rect 22959 16216 22983 16224
rect 23035 16224 23101 16232
rect 23035 16216 23059 16224
rect 22959 15672 22967 16216
rect 23051 15672 23059 16216
rect 22959 15664 22983 15672
rect 22917 15656 22983 15664
rect 23035 15664 23059 15672
rect 23077 16216 23101 16224
rect 23153 16224 23219 16232
rect 23153 16216 23177 16224
rect 23077 15672 23085 16216
rect 23169 15672 23177 16216
rect 23077 15664 23101 15672
rect 23035 15656 23101 15664
rect 23153 15664 23177 15672
rect 23195 16216 23219 16224
rect 23271 16224 23337 16232
rect 23271 16216 23295 16224
rect 23195 15672 23203 16216
rect 23287 15672 23295 16216
rect 23195 15664 23219 15672
rect 23153 15656 23219 15664
rect 23271 15664 23295 15672
rect 23313 16216 23337 16224
rect 23389 16224 23455 16232
rect 23389 16216 23413 16224
rect 23313 15672 23321 16216
rect 23405 15672 23413 16216
rect 23313 15664 23337 15672
rect 23271 15656 23337 15664
rect 23389 15664 23413 15672
rect 23431 16216 23455 16224
rect 23507 16224 23573 16232
rect 23507 16216 23531 16224
rect 23431 15672 23439 16216
rect 23523 15672 23531 16216
rect 23431 15664 23455 15672
rect 23389 15656 23455 15664
rect 23507 15664 23531 15672
rect 23549 16216 23573 16224
rect 23625 16224 23691 16232
rect 23625 16216 23649 16224
rect 23549 15672 23557 16216
rect 23641 15672 23649 16216
rect 23549 15664 23573 15672
rect 23507 15656 23573 15664
rect 23625 15664 23649 15672
rect 23667 16216 23691 16224
rect 23743 16224 23809 16232
rect 23743 16216 23767 16224
rect 23667 15672 23675 16216
rect 23759 15672 23767 16216
rect 23667 15664 23691 15672
rect 23625 15656 23691 15664
rect 23743 15664 23767 15672
rect 23785 16216 23809 16224
rect 23861 16224 23927 16232
rect 23861 16216 23885 16224
rect 23785 15672 23793 16216
rect 23877 15672 23885 16216
rect 23785 15664 23809 15672
rect 23743 15656 23809 15664
rect 23861 15664 23885 15672
rect 23903 16216 23927 16224
rect 23979 16224 24045 16232
rect 23979 16216 24003 16224
rect 23903 15672 23911 16216
rect 23995 15672 24003 16216
rect 23903 15664 23927 15672
rect 23861 15656 23927 15664
rect 23979 15664 24003 15672
rect 24021 16216 24045 16224
rect 24097 16224 24163 16232
rect 24097 16216 24121 16224
rect 24021 15672 24029 16216
rect 24113 15672 24121 16216
rect 24021 15664 24045 15672
rect 23979 15656 24045 15664
rect 24097 15664 24121 15672
rect 24139 16216 24163 16224
rect 24215 16224 24281 16232
rect 24215 16216 24239 16224
rect 24139 15672 24147 16216
rect 24231 15672 24239 16216
rect 24139 15664 24163 15672
rect 24097 15656 24163 15664
rect 24215 15664 24239 15672
rect 24257 16216 24281 16224
rect 25860 16224 25926 16232
rect 25860 16216 25884 16224
rect 24257 15672 24265 16216
rect 25876 15672 25884 16216
rect 24257 15664 24281 15672
rect 24215 15656 24281 15664
rect 25860 15664 25884 15672
rect 25902 16216 25926 16224
rect 25978 16224 26044 16232
rect 25978 16216 26002 16224
rect 25902 15672 25910 16216
rect 25994 15672 26002 16216
rect 25902 15664 25926 15672
rect 25860 15656 25926 15664
rect 25978 15664 26002 15672
rect 26020 16216 26044 16224
rect 26096 16224 26162 16232
rect 26096 16216 26120 16224
rect 26020 15672 26028 16216
rect 26112 15672 26120 16216
rect 26020 15664 26044 15672
rect 25978 15656 26044 15664
rect 26096 15664 26120 15672
rect 26138 16216 26162 16224
rect 26214 16224 26280 16232
rect 26214 16216 26238 16224
rect 26138 15672 26146 16216
rect 26230 15672 26238 16216
rect 26138 15664 26162 15672
rect 26096 15656 26162 15664
rect 26214 15664 26238 15672
rect 26256 16216 26280 16224
rect 26332 16224 26398 16232
rect 26332 16216 26356 16224
rect 26256 15672 26264 16216
rect 26348 15672 26356 16216
rect 26256 15664 26280 15672
rect 26214 15656 26280 15664
rect 26332 15664 26356 15672
rect 26374 16216 26398 16224
rect 26450 16224 26516 16232
rect 26450 16216 26474 16224
rect 26374 15672 26382 16216
rect 26466 15672 26474 16216
rect 26374 15664 26398 15672
rect 26332 15656 26398 15664
rect 26450 15664 26474 15672
rect 26492 16216 26516 16224
rect 26568 16224 26634 16232
rect 26568 16216 26592 16224
rect 26492 15672 26500 16216
rect 26584 15672 26592 16216
rect 26492 15664 26516 15672
rect 26450 15656 26516 15664
rect 26568 15664 26592 15672
rect 26610 16216 26634 16224
rect 26686 16224 26752 16232
rect 26686 16216 26710 16224
rect 26610 15672 26618 16216
rect 26702 15672 26710 16216
rect 26610 15664 26634 15672
rect 26568 15656 26634 15664
rect 26686 15664 26710 15672
rect 26728 16216 26752 16224
rect 26804 16224 26870 16232
rect 26804 16216 26828 16224
rect 26728 15672 26736 16216
rect 26820 15672 26828 16216
rect 26728 15664 26752 15672
rect 26686 15656 26752 15664
rect 26804 15664 26828 15672
rect 26846 16216 26870 16224
rect 26922 16224 26988 16232
rect 26922 16216 26946 16224
rect 26846 15672 26854 16216
rect 26938 15672 26946 16216
rect 26846 15664 26870 15672
rect 26804 15656 26870 15664
rect 26922 15664 26946 15672
rect 26964 16216 26988 16224
rect 27040 16224 27106 16232
rect 27040 16216 27064 16224
rect 26964 15672 26972 16216
rect 27056 15672 27064 16216
rect 26964 15664 26988 15672
rect 26922 15656 26988 15664
rect 27040 15664 27064 15672
rect 27082 16216 27106 16224
rect 27158 16224 27224 16232
rect 27158 16216 27182 16224
rect 27082 15672 27090 16216
rect 27174 15672 27182 16216
rect 27082 15664 27106 15672
rect 27040 15656 27106 15664
rect 27158 15664 27182 15672
rect 27200 16216 27224 16224
rect 27276 16224 27342 16232
rect 27276 16216 27300 16224
rect 27200 15672 27208 16216
rect 27292 15672 27300 16216
rect 27200 15664 27224 15672
rect 27158 15656 27224 15664
rect 27276 15664 27300 15672
rect 27318 16216 27342 16224
rect 27394 16224 27460 16232
rect 27394 16216 27418 16224
rect 27318 15672 27326 16216
rect 27410 15672 27418 16216
rect 27318 15664 27342 15672
rect 27276 15656 27342 15664
rect 27394 15664 27418 15672
rect 27436 16216 27460 16224
rect 27512 16224 27578 16232
rect 27512 16216 27536 16224
rect 27436 15672 27444 16216
rect 27528 15672 27536 16216
rect 27436 15664 27460 15672
rect 27394 15656 27460 15664
rect 27512 15664 27536 15672
rect 27554 16216 27578 16224
rect 27630 16224 27696 16232
rect 27630 16216 27654 16224
rect 27554 15672 27562 16216
rect 27646 15672 27654 16216
rect 27554 15664 27578 15672
rect 27512 15656 27578 15664
rect 27630 15664 27654 15672
rect 27672 16216 27696 16224
rect 27748 16224 27814 16232
rect 27748 16216 27772 16224
rect 27672 15672 27680 16216
rect 27764 15672 27772 16216
rect 27672 15664 27696 15672
rect 27630 15656 27696 15664
rect 27748 15664 27772 15672
rect 27790 16216 27814 16224
rect 27866 16224 27932 16232
rect 27866 16216 27890 16224
rect 27790 15672 27798 16216
rect 27882 15672 27890 16216
rect 27790 15664 27814 15672
rect 27748 15656 27814 15664
rect 27866 15664 27890 15672
rect 27908 16216 27932 16224
rect 27984 16224 28050 16232
rect 27984 16216 28008 16224
rect 27908 15672 27916 16216
rect 28000 15672 28008 16216
rect 27908 15664 27932 15672
rect 27866 15656 27932 15664
rect 27984 15664 28008 15672
rect 28026 16216 28050 16224
rect 28102 16224 28168 16232
rect 28102 16216 28126 16224
rect 28026 15672 28034 16216
rect 28118 15672 28126 16216
rect 28026 15664 28050 15672
rect 27984 15656 28050 15664
rect 28102 15664 28126 15672
rect 28144 16216 28168 16224
rect 28220 16224 28286 16232
rect 28220 16216 28244 16224
rect 28144 15672 28152 16216
rect 28236 15672 28244 16216
rect 28144 15664 28168 15672
rect 28102 15656 28168 15664
rect 28220 15664 28244 15672
rect 28262 16216 28286 16224
rect 28338 16224 28404 16232
rect 28338 16216 28362 16224
rect 28262 15672 28270 16216
rect 28354 15672 28362 16216
rect 28262 15664 28286 15672
rect 28220 15656 28286 15664
rect 28338 15664 28362 15672
rect 28380 16216 28404 16224
rect 29983 16224 30049 16232
rect 29983 16216 30007 16224
rect 28380 15672 28388 16216
rect 29999 15672 30007 16216
rect 28380 15664 28404 15672
rect 28338 15656 28404 15664
rect 29983 15664 30007 15672
rect 30025 16216 30049 16224
rect 30101 16224 30167 16232
rect 30101 16216 30125 16224
rect 30025 15672 30033 16216
rect 30117 15672 30125 16216
rect 30025 15664 30049 15672
rect 29983 15656 30049 15664
rect 30101 15664 30125 15672
rect 30143 16216 30167 16224
rect 30219 16224 30285 16232
rect 30219 16216 30243 16224
rect 30143 15672 30151 16216
rect 30235 15672 30243 16216
rect 30143 15664 30167 15672
rect 30101 15656 30167 15664
rect 30219 15664 30243 15672
rect 30261 16216 30285 16224
rect 30337 16224 30403 16232
rect 30337 16216 30361 16224
rect 30261 15672 30269 16216
rect 30353 15672 30361 16216
rect 30261 15664 30285 15672
rect 30219 15656 30285 15664
rect 30337 15664 30361 15672
rect 30379 16216 30403 16224
rect 30455 16224 30521 16232
rect 30455 16216 30479 16224
rect 30379 15672 30387 16216
rect 30471 15672 30479 16216
rect 30379 15664 30403 15672
rect 30337 15656 30403 15664
rect 30455 15664 30479 15672
rect 30497 16216 30521 16224
rect 30573 16224 30639 16232
rect 30573 16216 30597 16224
rect 30497 15672 30505 16216
rect 30589 15672 30597 16216
rect 30497 15664 30521 15672
rect 30455 15656 30521 15664
rect 30573 15664 30597 15672
rect 30615 16216 30639 16224
rect 30691 16224 30757 16232
rect 30691 16216 30715 16224
rect 30615 15672 30623 16216
rect 30707 15672 30715 16216
rect 30615 15664 30639 15672
rect 30573 15656 30639 15664
rect 30691 15664 30715 15672
rect 30733 16216 30757 16224
rect 30809 16224 30875 16232
rect 30809 16216 30833 16224
rect 30733 15672 30741 16216
rect 30825 15672 30833 16216
rect 30733 15664 30757 15672
rect 30691 15656 30757 15664
rect 30809 15664 30833 15672
rect 30851 16216 30875 16224
rect 30927 16224 30993 16232
rect 30927 16216 30951 16224
rect 30851 15672 30859 16216
rect 30943 15672 30951 16216
rect 30851 15664 30875 15672
rect 30809 15656 30875 15664
rect 30927 15664 30951 15672
rect 30969 16216 30993 16224
rect 31045 16224 31111 16232
rect 31045 16216 31069 16224
rect 30969 15672 30977 16216
rect 31061 15672 31069 16216
rect 30969 15664 30993 15672
rect 30927 15656 30993 15664
rect 31045 15664 31069 15672
rect 31087 16216 31111 16224
rect 31163 16224 31229 16232
rect 31163 16216 31187 16224
rect 31087 15672 31095 16216
rect 31179 15672 31187 16216
rect 31087 15664 31111 15672
rect 31045 15656 31111 15664
rect 31163 15664 31187 15672
rect 31205 16216 31229 16224
rect 31281 16224 31347 16232
rect 31281 16216 31305 16224
rect 31205 15672 31213 16216
rect 31297 15672 31305 16216
rect 31205 15664 31229 15672
rect 31163 15656 31229 15664
rect 31281 15664 31305 15672
rect 31323 16216 31347 16224
rect 31399 16224 31465 16232
rect 31399 16216 31423 16224
rect 31323 15672 31331 16216
rect 31415 15672 31423 16216
rect 31323 15664 31347 15672
rect 31281 15656 31347 15664
rect 31399 15664 31423 15672
rect 31441 16216 31465 16224
rect 31517 16224 31583 16232
rect 31517 16216 31541 16224
rect 31441 15672 31449 16216
rect 31533 15672 31541 16216
rect 31441 15664 31465 15672
rect 31399 15656 31465 15664
rect 31517 15664 31541 15672
rect 31559 16216 31583 16224
rect 31635 16224 31701 16232
rect 31635 16216 31659 16224
rect 31559 15672 31567 16216
rect 31651 15672 31659 16216
rect 31559 15664 31583 15672
rect 31517 15656 31583 15664
rect 31635 15664 31659 15672
rect 31677 16216 31701 16224
rect 31753 16224 31819 16232
rect 31753 16216 31777 16224
rect 31677 15672 31685 16216
rect 31769 15672 31777 16216
rect 31677 15664 31701 15672
rect 31635 15656 31701 15664
rect 31753 15664 31777 15672
rect 31795 16216 31819 16224
rect 31871 16224 31937 16232
rect 31871 16216 31895 16224
rect 31795 15672 31803 16216
rect 31887 15672 31895 16216
rect 31795 15664 31819 15672
rect 31753 15656 31819 15664
rect 31871 15664 31895 15672
rect 31913 16216 31937 16224
rect 31989 16224 32055 16232
rect 31989 16216 32013 16224
rect 31913 15672 31921 16216
rect 32005 15672 32013 16216
rect 31913 15664 31937 15672
rect 31871 15656 31937 15664
rect 31989 15664 32013 15672
rect 32031 16216 32055 16224
rect 32107 16224 32173 16232
rect 32107 16216 32131 16224
rect 32031 15672 32039 16216
rect 32123 15672 32131 16216
rect 32031 15664 32055 15672
rect 31989 15656 32055 15664
rect 32107 15664 32131 15672
rect 32149 16216 32173 16224
rect 32225 16224 32291 16232
rect 32225 16216 32249 16224
rect 32149 15672 32157 16216
rect 32241 15672 32249 16216
rect 32149 15664 32173 15672
rect 32107 15656 32173 15664
rect 32225 15664 32249 15672
rect 32267 16216 32291 16224
rect 32343 16224 32409 16232
rect 32343 16216 32367 16224
rect 32267 15672 32275 16216
rect 32359 15672 32367 16216
rect 32267 15664 32291 15672
rect 32225 15656 32291 15664
rect 32343 15664 32367 15672
rect 32385 16216 32409 16224
rect 32461 16224 32527 16232
rect 32461 16216 32485 16224
rect 32385 15672 32393 16216
rect 32477 15672 32485 16216
rect 32385 15664 32409 15672
rect 32343 15656 32409 15664
rect 32461 15664 32485 15672
rect 32503 16216 32527 16224
rect 32503 15672 32511 16216
rect 32503 15664 32527 15672
rect 32461 15656 32527 15664
rect 21753 15640 21769 15656
rect 21771 15640 21787 15656
rect 21871 15640 21887 15656
rect 21889 15640 21905 15656
rect 21989 15640 22005 15656
rect 22007 15640 22023 15656
rect 22107 15640 22123 15656
rect 22125 15640 22141 15656
rect 22225 15640 22241 15656
rect 22243 15640 22259 15656
rect 22343 15640 22359 15656
rect 22361 15640 22377 15656
rect 22461 15640 22477 15656
rect 22479 15640 22495 15656
rect 22579 15640 22595 15656
rect 22597 15640 22613 15656
rect 22697 15640 22713 15656
rect 22715 15640 22731 15656
rect 22815 15640 22831 15656
rect 22833 15640 22849 15656
rect 22933 15640 22949 15656
rect 22951 15640 22967 15656
rect 23051 15640 23067 15656
rect 23069 15640 23085 15656
rect 23169 15640 23185 15656
rect 23187 15640 23203 15656
rect 23287 15640 23303 15656
rect 23305 15640 23321 15656
rect 23405 15640 23421 15656
rect 23423 15640 23439 15656
rect 23523 15640 23539 15656
rect 23541 15640 23557 15656
rect 23641 15640 23657 15656
rect 23659 15640 23675 15656
rect 23759 15640 23775 15656
rect 23777 15640 23793 15656
rect 23877 15640 23893 15656
rect 23895 15640 23911 15656
rect 23995 15640 24011 15656
rect 24013 15640 24029 15656
rect 24113 15640 24129 15656
rect 24131 15640 24147 15656
rect 24231 15640 24247 15656
rect 24249 15640 24265 15656
rect 25876 15640 25892 15656
rect 25894 15640 25910 15656
rect 25994 15640 26010 15656
rect 26012 15640 26028 15656
rect 26112 15640 26128 15656
rect 26130 15640 26146 15656
rect 26230 15640 26246 15656
rect 26248 15640 26264 15656
rect 26348 15640 26364 15656
rect 26366 15640 26382 15656
rect 26466 15640 26482 15656
rect 26484 15640 26500 15656
rect 26584 15640 26600 15656
rect 26602 15640 26618 15656
rect 26702 15640 26718 15656
rect 26720 15640 26736 15656
rect 26820 15640 26836 15656
rect 26838 15640 26854 15656
rect 26938 15640 26954 15656
rect 26956 15640 26972 15656
rect 27056 15640 27072 15656
rect 27074 15640 27090 15656
rect 27174 15640 27190 15656
rect 27192 15640 27208 15656
rect 27292 15640 27308 15656
rect 27310 15640 27326 15656
rect 27410 15640 27426 15656
rect 27428 15640 27444 15656
rect 27528 15640 27544 15656
rect 27546 15640 27562 15656
rect 27646 15640 27662 15656
rect 27664 15640 27680 15656
rect 27764 15640 27780 15656
rect 27782 15640 27798 15656
rect 27882 15640 27898 15656
rect 27900 15640 27916 15656
rect 28000 15640 28016 15656
rect 28018 15640 28034 15656
rect 28118 15640 28134 15656
rect 28136 15640 28152 15656
rect 28236 15640 28252 15656
rect 28254 15640 28270 15656
rect 28354 15640 28370 15656
rect 28372 15640 28388 15656
rect 29999 15640 30015 15656
rect 30017 15640 30033 15656
rect 30117 15640 30133 15656
rect 30135 15640 30151 15656
rect 30235 15640 30251 15656
rect 30253 15640 30269 15656
rect 30353 15640 30369 15656
rect 30371 15640 30387 15656
rect 30471 15640 30487 15656
rect 30489 15640 30505 15656
rect 30589 15640 30605 15656
rect 30607 15640 30623 15656
rect 30707 15640 30723 15656
rect 30725 15640 30741 15656
rect 30825 15640 30841 15656
rect 30843 15640 30859 15656
rect 30943 15640 30959 15656
rect 30961 15640 30977 15656
rect 31061 15640 31077 15656
rect 31079 15640 31095 15656
rect 31179 15640 31195 15656
rect 31197 15640 31213 15656
rect 31297 15640 31313 15656
rect 31315 15640 31331 15656
rect 31415 15640 31431 15656
rect 31433 15640 31449 15656
rect 31533 15640 31549 15656
rect 31551 15640 31567 15656
rect 31651 15640 31667 15656
rect 31669 15640 31685 15656
rect 31769 15640 31785 15656
rect 31787 15640 31803 15656
rect 31887 15640 31903 15656
rect 31905 15640 31921 15656
rect 32005 15640 32021 15656
rect 32023 15640 32039 15656
rect 32123 15640 32139 15656
rect 32141 15640 32157 15656
rect 32241 15640 32257 15656
rect 32259 15640 32275 15656
rect 32359 15640 32375 15656
rect 32377 15640 32393 15656
rect 32477 15640 32493 15656
rect 32495 15640 32511 15656
rect 13650 15564 13684 15598
rect 13768 15564 13802 15598
rect 13886 15564 13920 15598
rect 14004 15564 14038 15598
rect 14122 15564 14156 15598
rect 14240 15564 14274 15598
rect 14358 15564 14392 15598
rect 14476 15564 14510 15598
rect 14594 15564 14628 15598
rect 14712 15564 14746 15598
rect 14830 15564 14864 15598
rect 14948 15564 14982 15598
rect 15066 15564 15100 15598
rect 15184 15564 15218 15598
rect 15302 15564 15336 15598
rect 15884 15564 15918 15598
rect 16002 15564 16036 15598
rect 16120 15564 16154 15598
rect 16238 15564 16272 15598
rect 16356 15564 16390 15598
rect 16474 15564 16508 15598
rect 21458 15597 21474 15613
rect 21476 15597 21492 15613
rect 25581 15597 25597 15613
rect 25599 15597 25615 15613
rect 29704 15597 29720 15613
rect 29722 15597 29738 15613
rect 21442 15593 21492 15597
rect 21442 15581 21458 15593
rect 21504 15581 21508 15597
rect 25565 15593 25615 15597
rect 25565 15581 25581 15593
rect 25627 15581 25631 15597
rect 29688 15593 29738 15597
rect 29688 15581 29704 15593
rect 29750 15581 29754 15597
rect 21446 15579 21458 15581
rect 25569 15579 25581 15581
rect 29692 15579 29704 15581
rect 21442 15563 21458 15579
rect 21504 15563 21508 15579
rect 25565 15563 25581 15579
rect 25627 15563 25631 15579
rect 29688 15563 29704 15579
rect 29750 15563 29754 15579
rect 21458 15547 21474 15563
rect 21476 15547 21492 15563
rect 25581 15547 25597 15563
rect 25599 15547 25615 15563
rect 29704 15547 29720 15563
rect 29722 15547 29738 15563
rect 21458 15489 21474 15505
rect 21476 15489 21492 15505
rect 25581 15489 25597 15505
rect 25599 15489 25615 15505
rect 29704 15489 29720 15505
rect 29722 15489 29738 15505
rect 21442 15473 21458 15489
rect 21504 15473 21508 15489
rect 25565 15473 25581 15489
rect 25627 15473 25631 15489
rect 29688 15473 29704 15489
rect 29750 15473 29754 15489
rect 21446 15471 21458 15473
rect 25569 15471 25581 15473
rect 29692 15471 29704 15473
rect 21442 15459 21458 15471
rect 21442 15455 21492 15459
rect 21504 15455 21508 15471
rect 25565 15459 25581 15471
rect 25565 15455 25615 15459
rect 25627 15455 25631 15471
rect 29688 15459 29704 15471
rect 29688 15455 29738 15459
rect 29750 15455 29754 15471
rect 21458 15439 21474 15455
rect 21476 15439 21492 15455
rect 25581 15439 25597 15455
rect 25599 15439 25615 15455
rect 29704 15439 29720 15455
rect 29722 15439 29738 15455
rect 21753 15396 21769 15412
rect 21771 15396 21787 15412
rect 21871 15396 21887 15412
rect 21889 15396 21905 15412
rect 21989 15396 22005 15412
rect 22007 15396 22023 15412
rect 22107 15396 22123 15412
rect 22125 15396 22141 15412
rect 22225 15396 22241 15412
rect 22243 15396 22259 15412
rect 22343 15396 22359 15412
rect 22361 15396 22377 15412
rect 22461 15396 22477 15412
rect 22479 15396 22495 15412
rect 22579 15396 22595 15412
rect 22597 15396 22613 15412
rect 22697 15396 22713 15412
rect 22715 15396 22731 15412
rect 22815 15396 22831 15412
rect 22833 15396 22849 15412
rect 22933 15396 22949 15412
rect 22951 15396 22967 15412
rect 23051 15396 23067 15412
rect 23069 15396 23085 15412
rect 23169 15396 23185 15412
rect 23187 15396 23203 15412
rect 23287 15396 23303 15412
rect 23305 15396 23321 15412
rect 23405 15396 23421 15412
rect 23423 15396 23439 15412
rect 23523 15396 23539 15412
rect 23541 15396 23557 15412
rect 23641 15396 23657 15412
rect 23659 15396 23675 15412
rect 23759 15396 23775 15412
rect 23777 15396 23793 15412
rect 23877 15396 23893 15412
rect 23895 15396 23911 15412
rect 23995 15396 24011 15412
rect 24013 15396 24029 15412
rect 24113 15396 24129 15412
rect 24131 15396 24147 15412
rect 24231 15396 24247 15412
rect 24249 15396 24265 15412
rect 25876 15396 25892 15412
rect 25894 15396 25910 15412
rect 25994 15396 26010 15412
rect 26012 15396 26028 15412
rect 26112 15396 26128 15412
rect 26130 15396 26146 15412
rect 26230 15396 26246 15412
rect 26248 15396 26264 15412
rect 26348 15396 26364 15412
rect 26366 15396 26382 15412
rect 26466 15396 26482 15412
rect 26484 15396 26500 15412
rect 26584 15396 26600 15412
rect 26602 15396 26618 15412
rect 26702 15396 26718 15412
rect 26720 15396 26736 15412
rect 26820 15396 26836 15412
rect 26838 15396 26854 15412
rect 26938 15396 26954 15412
rect 26956 15396 26972 15412
rect 27056 15396 27072 15412
rect 27074 15396 27090 15412
rect 27174 15396 27190 15412
rect 27192 15396 27208 15412
rect 27292 15396 27308 15412
rect 27310 15396 27326 15412
rect 27410 15396 27426 15412
rect 27428 15396 27444 15412
rect 27528 15396 27544 15412
rect 27546 15396 27562 15412
rect 27646 15396 27662 15412
rect 27664 15396 27680 15412
rect 27764 15396 27780 15412
rect 27782 15396 27798 15412
rect 27882 15396 27898 15412
rect 27900 15396 27916 15412
rect 28000 15396 28016 15412
rect 28018 15396 28034 15412
rect 28118 15396 28134 15412
rect 28136 15396 28152 15412
rect 28236 15396 28252 15412
rect 28254 15396 28270 15412
rect 28354 15396 28370 15412
rect 28372 15396 28388 15412
rect 29999 15396 30015 15412
rect 30017 15396 30033 15412
rect 30117 15396 30133 15412
rect 30135 15396 30151 15412
rect 30235 15396 30251 15412
rect 30253 15396 30269 15412
rect 30353 15396 30369 15412
rect 30371 15396 30387 15412
rect 30471 15396 30487 15412
rect 30489 15396 30505 15412
rect 30589 15396 30605 15412
rect 30607 15396 30623 15412
rect 30707 15396 30723 15412
rect 30725 15396 30741 15412
rect 30825 15396 30841 15412
rect 30843 15396 30859 15412
rect 30943 15396 30959 15412
rect 30961 15396 30977 15412
rect 31061 15396 31077 15412
rect 31079 15396 31095 15412
rect 31179 15396 31195 15412
rect 31197 15396 31213 15412
rect 31297 15396 31313 15412
rect 31315 15396 31331 15412
rect 31415 15396 31431 15412
rect 31433 15396 31449 15412
rect 31533 15396 31549 15412
rect 31551 15396 31567 15412
rect 31651 15396 31667 15412
rect 31669 15396 31685 15412
rect 31769 15396 31785 15412
rect 31787 15396 31803 15412
rect 31887 15396 31903 15412
rect 31905 15396 31921 15412
rect 32005 15396 32021 15412
rect 32023 15396 32039 15412
rect 32123 15396 32139 15412
rect 32141 15396 32157 15412
rect 32241 15396 32257 15412
rect 32259 15396 32275 15412
rect 32359 15396 32375 15412
rect 32377 15396 32393 15412
rect 32477 15396 32493 15412
rect 32495 15396 32511 15412
rect 21737 15388 21803 15396
rect 21737 15380 21761 15388
rect 13387 7120 13392 15328
rect 13415 7120 13420 15328
rect 13475 14849 13479 15156
rect 13503 15021 13507 15128
rect 13554 15053 13575 15128
rect 13582 15127 13588 15133
rect 13628 15127 13634 15133
rect 13818 15127 13824 15133
rect 13864 15127 13870 15133
rect 14054 15127 14060 15133
rect 14100 15127 14106 15133
rect 14290 15127 14296 15133
rect 14336 15127 14342 15133
rect 14526 15127 14532 15133
rect 14572 15127 14578 15133
rect 14762 15127 14768 15133
rect 14808 15127 14814 15133
rect 14998 15127 15004 15133
rect 15044 15127 15050 15133
rect 15234 15127 15240 15133
rect 15280 15127 15286 15133
rect 15470 15127 15476 15133
rect 15516 15127 15522 15133
rect 15706 15127 15712 15133
rect 15752 15127 15758 15133
rect 15942 15127 15948 15133
rect 15988 15127 15994 15133
rect 16178 15127 16184 15133
rect 16224 15127 16230 15133
rect 16414 15127 16420 15133
rect 16460 15127 16466 15133
rect 16650 15127 16656 15133
rect 16696 15127 16702 15133
rect 16886 15127 16892 15133
rect 16932 15127 16938 15133
rect 17122 15127 17128 15133
rect 17168 15127 17174 15133
rect 17358 15127 17364 15133
rect 17404 15127 17410 15133
rect 17594 15127 17600 15133
rect 17640 15127 17646 15133
rect 17830 15127 17836 15133
rect 17876 15127 17882 15133
rect 18066 15127 18072 15133
rect 18112 15127 18118 15133
rect 18302 15127 18308 15133
rect 18348 15127 18354 15133
rect 18538 15127 18544 15133
rect 18584 15127 18590 15133
rect 18774 15127 18780 15133
rect 18820 15127 18826 15133
rect 19010 15127 19016 15133
rect 19056 15127 19062 15133
rect 19246 15127 19252 15133
rect 19292 15127 19298 15133
rect 19482 15127 19488 15133
rect 19528 15127 19534 15133
rect 13576 15121 13603 15127
rect 13634 15121 13640 15127
rect 13812 15121 13818 15127
rect 13870 15121 13876 15127
rect 14048 15121 14054 15127
rect 14106 15121 14112 15127
rect 14284 15121 14290 15127
rect 14342 15121 14348 15127
rect 14520 15121 14526 15127
rect 14578 15121 14584 15127
rect 14756 15121 14762 15127
rect 14814 15121 14820 15127
rect 14992 15121 14998 15127
rect 15050 15121 15056 15127
rect 15228 15121 15234 15127
rect 15286 15121 15292 15127
rect 15464 15121 15470 15127
rect 15522 15121 15528 15127
rect 15700 15121 15706 15127
rect 15758 15121 15764 15127
rect 15936 15121 15942 15127
rect 15994 15121 16000 15127
rect 16172 15121 16178 15127
rect 16230 15121 16236 15127
rect 16408 15121 16414 15127
rect 16466 15121 16472 15127
rect 16644 15121 16650 15127
rect 16702 15121 16708 15127
rect 16880 15121 16886 15127
rect 16938 15121 16944 15127
rect 17116 15121 17122 15127
rect 17174 15121 17180 15127
rect 17352 15121 17358 15127
rect 17410 15121 17416 15127
rect 17588 15121 17594 15127
rect 17646 15121 17652 15127
rect 17824 15121 17830 15127
rect 17882 15121 17888 15127
rect 18060 15121 18066 15127
rect 18118 15121 18124 15127
rect 18296 15121 18302 15127
rect 18354 15121 18360 15127
rect 18532 15121 18538 15127
rect 18590 15121 18596 15127
rect 18768 15121 18774 15127
rect 18826 15121 18832 15127
rect 19004 15121 19010 15127
rect 19062 15121 19068 15127
rect 19240 15121 19246 15127
rect 19298 15121 19304 15127
rect 19476 15121 19482 15127
rect 19534 15121 19540 15127
rect 13582 15053 13603 15121
rect 13491 15019 13533 15021
rect 13503 14877 13507 15019
rect 13812 14877 13818 14883
rect 13870 14877 13876 14883
rect 14048 14877 14054 14883
rect 14106 14877 14112 14883
rect 14284 14877 14290 14883
rect 14342 14877 14348 14883
rect 14520 14877 14526 14883
rect 14578 14877 14584 14883
rect 14756 14877 14762 14883
rect 14814 14877 14820 14883
rect 14992 14877 14998 14883
rect 15050 14877 15056 14883
rect 15228 14877 15234 14883
rect 15286 14877 15292 14883
rect 15464 14877 15470 14883
rect 15522 14877 15528 14883
rect 15700 14877 15706 14883
rect 15758 14877 15764 14883
rect 15936 14877 15942 14883
rect 15994 14877 16000 14883
rect 16172 14877 16178 14883
rect 16230 14877 16236 14883
rect 16408 14877 16414 14883
rect 16466 14877 16472 14883
rect 16644 14877 16650 14883
rect 16702 14877 16708 14883
rect 16880 14877 16886 14883
rect 16938 14877 16944 14883
rect 17116 14877 17122 14883
rect 17174 14877 17180 14883
rect 17352 14877 17358 14883
rect 17410 14877 17416 14883
rect 17588 14877 17594 14883
rect 17646 14877 17652 14883
rect 17824 14877 17830 14883
rect 17882 14877 17888 14883
rect 18060 14877 18066 14883
rect 18118 14877 18124 14883
rect 18296 14877 18302 14883
rect 18354 14877 18360 14883
rect 18532 14877 18538 14883
rect 18590 14877 18596 14883
rect 18768 14877 18774 14883
rect 18826 14877 18832 14883
rect 19004 14877 19010 14883
rect 19062 14877 19068 14883
rect 19240 14877 19246 14883
rect 19298 14877 19304 14883
rect 19476 14877 19482 14883
rect 19534 14877 19540 14883
rect 13818 14871 13824 14877
rect 13864 14871 13870 14877
rect 14054 14871 14060 14877
rect 14100 14871 14106 14877
rect 14290 14871 14296 14877
rect 14336 14871 14342 14877
rect 14526 14871 14532 14877
rect 14572 14871 14578 14877
rect 14762 14871 14768 14877
rect 14808 14871 14814 14877
rect 14998 14871 15004 14877
rect 15044 14871 15050 14877
rect 15234 14871 15240 14877
rect 15280 14871 15286 14877
rect 15470 14871 15476 14877
rect 15516 14871 15522 14877
rect 15706 14871 15712 14877
rect 15752 14871 15758 14877
rect 15942 14871 15948 14877
rect 15988 14871 15994 14877
rect 16178 14871 16184 14877
rect 16224 14871 16230 14877
rect 16414 14871 16420 14877
rect 16460 14871 16466 14877
rect 16650 14871 16656 14877
rect 16696 14871 16702 14877
rect 16886 14871 16892 14877
rect 16932 14871 16938 14877
rect 17122 14871 17128 14877
rect 17168 14871 17174 14877
rect 17358 14871 17364 14877
rect 17404 14871 17410 14877
rect 17594 14871 17600 14877
rect 17640 14871 17646 14877
rect 17830 14871 17836 14877
rect 17876 14871 17882 14877
rect 18066 14871 18072 14877
rect 18112 14871 18118 14877
rect 18302 14871 18308 14877
rect 18348 14871 18354 14877
rect 18538 14871 18544 14877
rect 18584 14871 18590 14877
rect 18774 14871 18780 14877
rect 18820 14871 18826 14877
rect 19010 14871 19016 14877
rect 19056 14871 19062 14877
rect 19246 14871 19252 14877
rect 19292 14871 19298 14877
rect 19482 14871 19488 14877
rect 19528 14871 19534 14877
rect 21753 14836 21761 15380
rect 21737 14828 21761 14836
rect 21779 15380 21803 15388
rect 21855 15388 21921 15396
rect 21855 15380 21879 15388
rect 21779 14836 21787 15380
rect 21871 14836 21879 15380
rect 21779 14828 21803 14836
rect 21737 14820 21803 14828
rect 21855 14828 21879 14836
rect 21897 15380 21921 15388
rect 21973 15388 22039 15396
rect 21973 15380 21997 15388
rect 21897 14836 21905 15380
rect 21989 14836 21997 15380
rect 21897 14828 21921 14836
rect 21855 14820 21921 14828
rect 21973 14828 21997 14836
rect 22015 15380 22039 15388
rect 22091 15388 22157 15396
rect 22091 15380 22115 15388
rect 22015 14836 22023 15380
rect 22107 14836 22115 15380
rect 22015 14828 22039 14836
rect 21973 14820 22039 14828
rect 22091 14828 22115 14836
rect 22133 15380 22157 15388
rect 22209 15388 22275 15396
rect 22209 15380 22233 15388
rect 22133 14836 22141 15380
rect 22225 14836 22233 15380
rect 22133 14828 22157 14836
rect 22091 14820 22157 14828
rect 22209 14828 22233 14836
rect 22251 15380 22275 15388
rect 22327 15388 22393 15396
rect 22327 15380 22351 15388
rect 22251 14836 22259 15380
rect 22343 14836 22351 15380
rect 22251 14828 22275 14836
rect 22209 14820 22275 14828
rect 22327 14828 22351 14836
rect 22369 15380 22393 15388
rect 22445 15388 22511 15396
rect 22445 15380 22469 15388
rect 22369 14836 22377 15380
rect 22461 14836 22469 15380
rect 22369 14828 22393 14836
rect 22327 14820 22393 14828
rect 22445 14828 22469 14836
rect 22487 15380 22511 15388
rect 22563 15388 22629 15396
rect 22563 15380 22587 15388
rect 22487 14836 22495 15380
rect 22579 14836 22587 15380
rect 22487 14828 22511 14836
rect 22445 14820 22511 14828
rect 22563 14828 22587 14836
rect 22605 15380 22629 15388
rect 22681 15388 22747 15396
rect 22681 15380 22705 15388
rect 22605 14836 22613 15380
rect 22697 14836 22705 15380
rect 22605 14828 22629 14836
rect 22563 14820 22629 14828
rect 22681 14828 22705 14836
rect 22723 15380 22747 15388
rect 22799 15388 22865 15396
rect 22799 15380 22823 15388
rect 22723 14836 22731 15380
rect 22815 14836 22823 15380
rect 22723 14828 22747 14836
rect 22681 14820 22747 14828
rect 22799 14828 22823 14836
rect 22841 15380 22865 15388
rect 22917 15388 22983 15396
rect 22917 15380 22941 15388
rect 22841 14836 22849 15380
rect 22933 14836 22941 15380
rect 22841 14828 22865 14836
rect 22799 14820 22865 14828
rect 22917 14828 22941 14836
rect 22959 15380 22983 15388
rect 23035 15388 23101 15396
rect 23035 15380 23059 15388
rect 22959 14836 22967 15380
rect 23051 14836 23059 15380
rect 22959 14828 22983 14836
rect 22917 14820 22983 14828
rect 23035 14828 23059 14836
rect 23077 15380 23101 15388
rect 23153 15388 23219 15396
rect 23153 15380 23177 15388
rect 23077 14836 23085 15380
rect 23169 14836 23177 15380
rect 23077 14828 23101 14836
rect 23035 14820 23101 14828
rect 23153 14828 23177 14836
rect 23195 15380 23219 15388
rect 23271 15388 23337 15396
rect 23271 15380 23295 15388
rect 23195 14836 23203 15380
rect 23287 14836 23295 15380
rect 23195 14828 23219 14836
rect 23153 14820 23219 14828
rect 23271 14828 23295 14836
rect 23313 15380 23337 15388
rect 23389 15388 23455 15396
rect 23389 15380 23413 15388
rect 23313 14836 23321 15380
rect 23405 14836 23413 15380
rect 23313 14828 23337 14836
rect 23271 14820 23337 14828
rect 23389 14828 23413 14836
rect 23431 15380 23455 15388
rect 23507 15388 23573 15396
rect 23507 15380 23531 15388
rect 23431 14836 23439 15380
rect 23523 14836 23531 15380
rect 23431 14828 23455 14836
rect 23389 14820 23455 14828
rect 23507 14828 23531 14836
rect 23549 15380 23573 15388
rect 23625 15388 23691 15396
rect 23625 15380 23649 15388
rect 23549 14836 23557 15380
rect 23641 14836 23649 15380
rect 23549 14828 23573 14836
rect 23507 14820 23573 14828
rect 23625 14828 23649 14836
rect 23667 15380 23691 15388
rect 23743 15388 23809 15396
rect 23743 15380 23767 15388
rect 23667 14836 23675 15380
rect 23759 14836 23767 15380
rect 23667 14828 23691 14836
rect 23625 14820 23691 14828
rect 23743 14828 23767 14836
rect 23785 15380 23809 15388
rect 23861 15388 23927 15396
rect 23861 15380 23885 15388
rect 23785 14836 23793 15380
rect 23877 14836 23885 15380
rect 23785 14828 23809 14836
rect 23743 14820 23809 14828
rect 23861 14828 23885 14836
rect 23903 15380 23927 15388
rect 23979 15388 24045 15396
rect 23979 15380 24003 15388
rect 23903 14836 23911 15380
rect 23995 14836 24003 15380
rect 23903 14828 23927 14836
rect 23861 14820 23927 14828
rect 23979 14828 24003 14836
rect 24021 15380 24045 15388
rect 24097 15388 24163 15396
rect 24097 15380 24121 15388
rect 24021 14836 24029 15380
rect 24113 14836 24121 15380
rect 24021 14828 24045 14836
rect 23979 14820 24045 14828
rect 24097 14828 24121 14836
rect 24139 15380 24163 15388
rect 24215 15388 24281 15396
rect 24215 15380 24239 15388
rect 24139 14836 24147 15380
rect 24231 14836 24239 15380
rect 24139 14828 24163 14836
rect 24097 14820 24163 14828
rect 24215 14828 24239 14836
rect 24257 15380 24281 15388
rect 25860 15388 25926 15396
rect 25860 15380 25884 15388
rect 24257 14836 24265 15380
rect 25876 14836 25884 15380
rect 24257 14828 24281 14836
rect 24215 14820 24281 14828
rect 25860 14828 25884 14836
rect 25902 15380 25926 15388
rect 25978 15388 26044 15396
rect 25978 15380 26002 15388
rect 25902 14836 25910 15380
rect 25994 14836 26002 15380
rect 25902 14828 25926 14836
rect 25860 14820 25926 14828
rect 25978 14828 26002 14836
rect 26020 15380 26044 15388
rect 26096 15388 26162 15396
rect 26096 15380 26120 15388
rect 26020 14836 26028 15380
rect 26112 14836 26120 15380
rect 26020 14828 26044 14836
rect 25978 14820 26044 14828
rect 26096 14828 26120 14836
rect 26138 15380 26162 15388
rect 26214 15388 26280 15396
rect 26214 15380 26238 15388
rect 26138 14836 26146 15380
rect 26230 14836 26238 15380
rect 26138 14828 26162 14836
rect 26096 14820 26162 14828
rect 26214 14828 26238 14836
rect 26256 15380 26280 15388
rect 26332 15388 26398 15396
rect 26332 15380 26356 15388
rect 26256 14836 26264 15380
rect 26348 14836 26356 15380
rect 26256 14828 26280 14836
rect 26214 14820 26280 14828
rect 26332 14828 26356 14836
rect 26374 15380 26398 15388
rect 26450 15388 26516 15396
rect 26450 15380 26474 15388
rect 26374 14836 26382 15380
rect 26466 14836 26474 15380
rect 26374 14828 26398 14836
rect 26332 14820 26398 14828
rect 26450 14828 26474 14836
rect 26492 15380 26516 15388
rect 26568 15388 26634 15396
rect 26568 15380 26592 15388
rect 26492 14836 26500 15380
rect 26584 14836 26592 15380
rect 26492 14828 26516 14836
rect 26450 14820 26516 14828
rect 26568 14828 26592 14836
rect 26610 15380 26634 15388
rect 26686 15388 26752 15396
rect 26686 15380 26710 15388
rect 26610 14836 26618 15380
rect 26702 14836 26710 15380
rect 26610 14828 26634 14836
rect 26568 14820 26634 14828
rect 26686 14828 26710 14836
rect 26728 15380 26752 15388
rect 26804 15388 26870 15396
rect 26804 15380 26828 15388
rect 26728 14836 26736 15380
rect 26820 14836 26828 15380
rect 26728 14828 26752 14836
rect 26686 14820 26752 14828
rect 26804 14828 26828 14836
rect 26846 15380 26870 15388
rect 26922 15388 26988 15396
rect 26922 15380 26946 15388
rect 26846 14836 26854 15380
rect 26938 14836 26946 15380
rect 26846 14828 26870 14836
rect 26804 14820 26870 14828
rect 26922 14828 26946 14836
rect 26964 15380 26988 15388
rect 27040 15388 27106 15396
rect 27040 15380 27064 15388
rect 26964 14836 26972 15380
rect 27056 14836 27064 15380
rect 26964 14828 26988 14836
rect 26922 14820 26988 14828
rect 27040 14828 27064 14836
rect 27082 15380 27106 15388
rect 27158 15388 27224 15396
rect 27158 15380 27182 15388
rect 27082 14836 27090 15380
rect 27174 14836 27182 15380
rect 27082 14828 27106 14836
rect 27040 14820 27106 14828
rect 27158 14828 27182 14836
rect 27200 15380 27224 15388
rect 27276 15388 27342 15396
rect 27276 15380 27300 15388
rect 27200 14836 27208 15380
rect 27292 14836 27300 15380
rect 27200 14828 27224 14836
rect 27158 14820 27224 14828
rect 27276 14828 27300 14836
rect 27318 15380 27342 15388
rect 27394 15388 27460 15396
rect 27394 15380 27418 15388
rect 27318 14836 27326 15380
rect 27410 14836 27418 15380
rect 27318 14828 27342 14836
rect 27276 14820 27342 14828
rect 27394 14828 27418 14836
rect 27436 15380 27460 15388
rect 27512 15388 27578 15396
rect 27512 15380 27536 15388
rect 27436 14836 27444 15380
rect 27528 14836 27536 15380
rect 27436 14828 27460 14836
rect 27394 14820 27460 14828
rect 27512 14828 27536 14836
rect 27554 15380 27578 15388
rect 27630 15388 27696 15396
rect 27630 15380 27654 15388
rect 27554 14836 27562 15380
rect 27646 14836 27654 15380
rect 27554 14828 27578 14836
rect 27512 14820 27578 14828
rect 27630 14828 27654 14836
rect 27672 15380 27696 15388
rect 27748 15388 27814 15396
rect 27748 15380 27772 15388
rect 27672 14836 27680 15380
rect 27764 14836 27772 15380
rect 27672 14828 27696 14836
rect 27630 14820 27696 14828
rect 27748 14828 27772 14836
rect 27790 15380 27814 15388
rect 27866 15388 27932 15396
rect 27866 15380 27890 15388
rect 27790 14836 27798 15380
rect 27882 14836 27890 15380
rect 27790 14828 27814 14836
rect 27748 14820 27814 14828
rect 27866 14828 27890 14836
rect 27908 15380 27932 15388
rect 27984 15388 28050 15396
rect 27984 15380 28008 15388
rect 27908 14836 27916 15380
rect 28000 14836 28008 15380
rect 27908 14828 27932 14836
rect 27866 14820 27932 14828
rect 27984 14828 28008 14836
rect 28026 15380 28050 15388
rect 28102 15388 28168 15396
rect 28102 15380 28126 15388
rect 28026 14836 28034 15380
rect 28118 14836 28126 15380
rect 28026 14828 28050 14836
rect 27984 14820 28050 14828
rect 28102 14828 28126 14836
rect 28144 15380 28168 15388
rect 28220 15388 28286 15396
rect 28220 15380 28244 15388
rect 28144 14836 28152 15380
rect 28236 14836 28244 15380
rect 28144 14828 28168 14836
rect 28102 14820 28168 14828
rect 28220 14828 28244 14836
rect 28262 15380 28286 15388
rect 28338 15388 28404 15396
rect 28338 15380 28362 15388
rect 28262 14836 28270 15380
rect 28354 14836 28362 15380
rect 28262 14828 28286 14836
rect 28220 14820 28286 14828
rect 28338 14828 28362 14836
rect 28380 15380 28404 15388
rect 29983 15388 30049 15396
rect 29983 15380 30007 15388
rect 28380 14836 28388 15380
rect 29999 14836 30007 15380
rect 28380 14828 28404 14836
rect 28338 14820 28404 14828
rect 29983 14828 30007 14836
rect 30025 15380 30049 15388
rect 30101 15388 30167 15396
rect 30101 15380 30125 15388
rect 30025 14836 30033 15380
rect 30117 14836 30125 15380
rect 30025 14828 30049 14836
rect 29983 14820 30049 14828
rect 30101 14828 30125 14836
rect 30143 15380 30167 15388
rect 30219 15388 30285 15396
rect 30219 15380 30243 15388
rect 30143 14836 30151 15380
rect 30235 14836 30243 15380
rect 30143 14828 30167 14836
rect 30101 14820 30167 14828
rect 30219 14828 30243 14836
rect 30261 15380 30285 15388
rect 30337 15388 30403 15396
rect 30337 15380 30361 15388
rect 30261 14836 30269 15380
rect 30353 14836 30361 15380
rect 30261 14828 30285 14836
rect 30219 14820 30285 14828
rect 30337 14828 30361 14836
rect 30379 15380 30403 15388
rect 30455 15388 30521 15396
rect 30455 15380 30479 15388
rect 30379 14836 30387 15380
rect 30471 14836 30479 15380
rect 30379 14828 30403 14836
rect 30337 14820 30403 14828
rect 30455 14828 30479 14836
rect 30497 15380 30521 15388
rect 30573 15388 30639 15396
rect 30573 15380 30597 15388
rect 30497 14836 30505 15380
rect 30589 14836 30597 15380
rect 30497 14828 30521 14836
rect 30455 14820 30521 14828
rect 30573 14828 30597 14836
rect 30615 15380 30639 15388
rect 30691 15388 30757 15396
rect 30691 15380 30715 15388
rect 30615 14836 30623 15380
rect 30707 14836 30715 15380
rect 30615 14828 30639 14836
rect 30573 14820 30639 14828
rect 30691 14828 30715 14836
rect 30733 15380 30757 15388
rect 30809 15388 30875 15396
rect 30809 15380 30833 15388
rect 30733 14836 30741 15380
rect 30825 14836 30833 15380
rect 30733 14828 30757 14836
rect 30691 14820 30757 14828
rect 30809 14828 30833 14836
rect 30851 15380 30875 15388
rect 30927 15388 30993 15396
rect 30927 15380 30951 15388
rect 30851 14836 30859 15380
rect 30943 14836 30951 15380
rect 30851 14828 30875 14836
rect 30809 14820 30875 14828
rect 30927 14828 30951 14836
rect 30969 15380 30993 15388
rect 31045 15388 31111 15396
rect 31045 15380 31069 15388
rect 30969 14836 30977 15380
rect 31061 14836 31069 15380
rect 30969 14828 30993 14836
rect 30927 14820 30993 14828
rect 31045 14828 31069 14836
rect 31087 15380 31111 15388
rect 31163 15388 31229 15396
rect 31163 15380 31187 15388
rect 31087 14836 31095 15380
rect 31179 14836 31187 15380
rect 31087 14828 31111 14836
rect 31045 14820 31111 14828
rect 31163 14828 31187 14836
rect 31205 15380 31229 15388
rect 31281 15388 31347 15396
rect 31281 15380 31305 15388
rect 31205 14836 31213 15380
rect 31297 14836 31305 15380
rect 31205 14828 31229 14836
rect 31163 14820 31229 14828
rect 31281 14828 31305 14836
rect 31323 15380 31347 15388
rect 31399 15388 31465 15396
rect 31399 15380 31423 15388
rect 31323 14836 31331 15380
rect 31415 14836 31423 15380
rect 31323 14828 31347 14836
rect 31281 14820 31347 14828
rect 31399 14828 31423 14836
rect 31441 15380 31465 15388
rect 31517 15388 31583 15396
rect 31517 15380 31541 15388
rect 31441 14836 31449 15380
rect 31533 14836 31541 15380
rect 31441 14828 31465 14836
rect 31399 14820 31465 14828
rect 31517 14828 31541 14836
rect 31559 15380 31583 15388
rect 31635 15388 31701 15396
rect 31635 15380 31659 15388
rect 31559 14836 31567 15380
rect 31651 14836 31659 15380
rect 31559 14828 31583 14836
rect 31517 14820 31583 14828
rect 31635 14828 31659 14836
rect 31677 15380 31701 15388
rect 31753 15388 31819 15396
rect 31753 15380 31777 15388
rect 31677 14836 31685 15380
rect 31769 14836 31777 15380
rect 31677 14828 31701 14836
rect 31635 14820 31701 14828
rect 31753 14828 31777 14836
rect 31795 15380 31819 15388
rect 31871 15388 31937 15396
rect 31871 15380 31895 15388
rect 31795 14836 31803 15380
rect 31887 14836 31895 15380
rect 31795 14828 31819 14836
rect 31753 14820 31819 14828
rect 31871 14828 31895 14836
rect 31913 15380 31937 15388
rect 31989 15388 32055 15396
rect 31989 15380 32013 15388
rect 31913 14836 31921 15380
rect 32005 14836 32013 15380
rect 31913 14828 31937 14836
rect 31871 14820 31937 14828
rect 31989 14828 32013 14836
rect 32031 15380 32055 15388
rect 32107 15388 32173 15396
rect 32107 15380 32131 15388
rect 32031 14836 32039 15380
rect 32123 14836 32131 15380
rect 32031 14828 32055 14836
rect 31989 14820 32055 14828
rect 32107 14828 32131 14836
rect 32149 15380 32173 15388
rect 32225 15388 32291 15396
rect 32225 15380 32249 15388
rect 32149 14836 32157 15380
rect 32241 14836 32249 15380
rect 32149 14828 32173 14836
rect 32107 14820 32173 14828
rect 32225 14828 32249 14836
rect 32267 15380 32291 15388
rect 32343 15388 32409 15396
rect 32343 15380 32367 15388
rect 32267 14836 32275 15380
rect 32359 14836 32367 15380
rect 32267 14828 32291 14836
rect 32225 14820 32291 14828
rect 32343 14828 32367 14836
rect 32385 15380 32409 15388
rect 32461 15388 32527 15396
rect 32461 15380 32485 15388
rect 32385 14836 32393 15380
rect 32477 14836 32485 15380
rect 32385 14828 32409 14836
rect 32343 14820 32409 14828
rect 32461 14828 32485 14836
rect 32503 15380 32527 15388
rect 32503 14836 32511 15380
rect 32503 14828 32527 14836
rect 32461 14820 32527 14828
rect 21753 14804 21769 14820
rect 21771 14804 21787 14820
rect 21871 14804 21887 14820
rect 21889 14804 21905 14820
rect 21989 14804 22005 14820
rect 22007 14804 22023 14820
rect 22107 14804 22123 14820
rect 22125 14804 22141 14820
rect 22225 14804 22241 14820
rect 22243 14804 22259 14820
rect 22343 14804 22359 14820
rect 22361 14804 22377 14820
rect 22461 14804 22477 14820
rect 22479 14804 22495 14820
rect 22579 14804 22595 14820
rect 22597 14804 22613 14820
rect 22697 14804 22713 14820
rect 22715 14804 22731 14820
rect 22815 14804 22831 14820
rect 22833 14804 22849 14820
rect 22933 14804 22949 14820
rect 22951 14804 22967 14820
rect 23051 14804 23067 14820
rect 23069 14804 23085 14820
rect 23169 14804 23185 14820
rect 23187 14804 23203 14820
rect 23287 14804 23303 14820
rect 23305 14804 23321 14820
rect 23405 14804 23421 14820
rect 23423 14804 23439 14820
rect 23523 14804 23539 14820
rect 23541 14804 23557 14820
rect 23641 14804 23657 14820
rect 23659 14804 23675 14820
rect 23759 14804 23775 14820
rect 23777 14804 23793 14820
rect 23877 14804 23893 14820
rect 23895 14804 23911 14820
rect 23995 14804 24011 14820
rect 24013 14804 24029 14820
rect 24113 14804 24129 14820
rect 24131 14804 24147 14820
rect 24231 14804 24247 14820
rect 24249 14804 24265 14820
rect 25876 14804 25892 14820
rect 25894 14804 25910 14820
rect 25994 14804 26010 14820
rect 26012 14804 26028 14820
rect 26112 14804 26128 14820
rect 26130 14804 26146 14820
rect 26230 14804 26246 14820
rect 26248 14804 26264 14820
rect 26348 14804 26364 14820
rect 26366 14804 26382 14820
rect 26466 14804 26482 14820
rect 26484 14804 26500 14820
rect 26584 14804 26600 14820
rect 26602 14804 26618 14820
rect 26702 14804 26718 14820
rect 26720 14804 26736 14820
rect 26820 14804 26836 14820
rect 26838 14804 26854 14820
rect 26938 14804 26954 14820
rect 26956 14804 26972 14820
rect 27056 14804 27072 14820
rect 27074 14804 27090 14820
rect 27174 14804 27190 14820
rect 27192 14804 27208 14820
rect 27292 14804 27308 14820
rect 27310 14804 27326 14820
rect 27410 14804 27426 14820
rect 27428 14804 27444 14820
rect 27528 14804 27544 14820
rect 27546 14804 27562 14820
rect 27646 14804 27662 14820
rect 27664 14804 27680 14820
rect 27764 14804 27780 14820
rect 27782 14804 27798 14820
rect 27882 14804 27898 14820
rect 27900 14804 27916 14820
rect 28000 14804 28016 14820
rect 28018 14804 28034 14820
rect 28118 14804 28134 14820
rect 28136 14804 28152 14820
rect 28236 14804 28252 14820
rect 28254 14804 28270 14820
rect 28354 14804 28370 14820
rect 28372 14804 28388 14820
rect 29999 14804 30015 14820
rect 30017 14804 30033 14820
rect 30117 14804 30133 14820
rect 30135 14804 30151 14820
rect 30235 14804 30251 14820
rect 30253 14804 30269 14820
rect 30353 14804 30369 14820
rect 30371 14804 30387 14820
rect 30471 14804 30487 14820
rect 30489 14804 30505 14820
rect 30589 14804 30605 14820
rect 30607 14804 30623 14820
rect 30707 14804 30723 14820
rect 30725 14804 30741 14820
rect 30825 14804 30841 14820
rect 30843 14804 30859 14820
rect 30943 14804 30959 14820
rect 30961 14804 30977 14820
rect 31061 14804 31077 14820
rect 31079 14804 31095 14820
rect 31179 14804 31195 14820
rect 31197 14804 31213 14820
rect 31297 14804 31313 14820
rect 31315 14804 31331 14820
rect 31415 14804 31431 14820
rect 31433 14804 31449 14820
rect 31533 14804 31549 14820
rect 31551 14804 31567 14820
rect 31651 14804 31667 14820
rect 31669 14804 31685 14820
rect 31769 14804 31785 14820
rect 31787 14804 31803 14820
rect 31887 14804 31903 14820
rect 31905 14804 31921 14820
rect 32005 14804 32021 14820
rect 32023 14804 32039 14820
rect 32123 14804 32139 14820
rect 32141 14804 32157 14820
rect 32241 14804 32257 14820
rect 32259 14804 32275 14820
rect 32359 14804 32375 14820
rect 32377 14804 32393 14820
rect 32477 14804 32493 14820
rect 32495 14804 32511 14820
rect 21260 14625 21294 14659
rect 26693 14317 26752 14480
rect 26753 14257 26812 14420
rect 27098 14230 27137 14420
rect 27158 14290 27197 14480
rect 30859 14314 30875 14512
rect 30919 14254 30935 14452
rect 13490 13075 13530 13079
rect 14063 12680 14097 12686
rect 14063 12672 14069 12680
rect 14091 12672 14097 12680
rect 14299 12680 14333 12686
rect 14299 12672 14305 12680
rect 14327 12672 14333 12680
rect 14535 12680 14569 12686
rect 14535 12672 14541 12680
rect 14563 12672 14569 12680
rect 14771 12680 14805 12686
rect 14771 12672 14777 12680
rect 14799 12672 14805 12680
rect 15007 12680 15041 12686
rect 15007 12672 15013 12680
rect 15035 12672 15041 12680
rect 15243 12680 15277 12686
rect 15243 12672 15249 12680
rect 15271 12672 15277 12680
rect 15479 12680 15513 12686
rect 15479 12672 15485 12680
rect 15507 12672 15513 12680
rect 15715 12680 15749 12686
rect 15715 12672 15721 12680
rect 15743 12672 15749 12680
rect 15951 12680 15985 12686
rect 15951 12672 15957 12680
rect 15979 12672 15985 12680
rect 16187 12680 16221 12686
rect 16187 12672 16193 12680
rect 16215 12672 16221 12680
rect 16423 12680 16457 12686
rect 16423 12672 16429 12680
rect 16451 12672 16457 12680
rect 16659 12680 16693 12686
rect 16659 12672 16665 12680
rect 16687 12672 16693 12680
rect 16895 12680 16929 12686
rect 16895 12672 16901 12680
rect 16923 12672 16929 12680
rect 17131 12680 17165 12686
rect 17131 12672 17137 12680
rect 17159 12672 17165 12680
rect 17367 12680 17401 12686
rect 17367 12672 17373 12680
rect 17395 12672 17401 12680
rect 17603 12680 17637 12686
rect 17603 12672 17609 12680
rect 17631 12672 17637 12680
rect 17839 12680 17873 12686
rect 17839 12672 17845 12680
rect 17867 12672 17873 12680
rect 18075 12680 18109 12686
rect 18075 12672 18081 12680
rect 18103 12672 18109 12680
rect 18311 12680 18345 12686
rect 18311 12672 18317 12680
rect 18339 12672 18345 12680
rect 18547 12680 18581 12686
rect 18547 12672 18553 12680
rect 18575 12672 18581 12680
rect 18783 12680 18817 12686
rect 18783 12672 18789 12680
rect 18811 12672 18817 12680
rect 19019 12680 19053 12686
rect 19019 12672 19025 12680
rect 19047 12672 19053 12680
rect 19255 12680 19289 12686
rect 19255 12672 19261 12680
rect 19283 12672 19289 12680
rect 19491 12680 19525 12686
rect 19491 12672 19497 12680
rect 19519 12672 19525 12680
rect 13484 11025 13524 11028
rect 13492 10937 13529 10941
rect 13490 8975 13529 9001
rect 13488 8887 13534 8891
rect 14535 8586 14551 8602
rect 14553 8586 14569 8602
rect 14653 8586 14669 8602
rect 14671 8586 14687 8602
rect 14771 8586 14787 8602
rect 14789 8586 14805 8602
rect 14889 8586 14905 8602
rect 14907 8586 14923 8602
rect 17839 8586 17855 8602
rect 17857 8586 17873 8602
rect 17957 8586 17973 8602
rect 17975 8586 17991 8602
rect 18075 8586 18091 8602
rect 18093 8586 18109 8602
rect 18193 8586 18209 8602
rect 18211 8586 18227 8602
rect 18311 8586 18327 8602
rect 18329 8586 18345 8602
rect 18429 8586 18445 8602
rect 18447 8586 18463 8602
rect 18547 8586 18563 8602
rect 18565 8586 18581 8602
rect 18665 8586 18681 8602
rect 18683 8586 18699 8602
rect 18783 8586 18799 8602
rect 18801 8586 18817 8602
rect 18901 8586 18917 8602
rect 18919 8586 18935 8602
rect 19019 8586 19035 8602
rect 19037 8586 19053 8602
rect 19137 8586 19153 8602
rect 19155 8586 19171 8602
rect 14519 8578 14585 8586
rect 14519 8570 14543 8578
rect 14535 8026 14543 8570
rect 14519 8018 14543 8026
rect 14561 8570 14585 8578
rect 14637 8578 14703 8586
rect 14637 8570 14661 8578
rect 14561 8026 14569 8570
rect 14653 8026 14661 8570
rect 14561 8018 14585 8026
rect 14519 8010 14585 8018
rect 14637 8018 14661 8026
rect 14679 8570 14703 8578
rect 14755 8578 14821 8586
rect 14755 8570 14779 8578
rect 14679 8026 14687 8570
rect 14771 8026 14779 8570
rect 14679 8018 14703 8026
rect 14637 8010 14703 8018
rect 14755 8018 14779 8026
rect 14797 8570 14821 8578
rect 14873 8578 14939 8586
rect 14873 8570 14897 8578
rect 14797 8026 14805 8570
rect 14889 8026 14897 8570
rect 14797 8018 14821 8026
rect 14755 8010 14821 8018
rect 14873 8018 14897 8026
rect 14915 8570 14939 8578
rect 17823 8578 17889 8586
rect 17823 8570 17847 8578
rect 14915 8026 14923 8570
rect 17839 8026 17847 8570
rect 14915 8018 14939 8026
rect 14873 8010 14939 8018
rect 17823 8018 17847 8026
rect 17865 8570 17889 8578
rect 17941 8578 18007 8586
rect 17941 8570 17965 8578
rect 17865 8026 17873 8570
rect 17957 8026 17965 8570
rect 17865 8018 17889 8026
rect 17823 8010 17889 8018
rect 17941 8018 17965 8026
rect 17983 8570 18007 8578
rect 18059 8578 18125 8586
rect 18059 8570 18083 8578
rect 17983 8026 17991 8570
rect 18075 8026 18083 8570
rect 17983 8018 18007 8026
rect 17941 8010 18007 8018
rect 18059 8018 18083 8026
rect 18101 8570 18125 8578
rect 18177 8578 18243 8586
rect 18177 8570 18201 8578
rect 18101 8026 18109 8570
rect 18193 8026 18201 8570
rect 18101 8018 18125 8026
rect 18059 8010 18125 8018
rect 18177 8018 18201 8026
rect 18219 8570 18243 8578
rect 18295 8578 18361 8586
rect 18295 8570 18319 8578
rect 18219 8026 18227 8570
rect 18311 8026 18319 8570
rect 18219 8018 18243 8026
rect 18177 8010 18243 8018
rect 18295 8018 18319 8026
rect 18337 8570 18361 8578
rect 18413 8578 18479 8586
rect 18413 8570 18437 8578
rect 18337 8026 18345 8570
rect 18429 8026 18437 8570
rect 18337 8018 18361 8026
rect 18295 8010 18361 8018
rect 18413 8018 18437 8026
rect 18455 8570 18479 8578
rect 18531 8578 18597 8586
rect 18531 8570 18555 8578
rect 18455 8026 18463 8570
rect 18547 8026 18555 8570
rect 18455 8018 18479 8026
rect 18413 8010 18479 8018
rect 18531 8018 18555 8026
rect 18573 8570 18597 8578
rect 18649 8578 18715 8586
rect 18649 8570 18673 8578
rect 18573 8026 18581 8570
rect 18665 8026 18673 8570
rect 18573 8018 18597 8026
rect 18531 8010 18597 8018
rect 18649 8018 18673 8026
rect 18691 8570 18715 8578
rect 18767 8578 18833 8586
rect 18767 8570 18791 8578
rect 18691 8026 18699 8570
rect 18783 8026 18791 8570
rect 18691 8018 18715 8026
rect 18649 8010 18715 8018
rect 18767 8018 18791 8026
rect 18809 8570 18833 8578
rect 18885 8578 18951 8586
rect 18885 8570 18909 8578
rect 18809 8026 18817 8570
rect 18901 8026 18909 8570
rect 18809 8018 18833 8026
rect 18767 8010 18833 8018
rect 18885 8018 18909 8026
rect 18927 8570 18951 8578
rect 19003 8578 19069 8586
rect 19003 8570 19027 8578
rect 18927 8026 18935 8570
rect 19019 8026 19027 8570
rect 18927 8018 18951 8026
rect 18885 8010 18951 8018
rect 19003 8018 19027 8026
rect 19045 8570 19069 8578
rect 19121 8578 19187 8586
rect 19121 8570 19145 8578
rect 19045 8026 19053 8570
rect 19137 8026 19145 8570
rect 19045 8018 19069 8026
rect 19003 8010 19069 8018
rect 19121 8018 19145 8026
rect 19163 8570 19187 8578
rect 19163 8026 19171 8570
rect 19163 8018 19187 8026
rect 19121 8010 19187 8018
rect 14535 7994 14551 8010
rect 14553 7994 14569 8010
rect 14653 7994 14669 8010
rect 14671 7994 14687 8010
rect 14771 7994 14787 8010
rect 14789 7994 14805 8010
rect 14889 7994 14905 8010
rect 14907 7994 14923 8010
rect 17839 7994 17855 8010
rect 17857 7994 17873 8010
rect 17957 7994 17973 8010
rect 17975 7994 17991 8010
rect 18075 7994 18091 8010
rect 18093 7994 18109 8010
rect 18193 7994 18209 8010
rect 18211 7994 18227 8010
rect 18311 7994 18327 8010
rect 18329 7994 18345 8010
rect 18429 7994 18445 8010
rect 18447 7994 18463 8010
rect 18547 7994 18563 8010
rect 18565 7994 18581 8010
rect 18665 7994 18681 8010
rect 18683 7994 18699 8010
rect 18783 7994 18799 8010
rect 18801 7994 18817 8010
rect 18901 7994 18917 8010
rect 18919 7994 18935 8010
rect 19019 7994 19035 8010
rect 19037 7994 19053 8010
rect 19137 7994 19153 8010
rect 19155 7994 19171 8010
rect 14535 7750 14551 7766
rect 14553 7750 14569 7766
rect 14653 7750 14669 7766
rect 14671 7750 14687 7766
rect 14771 7750 14787 7766
rect 14789 7750 14805 7766
rect 14889 7750 14905 7766
rect 14907 7750 14923 7766
rect 17839 7750 17855 7766
rect 17857 7750 17873 7766
rect 17957 7750 17973 7766
rect 17975 7750 17991 7766
rect 18075 7750 18091 7766
rect 18093 7750 18109 7766
rect 18193 7750 18209 7766
rect 18211 7750 18227 7766
rect 18311 7750 18327 7766
rect 18329 7750 18345 7766
rect 18429 7750 18445 7766
rect 18447 7750 18463 7766
rect 18547 7750 18563 7766
rect 18565 7750 18581 7766
rect 18665 7750 18681 7766
rect 18683 7750 18699 7766
rect 18783 7750 18799 7766
rect 18801 7750 18817 7766
rect 18901 7750 18917 7766
rect 18919 7750 18935 7766
rect 19019 7750 19035 7766
rect 19037 7750 19053 7766
rect 19137 7750 19153 7766
rect 19155 7750 19171 7766
rect 14519 7742 14585 7750
rect 14519 7734 14543 7742
rect 14535 7190 14543 7734
rect 14519 7182 14543 7190
rect 14561 7734 14585 7742
rect 14637 7742 14703 7750
rect 14637 7734 14661 7742
rect 14561 7190 14569 7734
rect 14653 7190 14661 7734
rect 14561 7182 14585 7190
rect 14519 7174 14585 7182
rect 14637 7182 14661 7190
rect 14679 7734 14703 7742
rect 14755 7742 14821 7750
rect 14755 7734 14779 7742
rect 14679 7190 14687 7734
rect 14771 7190 14779 7734
rect 14679 7182 14703 7190
rect 14637 7174 14703 7182
rect 14755 7182 14779 7190
rect 14797 7734 14821 7742
rect 14873 7742 14939 7750
rect 14873 7734 14897 7742
rect 14797 7190 14805 7734
rect 14889 7190 14897 7734
rect 14797 7182 14821 7190
rect 14755 7174 14821 7182
rect 14873 7182 14897 7190
rect 14915 7734 14939 7742
rect 17823 7742 17889 7750
rect 17823 7734 17847 7742
rect 14915 7190 14923 7734
rect 17839 7190 17847 7734
rect 14915 7182 14939 7190
rect 14873 7174 14939 7182
rect 17823 7182 17847 7190
rect 17865 7734 17889 7742
rect 17941 7742 18007 7750
rect 17941 7734 17965 7742
rect 17865 7190 17873 7734
rect 17957 7190 17965 7734
rect 17865 7182 17889 7190
rect 17823 7174 17889 7182
rect 17941 7182 17965 7190
rect 17983 7734 18007 7742
rect 18059 7742 18125 7750
rect 18059 7734 18083 7742
rect 17983 7190 17991 7734
rect 18075 7190 18083 7734
rect 17983 7182 18007 7190
rect 17941 7174 18007 7182
rect 18059 7182 18083 7190
rect 18101 7734 18125 7742
rect 18177 7742 18243 7750
rect 18177 7734 18201 7742
rect 18101 7190 18109 7734
rect 18193 7190 18201 7734
rect 18101 7182 18125 7190
rect 18059 7174 18125 7182
rect 18177 7182 18201 7190
rect 18219 7734 18243 7742
rect 18295 7742 18361 7750
rect 18295 7734 18319 7742
rect 18219 7190 18227 7734
rect 18311 7190 18319 7734
rect 18219 7182 18243 7190
rect 18177 7174 18243 7182
rect 18295 7182 18319 7190
rect 18337 7734 18361 7742
rect 18413 7742 18479 7750
rect 18413 7734 18437 7742
rect 18337 7190 18345 7734
rect 18429 7190 18437 7734
rect 18337 7182 18361 7190
rect 18295 7174 18361 7182
rect 18413 7182 18437 7190
rect 18455 7734 18479 7742
rect 18531 7742 18597 7750
rect 18531 7734 18555 7742
rect 18455 7190 18463 7734
rect 18547 7190 18555 7734
rect 18455 7182 18479 7190
rect 18413 7174 18479 7182
rect 18531 7182 18555 7190
rect 18573 7734 18597 7742
rect 18649 7742 18715 7750
rect 18649 7734 18673 7742
rect 18573 7190 18581 7734
rect 18665 7190 18673 7734
rect 18573 7182 18597 7190
rect 18531 7174 18597 7182
rect 18649 7182 18673 7190
rect 18691 7734 18715 7742
rect 18767 7742 18833 7750
rect 18767 7734 18791 7742
rect 18691 7190 18699 7734
rect 18783 7190 18791 7734
rect 18691 7182 18715 7190
rect 18649 7174 18715 7182
rect 18767 7182 18791 7190
rect 18809 7734 18833 7742
rect 18885 7742 18951 7750
rect 18885 7734 18909 7742
rect 18809 7190 18817 7734
rect 18901 7190 18909 7734
rect 18809 7182 18833 7190
rect 18767 7174 18833 7182
rect 18885 7182 18909 7190
rect 18927 7734 18951 7742
rect 19003 7742 19069 7750
rect 19003 7734 19027 7742
rect 18927 7190 18935 7734
rect 19019 7190 19027 7734
rect 18927 7182 18951 7190
rect 18885 7174 18951 7182
rect 19003 7182 19027 7190
rect 19045 7734 19069 7742
rect 19121 7742 19187 7750
rect 19121 7734 19145 7742
rect 19045 7190 19053 7734
rect 19137 7190 19145 7734
rect 19045 7182 19069 7190
rect 19003 7174 19069 7182
rect 19121 7182 19145 7190
rect 19163 7734 19187 7742
rect 19163 7190 19171 7734
rect 19163 7182 19187 7190
rect 19121 7174 19187 7182
rect 14535 7158 14551 7174
rect 14553 7158 14569 7174
rect 14653 7158 14669 7174
rect 14671 7158 14687 7174
rect 14771 7158 14787 7174
rect 14789 7158 14805 7174
rect 14889 7158 14905 7174
rect 14907 7158 14923 7174
rect 17839 7158 17855 7174
rect 17857 7158 17873 7174
rect 17957 7158 17973 7174
rect 17975 7158 17991 7174
rect 18075 7158 18091 7174
rect 18093 7158 18109 7174
rect 18193 7158 18209 7174
rect 18211 7158 18227 7174
rect 18311 7158 18327 7174
rect 18329 7158 18345 7174
rect 18429 7158 18445 7174
rect 18447 7158 18463 7174
rect 18547 7158 18563 7174
rect 18565 7158 18581 7174
rect 18665 7158 18681 7174
rect 18683 7158 18699 7174
rect 18783 7158 18799 7174
rect 18801 7158 18817 7174
rect 18901 7158 18917 7174
rect 18919 7158 18935 7174
rect 19019 7158 19035 7174
rect 19037 7158 19053 7174
rect 19137 7158 19153 7174
rect 19155 7158 19171 7174
rect 13419 7048 13437 7102
rect 13447 7048 13465 7102
rect 13456 7020 13465 7048
rect 13818 7033 13824 7039
rect 13864 7033 13870 7039
rect 14054 7033 14060 7039
rect 14100 7033 14106 7039
rect 14290 7033 14296 7039
rect 14336 7033 14342 7039
rect 14526 7033 14532 7039
rect 14572 7033 14578 7039
rect 14762 7033 14768 7039
rect 14808 7033 14814 7039
rect 14998 7033 15004 7039
rect 15044 7033 15050 7039
rect 15234 7033 15240 7039
rect 15280 7033 15286 7039
rect 15470 7033 15476 7039
rect 15516 7033 15522 7039
rect 15706 7033 15712 7039
rect 15752 7033 15758 7039
rect 15942 7033 15948 7039
rect 15988 7033 15994 7039
rect 16178 7033 16184 7039
rect 16224 7033 16230 7039
rect 16414 7033 16420 7039
rect 16460 7033 16466 7039
rect 16650 7033 16656 7039
rect 16696 7033 16702 7039
rect 16886 7033 16892 7039
rect 16932 7033 16938 7039
rect 17122 7033 17128 7039
rect 17168 7033 17174 7039
rect 17358 7033 17364 7039
rect 17404 7033 17410 7039
rect 17594 7033 17600 7039
rect 17640 7033 17646 7039
rect 17830 7033 17836 7039
rect 17876 7033 17882 7039
rect 18066 7033 18072 7039
rect 18112 7033 18118 7039
rect 18302 7033 18308 7039
rect 18348 7033 18354 7039
rect 18538 7033 18544 7039
rect 18584 7033 18590 7039
rect 18774 7033 18780 7039
rect 18820 7033 18826 7039
rect 19010 7033 19016 7039
rect 19056 7033 19062 7039
rect 19246 7033 19252 7039
rect 19292 7033 19298 7039
rect 19482 7033 19488 7039
rect 19528 7033 19534 7039
rect 13812 7027 13818 7033
rect 13870 7027 13876 7033
rect 14048 7027 14054 7033
rect 14106 7027 14112 7033
rect 14284 7027 14290 7033
rect 14342 7027 14348 7033
rect 14520 7027 14526 7033
rect 14578 7027 14584 7033
rect 14756 7027 14762 7033
rect 14814 7027 14820 7033
rect 14992 7027 14998 7033
rect 15050 7027 15056 7033
rect 15228 7027 15234 7033
rect 15286 7027 15292 7033
rect 15464 7027 15470 7033
rect 15522 7027 15528 7033
rect 15700 7027 15706 7033
rect 15758 7027 15764 7033
rect 15936 7027 15942 7033
rect 15994 7027 16000 7033
rect 16172 7027 16178 7033
rect 16230 7027 16236 7033
rect 16408 7027 16414 7033
rect 16466 7027 16472 7033
rect 16644 7027 16650 7033
rect 16702 7027 16708 7033
rect 16880 7027 16886 7033
rect 16938 7027 16944 7033
rect 17116 7027 17122 7033
rect 17174 7027 17180 7033
rect 17352 7027 17358 7033
rect 17410 7027 17416 7033
rect 17588 7027 17594 7033
rect 17646 7027 17652 7033
rect 17824 7027 17830 7033
rect 17882 7027 17888 7033
rect 18060 7027 18066 7033
rect 18118 7027 18124 7033
rect 18296 7027 18302 7033
rect 18354 7027 18360 7033
rect 18532 7027 18538 7033
rect 18590 7027 18596 7033
rect 18768 7027 18774 7033
rect 18826 7027 18832 7033
rect 19004 7027 19010 7033
rect 19062 7027 19068 7033
rect 19240 7027 19246 7033
rect 19298 7027 19304 7033
rect 19476 7027 19482 7033
rect 19534 7027 19540 7033
rect 13813 6948 19603 6961
rect 13777 6912 19567 6925
rect 26214 6815 26238 6901
rect 26550 6817 26576 6901
rect 13812 6783 13818 6789
rect 13870 6783 13876 6789
rect 14048 6783 14054 6789
rect 14106 6783 14112 6789
rect 14284 6783 14290 6789
rect 14342 6783 14348 6789
rect 14520 6783 14526 6789
rect 14578 6783 14584 6789
rect 14756 6783 14762 6789
rect 14814 6783 14820 6789
rect 14992 6783 14998 6789
rect 15050 6783 15056 6789
rect 15228 6783 15234 6789
rect 15286 6783 15292 6789
rect 15464 6783 15470 6789
rect 15522 6783 15528 6789
rect 15700 6783 15706 6789
rect 15758 6783 15764 6789
rect 15936 6783 15942 6789
rect 15994 6783 16000 6789
rect 16172 6783 16178 6789
rect 16230 6783 16236 6789
rect 16408 6783 16414 6789
rect 16466 6783 16472 6789
rect 16644 6783 16650 6789
rect 16702 6783 16708 6789
rect 16880 6783 16886 6789
rect 16938 6783 16944 6789
rect 17116 6783 17122 6789
rect 17174 6783 17180 6789
rect 17352 6783 17358 6789
rect 17410 6783 17416 6789
rect 17588 6783 17594 6789
rect 17646 6783 17652 6789
rect 17824 6783 17830 6789
rect 17882 6783 17888 6789
rect 18060 6783 18066 6789
rect 18118 6783 18124 6789
rect 18296 6783 18302 6789
rect 18354 6783 18360 6789
rect 18532 6783 18538 6789
rect 18590 6783 18596 6789
rect 18768 6783 18774 6789
rect 18826 6783 18832 6789
rect 19004 6783 19010 6789
rect 19062 6783 19068 6789
rect 19240 6783 19246 6789
rect 19298 6783 19304 6789
rect 19476 6783 19482 6789
rect 19534 6783 19540 6789
rect 13818 6777 13824 6783
rect 13864 6777 13870 6783
rect 14054 6777 14060 6783
rect 14100 6777 14106 6783
rect 14290 6777 14296 6783
rect 14336 6777 14342 6783
rect 14526 6777 14532 6783
rect 14572 6777 14578 6783
rect 14762 6777 14768 6783
rect 14808 6777 14814 6783
rect 14998 6777 15004 6783
rect 15044 6777 15050 6783
rect 15234 6777 15240 6783
rect 15280 6777 15286 6783
rect 15470 6777 15476 6783
rect 15516 6777 15522 6783
rect 15706 6777 15712 6783
rect 15752 6777 15758 6783
rect 15942 6777 15948 6783
rect 15988 6777 15994 6783
rect 16178 6777 16184 6783
rect 16224 6777 16230 6783
rect 16414 6777 16420 6783
rect 16460 6777 16466 6783
rect 16650 6777 16656 6783
rect 16696 6777 16702 6783
rect 16886 6777 16892 6783
rect 16932 6777 16938 6783
rect 17122 6777 17128 6783
rect 17168 6777 17174 6783
rect 17358 6777 17364 6783
rect 17404 6777 17410 6783
rect 17594 6777 17600 6783
rect 17640 6777 17646 6783
rect 17830 6777 17836 6783
rect 17876 6777 17882 6783
rect 18066 6777 18072 6783
rect 18112 6777 18118 6783
rect 18302 6777 18308 6783
rect 18348 6777 18354 6783
rect 18538 6777 18544 6783
rect 18584 6777 18590 6783
rect 18774 6777 18780 6783
rect 18820 6777 18826 6783
rect 19010 6777 19016 6783
rect 19056 6777 19062 6783
rect 19246 6777 19252 6783
rect 19292 6777 19298 6783
rect 19482 6777 19488 6783
rect 19528 6777 19534 6783
rect 15129 6343 15145 6359
rect 15147 6343 15163 6359
rect 15247 6343 15263 6359
rect 15265 6343 15281 6359
rect 15365 6343 15381 6359
rect 15383 6343 15399 6359
rect 15483 6343 15499 6359
rect 15501 6343 15517 6359
rect 16655 6343 16671 6359
rect 16673 6343 16689 6359
rect 16773 6343 16789 6359
rect 16791 6343 16807 6359
rect 16891 6343 16907 6359
rect 16909 6343 16925 6359
rect 17009 6343 17025 6359
rect 17027 6343 17043 6359
rect 17127 6343 17143 6359
rect 17145 6343 17161 6359
rect 17245 6343 17261 6359
rect 17263 6343 17279 6359
rect 17363 6343 17379 6359
rect 17381 6343 17397 6359
rect 17481 6343 17497 6359
rect 17499 6343 17515 6359
rect 17599 6343 17615 6359
rect 17617 6343 17633 6359
rect 17717 6343 17733 6359
rect 17735 6343 17751 6359
rect 17835 6343 17851 6359
rect 17853 6343 17869 6359
rect 17953 6343 17969 6359
rect 17971 6343 17987 6359
rect 18071 6343 18087 6359
rect 18089 6343 18105 6359
rect 18189 6343 18205 6359
rect 18207 6343 18223 6359
rect 18307 6343 18323 6359
rect 18325 6343 18341 6359
rect 18425 6343 18441 6359
rect 18443 6343 18459 6359
rect 15113 6335 15179 6343
rect 15113 6327 15137 6335
rect 15129 5783 15137 6327
rect 15113 5775 15137 5783
rect 15155 6327 15179 6335
rect 15231 6335 15297 6343
rect 15231 6327 15255 6335
rect 15155 5783 15163 6327
rect 15247 5783 15255 6327
rect 15155 5775 15179 5783
rect 15113 5767 15179 5775
rect 15231 5775 15255 5783
rect 15273 6327 15297 6335
rect 15349 6335 15415 6343
rect 15349 6327 15373 6335
rect 15273 5783 15281 6327
rect 15365 5783 15373 6327
rect 15273 5775 15297 5783
rect 15231 5767 15297 5775
rect 15349 5775 15373 5783
rect 15391 6327 15415 6335
rect 15467 6335 15533 6343
rect 15467 6327 15491 6335
rect 15391 5783 15399 6327
rect 15483 5783 15491 6327
rect 15391 5775 15415 5783
rect 15349 5767 15415 5775
rect 15467 5775 15491 5783
rect 15509 6327 15533 6335
rect 16639 6335 16705 6343
rect 16639 6327 16663 6335
rect 15509 5783 15517 6327
rect 16655 5783 16663 6327
rect 15509 5775 15533 5783
rect 15467 5767 15533 5775
rect 16639 5775 16663 5783
rect 16681 6327 16705 6335
rect 16757 6335 16823 6343
rect 16757 6327 16781 6335
rect 16681 5783 16689 6327
rect 16773 5783 16781 6327
rect 16681 5775 16705 5783
rect 16639 5767 16705 5775
rect 16757 5775 16781 5783
rect 16799 6327 16823 6335
rect 16875 6335 16941 6343
rect 16875 6327 16899 6335
rect 16799 5783 16807 6327
rect 16891 5783 16899 6327
rect 16799 5775 16823 5783
rect 16757 5767 16823 5775
rect 16875 5775 16899 5783
rect 16917 6327 16941 6335
rect 16993 6335 17059 6343
rect 16993 6327 17017 6335
rect 16917 5783 16925 6327
rect 17009 5783 17017 6327
rect 16917 5775 16941 5783
rect 16875 5767 16941 5775
rect 16993 5775 17017 5783
rect 17035 6327 17059 6335
rect 17111 6335 17177 6343
rect 17111 6327 17135 6335
rect 17035 5783 17043 6327
rect 17127 5783 17135 6327
rect 17035 5775 17059 5783
rect 16993 5767 17059 5775
rect 17111 5775 17135 5783
rect 17153 6327 17177 6335
rect 17229 6335 17295 6343
rect 17229 6327 17253 6335
rect 17153 5783 17161 6327
rect 17245 5783 17253 6327
rect 17153 5775 17177 5783
rect 17111 5767 17177 5775
rect 17229 5775 17253 5783
rect 17271 6327 17295 6335
rect 17347 6335 17413 6343
rect 17347 6327 17371 6335
rect 17271 5783 17279 6327
rect 17363 5783 17371 6327
rect 17271 5775 17295 5783
rect 17229 5767 17295 5775
rect 17347 5775 17371 5783
rect 17389 6327 17413 6335
rect 17465 6335 17531 6343
rect 17465 6327 17489 6335
rect 17389 5783 17397 6327
rect 17481 5783 17489 6327
rect 17389 5775 17413 5783
rect 17347 5767 17413 5775
rect 17465 5775 17489 5783
rect 17507 6327 17531 6335
rect 17583 6335 17649 6343
rect 17583 6327 17607 6335
rect 17507 5783 17515 6327
rect 17599 5783 17607 6327
rect 17507 5775 17531 5783
rect 17465 5767 17531 5775
rect 17583 5775 17607 5783
rect 17625 6327 17649 6335
rect 17701 6335 17767 6343
rect 17701 6327 17725 6335
rect 17625 5783 17633 6327
rect 17717 5783 17725 6327
rect 17625 5775 17649 5783
rect 17583 5767 17649 5775
rect 17701 5775 17725 5783
rect 17743 6327 17767 6335
rect 17819 6335 17885 6343
rect 17819 6327 17843 6335
rect 17743 5783 17751 6327
rect 17835 5783 17843 6327
rect 17743 5775 17767 5783
rect 17701 5767 17767 5775
rect 17819 5775 17843 5783
rect 17861 6327 17885 6335
rect 17937 6335 18003 6343
rect 17937 6327 17961 6335
rect 17861 5783 17869 6327
rect 17953 5783 17961 6327
rect 17861 5775 17885 5783
rect 17819 5767 17885 5775
rect 17937 5775 17961 5783
rect 17979 6327 18003 6335
rect 18055 6335 18121 6343
rect 18055 6327 18079 6335
rect 17979 5783 17987 6327
rect 18071 5783 18079 6327
rect 17979 5775 18003 5783
rect 17937 5767 18003 5775
rect 18055 5775 18079 5783
rect 18097 6327 18121 6335
rect 18173 6335 18239 6343
rect 18173 6327 18197 6335
rect 18097 5783 18105 6327
rect 18189 5783 18197 6327
rect 18097 5775 18121 5783
rect 18055 5767 18121 5775
rect 18173 5775 18197 5783
rect 18215 6327 18239 6335
rect 18291 6335 18357 6343
rect 18291 6327 18315 6335
rect 18215 5783 18223 6327
rect 18307 5783 18315 6327
rect 18215 5775 18239 5783
rect 18173 5767 18239 5775
rect 18291 5775 18315 5783
rect 18333 6327 18357 6335
rect 18409 6335 18475 6343
rect 18409 6327 18433 6335
rect 18333 5783 18341 6327
rect 18425 5783 18433 6327
rect 18333 5775 18357 5783
rect 18291 5767 18357 5775
rect 18409 5775 18433 5783
rect 18451 6327 18475 6335
rect 19202 6333 19236 6367
rect 22499 6343 22515 6359
rect 22517 6343 22533 6359
rect 22647 6343 22663 6359
rect 22665 6343 22681 6359
rect 22795 6343 22811 6359
rect 22813 6343 22829 6359
rect 22943 6343 22959 6359
rect 22961 6343 22977 6359
rect 23091 6343 23107 6359
rect 23109 6343 23125 6359
rect 23239 6343 23255 6359
rect 23257 6343 23273 6359
rect 23387 6343 23403 6359
rect 23405 6343 23421 6359
rect 23535 6343 23551 6359
rect 23553 6343 23569 6359
rect 23683 6343 23699 6359
rect 23701 6343 23717 6359
rect 23831 6343 23847 6359
rect 23849 6343 23865 6359
rect 23979 6343 23995 6359
rect 23997 6343 24013 6359
rect 24127 6343 24143 6359
rect 24145 6343 24161 6359
rect 24275 6343 24291 6359
rect 24293 6343 24309 6359
rect 24423 6343 24439 6359
rect 24441 6343 24457 6359
rect 24571 6343 24587 6359
rect 24589 6343 24605 6359
rect 24719 6343 24735 6359
rect 24737 6343 24753 6359
rect 24867 6343 24883 6359
rect 24885 6343 24901 6359
rect 25015 6343 25031 6359
rect 25033 6343 25049 6359
rect 25163 6343 25179 6359
rect 25181 6343 25197 6359
rect 25311 6343 25327 6359
rect 25329 6343 25345 6359
rect 25459 6343 25475 6359
rect 25477 6343 25493 6359
rect 25607 6343 25623 6359
rect 25625 6343 25641 6359
rect 25755 6343 25771 6359
rect 25773 6343 25789 6359
rect 25903 6343 25919 6359
rect 25921 6343 25937 6359
rect 26051 6343 26067 6359
rect 26069 6343 26085 6359
rect 26199 6343 26215 6359
rect 26217 6343 26233 6359
rect 26347 6343 26363 6359
rect 26365 6343 26381 6359
rect 26495 6343 26511 6359
rect 26513 6343 26529 6359
rect 26643 6343 26659 6359
rect 26661 6343 26677 6359
rect 26791 6343 26807 6359
rect 26809 6343 26825 6359
rect 26939 6343 26955 6359
rect 26957 6343 26973 6359
rect 27087 6343 27103 6359
rect 27105 6343 27121 6359
rect 27235 6343 27251 6359
rect 27253 6343 27269 6359
rect 27383 6343 27399 6359
rect 27401 6343 27417 6359
rect 27531 6343 27547 6359
rect 27549 6343 27565 6359
rect 27679 6343 27695 6359
rect 27697 6343 27713 6359
rect 27827 6343 27843 6359
rect 27845 6343 27861 6359
rect 27975 6343 27991 6359
rect 27993 6343 28009 6359
rect 28123 6343 28139 6359
rect 28141 6343 28157 6359
rect 28271 6343 28287 6359
rect 28289 6343 28305 6359
rect 28419 6343 28435 6359
rect 28437 6343 28453 6359
rect 28567 6343 28583 6359
rect 28585 6343 28601 6359
rect 28715 6343 28731 6359
rect 28733 6343 28749 6359
rect 28863 6343 28879 6359
rect 28881 6343 28897 6359
rect 29011 6343 29027 6359
rect 29029 6343 29045 6359
rect 29159 6343 29175 6359
rect 29177 6343 29193 6359
rect 29307 6343 29323 6359
rect 29325 6343 29341 6359
rect 29455 6343 29471 6359
rect 29473 6343 29489 6359
rect 29603 6343 29619 6359
rect 29621 6343 29637 6359
rect 29751 6343 29767 6359
rect 29769 6343 29785 6359
rect 29899 6343 29915 6359
rect 29917 6343 29933 6359
rect 30047 6343 30063 6359
rect 30065 6343 30081 6359
rect 30195 6343 30211 6359
rect 30213 6343 30229 6359
rect 30343 6343 30359 6359
rect 30361 6343 30377 6359
rect 30491 6343 30507 6359
rect 30509 6343 30525 6359
rect 30639 6343 30655 6359
rect 30657 6343 30660 6359
rect 22483 6335 22549 6343
rect 22483 6327 22507 6335
rect 18451 5783 18459 6327
rect 19202 6299 19236 6324
rect 19708 6043 19732 6193
rect 20024 6043 20048 6193
rect 20340 6043 20364 6193
rect 20656 6043 20680 6193
rect 20972 6043 20996 6193
rect 19202 5918 19236 5957
rect 19518 5943 19552 5957
rect 19494 5909 19552 5943
rect 19834 5909 19868 5957
rect 20150 5909 20184 5957
rect 20466 5909 20500 5957
rect 20782 5909 20816 5957
rect 21098 5909 21132 5957
rect 19528 5903 19552 5909
rect 19275 5869 19309 5903
rect 19348 5869 19382 5903
rect 19421 5869 19455 5903
rect 19567 5869 19601 5903
rect 19640 5869 19674 5903
rect 19713 5869 19747 5903
rect 19786 5869 19820 5903
rect 19859 5869 19893 5903
rect 19932 5869 19966 5903
rect 20005 5869 20039 5903
rect 20078 5869 20112 5903
rect 20151 5869 20185 5903
rect 20224 5869 20258 5903
rect 20297 5869 20331 5903
rect 20370 5869 20404 5903
rect 20443 5869 20477 5903
rect 20516 5869 20550 5903
rect 20589 5869 20623 5903
rect 20662 5869 20696 5903
rect 20735 5869 20769 5903
rect 20808 5869 20842 5903
rect 20881 5869 20915 5903
rect 20954 5869 20988 5903
rect 21027 5869 21061 5903
rect 21100 5869 21134 5903
rect 18451 5775 18475 5783
rect 18409 5767 18475 5775
rect 15129 5751 15145 5767
rect 15147 5751 15163 5767
rect 15247 5751 15263 5767
rect 15265 5751 15281 5767
rect 15365 5751 15381 5767
rect 15383 5751 15399 5767
rect 15483 5751 15499 5767
rect 15501 5751 15517 5767
rect 16655 5751 16671 5767
rect 16673 5751 16689 5767
rect 16773 5751 16789 5767
rect 16791 5751 16807 5767
rect 16891 5751 16907 5767
rect 16909 5751 16925 5767
rect 17009 5751 17025 5767
rect 17027 5751 17043 5767
rect 17127 5751 17143 5767
rect 17145 5751 17161 5767
rect 17245 5751 17261 5767
rect 17263 5751 17279 5767
rect 17363 5751 17379 5767
rect 17381 5751 17397 5767
rect 17481 5751 17497 5767
rect 17499 5751 17515 5767
rect 17599 5751 17615 5767
rect 17617 5751 17633 5767
rect 17717 5751 17733 5767
rect 17735 5751 17751 5767
rect 17835 5751 17851 5767
rect 17853 5751 17869 5767
rect 17953 5751 17969 5767
rect 17971 5751 17987 5767
rect 18071 5751 18087 5767
rect 18089 5751 18105 5767
rect 18189 5751 18205 5767
rect 18207 5751 18223 5767
rect 18307 5751 18323 5767
rect 18325 5751 18341 5767
rect 18425 5751 18441 5767
rect 18443 5751 18459 5767
rect 16684 5733 16778 5747
rect 16684 5717 16698 5733
rect 16714 5717 16748 5725
rect 16714 5683 16728 5717
rect 16748 5683 16756 5717
rect 16764 5683 16778 5733
rect 16802 5733 16896 5747
rect 16802 5717 16816 5733
rect 16832 5717 16866 5725
rect 16832 5683 16846 5717
rect 16866 5683 16874 5717
rect 16882 5683 16896 5733
rect 16920 5733 17014 5747
rect 16920 5717 16934 5733
rect 16950 5717 16984 5725
rect 16950 5683 16964 5717
rect 16984 5683 16992 5717
rect 17000 5683 17014 5733
rect 17038 5733 17132 5747
rect 17038 5717 17052 5733
rect 17068 5717 17102 5725
rect 17068 5683 17082 5717
rect 17102 5683 17110 5717
rect 17118 5683 17132 5733
rect 17156 5733 17250 5747
rect 17156 5717 17170 5733
rect 17186 5717 17220 5725
rect 17186 5683 17200 5717
rect 17220 5683 17228 5717
rect 17236 5683 17250 5733
rect 17274 5733 17368 5747
rect 17274 5717 17288 5733
rect 17304 5717 17338 5725
rect 17304 5683 17318 5717
rect 17338 5683 17346 5717
rect 17354 5683 17368 5733
rect 17392 5733 17486 5747
rect 17392 5717 17406 5733
rect 17422 5717 17456 5725
rect 17422 5683 17436 5717
rect 17456 5683 17464 5717
rect 17472 5683 17486 5733
rect 17510 5733 17604 5747
rect 17510 5717 17524 5733
rect 17540 5717 17574 5725
rect 17540 5683 17554 5717
rect 17574 5683 17582 5717
rect 17590 5683 17604 5733
rect 17628 5733 17722 5747
rect 17628 5717 17642 5733
rect 17658 5717 17692 5725
rect 17658 5683 17672 5717
rect 17692 5683 17700 5717
rect 17708 5683 17722 5733
rect 17746 5733 17840 5747
rect 17746 5717 17760 5733
rect 17776 5717 17810 5725
rect 17776 5683 17790 5717
rect 17810 5683 17818 5717
rect 17826 5683 17840 5733
rect 17864 5733 17958 5747
rect 17864 5717 17878 5733
rect 17894 5717 17928 5725
rect 17894 5683 17908 5717
rect 17928 5683 17936 5717
rect 17944 5683 17958 5733
rect 17982 5733 18076 5747
rect 17982 5717 17996 5733
rect 18012 5717 18046 5725
rect 18012 5683 18026 5717
rect 18046 5683 18054 5717
rect 18062 5683 18076 5733
rect 18100 5733 18194 5747
rect 18100 5717 18114 5733
rect 18130 5717 18164 5725
rect 18130 5683 18144 5717
rect 18164 5683 18172 5717
rect 18180 5683 18194 5733
rect 18218 5733 18312 5747
rect 18218 5717 18232 5733
rect 18248 5717 18282 5725
rect 18248 5683 18262 5717
rect 18282 5683 18290 5717
rect 18298 5683 18312 5733
rect 18336 5733 18430 5747
rect 18336 5717 18350 5733
rect 18366 5717 18400 5725
rect 18366 5683 18380 5717
rect 18400 5683 18408 5717
rect 18416 5683 18430 5733
rect 16684 5609 16698 5639
rect 16714 5609 16748 5617
rect 16714 5589 16728 5609
rect 16748 5589 16756 5609
rect 16714 5575 16756 5589
rect 16764 5575 16778 5639
rect 16802 5609 16816 5639
rect 16832 5609 16866 5617
rect 16832 5589 16846 5609
rect 16866 5589 16874 5609
rect 16832 5575 16874 5589
rect 16882 5575 16896 5639
rect 16920 5609 16934 5639
rect 16950 5609 16984 5617
rect 16950 5589 16964 5609
rect 16984 5589 16992 5609
rect 16950 5575 16992 5589
rect 17000 5575 17014 5639
rect 17038 5609 17052 5639
rect 17068 5609 17102 5617
rect 17068 5589 17082 5609
rect 17102 5589 17110 5609
rect 17068 5575 17110 5589
rect 17118 5575 17132 5639
rect 17156 5609 17170 5639
rect 17186 5609 17220 5617
rect 17186 5589 17200 5609
rect 17220 5589 17228 5609
rect 17186 5575 17228 5589
rect 17236 5575 17250 5639
rect 17274 5609 17288 5639
rect 17304 5609 17338 5617
rect 17304 5589 17318 5609
rect 17338 5589 17346 5609
rect 17304 5575 17346 5589
rect 17354 5575 17368 5639
rect 17392 5609 17406 5639
rect 17422 5609 17456 5617
rect 17422 5589 17436 5609
rect 17456 5589 17464 5609
rect 17422 5575 17464 5589
rect 17472 5575 17486 5639
rect 17510 5609 17524 5639
rect 17540 5609 17574 5617
rect 17540 5589 17554 5609
rect 17574 5589 17582 5609
rect 17540 5575 17582 5589
rect 17590 5575 17604 5639
rect 17628 5609 17642 5639
rect 17658 5609 17692 5617
rect 17658 5589 17672 5609
rect 17692 5589 17700 5609
rect 17658 5575 17700 5589
rect 17708 5575 17722 5639
rect 17746 5609 17760 5639
rect 17776 5609 17810 5617
rect 17776 5589 17790 5609
rect 17810 5589 17818 5609
rect 17776 5575 17818 5589
rect 17826 5575 17840 5639
rect 17864 5609 17878 5639
rect 17894 5609 17928 5617
rect 17894 5589 17908 5609
rect 17928 5589 17936 5609
rect 17894 5575 17936 5589
rect 17944 5575 17958 5639
rect 17982 5609 17996 5639
rect 18012 5609 18046 5617
rect 18012 5589 18026 5609
rect 18046 5589 18054 5609
rect 18012 5575 18054 5589
rect 18062 5575 18076 5639
rect 18100 5609 18114 5639
rect 18130 5609 18164 5617
rect 18130 5589 18144 5609
rect 18164 5589 18172 5609
rect 18130 5575 18172 5589
rect 18180 5575 18194 5639
rect 18218 5609 18232 5639
rect 18248 5609 18282 5617
rect 18248 5589 18262 5609
rect 18282 5589 18290 5609
rect 18248 5575 18290 5589
rect 18298 5575 18312 5639
rect 18336 5609 18350 5639
rect 18366 5609 18400 5617
rect 18366 5589 18380 5609
rect 18400 5589 18408 5609
rect 18366 5575 18408 5589
rect 18416 5575 18430 5639
rect 15129 5525 15145 5541
rect 15147 5525 15163 5541
rect 15247 5525 15263 5541
rect 15265 5525 15281 5541
rect 15365 5525 15381 5541
rect 15383 5525 15399 5541
rect 15483 5525 15499 5541
rect 15501 5525 15517 5541
rect 16655 5525 16671 5541
rect 16673 5525 16689 5541
rect 16773 5525 16789 5541
rect 16791 5525 16807 5541
rect 16891 5525 16907 5541
rect 16909 5525 16925 5541
rect 17009 5525 17025 5541
rect 17027 5525 17043 5541
rect 17127 5525 17143 5541
rect 17145 5525 17161 5541
rect 17245 5525 17261 5541
rect 17263 5525 17279 5541
rect 17363 5525 17379 5541
rect 17381 5525 17397 5541
rect 17481 5525 17497 5541
rect 17499 5525 17515 5541
rect 17599 5525 17615 5541
rect 17617 5525 17633 5541
rect 17717 5525 17733 5541
rect 17735 5525 17751 5541
rect 17835 5525 17851 5541
rect 17853 5525 17869 5541
rect 17953 5525 17969 5541
rect 17971 5525 17987 5541
rect 18071 5525 18087 5541
rect 18089 5525 18105 5541
rect 18189 5525 18205 5541
rect 18207 5525 18223 5541
rect 18307 5525 18323 5541
rect 18325 5525 18341 5541
rect 18425 5525 18441 5541
rect 18443 5525 18459 5541
rect 15113 5517 15179 5525
rect 15113 5509 15137 5517
rect 15129 5170 15137 5509
rect 15155 5509 15179 5517
rect 15231 5517 15297 5525
rect 15231 5509 15255 5517
rect 15155 5170 15163 5509
rect 15247 5170 15255 5509
rect 15273 5509 15297 5517
rect 15349 5517 15415 5525
rect 15349 5509 15373 5517
rect 15273 5170 15281 5509
rect 15365 5170 15373 5509
rect 15391 5509 15415 5517
rect 15467 5517 15533 5525
rect 15467 5509 15491 5517
rect 15391 5170 15399 5509
rect 15483 5170 15491 5509
rect 15509 5509 15533 5517
rect 16639 5517 16705 5525
rect 16639 5509 16663 5517
rect 15509 5170 15517 5509
rect 16655 5170 16663 5509
rect 16681 5509 16705 5517
rect 16757 5517 16823 5525
rect 16757 5509 16781 5517
rect 16681 5170 16689 5509
rect 16773 5170 16781 5509
rect 16799 5509 16823 5517
rect 16875 5517 16941 5525
rect 16875 5509 16899 5517
rect 16799 5170 16807 5509
rect 16891 5170 16899 5509
rect 16917 5509 16941 5517
rect 16993 5517 17059 5525
rect 16993 5509 17017 5517
rect 16917 5170 16925 5509
rect 17009 5170 17017 5509
rect 17035 5509 17059 5517
rect 17111 5517 17177 5525
rect 17111 5509 17135 5517
rect 17035 5170 17043 5509
rect 17127 5170 17135 5509
rect 17153 5509 17177 5517
rect 17229 5517 17295 5525
rect 17229 5509 17253 5517
rect 17153 5170 17161 5509
rect 17245 5170 17253 5509
rect 17271 5509 17295 5517
rect 17347 5517 17413 5525
rect 17347 5509 17371 5517
rect 17271 5170 17279 5509
rect 17363 5170 17371 5509
rect 17389 5509 17413 5517
rect 17465 5517 17531 5525
rect 17465 5509 17489 5517
rect 17389 5170 17397 5509
rect 17481 5170 17489 5509
rect 17507 5509 17531 5517
rect 17583 5517 17649 5525
rect 17583 5509 17607 5517
rect 17507 5170 17515 5509
rect 17599 5170 17607 5509
rect 17625 5509 17649 5517
rect 17701 5517 17767 5525
rect 17701 5509 17725 5517
rect 17625 5170 17633 5509
rect 17717 5170 17725 5509
rect 17743 5509 17767 5517
rect 17819 5517 17885 5525
rect 17819 5509 17843 5517
rect 17743 5170 17751 5509
rect 17835 5170 17843 5509
rect 17861 5509 17885 5517
rect 17937 5517 18003 5525
rect 17937 5509 17961 5517
rect 17861 5170 17869 5509
rect 17953 5170 17961 5509
rect 17979 5509 18003 5517
rect 18055 5517 18121 5525
rect 18055 5509 18079 5517
rect 17979 5170 17987 5509
rect 18071 5170 18079 5509
rect 18097 5509 18121 5517
rect 18173 5517 18239 5525
rect 18173 5509 18197 5517
rect 18097 5170 18105 5509
rect 18189 5170 18197 5509
rect 18215 5509 18239 5517
rect 18291 5517 18357 5525
rect 18291 5509 18315 5517
rect 18215 5170 18223 5509
rect 18307 5170 18315 5509
rect 18333 5509 18357 5517
rect 18409 5517 18475 5525
rect 18409 5509 18433 5517
rect 18333 5170 18341 5509
rect 18425 5170 18433 5509
rect 18451 5509 18475 5517
rect 18451 5170 18459 5509
rect 22499 5483 22507 6327
rect 22483 5475 22507 5483
rect 22525 6327 22549 6335
rect 22631 6335 22697 6343
rect 22631 6327 22655 6335
rect 22525 5483 22533 6327
rect 22647 5483 22655 6327
rect 22525 5475 22549 5483
rect 22483 5467 22549 5475
rect 22631 5475 22655 5483
rect 22673 6327 22697 6335
rect 22779 6335 22845 6343
rect 22779 6327 22803 6335
rect 22673 5483 22681 6327
rect 22795 5483 22803 6327
rect 22673 5475 22697 5483
rect 22631 5467 22697 5475
rect 22779 5475 22803 5483
rect 22821 6327 22845 6335
rect 22927 6335 22993 6343
rect 22927 6327 22951 6335
rect 22821 5483 22829 6327
rect 22943 5483 22951 6327
rect 22821 5475 22845 5483
rect 22779 5467 22845 5475
rect 22927 5475 22951 5483
rect 22969 6327 22993 6335
rect 23075 6335 23141 6343
rect 23075 6327 23099 6335
rect 22969 5483 22977 6327
rect 23091 5483 23099 6327
rect 22969 5475 22993 5483
rect 22927 5467 22993 5475
rect 23075 5475 23099 5483
rect 23117 6327 23141 6335
rect 23223 6335 23289 6343
rect 23223 6327 23247 6335
rect 23117 5483 23125 6327
rect 23239 5483 23247 6327
rect 23117 5475 23141 5483
rect 23075 5467 23141 5475
rect 23223 5475 23247 5483
rect 23265 6327 23289 6335
rect 23371 6335 23437 6343
rect 23371 6327 23395 6335
rect 23265 5483 23273 6327
rect 23387 5483 23395 6327
rect 23265 5475 23289 5483
rect 23223 5467 23289 5475
rect 23371 5475 23395 5483
rect 23413 6327 23437 6335
rect 23519 6335 23585 6343
rect 23519 6327 23543 6335
rect 23413 5483 23421 6327
rect 23535 5483 23543 6327
rect 23413 5475 23437 5483
rect 23371 5467 23437 5475
rect 23519 5475 23543 5483
rect 23561 6327 23585 6335
rect 23667 6335 23733 6343
rect 23667 6327 23691 6335
rect 23561 5483 23569 6327
rect 23683 5483 23691 6327
rect 23561 5475 23585 5483
rect 23519 5467 23585 5475
rect 23667 5475 23691 5483
rect 23709 6327 23733 6335
rect 23815 6335 23881 6343
rect 23815 6327 23839 6335
rect 23709 5483 23717 6327
rect 23831 5483 23839 6327
rect 23709 5475 23733 5483
rect 23667 5467 23733 5475
rect 23815 5475 23839 5483
rect 23857 6327 23881 6335
rect 23963 6335 24029 6343
rect 23963 6327 23987 6335
rect 23857 5483 23865 6327
rect 23979 5483 23987 6327
rect 23857 5475 23881 5483
rect 23815 5467 23881 5475
rect 23963 5475 23987 5483
rect 24005 6327 24029 6335
rect 24111 6335 24177 6343
rect 24111 6327 24135 6335
rect 24005 5483 24013 6327
rect 24127 5483 24135 6327
rect 24005 5475 24029 5483
rect 23963 5467 24029 5475
rect 24111 5475 24135 5483
rect 24153 6327 24177 6335
rect 24259 6335 24325 6343
rect 24259 6327 24283 6335
rect 24153 5483 24161 6327
rect 24275 5483 24283 6327
rect 24153 5475 24177 5483
rect 24111 5467 24177 5475
rect 24259 5475 24283 5483
rect 24301 6327 24325 6335
rect 24407 6335 24473 6343
rect 24407 6327 24431 6335
rect 24301 5483 24309 6327
rect 24423 5483 24431 6327
rect 24301 5475 24325 5483
rect 24259 5467 24325 5475
rect 24407 5475 24431 5483
rect 24449 6327 24473 6335
rect 24555 6335 24621 6343
rect 24555 6327 24579 6335
rect 24449 5483 24457 6327
rect 24571 5483 24579 6327
rect 24449 5475 24473 5483
rect 24407 5467 24473 5475
rect 24555 5475 24579 5483
rect 24597 6327 24621 6335
rect 24703 6335 24769 6343
rect 24703 6327 24727 6335
rect 24597 5483 24605 6327
rect 24719 5483 24727 6327
rect 24597 5475 24621 5483
rect 24555 5467 24621 5475
rect 24703 5475 24727 5483
rect 24745 6327 24769 6335
rect 24851 6335 24917 6343
rect 24851 6327 24875 6335
rect 24745 5483 24753 6327
rect 24867 5483 24875 6327
rect 24745 5475 24769 5483
rect 24703 5467 24769 5475
rect 24851 5475 24875 5483
rect 24893 6327 24917 6335
rect 24999 6335 25065 6343
rect 24999 6327 25023 6335
rect 24893 5483 24901 6327
rect 25015 5483 25023 6327
rect 24893 5475 24917 5483
rect 24851 5467 24917 5475
rect 24999 5475 25023 5483
rect 25041 6327 25065 6335
rect 25147 6335 25213 6343
rect 25147 6327 25171 6335
rect 25041 5483 25049 6327
rect 25163 5483 25171 6327
rect 25041 5475 25065 5483
rect 24999 5467 25065 5475
rect 25147 5475 25171 5483
rect 25189 6327 25213 6335
rect 25295 6335 25361 6343
rect 25295 6327 25319 6335
rect 25189 5483 25197 6327
rect 25311 5483 25319 6327
rect 25189 5475 25213 5483
rect 25147 5467 25213 5475
rect 25295 5475 25319 5483
rect 25337 6327 25361 6335
rect 25443 6335 25509 6343
rect 25443 6327 25467 6335
rect 25337 5483 25345 6327
rect 25459 5483 25467 6327
rect 25337 5475 25361 5483
rect 25295 5467 25361 5475
rect 25443 5475 25467 5483
rect 25485 6327 25509 6335
rect 25591 6335 25657 6343
rect 25591 6327 25615 6335
rect 25485 5483 25493 6327
rect 25607 5483 25615 6327
rect 25485 5475 25509 5483
rect 25443 5467 25509 5475
rect 25591 5475 25615 5483
rect 25633 6327 25657 6335
rect 25739 6335 25805 6343
rect 25739 6327 25763 6335
rect 25633 5483 25641 6327
rect 25755 5483 25763 6327
rect 25633 5475 25657 5483
rect 25591 5467 25657 5475
rect 25739 5475 25763 5483
rect 25781 6327 25805 6335
rect 25887 6335 25953 6343
rect 25887 6327 25911 6335
rect 25781 5483 25789 6327
rect 25903 5483 25911 6327
rect 25781 5475 25805 5483
rect 25739 5467 25805 5475
rect 25887 5475 25911 5483
rect 25929 6327 25953 6335
rect 26035 6335 26101 6343
rect 26035 6327 26059 6335
rect 25929 5483 25937 6327
rect 26051 5483 26059 6327
rect 25929 5475 25953 5483
rect 25887 5467 25953 5475
rect 26035 5475 26059 5483
rect 26077 6327 26101 6335
rect 26183 6335 26249 6343
rect 26183 6327 26207 6335
rect 26077 5483 26085 6327
rect 26199 5483 26207 6327
rect 26077 5475 26101 5483
rect 26035 5467 26101 5475
rect 26183 5475 26207 5483
rect 26225 6327 26249 6335
rect 26331 6335 26397 6343
rect 26331 6327 26355 6335
rect 26225 5483 26233 6327
rect 26347 5483 26355 6327
rect 26225 5475 26249 5483
rect 26183 5467 26249 5475
rect 26331 5475 26355 5483
rect 26373 6327 26397 6335
rect 26479 6335 26545 6343
rect 26479 6327 26503 6335
rect 26373 5483 26381 6327
rect 26495 5483 26503 6327
rect 26373 5475 26397 5483
rect 26331 5467 26397 5475
rect 26479 5475 26503 5483
rect 26521 6327 26545 6335
rect 26627 6335 26693 6343
rect 26627 6327 26651 6335
rect 26521 5483 26529 6327
rect 26643 5483 26651 6327
rect 26521 5475 26545 5483
rect 26479 5467 26545 5475
rect 26627 5475 26651 5483
rect 26669 6327 26693 6335
rect 26775 6335 26841 6343
rect 26775 6327 26799 6335
rect 26669 5483 26677 6327
rect 26791 5483 26799 6327
rect 26669 5475 26693 5483
rect 26627 5467 26693 5475
rect 26775 5475 26799 5483
rect 26817 6327 26841 6335
rect 26923 6335 26989 6343
rect 26923 6327 26947 6335
rect 26817 5483 26825 6327
rect 26939 5483 26947 6327
rect 26817 5475 26841 5483
rect 26775 5467 26841 5475
rect 26923 5475 26947 5483
rect 26965 6327 26989 6335
rect 27071 6335 27137 6343
rect 27071 6327 27095 6335
rect 26965 5483 26973 6327
rect 27087 5483 27095 6327
rect 26965 5475 26989 5483
rect 26923 5467 26989 5475
rect 27071 5475 27095 5483
rect 27113 6327 27137 6335
rect 27219 6335 27285 6343
rect 27219 6327 27243 6335
rect 27113 5483 27121 6327
rect 27235 5483 27243 6327
rect 27113 5475 27137 5483
rect 27071 5467 27137 5475
rect 27219 5475 27243 5483
rect 27261 6327 27285 6335
rect 27367 6335 27433 6343
rect 27367 6327 27391 6335
rect 27261 5483 27269 6327
rect 27383 5483 27391 6327
rect 27261 5475 27285 5483
rect 27219 5467 27285 5475
rect 27367 5475 27391 5483
rect 27409 6327 27433 6335
rect 27515 6335 27581 6343
rect 27515 6327 27539 6335
rect 27409 5483 27417 6327
rect 27531 5483 27539 6327
rect 27409 5475 27433 5483
rect 27367 5467 27433 5475
rect 27515 5475 27539 5483
rect 27557 6327 27581 6335
rect 27663 6335 27729 6343
rect 27663 6327 27687 6335
rect 27557 5483 27565 6327
rect 27679 5483 27687 6327
rect 27557 5475 27581 5483
rect 27515 5467 27581 5475
rect 27663 5475 27687 5483
rect 27705 6327 27729 6335
rect 27811 6335 27877 6343
rect 27811 6327 27835 6335
rect 27705 5483 27713 6327
rect 27827 5483 27835 6327
rect 27705 5475 27729 5483
rect 27663 5467 27729 5475
rect 27811 5475 27835 5483
rect 27853 6327 27877 6335
rect 27959 6335 28025 6343
rect 27959 6327 27983 6335
rect 27853 5483 27861 6327
rect 27975 5483 27983 6327
rect 27853 5475 27877 5483
rect 27811 5467 27877 5475
rect 27959 5475 27983 5483
rect 28001 6327 28025 6335
rect 28107 6335 28173 6343
rect 28107 6327 28131 6335
rect 28001 5483 28009 6327
rect 28123 5483 28131 6327
rect 28001 5475 28025 5483
rect 27959 5467 28025 5475
rect 28107 5475 28131 5483
rect 28149 6327 28173 6335
rect 28255 6335 28321 6343
rect 28255 6327 28279 6335
rect 28149 5483 28157 6327
rect 28271 5483 28279 6327
rect 28149 5475 28173 5483
rect 28107 5467 28173 5475
rect 28255 5475 28279 5483
rect 28297 6327 28321 6335
rect 28403 6335 28469 6343
rect 28403 6327 28427 6335
rect 28297 5483 28305 6327
rect 28419 5483 28427 6327
rect 28297 5475 28321 5483
rect 28255 5467 28321 5475
rect 28403 5475 28427 5483
rect 28445 6327 28469 6335
rect 28551 6335 28617 6343
rect 28551 6327 28575 6335
rect 28445 5483 28453 6327
rect 28567 5483 28575 6327
rect 28445 5475 28469 5483
rect 28403 5467 28469 5475
rect 28551 5475 28575 5483
rect 28593 6327 28617 6335
rect 28699 6335 28765 6343
rect 28699 6327 28723 6335
rect 28593 5483 28601 6327
rect 28715 5483 28723 6327
rect 28593 5475 28617 5483
rect 28551 5467 28617 5475
rect 28699 5475 28723 5483
rect 28741 6327 28765 6335
rect 28847 6335 28913 6343
rect 28847 6327 28871 6335
rect 28741 5483 28749 6327
rect 28863 5483 28871 6327
rect 28741 5475 28765 5483
rect 28699 5467 28765 5475
rect 28847 5475 28871 5483
rect 28889 6327 28913 6335
rect 28995 6335 29061 6343
rect 28995 6327 29019 6335
rect 28889 5483 28897 6327
rect 29011 5483 29019 6327
rect 28889 5475 28913 5483
rect 28847 5467 28913 5475
rect 28995 5475 29019 5483
rect 29037 6327 29061 6335
rect 29143 6335 29209 6343
rect 29143 6327 29167 6335
rect 29037 5483 29045 6327
rect 29159 5483 29167 6327
rect 29037 5475 29061 5483
rect 28995 5467 29061 5475
rect 29143 5475 29167 5483
rect 29185 6327 29209 6335
rect 29291 6335 29357 6343
rect 29291 6327 29315 6335
rect 29185 5483 29193 6327
rect 29307 5483 29315 6327
rect 29185 5475 29209 5483
rect 29143 5467 29209 5475
rect 29291 5475 29315 5483
rect 29333 6327 29357 6335
rect 29439 6335 29505 6343
rect 29439 6327 29463 6335
rect 29333 5483 29341 6327
rect 29455 5483 29463 6327
rect 29333 5475 29357 5483
rect 29291 5467 29357 5475
rect 29439 5475 29463 5483
rect 29481 6327 29505 6335
rect 29587 6335 29653 6343
rect 29587 6327 29611 6335
rect 29481 5483 29489 6327
rect 29603 5483 29611 6327
rect 29481 5475 29505 5483
rect 29439 5467 29505 5475
rect 29587 5475 29611 5483
rect 29629 6327 29653 6335
rect 29735 6335 29801 6343
rect 29735 6327 29759 6335
rect 29629 5483 29637 6327
rect 29751 5483 29759 6327
rect 29629 5475 29653 5483
rect 29587 5467 29653 5475
rect 29735 5475 29759 5483
rect 29777 6327 29801 6335
rect 29883 6335 29949 6343
rect 29883 6327 29907 6335
rect 29777 5483 29785 6327
rect 29899 5483 29907 6327
rect 29777 5475 29801 5483
rect 29735 5467 29801 5475
rect 29883 5475 29907 5483
rect 29925 6327 29949 6335
rect 30031 6335 30097 6343
rect 30031 6327 30055 6335
rect 29925 5483 29933 6327
rect 30047 5483 30055 6327
rect 29925 5475 29949 5483
rect 29883 5467 29949 5475
rect 30031 5475 30055 5483
rect 30073 6327 30097 6335
rect 30179 6335 30245 6343
rect 30179 6327 30203 6335
rect 30073 5483 30081 6327
rect 30195 5483 30203 6327
rect 30073 5475 30097 5483
rect 30031 5467 30097 5475
rect 30179 5475 30203 5483
rect 30221 6327 30245 6335
rect 30327 6335 30393 6343
rect 30327 6327 30351 6335
rect 30221 5483 30229 6327
rect 30343 5483 30351 6327
rect 30221 5475 30245 5483
rect 30179 5467 30245 5475
rect 30327 5475 30351 5483
rect 30369 6327 30393 6335
rect 30475 6335 30541 6343
rect 30475 6327 30499 6335
rect 30369 5483 30377 6327
rect 30491 5483 30499 6327
rect 30369 5475 30393 5483
rect 30327 5467 30393 5475
rect 30475 5475 30499 5483
rect 30517 6327 30541 6335
rect 30623 6335 30660 6343
rect 30623 6327 30647 6335
rect 30517 5483 30525 6327
rect 30639 5483 30647 6327
rect 30517 5475 30541 5483
rect 30475 5467 30541 5475
rect 30623 5475 30647 5483
rect 30623 5467 30660 5475
rect 22499 5451 22515 5467
rect 22517 5451 22533 5467
rect 22647 5451 22663 5467
rect 22665 5451 22681 5467
rect 22795 5451 22811 5467
rect 22813 5451 22829 5467
rect 22943 5451 22959 5467
rect 22961 5451 22977 5467
rect 23091 5451 23107 5467
rect 23109 5451 23125 5467
rect 23239 5451 23255 5467
rect 23257 5451 23273 5467
rect 23387 5451 23403 5467
rect 23405 5451 23421 5467
rect 23535 5451 23551 5467
rect 23553 5451 23569 5467
rect 23683 5451 23699 5467
rect 23701 5451 23717 5467
rect 23831 5451 23847 5467
rect 23849 5451 23865 5467
rect 23979 5451 23995 5467
rect 23997 5451 24013 5467
rect 24127 5451 24143 5467
rect 24145 5451 24161 5467
rect 24275 5451 24291 5467
rect 24293 5451 24309 5467
rect 24423 5451 24439 5467
rect 24441 5451 24457 5467
rect 24571 5451 24587 5467
rect 24589 5451 24605 5467
rect 24719 5451 24735 5467
rect 24737 5451 24753 5467
rect 24867 5451 24883 5467
rect 24885 5451 24901 5467
rect 25015 5451 25031 5467
rect 25033 5451 25049 5467
rect 25163 5451 25179 5467
rect 25181 5451 25197 5467
rect 25311 5451 25327 5467
rect 25329 5451 25345 5467
rect 25459 5451 25475 5467
rect 25477 5451 25493 5467
rect 25607 5451 25623 5467
rect 25625 5451 25641 5467
rect 25755 5451 25771 5467
rect 25773 5451 25789 5467
rect 25903 5451 25919 5467
rect 25921 5451 25937 5467
rect 26051 5451 26067 5467
rect 26069 5451 26085 5467
rect 26199 5451 26215 5467
rect 26217 5451 26233 5467
rect 26347 5451 26363 5467
rect 26365 5451 26381 5467
rect 26495 5451 26511 5467
rect 26513 5451 26529 5467
rect 26643 5451 26659 5467
rect 26661 5451 26677 5467
rect 26791 5451 26807 5467
rect 26809 5451 26825 5467
rect 26939 5451 26955 5467
rect 26957 5451 26973 5467
rect 27087 5451 27103 5467
rect 27105 5451 27121 5467
rect 27235 5451 27251 5467
rect 27253 5451 27269 5467
rect 27383 5451 27399 5467
rect 27401 5451 27417 5467
rect 27531 5451 27547 5467
rect 27549 5451 27565 5467
rect 27679 5451 27695 5467
rect 27697 5451 27713 5467
rect 27827 5451 27843 5467
rect 27845 5451 27861 5467
rect 27975 5451 27991 5467
rect 27993 5451 28009 5467
rect 28123 5451 28139 5467
rect 28141 5451 28157 5467
rect 28271 5451 28287 5467
rect 28289 5451 28305 5467
rect 28419 5451 28435 5467
rect 28437 5451 28453 5467
rect 28567 5451 28583 5467
rect 28585 5451 28601 5467
rect 28715 5451 28731 5467
rect 28733 5451 28749 5467
rect 28863 5451 28879 5467
rect 28881 5451 28897 5467
rect 29011 5451 29027 5467
rect 29029 5451 29045 5467
rect 29159 5451 29175 5467
rect 29177 5451 29193 5467
rect 29307 5451 29323 5467
rect 29325 5451 29341 5467
rect 29455 5451 29471 5467
rect 29473 5451 29489 5467
rect 29603 5451 29619 5467
rect 29621 5451 29637 5467
rect 29751 5451 29767 5467
rect 29769 5451 29785 5467
rect 29899 5451 29915 5467
rect 29917 5451 29933 5467
rect 30047 5451 30063 5467
rect 30065 5451 30081 5467
rect 30195 5451 30211 5467
rect 30213 5451 30229 5467
rect 30343 5451 30359 5467
rect 30361 5451 30377 5467
rect 30491 5451 30507 5467
rect 30509 5451 30525 5467
rect 30639 5451 30655 5467
rect 30657 5451 30660 5467
rect 23419 5433 23537 5447
rect 23419 5417 23433 5433
rect 23449 5417 23507 5425
rect 23449 5383 23463 5417
rect 23523 5383 23537 5433
rect 23567 5433 23685 5447
rect 23567 5417 23581 5433
rect 23597 5417 23655 5425
rect 23597 5383 23611 5417
rect 23671 5383 23685 5433
rect 23715 5433 23833 5447
rect 23715 5417 23729 5433
rect 23745 5417 23803 5425
rect 23745 5383 23759 5417
rect 23819 5383 23833 5433
rect 23863 5433 23981 5447
rect 23863 5417 23877 5433
rect 23893 5417 23951 5425
rect 23893 5383 23907 5417
rect 23967 5383 23981 5433
rect 24011 5433 24129 5447
rect 24011 5417 24025 5433
rect 24041 5417 24099 5425
rect 24041 5383 24055 5417
rect 24115 5383 24129 5433
rect 24159 5433 24277 5447
rect 24159 5417 24173 5433
rect 24189 5417 24247 5425
rect 24189 5383 24203 5417
rect 24263 5383 24277 5433
rect 27267 5433 27385 5447
rect 27267 5417 27281 5433
rect 27297 5417 27355 5425
rect 27297 5383 27311 5417
rect 27371 5383 27385 5433
rect 27415 5433 27533 5447
rect 27415 5417 27429 5433
rect 27445 5417 27503 5425
rect 27445 5383 27459 5417
rect 27519 5383 27533 5433
rect 27563 5433 27681 5447
rect 27563 5417 27577 5433
rect 27593 5417 27651 5425
rect 27593 5383 27607 5417
rect 27667 5383 27681 5433
rect 27711 5433 27829 5447
rect 27711 5417 27725 5433
rect 27741 5417 27799 5425
rect 27741 5383 27755 5417
rect 27815 5383 27829 5433
rect 27859 5433 27977 5447
rect 27859 5417 27873 5433
rect 27889 5417 27947 5425
rect 27889 5383 27903 5417
rect 27963 5383 27977 5433
rect 28599 5433 28717 5447
rect 28599 5417 28613 5433
rect 28629 5417 28687 5425
rect 28629 5383 28643 5417
rect 28703 5383 28717 5433
rect 28747 5433 28865 5447
rect 28747 5417 28761 5433
rect 28777 5417 28835 5425
rect 28777 5383 28791 5417
rect 28851 5383 28865 5433
rect 28895 5433 29013 5447
rect 28895 5417 28909 5433
rect 28925 5417 28983 5425
rect 28925 5383 28939 5417
rect 28999 5383 29013 5433
rect 29043 5433 29161 5447
rect 29043 5417 29057 5433
rect 29073 5417 29131 5425
rect 29073 5383 29087 5417
rect 29147 5383 29161 5433
rect 29191 5433 29309 5447
rect 29191 5417 29205 5433
rect 29221 5417 29279 5425
rect 29221 5383 29235 5417
rect 29295 5383 29309 5433
rect 29339 5433 29457 5447
rect 29339 5417 29353 5433
rect 29369 5417 29427 5425
rect 29369 5383 29383 5417
rect 29443 5383 29457 5433
rect 29487 5433 29605 5447
rect 29487 5417 29501 5433
rect 29517 5417 29575 5425
rect 29517 5383 29531 5417
rect 29591 5383 29605 5433
rect 29635 5433 29753 5447
rect 29635 5417 29649 5433
rect 29665 5417 29723 5425
rect 29665 5383 29679 5417
rect 29739 5383 29753 5433
rect 29783 5433 29901 5447
rect 29783 5417 29797 5433
rect 29813 5417 29871 5425
rect 29813 5383 29827 5417
rect 29887 5383 29901 5433
rect 29931 5433 30049 5447
rect 29931 5417 29945 5433
rect 29961 5417 30019 5425
rect 29961 5383 29975 5417
rect 30035 5383 30049 5433
rect 30079 5433 30197 5447
rect 30079 5417 30093 5433
rect 30109 5417 30167 5425
rect 30109 5383 30123 5417
rect 30183 5383 30197 5433
rect 30227 5433 30345 5447
rect 30227 5417 30241 5433
rect 30257 5417 30315 5425
rect 30257 5383 30271 5417
rect 30331 5383 30345 5433
rect 30375 5433 30493 5447
rect 30375 5417 30389 5433
rect 30405 5417 30463 5425
rect 30405 5383 30419 5417
rect 30479 5383 30493 5433
rect 30523 5433 30641 5447
rect 30523 5417 30537 5433
rect 30553 5417 30611 5425
rect 30553 5383 30567 5417
rect 30627 5383 30641 5433
rect 23419 5309 23433 5339
rect 23449 5309 23507 5317
rect 23449 5289 23463 5309
rect 23449 5275 23507 5289
rect 23523 5275 23537 5339
rect 23567 5309 23581 5339
rect 23597 5309 23655 5317
rect 23597 5289 23611 5309
rect 23597 5275 23655 5289
rect 23671 5275 23685 5339
rect 23715 5309 23729 5339
rect 23745 5309 23803 5317
rect 23745 5289 23759 5309
rect 23745 5275 23803 5289
rect 23819 5275 23833 5339
rect 23863 5309 23877 5339
rect 23893 5309 23951 5317
rect 23893 5289 23907 5309
rect 23893 5275 23951 5289
rect 23967 5275 23981 5339
rect 24011 5309 24025 5339
rect 24041 5309 24099 5317
rect 24041 5289 24055 5309
rect 24041 5275 24099 5289
rect 24115 5275 24129 5339
rect 24159 5309 24173 5339
rect 24189 5309 24247 5317
rect 24189 5289 24203 5309
rect 24189 5275 24247 5289
rect 24263 5275 24277 5339
rect 27267 5309 27281 5339
rect 27297 5309 27355 5317
rect 27297 5289 27311 5309
rect 27297 5275 27355 5289
rect 27371 5275 27385 5339
rect 27415 5309 27429 5339
rect 27445 5309 27503 5317
rect 27445 5289 27459 5309
rect 27445 5275 27503 5289
rect 27519 5275 27533 5339
rect 27563 5309 27577 5339
rect 27593 5309 27651 5317
rect 27593 5289 27607 5309
rect 27593 5275 27651 5289
rect 27667 5275 27681 5339
rect 27711 5309 27725 5339
rect 27741 5309 27799 5317
rect 27741 5289 27755 5309
rect 27741 5275 27799 5289
rect 27815 5275 27829 5339
rect 27859 5309 27873 5339
rect 27889 5309 27947 5317
rect 27889 5289 27903 5309
rect 27889 5275 27947 5289
rect 27963 5275 27977 5339
rect 28599 5309 28613 5339
rect 28629 5309 28687 5317
rect 28629 5289 28643 5309
rect 28629 5275 28687 5289
rect 28703 5275 28717 5339
rect 28747 5309 28761 5339
rect 28777 5309 28835 5317
rect 28777 5289 28791 5309
rect 28777 5275 28835 5289
rect 28851 5275 28865 5339
rect 28895 5309 28909 5339
rect 28925 5309 28983 5317
rect 28925 5289 28939 5309
rect 28925 5275 28983 5289
rect 28999 5275 29013 5339
rect 29043 5309 29057 5339
rect 29073 5309 29131 5317
rect 29073 5289 29087 5309
rect 29073 5275 29131 5289
rect 29147 5275 29161 5339
rect 29191 5309 29205 5339
rect 29221 5309 29279 5317
rect 29221 5289 29235 5309
rect 29221 5275 29279 5289
rect 29295 5275 29309 5339
rect 29339 5309 29353 5339
rect 29369 5309 29427 5317
rect 29369 5289 29383 5309
rect 29369 5275 29427 5289
rect 29443 5275 29457 5339
rect 29487 5309 29501 5339
rect 29517 5309 29575 5317
rect 29517 5289 29531 5309
rect 29517 5275 29575 5289
rect 29591 5275 29605 5339
rect 29635 5309 29649 5339
rect 29665 5309 29723 5317
rect 29665 5289 29679 5309
rect 29665 5275 29723 5289
rect 29739 5275 29753 5339
rect 29783 5309 29797 5339
rect 29813 5309 29871 5317
rect 29813 5289 29827 5309
rect 29813 5275 29871 5289
rect 29887 5275 29901 5339
rect 29931 5309 29945 5339
rect 29961 5309 30019 5317
rect 29961 5289 29975 5309
rect 29961 5275 30019 5289
rect 30035 5275 30049 5339
rect 30079 5309 30093 5339
rect 30109 5309 30167 5317
rect 30109 5289 30123 5309
rect 30109 5275 30167 5289
rect 30183 5275 30197 5339
rect 30227 5309 30241 5339
rect 30257 5309 30315 5317
rect 30257 5289 30271 5309
rect 30257 5275 30315 5289
rect 30331 5275 30345 5339
rect 30375 5309 30389 5339
rect 30405 5309 30463 5317
rect 30405 5289 30419 5309
rect 30405 5275 30463 5289
rect 30479 5275 30493 5339
rect 30523 5309 30537 5339
rect 30553 5309 30611 5317
rect 30553 5289 30567 5309
rect 30553 5275 30611 5289
rect 30627 5275 30641 5339
rect 30195 5225 30211 5241
rect 30213 5225 30229 5241
rect 30343 5225 30359 5241
rect 30361 5225 30377 5241
rect 30491 5225 30507 5241
rect 30509 5225 30525 5241
rect 30639 5225 30655 5241
rect 30657 5225 30660 5241
rect 30179 5217 30245 5225
rect 30179 5209 30203 5217
rect 30195 5170 30203 5209
rect 30221 5209 30245 5217
rect 30327 5217 30393 5225
rect 30327 5209 30351 5217
rect 30221 5170 30229 5209
rect 30343 5170 30351 5209
rect 30369 5209 30393 5217
rect 30475 5217 30541 5225
rect 30475 5209 30499 5217
rect 30369 5170 30377 5209
rect 30491 5170 30499 5209
rect 30517 5209 30541 5217
rect 30623 5217 30660 5225
rect 30623 5209 30647 5217
rect 30517 5170 30525 5209
rect 30639 5170 30647 5209
rect 12837 4703 12861 4708
rect 12895 4703 12933 4708
rect 12967 4703 13015 4708
rect 13049 4703 13087 4708
rect 13121 4703 13169 4708
rect 13203 4703 13241 4708
rect 13275 4703 13323 4708
rect 13357 4703 13395 4708
rect 13429 4703 13477 4708
rect 13511 4703 13549 4708
rect 13583 4703 13631 4708
rect 13665 4703 13703 4708
rect 13737 4703 13785 4708
rect 13819 4703 13857 4708
rect 13891 4703 13939 4708
rect 13973 4703 14011 4708
rect 14045 4703 14093 4708
rect 14127 4703 14165 4708
rect 14199 4703 14247 4708
rect 12837 4687 12877 4703
rect 12879 4687 12949 4703
rect 12951 4687 13031 4703
rect 13033 4687 13103 4703
rect 13105 4687 13185 4703
rect 13187 4687 13257 4703
rect 13259 4687 13339 4703
rect 13341 4687 13411 4703
rect 13413 4687 13493 4703
rect 13495 4687 13565 4703
rect 13567 4687 13647 4703
rect 13649 4687 13719 4703
rect 13721 4687 13801 4703
rect 13803 4687 13873 4703
rect 13875 4687 13955 4703
rect 13957 4687 14027 4703
rect 14029 4687 14109 4703
rect 14111 4687 14181 4703
rect 14183 4687 14260 4703
rect 12837 4682 14260 4687
rect 12845 4680 12911 4682
rect 12917 4680 12983 4682
rect 12999 4680 13065 4682
rect 13071 4680 13137 4682
rect 13153 4680 13219 4682
rect 13225 4680 13291 4682
rect 13307 4680 13373 4682
rect 13379 4680 13445 4682
rect 13461 4680 13527 4682
rect 13533 4680 13599 4682
rect 13615 4680 13681 4682
rect 13687 4680 13753 4682
rect 13769 4680 13835 4682
rect 13841 4680 13907 4682
rect 13923 4680 13989 4682
rect 13995 4680 14061 4682
rect 14077 4680 14143 4682
rect 14149 4680 14215 4682
rect 14231 4680 14260 4682
rect 12837 4654 14260 4680
rect 12845 4653 12911 4654
rect 12917 4653 12983 4654
rect 12999 4653 13065 4654
rect 13071 4653 13137 4654
rect 13153 4653 13219 4654
rect 13225 4653 13291 4654
rect 13307 4653 13373 4654
rect 13379 4653 13445 4654
rect 13461 4653 13527 4654
rect 13533 4653 13599 4654
rect 13615 4653 13681 4654
rect 13687 4653 13753 4654
rect 13769 4653 13835 4654
rect 13841 4653 13907 4654
rect 13923 4653 13989 4654
rect 13995 4653 14061 4654
rect 14077 4653 14143 4654
rect 14149 4653 14215 4654
rect 14231 4653 14260 4654
rect 12861 4637 12877 4653
rect 12879 4637 12895 4653
rect 12933 4637 12949 4653
rect 12951 4637 12967 4653
rect 13015 4637 13031 4653
rect 13033 4637 13049 4653
rect 13087 4637 13103 4653
rect 13105 4637 13121 4653
rect 13169 4637 13185 4653
rect 13187 4637 13203 4653
rect 13241 4637 13257 4653
rect 13259 4637 13275 4653
rect 13323 4637 13339 4653
rect 13341 4637 13357 4653
rect 13395 4637 13411 4653
rect 13413 4637 13429 4653
rect 13477 4637 13493 4653
rect 13495 4637 13511 4653
rect 13549 4637 13565 4653
rect 13567 4637 13583 4653
rect 13631 4637 13647 4653
rect 13649 4637 13665 4653
rect 13703 4637 13719 4653
rect 13721 4637 13737 4653
rect 13785 4637 13801 4653
rect 13803 4637 13819 4653
rect 13857 4637 13873 4653
rect 13875 4637 13891 4653
rect 13939 4637 13955 4653
rect 13957 4637 13973 4653
rect 14011 4637 14027 4653
rect 14029 4637 14045 4653
rect 14093 4637 14109 4653
rect 14111 4637 14127 4653
rect 14165 4637 14181 4653
rect 14183 4637 14199 4653
rect 14247 4637 14260 4653
rect 12861 4613 12877 4629
rect 12879 4613 12895 4629
rect 12933 4613 12949 4629
rect 12951 4613 12967 4629
rect 13015 4613 13031 4629
rect 13033 4613 13049 4629
rect 13087 4613 13103 4629
rect 13105 4613 13121 4629
rect 13169 4613 13185 4629
rect 13187 4613 13203 4629
rect 13241 4613 13257 4629
rect 13259 4613 13275 4629
rect 13323 4613 13339 4629
rect 13341 4613 13357 4629
rect 13395 4613 13411 4629
rect 13413 4613 13429 4629
rect 13477 4613 13493 4629
rect 13495 4613 13511 4629
rect 13549 4613 13565 4629
rect 13567 4613 13583 4629
rect 13631 4613 13647 4629
rect 13649 4613 13665 4629
rect 13703 4613 13719 4629
rect 13721 4613 13737 4629
rect 13785 4613 13801 4629
rect 13803 4613 13819 4629
rect 13857 4613 13873 4629
rect 13875 4613 13891 4629
rect 13939 4613 13955 4629
rect 13957 4613 13973 4629
rect 14011 4613 14027 4629
rect 14029 4613 14045 4629
rect 14093 4613 14109 4629
rect 14111 4613 14127 4629
rect 14165 4613 14181 4629
rect 14183 4613 14199 4629
rect 14247 4613 14260 4629
rect 12845 4597 12911 4613
rect 12917 4597 12983 4613
rect 12999 4597 13065 4613
rect 13071 4597 13137 4613
rect 13153 4597 13219 4613
rect 13225 4597 13291 4613
rect 13307 4597 13373 4613
rect 13379 4597 13445 4613
rect 13461 4597 13527 4613
rect 13533 4597 13599 4613
rect 13615 4597 13681 4613
rect 13687 4597 13753 4613
rect 13769 4597 13835 4613
rect 13841 4597 13907 4613
rect 13923 4597 13989 4613
rect 13995 4597 14061 4613
rect 14077 4597 14143 4613
rect 14149 4597 14215 4613
rect 14231 4597 14260 4613
rect 12861 4595 12895 4597
rect 12933 4595 12967 4597
rect 13015 4595 13049 4597
rect 13087 4595 13121 4597
rect 13169 4595 13203 4597
rect 13241 4595 13275 4597
rect 13323 4595 13357 4597
rect 13395 4595 13429 4597
rect 13477 4595 13511 4597
rect 13549 4595 13583 4597
rect 13631 4595 13665 4597
rect 13703 4595 13737 4597
rect 13785 4595 13819 4597
rect 13857 4595 13891 4597
rect 13939 4595 13973 4597
rect 14011 4595 14045 4597
rect 14093 4595 14127 4597
rect 14165 4595 14199 4597
rect 14247 4595 14260 4597
rect 12845 4579 12911 4595
rect 12917 4579 12983 4595
rect 12999 4579 13065 4595
rect 13071 4579 13137 4595
rect 13153 4579 13219 4595
rect 13225 4579 13291 4595
rect 13307 4579 13373 4595
rect 13379 4579 13445 4595
rect 13461 4579 13527 4595
rect 13533 4579 13599 4595
rect 13615 4579 13681 4595
rect 13687 4579 13753 4595
rect 13769 4579 13835 4595
rect 13841 4579 13907 4595
rect 13923 4579 13989 4595
rect 13995 4579 14061 4595
rect 14077 4579 14143 4595
rect 14149 4579 14215 4595
rect 14231 4579 14260 4595
rect 12861 4563 12877 4579
rect 12879 4563 12895 4579
rect 12933 4563 12949 4579
rect 12951 4563 12967 4579
rect 13015 4563 13031 4579
rect 13033 4563 13049 4579
rect 13087 4563 13103 4579
rect 13105 4563 13121 4579
rect 13169 4563 13185 4579
rect 13187 4563 13203 4579
rect 13241 4563 13257 4579
rect 13259 4563 13275 4579
rect 13323 4563 13339 4579
rect 13341 4563 13357 4579
rect 13395 4563 13411 4579
rect 13413 4563 13429 4579
rect 13477 4563 13493 4579
rect 13495 4563 13511 4579
rect 13549 4563 13565 4579
rect 13567 4563 13583 4579
rect 13631 4563 13647 4579
rect 13649 4563 13665 4579
rect 13703 4563 13719 4579
rect 13721 4563 13737 4579
rect 13785 4563 13801 4579
rect 13803 4563 13819 4579
rect 13857 4563 13873 4579
rect 13875 4563 13891 4579
rect 13939 4563 13955 4579
rect 13957 4563 13973 4579
rect 14011 4563 14027 4579
rect 14029 4563 14045 4579
rect 14093 4563 14109 4579
rect 14111 4563 14127 4579
rect 14165 4563 14181 4579
rect 14183 4563 14199 4579
rect 14247 4563 14260 4579
rect 12861 4539 12877 4555
rect 12879 4539 12895 4555
rect 12933 4539 12949 4555
rect 12951 4539 12967 4555
rect 13015 4539 13031 4555
rect 13033 4539 13049 4555
rect 13087 4539 13103 4555
rect 13105 4539 13121 4555
rect 13169 4539 13185 4555
rect 13187 4539 13203 4555
rect 13241 4539 13257 4555
rect 13259 4539 13275 4555
rect 13323 4539 13339 4555
rect 13341 4539 13357 4555
rect 13395 4539 13411 4555
rect 13413 4539 13429 4555
rect 13477 4539 13493 4555
rect 13495 4539 13511 4555
rect 13549 4539 13565 4555
rect 13567 4539 13583 4555
rect 13631 4539 13647 4555
rect 13649 4539 13665 4555
rect 13703 4539 13719 4555
rect 13721 4539 13737 4555
rect 13785 4539 13801 4555
rect 13803 4539 13819 4555
rect 13857 4539 13873 4555
rect 13875 4539 13891 4555
rect 13939 4539 13955 4555
rect 13957 4539 13973 4555
rect 14011 4539 14027 4555
rect 14029 4539 14045 4555
rect 14093 4539 14109 4555
rect 14111 4539 14127 4555
rect 14165 4539 14181 4555
rect 14183 4539 14199 4555
rect 14247 4539 14260 4555
rect 12845 4523 12911 4539
rect 12917 4523 12983 4539
rect 12999 4523 13065 4539
rect 13071 4523 13137 4539
rect 13153 4523 13219 4539
rect 13225 4523 13291 4539
rect 13307 4523 13373 4539
rect 13379 4523 13445 4539
rect 13461 4523 13527 4539
rect 13533 4523 13599 4539
rect 13615 4523 13681 4539
rect 13687 4523 13753 4539
rect 13769 4523 13835 4539
rect 13841 4523 13907 4539
rect 13923 4523 13989 4539
rect 13995 4523 14061 4539
rect 14077 4523 14143 4539
rect 14149 4523 14215 4539
rect 14231 4523 14260 4539
rect 12861 4521 12895 4523
rect 12933 4521 12967 4523
rect 13015 4521 13049 4523
rect 13087 4521 13121 4523
rect 13169 4521 13203 4523
rect 13241 4521 13275 4523
rect 13323 4521 13357 4523
rect 13395 4521 13429 4523
rect 13477 4521 13511 4523
rect 13549 4521 13583 4523
rect 13631 4521 13665 4523
rect 13703 4521 13737 4523
rect 13785 4521 13819 4523
rect 13857 4521 13891 4523
rect 13939 4521 13973 4523
rect 14011 4521 14045 4523
rect 14093 4521 14127 4523
rect 14165 4521 14199 4523
rect 14247 4521 14260 4523
rect 12845 4505 12911 4521
rect 12917 4505 12983 4521
rect 12999 4505 13065 4521
rect 13071 4505 13137 4521
rect 13153 4505 13219 4521
rect 13225 4505 13291 4521
rect 13307 4505 13373 4521
rect 13379 4505 13445 4521
rect 13461 4505 13527 4521
rect 13533 4505 13599 4521
rect 13615 4505 13681 4521
rect 13687 4505 13753 4521
rect 13769 4505 13835 4521
rect 13841 4505 13907 4521
rect 13923 4505 13989 4521
rect 13995 4505 14061 4521
rect 14077 4505 14143 4521
rect 14149 4505 14215 4521
rect 14231 4505 14260 4521
rect 12861 4489 12877 4505
rect 12879 4489 12895 4505
rect 12933 4489 12949 4505
rect 12951 4489 12967 4505
rect 13015 4489 13031 4505
rect 13033 4489 13049 4505
rect 13087 4489 13103 4505
rect 13105 4489 13121 4505
rect 13169 4489 13185 4505
rect 13187 4489 13203 4505
rect 13241 4489 13257 4505
rect 13259 4489 13275 4505
rect 13323 4489 13339 4505
rect 13341 4489 13357 4505
rect 13395 4489 13411 4505
rect 13413 4489 13429 4505
rect 13477 4489 13493 4505
rect 13495 4489 13511 4505
rect 13549 4489 13565 4505
rect 13567 4489 13583 4505
rect 13631 4489 13647 4505
rect 13649 4489 13665 4505
rect 13703 4489 13719 4505
rect 13721 4489 13737 4505
rect 13785 4489 13801 4505
rect 13803 4489 13819 4505
rect 13857 4489 13873 4505
rect 13875 4489 13891 4505
rect 13939 4489 13955 4505
rect 13957 4489 13973 4505
rect 14011 4489 14027 4505
rect 14029 4489 14045 4505
rect 14093 4489 14109 4505
rect 14111 4489 14127 4505
rect 14165 4489 14181 4505
rect 14183 4489 14199 4505
rect 14247 4489 14260 4505
rect 12861 4465 12877 4481
rect 12879 4465 12895 4481
rect 12933 4465 12949 4481
rect 12951 4465 12967 4481
rect 13015 4465 13031 4481
rect 13033 4465 13049 4481
rect 13087 4465 13103 4481
rect 13105 4465 13121 4481
rect 13169 4465 13185 4481
rect 13187 4465 13203 4481
rect 13241 4465 13257 4481
rect 13259 4465 13275 4481
rect 13323 4465 13339 4481
rect 13341 4465 13357 4481
rect 13395 4465 13411 4481
rect 13413 4465 13429 4481
rect 13477 4465 13493 4481
rect 13495 4465 13511 4481
rect 13549 4465 13565 4481
rect 13567 4465 13583 4481
rect 13631 4465 13647 4481
rect 13649 4465 13665 4481
rect 13703 4465 13719 4481
rect 13721 4465 13737 4481
rect 13785 4465 13801 4481
rect 13803 4465 13819 4481
rect 13857 4465 13873 4481
rect 13875 4465 13891 4481
rect 13939 4465 13955 4481
rect 13957 4465 13973 4481
rect 14011 4465 14027 4481
rect 14029 4465 14045 4481
rect 14093 4465 14109 4481
rect 14111 4465 14127 4481
rect 14165 4465 14181 4481
rect 14183 4465 14199 4481
rect 14247 4465 14260 4481
rect 12845 4449 12911 4465
rect 12917 4449 12983 4465
rect 12999 4449 13065 4465
rect 13071 4449 13137 4465
rect 13153 4449 13219 4465
rect 13225 4449 13291 4465
rect 13307 4449 13373 4465
rect 13379 4449 13445 4465
rect 13461 4449 13527 4465
rect 13533 4449 13599 4465
rect 13615 4449 13681 4465
rect 13687 4449 13753 4465
rect 13769 4449 13835 4465
rect 13841 4449 13907 4465
rect 13923 4449 13989 4465
rect 13995 4449 14061 4465
rect 14077 4449 14143 4465
rect 14149 4449 14215 4465
rect 14231 4449 14260 4465
rect 12861 4447 12895 4449
rect 12933 4447 12967 4449
rect 13015 4447 13049 4449
rect 13087 4447 13121 4449
rect 13169 4447 13203 4449
rect 13241 4447 13275 4449
rect 13323 4447 13357 4449
rect 13395 4447 13429 4449
rect 13477 4447 13511 4449
rect 13549 4447 13583 4449
rect 13631 4447 13665 4449
rect 13703 4447 13737 4449
rect 13785 4447 13819 4449
rect 13857 4447 13891 4449
rect 13939 4447 13973 4449
rect 14011 4447 14045 4449
rect 14093 4447 14127 4449
rect 14165 4447 14199 4449
rect 14247 4447 14260 4449
rect 12845 4431 12911 4447
rect 12917 4431 12983 4447
rect 12999 4431 13065 4447
rect 13071 4431 13137 4447
rect 13153 4431 13219 4447
rect 13225 4431 13291 4447
rect 13307 4431 13373 4447
rect 13379 4431 13445 4447
rect 13461 4431 13527 4447
rect 13533 4431 13599 4447
rect 13615 4431 13681 4447
rect 13687 4431 13753 4447
rect 13769 4431 13835 4447
rect 13841 4431 13907 4447
rect 13923 4431 13989 4447
rect 13995 4431 14061 4447
rect 14077 4431 14143 4447
rect 14149 4431 14215 4447
rect 14231 4431 14260 4447
rect 12861 4415 12877 4431
rect 12879 4415 12895 4431
rect 12933 4415 12949 4431
rect 12951 4415 12967 4431
rect 13015 4415 13031 4431
rect 13033 4415 13049 4431
rect 13087 4415 13103 4431
rect 13105 4415 13121 4431
rect 13169 4415 13185 4431
rect 13187 4415 13203 4431
rect 13241 4415 13257 4431
rect 13259 4415 13275 4431
rect 13323 4415 13339 4431
rect 13341 4415 13357 4431
rect 13395 4415 13411 4431
rect 13413 4415 13429 4431
rect 13477 4415 13493 4431
rect 13495 4415 13511 4431
rect 13549 4415 13565 4431
rect 13567 4415 13583 4431
rect 13631 4415 13647 4431
rect 13649 4415 13665 4431
rect 13703 4415 13719 4431
rect 13721 4415 13737 4431
rect 13785 4415 13801 4431
rect 13803 4415 13819 4431
rect 13857 4415 13873 4431
rect 13875 4415 13891 4431
rect 13939 4415 13955 4431
rect 13957 4415 13973 4431
rect 14011 4415 14027 4431
rect 14029 4415 14045 4431
rect 14093 4415 14109 4431
rect 14111 4415 14127 4431
rect 14165 4415 14181 4431
rect 14183 4415 14199 4431
rect 14247 4415 14260 4431
rect 12861 4391 12877 4407
rect 12879 4391 12895 4407
rect 12933 4391 12949 4407
rect 12951 4391 12967 4407
rect 13015 4391 13031 4407
rect 13033 4391 13049 4407
rect 13087 4391 13103 4407
rect 13105 4391 13121 4407
rect 13169 4391 13185 4407
rect 13187 4391 13203 4407
rect 13241 4391 13257 4407
rect 13259 4391 13275 4407
rect 13323 4391 13339 4407
rect 13341 4391 13357 4407
rect 13395 4391 13411 4407
rect 13413 4391 13429 4407
rect 13477 4391 13493 4407
rect 13495 4391 13511 4407
rect 13549 4391 13565 4407
rect 13567 4391 13583 4407
rect 13631 4391 13647 4407
rect 13649 4391 13665 4407
rect 13703 4391 13719 4407
rect 13721 4391 13737 4407
rect 13785 4391 13801 4407
rect 13803 4391 13819 4407
rect 13857 4391 13873 4407
rect 13875 4391 13891 4407
rect 13939 4391 13955 4407
rect 13957 4391 13973 4407
rect 14011 4391 14027 4407
rect 14029 4391 14045 4407
rect 14093 4391 14109 4407
rect 14111 4391 14127 4407
rect 14165 4391 14181 4407
rect 14183 4391 14199 4407
rect 14247 4391 14260 4407
rect 12845 4375 12911 4391
rect 12917 4375 12983 4391
rect 12999 4375 13065 4391
rect 13071 4375 13137 4391
rect 13153 4375 13219 4391
rect 13225 4375 13291 4391
rect 13307 4375 13373 4391
rect 13379 4375 13445 4391
rect 13461 4375 13527 4391
rect 13533 4375 13599 4391
rect 13615 4375 13681 4391
rect 13687 4375 13753 4391
rect 13769 4375 13835 4391
rect 13841 4375 13907 4391
rect 13923 4375 13989 4391
rect 13995 4375 14061 4391
rect 14077 4375 14143 4391
rect 14149 4375 14215 4391
rect 14231 4375 14260 4391
rect 12861 4373 12895 4375
rect 12933 4373 12967 4375
rect 13015 4373 13049 4375
rect 13087 4373 13121 4375
rect 13169 4373 13203 4375
rect 13241 4373 13275 4375
rect 13323 4373 13357 4375
rect 13395 4373 13429 4375
rect 13477 4373 13511 4375
rect 13549 4373 13583 4375
rect 13631 4373 13665 4375
rect 13703 4373 13737 4375
rect 13785 4373 13819 4375
rect 13857 4373 13891 4375
rect 13939 4373 13973 4375
rect 14011 4373 14045 4375
rect 14093 4373 14127 4375
rect 14165 4373 14199 4375
rect 14247 4373 14260 4375
rect 12845 4357 12911 4373
rect 12917 4357 12983 4373
rect 12999 4357 13065 4373
rect 13071 4357 13137 4373
rect 13153 4357 13219 4373
rect 13225 4357 13291 4373
rect 13307 4357 13373 4373
rect 13379 4357 13445 4373
rect 13461 4357 13527 4373
rect 13533 4357 13599 4373
rect 13615 4357 13681 4373
rect 13687 4357 13753 4373
rect 13769 4357 13835 4373
rect 13841 4357 13907 4373
rect 13923 4357 13989 4373
rect 13995 4357 14061 4373
rect 14077 4357 14143 4373
rect 14149 4357 14215 4373
rect 14231 4357 14260 4373
rect 12861 4341 12877 4357
rect 12879 4341 12895 4357
rect 12933 4341 12949 4357
rect 12951 4341 12967 4357
rect 13015 4341 13031 4357
rect 13033 4341 13049 4357
rect 13087 4341 13103 4357
rect 13105 4341 13121 4357
rect 13169 4341 13185 4357
rect 13187 4341 13203 4357
rect 13241 4341 13257 4357
rect 13259 4341 13275 4357
rect 13323 4341 13339 4357
rect 13341 4341 13357 4357
rect 13395 4341 13411 4357
rect 13413 4341 13429 4357
rect 13477 4341 13493 4357
rect 13495 4341 13511 4357
rect 13549 4341 13565 4357
rect 13567 4341 13583 4357
rect 13631 4341 13647 4357
rect 13649 4341 13665 4357
rect 13703 4341 13719 4357
rect 13721 4341 13737 4357
rect 13785 4341 13801 4357
rect 13803 4341 13819 4357
rect 13857 4341 13873 4357
rect 13875 4341 13891 4357
rect 13939 4341 13955 4357
rect 13957 4341 13973 4357
rect 14011 4341 14027 4357
rect 14029 4341 14045 4357
rect 14093 4341 14109 4357
rect 14111 4341 14127 4357
rect 14165 4341 14181 4357
rect 14183 4341 14199 4357
rect 14247 4341 14260 4357
rect 12861 4317 12877 4333
rect 12879 4317 12895 4333
rect 12933 4317 12949 4333
rect 12951 4317 12967 4333
rect 13015 4317 13031 4333
rect 13033 4317 13049 4333
rect 13087 4317 13103 4333
rect 13105 4317 13121 4333
rect 13169 4317 13185 4333
rect 13187 4317 13203 4333
rect 13241 4317 13257 4333
rect 13259 4317 13275 4333
rect 13323 4317 13339 4333
rect 13341 4317 13357 4333
rect 13395 4317 13411 4333
rect 13413 4317 13429 4333
rect 13477 4317 13493 4333
rect 13495 4317 13511 4333
rect 13549 4317 13565 4333
rect 13567 4317 13583 4333
rect 13631 4317 13647 4333
rect 13649 4317 13665 4333
rect 13703 4317 13719 4333
rect 13721 4317 13737 4333
rect 13785 4317 13801 4333
rect 13803 4317 13819 4333
rect 13857 4317 13873 4333
rect 13875 4317 13891 4333
rect 13939 4317 13955 4333
rect 13957 4317 13973 4333
rect 14011 4317 14027 4333
rect 14029 4317 14045 4333
rect 14093 4317 14109 4333
rect 14111 4317 14127 4333
rect 14165 4317 14181 4333
rect 14183 4317 14199 4333
rect 14247 4317 14260 4333
rect 12845 4301 12911 4317
rect 12917 4301 12983 4317
rect 12999 4301 13065 4317
rect 13071 4301 13137 4317
rect 13153 4301 13219 4317
rect 13225 4301 13291 4317
rect 13307 4301 13373 4317
rect 13379 4301 13445 4317
rect 13461 4301 13527 4317
rect 13533 4301 13599 4317
rect 13615 4301 13681 4317
rect 13687 4301 13753 4317
rect 13769 4301 13835 4317
rect 13841 4301 13907 4317
rect 13923 4301 13989 4317
rect 13995 4301 14061 4317
rect 14077 4301 14143 4317
rect 14149 4301 14215 4317
rect 14231 4301 14260 4317
rect 12861 4299 12895 4301
rect 12933 4299 12967 4301
rect 13015 4299 13049 4301
rect 13087 4299 13121 4301
rect 13169 4299 13203 4301
rect 13241 4299 13275 4301
rect 13323 4299 13357 4301
rect 13395 4299 13429 4301
rect 13477 4299 13511 4301
rect 13549 4299 13583 4301
rect 13631 4299 13665 4301
rect 13703 4299 13737 4301
rect 13785 4299 13819 4301
rect 13857 4299 13891 4301
rect 13939 4299 13973 4301
rect 14011 4299 14045 4301
rect 14093 4299 14127 4301
rect 14165 4299 14199 4301
rect 14247 4299 14260 4301
rect 12845 4283 12911 4299
rect 12917 4283 12983 4299
rect 12999 4283 13065 4299
rect 13071 4283 13137 4299
rect 13153 4283 13219 4299
rect 13225 4283 13291 4299
rect 13307 4283 13373 4299
rect 13379 4283 13445 4299
rect 13461 4283 13527 4299
rect 13533 4283 13599 4299
rect 13615 4283 13681 4299
rect 13687 4283 13753 4299
rect 13769 4283 13835 4299
rect 13841 4283 13907 4299
rect 13923 4283 13989 4299
rect 13995 4283 14061 4299
rect 14077 4283 14143 4299
rect 14149 4283 14215 4299
rect 14231 4283 14260 4299
rect 12861 4267 12877 4283
rect 12879 4267 12895 4283
rect 12933 4267 12949 4283
rect 12951 4267 12967 4283
rect 13015 4267 13031 4283
rect 13033 4267 13049 4283
rect 13087 4267 13103 4283
rect 13105 4267 13121 4283
rect 13169 4267 13185 4283
rect 13187 4267 13203 4283
rect 13241 4267 13257 4283
rect 13259 4267 13275 4283
rect 13323 4267 13339 4283
rect 13341 4267 13357 4283
rect 13395 4267 13411 4283
rect 13413 4267 13429 4283
rect 13477 4267 13493 4283
rect 13495 4267 13511 4283
rect 13549 4267 13565 4283
rect 13567 4267 13583 4283
rect 13631 4267 13647 4283
rect 13649 4267 13665 4283
rect 13703 4267 13719 4283
rect 13721 4267 13737 4283
rect 13785 4267 13801 4283
rect 13803 4267 13819 4283
rect 13857 4267 13873 4283
rect 13875 4267 13891 4283
rect 13939 4267 13955 4283
rect 13957 4267 13973 4283
rect 14011 4267 14027 4283
rect 14029 4267 14045 4283
rect 14093 4267 14109 4283
rect 14111 4267 14127 4283
rect 14165 4267 14181 4283
rect 14183 4267 14199 4283
rect 14247 4267 14260 4283
rect 12861 4243 12877 4259
rect 12879 4243 12895 4259
rect 12933 4243 12949 4259
rect 12951 4243 12967 4259
rect 13015 4243 13031 4259
rect 13033 4243 13049 4259
rect 13087 4243 13103 4259
rect 13105 4243 13121 4259
rect 13169 4243 13185 4259
rect 13187 4243 13203 4259
rect 13241 4243 13257 4259
rect 13259 4243 13275 4259
rect 13323 4243 13339 4259
rect 13341 4243 13357 4259
rect 13395 4243 13411 4259
rect 13413 4243 13429 4259
rect 13477 4243 13493 4259
rect 13495 4243 13511 4259
rect 13549 4243 13565 4259
rect 13567 4243 13583 4259
rect 13631 4243 13647 4259
rect 13649 4243 13665 4259
rect 13703 4243 13719 4259
rect 13721 4243 13737 4259
rect 13785 4243 13801 4259
rect 13803 4243 13819 4259
rect 13857 4243 13873 4259
rect 13875 4243 13891 4259
rect 13939 4243 13955 4259
rect 13957 4243 13973 4259
rect 14011 4243 14027 4259
rect 14029 4243 14045 4259
rect 14093 4243 14109 4259
rect 14111 4243 14127 4259
rect 14165 4243 14181 4259
rect 14183 4243 14199 4259
rect 14247 4243 14260 4259
rect 12845 4227 12911 4243
rect 12917 4227 12983 4243
rect 12999 4227 13065 4243
rect 13071 4227 13137 4243
rect 13153 4227 13219 4243
rect 13225 4227 13291 4243
rect 13307 4227 13373 4243
rect 13379 4227 13445 4243
rect 13461 4227 13527 4243
rect 13533 4227 13599 4243
rect 13615 4227 13681 4243
rect 13687 4227 13753 4243
rect 13769 4227 13835 4243
rect 13841 4227 13907 4243
rect 13923 4227 13989 4243
rect 13995 4227 14061 4243
rect 14077 4227 14143 4243
rect 14149 4227 14215 4243
rect 14231 4227 14260 4243
rect 12861 4225 12895 4227
rect 12933 4225 12967 4227
rect 13015 4225 13049 4227
rect 13087 4225 13121 4227
rect 13169 4225 13203 4227
rect 13241 4225 13275 4227
rect 13323 4225 13357 4227
rect 13395 4225 13429 4227
rect 13477 4225 13511 4227
rect 13549 4225 13583 4227
rect 13631 4225 13665 4227
rect 13703 4225 13737 4227
rect 13785 4225 13819 4227
rect 13857 4225 13891 4227
rect 13939 4225 13973 4227
rect 14011 4225 14045 4227
rect 14093 4225 14127 4227
rect 14165 4225 14199 4227
rect 14247 4225 14260 4227
rect 12845 4209 12911 4225
rect 12917 4209 12983 4225
rect 12999 4209 13065 4225
rect 13071 4209 13137 4225
rect 13153 4209 13219 4225
rect 13225 4209 13291 4225
rect 13307 4209 13373 4225
rect 13379 4209 13445 4225
rect 13461 4209 13527 4225
rect 13533 4209 13599 4225
rect 13615 4209 13681 4225
rect 13687 4209 13753 4225
rect 13769 4209 13835 4225
rect 13841 4209 13907 4225
rect 13923 4209 13989 4225
rect 13995 4209 14061 4225
rect 14077 4209 14143 4225
rect 14149 4209 14215 4225
rect 14231 4209 14260 4225
rect 12861 4193 12877 4209
rect 12879 4193 12895 4209
rect 12933 4193 12949 4209
rect 12951 4193 12967 4209
rect 13015 4193 13031 4209
rect 13033 4193 13049 4209
rect 13087 4193 13103 4209
rect 13105 4193 13121 4209
rect 13169 4193 13185 4209
rect 13187 4193 13203 4209
rect 13241 4193 13257 4209
rect 13259 4193 13275 4209
rect 13323 4193 13339 4209
rect 13341 4193 13357 4209
rect 13395 4193 13411 4209
rect 13413 4193 13429 4209
rect 13477 4193 13493 4209
rect 13495 4193 13511 4209
rect 13549 4193 13565 4209
rect 13567 4193 13583 4209
rect 13631 4193 13647 4209
rect 13649 4193 13665 4209
rect 13703 4193 13719 4209
rect 13721 4193 13737 4209
rect 13785 4193 13801 4209
rect 13803 4193 13819 4209
rect 13857 4193 13873 4209
rect 13875 4193 13891 4209
rect 13939 4193 13955 4209
rect 13957 4193 13973 4209
rect 14011 4193 14027 4209
rect 14029 4193 14045 4209
rect 14093 4193 14109 4209
rect 14111 4193 14127 4209
rect 14165 4193 14181 4209
rect 14183 4193 14199 4209
rect 14247 4193 14260 4209
rect 12861 4169 12877 4185
rect 12879 4169 12895 4185
rect 12933 4169 12949 4185
rect 12951 4169 12967 4185
rect 13015 4169 13031 4185
rect 13033 4169 13049 4185
rect 13087 4169 13103 4185
rect 13105 4169 13121 4185
rect 13169 4169 13185 4185
rect 13187 4169 13203 4185
rect 13241 4169 13257 4185
rect 13259 4169 13275 4185
rect 13323 4169 13339 4185
rect 13341 4169 13357 4185
rect 13395 4169 13411 4185
rect 13413 4169 13429 4185
rect 13477 4169 13493 4185
rect 13495 4169 13511 4185
rect 13549 4169 13565 4185
rect 13567 4169 13583 4185
rect 13631 4169 13647 4185
rect 13649 4169 13665 4185
rect 13703 4169 13719 4185
rect 13721 4169 13737 4185
rect 13785 4169 13801 4185
rect 13803 4169 13819 4185
rect 13857 4169 13873 4185
rect 13875 4169 13891 4185
rect 13939 4169 13955 4185
rect 13957 4169 13973 4185
rect 14011 4169 14027 4185
rect 14029 4169 14045 4185
rect 14093 4169 14109 4185
rect 14111 4169 14127 4185
rect 14165 4169 14181 4185
rect 14183 4169 14199 4185
rect 14247 4169 14260 4185
rect 12845 4153 12911 4169
rect 12917 4153 12983 4169
rect 12999 4153 13065 4169
rect 13071 4153 13137 4169
rect 13153 4153 13219 4169
rect 13225 4153 13291 4169
rect 13307 4153 13373 4169
rect 13379 4153 13445 4169
rect 13461 4153 13527 4169
rect 13533 4153 13599 4169
rect 13615 4153 13681 4169
rect 13687 4153 13753 4169
rect 13769 4153 13835 4169
rect 13841 4153 13907 4169
rect 13923 4153 13989 4169
rect 13995 4153 14061 4169
rect 14077 4153 14143 4169
rect 14149 4153 14215 4169
rect 14231 4153 14260 4169
rect 12861 4151 12895 4153
rect 12933 4151 12967 4153
rect 13015 4151 13049 4153
rect 13087 4151 13121 4153
rect 13169 4151 13203 4153
rect 13241 4151 13275 4153
rect 13323 4151 13357 4153
rect 13395 4151 13429 4153
rect 13477 4151 13511 4153
rect 13549 4151 13583 4153
rect 13631 4151 13665 4153
rect 13703 4151 13737 4153
rect 13785 4151 13819 4153
rect 13857 4151 13891 4153
rect 13939 4151 13973 4153
rect 14011 4151 14045 4153
rect 14093 4151 14127 4153
rect 14165 4151 14199 4153
rect 14247 4151 14260 4153
rect 12845 4135 12911 4151
rect 12917 4135 12983 4151
rect 12999 4135 13065 4151
rect 13071 4135 13137 4151
rect 13153 4135 13219 4151
rect 13225 4135 13291 4151
rect 13307 4135 13373 4151
rect 13379 4135 13445 4151
rect 13461 4135 13527 4151
rect 13533 4135 13599 4151
rect 13615 4135 13681 4151
rect 13687 4135 13753 4151
rect 13769 4135 13835 4151
rect 13841 4135 13907 4151
rect 13923 4135 13989 4151
rect 13995 4135 14061 4151
rect 14077 4135 14143 4151
rect 14149 4135 14215 4151
rect 14231 4135 14260 4151
rect 12861 4119 12877 4135
rect 12879 4119 12895 4135
rect 12933 4119 12949 4135
rect 12951 4119 12967 4135
rect 13015 4119 13031 4135
rect 13033 4119 13049 4135
rect 13087 4119 13103 4135
rect 13105 4119 13121 4135
rect 13169 4119 13185 4135
rect 13187 4119 13203 4135
rect 13241 4119 13257 4135
rect 13259 4119 13275 4135
rect 13323 4119 13339 4135
rect 13341 4119 13357 4135
rect 13395 4119 13411 4135
rect 13413 4119 13429 4135
rect 13477 4119 13493 4135
rect 13495 4119 13511 4135
rect 13549 4119 13565 4135
rect 13567 4119 13583 4135
rect 13631 4119 13647 4135
rect 13649 4119 13665 4135
rect 13703 4119 13719 4135
rect 13721 4119 13737 4135
rect 13785 4119 13801 4135
rect 13803 4119 13819 4135
rect 13857 4119 13873 4135
rect 13875 4119 13891 4135
rect 13939 4119 13955 4135
rect 13957 4119 13973 4135
rect 14011 4119 14027 4135
rect 14029 4119 14045 4135
rect 14093 4119 14109 4135
rect 14111 4119 14127 4135
rect 14165 4119 14181 4135
rect 14183 4119 14199 4135
rect 14247 4119 14260 4135
rect 12907 3890 12932 3900
rect 12981 3890 13006 3900
rect 13052 3881 13080 3900
rect 13044 3875 13050 3881
rect 13052 3875 13085 3881
rect 13125 3875 13126 3881
rect 13129 3875 13154 3900
rect 13160 3875 13166 3881
rect 13203 3875 13228 3900
rect 13241 3875 13247 3881
rect 13277 3875 13302 3900
rect 13322 3875 13328 3881
rect 13351 3875 13376 3900
rect 13425 3881 13450 3900
rect 13404 3875 13410 3881
rect 13425 3875 13456 3881
rect 13485 3875 13491 3881
rect 13499 3875 13524 3900
rect 13531 3875 13537 3881
rect 13566 3875 13570 3881
rect 13573 3875 13598 3900
rect 13612 3875 13618 3881
rect 13644 3875 13646 3900
rect 13647 3875 13672 3900
rect 13693 3875 13699 3881
rect 13718 3875 13746 3900
rect 13774 3875 13780 3881
rect 13792 3875 13820 3900
rect 13866 3881 13894 3900
rect 13855 3875 13861 3881
rect 13866 3875 13896 3881
rect 13936 3875 13940 3881
rect 13943 3875 13968 3900
rect 13972 3875 13978 3881
rect 14017 3875 14042 3900
rect 14053 3875 14059 3881
rect 14091 3875 14116 3900
rect 14134 3875 14140 3881
rect 14165 3875 14190 3900
rect 14215 3875 14221 3881
rect 14239 3875 14260 3900
rect 33770 3875 33772 3881
rect 33775 3875 33800 3900
rect 33816 3875 33822 3881
rect 33846 3875 33874 3900
rect 33897 3875 33903 3881
rect 33920 3875 33948 3900
rect 33978 3875 33984 3881
rect 33994 3875 34022 3900
rect 34068 3881 34096 3900
rect 34059 3875 34065 3881
rect 34068 3875 34100 3881
rect 34140 3875 34142 3881
rect 34145 3875 34170 3900
rect 34175 3875 34181 3881
rect 34219 3875 34244 3900
rect 34256 3875 34262 3881
rect 34293 3875 34318 3900
rect 34338 3875 34344 3881
rect 34367 3875 34392 3900
rect 34441 3881 34466 3900
rect 34419 3875 34425 3881
rect 34441 3875 34471 3881
rect 34500 3875 34506 3881
rect 34515 3875 34540 3900
rect 34546 3875 34552 3881
rect 34581 3875 34586 3881
rect 34589 3875 34614 3900
rect 34627 3875 34633 3881
rect 34660 3875 34661 3900
rect 34663 3875 34688 3900
rect 34708 3875 34714 3881
rect 34734 3875 34762 3900
rect 34789 3875 34795 3881
rect 34808 3875 34836 3900
rect 34882 3881 34910 3900
rect 34870 3875 34876 3881
rect 34882 3875 34912 3881
rect 34952 3875 34956 3881
rect 34959 3875 34984 3900
rect 34987 3875 34993 3881
rect 13024 3869 13083 3875
rect 13131 3869 13137 3875
rect 13154 3869 13160 3875
rect 13212 3869 13218 3875
rect 13235 3869 13241 3875
rect 13293 3869 13299 3875
rect 13316 3869 13322 3875
rect 13374 3869 13380 3875
rect 13398 3869 13404 3875
rect 13456 3869 13462 3875
rect 13479 3869 13485 3875
rect 13537 3869 13543 3875
rect 13560 3869 13566 3875
rect 13616 3869 13624 3875
rect 13641 3869 13646 3875
rect 13024 3829 13050 3869
rect 13052 3829 13083 3869
rect 13024 3823 13083 3829
rect 13131 3829 13154 3851
rect 13131 3823 13160 3829
rect 13212 3823 13228 3851
rect 13235 3823 13241 3829
rect 13293 3823 13302 3851
rect 13374 3829 13376 3851
rect 13316 3823 13322 3829
rect 13374 3823 13380 3829
rect 13397 3823 13404 3851
rect 13456 3823 13462 3829
rect 13471 3823 13485 3851
rect 13537 3823 13543 3829
rect 13545 3823 13566 3851
rect 13616 3829 13618 3869
rect 13644 3851 13646 3869
rect 13619 3829 13646 3851
rect 13616 3823 13646 3829
rect 13690 3869 13705 3875
rect 13718 3869 13786 3875
rect 13792 3869 13897 3875
rect 13943 3869 13946 3875
rect 13966 3869 13972 3875
rect 14024 3869 14030 3875
rect 14047 3869 14053 3875
rect 14105 3869 14111 3875
rect 14128 3869 14134 3875
rect 14186 3869 14192 3875
rect 14209 3869 14215 3875
rect 33818 3869 33828 3875
rect 33845 3869 33909 3875
rect 33920 3869 33990 3875
rect 33994 3869 34099 3875
rect 34146 3869 34152 3875
rect 34169 3869 34175 3875
rect 34227 3869 34233 3875
rect 34250 3869 34256 3875
rect 34308 3869 34314 3875
rect 34332 3869 34338 3875
rect 34390 3869 34396 3875
rect 34413 3869 34419 3875
rect 34471 3869 34477 3875
rect 34494 3869 34500 3875
rect 34552 3869 34558 3875
rect 34575 3869 34581 3875
rect 34632 3869 34639 3875
rect 34657 3869 34661 3875
rect 13690 3829 13699 3869
rect 13718 3829 13780 3869
rect 13792 3829 13861 3869
rect 13866 3829 13897 3869
rect 13690 3823 13705 3829
rect 13718 3823 13786 3829
rect 13792 3823 13897 3829
rect 13943 3829 13968 3851
rect 13943 3823 13972 3829
rect 14024 3823 14042 3851
rect 14047 3823 14053 3829
rect 14105 3823 14116 3851
rect 14186 3829 14190 3851
rect 14211 3829 14215 3851
rect 14128 3823 14134 3829
rect 14186 3823 14192 3829
rect 14209 3823 14215 3829
rect 33818 3829 33822 3869
rect 33846 3829 33903 3869
rect 33920 3829 33984 3869
rect 33994 3829 34065 3869
rect 34068 3829 34099 3869
rect 33818 3823 33828 3829
rect 33845 3823 33909 3829
rect 33920 3823 33990 3829
rect 33994 3823 34099 3829
rect 34146 3829 34170 3851
rect 34146 3823 34175 3829
rect 34227 3823 34244 3851
rect 34250 3823 34256 3829
rect 34308 3823 34318 3851
rect 34390 3829 34392 3851
rect 34332 3823 34338 3829
rect 34390 3823 34396 3829
rect 34413 3823 34419 3851
rect 34471 3823 34477 3829
rect 34487 3823 34500 3851
rect 34552 3823 34558 3829
rect 34561 3823 34581 3851
rect 34632 3829 34633 3869
rect 34660 3851 34661 3869
rect 34635 3829 34661 3851
rect 34632 3823 34661 3829
rect 34706 3869 34720 3875
rect 34734 3869 34801 3875
rect 34808 3869 34913 3875
rect 34959 3869 34962 3875
rect 34981 3869 34987 3875
rect 34706 3829 34714 3869
rect 34734 3829 34795 3869
rect 34808 3829 34876 3869
rect 34882 3829 34913 3869
rect 34706 3823 34720 3829
rect 34734 3823 34801 3829
rect 34808 3823 34913 3829
rect 34959 3829 34984 3851
rect 34959 3823 34987 3829
rect 13044 3817 13050 3823
rect 13052 3817 13085 3823
rect 13125 3817 13126 3823
rect 13052 3777 13080 3817
rect 13044 3771 13050 3777
rect 13052 3771 13085 3777
rect 13125 3771 13126 3777
rect 13129 3771 13154 3823
rect 13160 3817 13166 3823
rect 13160 3771 13166 3777
rect 13203 3771 13228 3823
rect 13241 3817 13247 3823
rect 13241 3771 13247 3777
rect 13277 3771 13302 3823
rect 13322 3817 13328 3823
rect 13322 3771 13328 3777
rect 13351 3771 13376 3823
rect 13404 3817 13410 3823
rect 13425 3817 13456 3823
rect 13485 3817 13491 3823
rect 13425 3777 13450 3817
rect 13404 3771 13410 3777
rect 13425 3771 13456 3777
rect 13485 3771 13491 3777
rect 13499 3771 13524 3823
rect 13531 3817 13537 3823
rect 13566 3817 13570 3823
rect 13531 3771 13537 3777
rect 13566 3771 13570 3777
rect 13573 3771 13598 3823
rect 13612 3817 13618 3823
rect 13612 3771 13618 3777
rect 13644 3771 13646 3823
rect 13647 3771 13672 3823
rect 13693 3817 13699 3823
rect 13693 3771 13699 3777
rect 13718 3771 13746 3823
rect 13774 3817 13780 3823
rect 13774 3771 13780 3777
rect 13792 3771 13820 3823
rect 13855 3817 13861 3823
rect 13866 3817 13896 3823
rect 13936 3817 13940 3823
rect 13866 3777 13894 3817
rect 13855 3771 13861 3777
rect 13866 3771 13896 3777
rect 13936 3771 13940 3777
rect 13943 3771 13968 3823
rect 13972 3817 13978 3823
rect 13972 3771 13978 3777
rect 14017 3771 14042 3823
rect 14053 3817 14059 3823
rect 14053 3771 14059 3777
rect 14091 3771 14116 3823
rect 14134 3817 14140 3823
rect 14134 3771 14140 3777
rect 14165 3771 14190 3823
rect 14215 3817 14221 3823
rect 14215 3771 14221 3777
rect 14239 3771 14260 3823
rect 33770 3817 33772 3823
rect 33770 3771 33772 3777
rect 33775 3771 33800 3823
rect 33816 3817 33822 3823
rect 33816 3771 33822 3777
rect 33846 3771 33874 3823
rect 33897 3817 33903 3823
rect 33897 3771 33903 3777
rect 33920 3771 33948 3823
rect 33978 3817 33984 3823
rect 33978 3771 33984 3777
rect 33994 3771 34022 3823
rect 34059 3817 34065 3823
rect 34068 3817 34100 3823
rect 34140 3817 34142 3823
rect 34068 3777 34096 3817
rect 34059 3771 34065 3777
rect 34068 3771 34100 3777
rect 34140 3771 34142 3777
rect 34145 3771 34170 3823
rect 34175 3817 34181 3823
rect 34175 3771 34181 3777
rect 34219 3771 34244 3823
rect 34256 3817 34262 3823
rect 34256 3771 34262 3777
rect 34293 3771 34318 3823
rect 34338 3817 34344 3823
rect 34338 3771 34344 3777
rect 34367 3771 34392 3823
rect 34419 3817 34425 3823
rect 34441 3817 34471 3823
rect 34500 3817 34506 3823
rect 34441 3777 34466 3817
rect 34419 3771 34425 3777
rect 34441 3771 34471 3777
rect 34500 3771 34506 3777
rect 34515 3771 34540 3823
rect 34546 3817 34552 3823
rect 34581 3817 34586 3823
rect 34546 3771 34552 3777
rect 34581 3771 34586 3777
rect 34589 3771 34614 3823
rect 34627 3817 34633 3823
rect 34627 3771 34633 3777
rect 34660 3771 34661 3823
rect 34663 3771 34688 3823
rect 34708 3817 34714 3823
rect 34708 3771 34714 3777
rect 34734 3771 34762 3823
rect 34789 3817 34795 3823
rect 34789 3771 34795 3777
rect 34808 3771 34836 3823
rect 34870 3817 34876 3823
rect 34882 3817 34912 3823
rect 34952 3817 34956 3823
rect 34882 3777 34910 3817
rect 34870 3771 34876 3777
rect 34882 3771 34912 3777
rect 34952 3771 34956 3777
rect 34959 3771 34984 3823
rect 34987 3817 34993 3823
rect 34987 3771 34993 3777
rect 13024 3765 13083 3771
rect 13131 3765 13137 3771
rect 13154 3765 13160 3771
rect 13212 3765 13218 3771
rect 13235 3765 13241 3771
rect 13293 3765 13299 3771
rect 13316 3765 13322 3771
rect 13374 3765 13380 3771
rect 13398 3765 13404 3771
rect 13456 3765 13462 3771
rect 13479 3765 13485 3771
rect 13537 3765 13543 3771
rect 13560 3765 13566 3771
rect 13616 3765 13624 3771
rect 13641 3765 13646 3771
rect 13024 3725 13050 3765
rect 13052 3725 13083 3765
rect 13024 3719 13083 3725
rect 13131 3725 13154 3747
rect 13131 3719 13160 3725
rect 13212 3719 13228 3747
rect 13235 3719 13241 3725
rect 13293 3719 13302 3747
rect 13374 3725 13376 3747
rect 13316 3719 13322 3725
rect 13374 3719 13380 3725
rect 13397 3719 13404 3747
rect 13456 3719 13462 3725
rect 13471 3719 13485 3747
rect 13537 3719 13543 3725
rect 13545 3719 13566 3747
rect 13616 3725 13618 3765
rect 13644 3747 13646 3765
rect 13619 3725 13646 3747
rect 13616 3719 13646 3725
rect 13690 3765 13705 3771
rect 13718 3765 13786 3771
rect 13792 3765 13897 3771
rect 13943 3765 13946 3771
rect 13966 3765 13972 3771
rect 14024 3765 14030 3771
rect 14047 3765 14053 3771
rect 14105 3765 14111 3771
rect 14128 3765 14134 3771
rect 14186 3765 14192 3771
rect 14209 3765 14215 3771
rect 33818 3765 33828 3771
rect 33845 3765 33909 3771
rect 33920 3765 33990 3771
rect 33994 3765 34099 3771
rect 34146 3765 34152 3771
rect 34169 3765 34175 3771
rect 34227 3765 34233 3771
rect 34250 3765 34256 3771
rect 34308 3765 34314 3771
rect 34332 3765 34338 3771
rect 34390 3765 34396 3771
rect 34413 3765 34419 3771
rect 34471 3765 34477 3771
rect 34494 3765 34500 3771
rect 34552 3765 34558 3771
rect 34575 3765 34581 3771
rect 34632 3765 34639 3771
rect 34657 3765 34661 3771
rect 13690 3725 13699 3765
rect 13718 3725 13780 3765
rect 13792 3725 13861 3765
rect 13866 3725 13897 3765
rect 13690 3719 13705 3725
rect 13718 3719 13786 3725
rect 13792 3719 13897 3725
rect 13943 3725 13968 3747
rect 13943 3719 13972 3725
rect 14024 3719 14042 3747
rect 14047 3719 14053 3725
rect 14105 3719 14116 3747
rect 14186 3725 14190 3747
rect 14211 3725 14215 3747
rect 14128 3719 14134 3725
rect 14186 3719 14192 3725
rect 14209 3719 14215 3725
rect 33818 3725 33822 3765
rect 33846 3725 33903 3765
rect 33920 3725 33984 3765
rect 33994 3725 34065 3765
rect 34068 3725 34099 3765
rect 33818 3719 33828 3725
rect 33845 3719 33909 3725
rect 33920 3719 33990 3725
rect 33994 3719 34099 3725
rect 34146 3725 34170 3747
rect 34146 3719 34175 3725
rect 34227 3719 34244 3747
rect 34250 3719 34256 3725
rect 34308 3719 34318 3747
rect 34390 3725 34392 3747
rect 34332 3719 34338 3725
rect 34390 3719 34396 3725
rect 34413 3719 34419 3747
rect 34471 3719 34477 3725
rect 34487 3719 34500 3747
rect 34552 3719 34558 3725
rect 34561 3719 34581 3747
rect 34632 3725 34633 3765
rect 34660 3747 34661 3765
rect 34635 3725 34661 3747
rect 34632 3719 34661 3725
rect 34706 3765 34720 3771
rect 34734 3765 34801 3771
rect 34808 3765 34913 3771
rect 34959 3765 34962 3771
rect 34981 3765 34987 3771
rect 34706 3725 34714 3765
rect 34734 3725 34795 3765
rect 34808 3725 34876 3765
rect 34882 3725 34913 3765
rect 34706 3719 34720 3725
rect 34734 3719 34801 3725
rect 34808 3719 34913 3725
rect 34959 3725 34984 3747
rect 34959 3719 34987 3725
rect 13044 3713 13050 3719
rect 13052 3713 13085 3719
rect 13125 3713 13126 3719
rect 13052 3673 13080 3713
rect 13044 3667 13050 3673
rect 13052 3667 13085 3673
rect 13125 3667 13126 3673
rect 13129 3667 13154 3719
rect 13160 3713 13166 3719
rect 13160 3667 13166 3673
rect 13203 3667 13228 3719
rect 13241 3713 13247 3719
rect 13241 3667 13247 3673
rect 13277 3667 13302 3719
rect 13322 3713 13328 3719
rect 13322 3667 13328 3673
rect 13351 3667 13376 3719
rect 13404 3713 13410 3719
rect 13425 3713 13456 3719
rect 13485 3713 13491 3719
rect 13425 3673 13450 3713
rect 13404 3667 13410 3673
rect 13425 3667 13456 3673
rect 13485 3667 13491 3673
rect 13499 3667 13524 3719
rect 13531 3713 13537 3719
rect 13566 3713 13570 3719
rect 13531 3667 13537 3673
rect 13566 3667 13570 3673
rect 13573 3667 13598 3719
rect 13612 3713 13618 3719
rect 13612 3667 13618 3673
rect 13644 3667 13646 3719
rect 13647 3667 13672 3719
rect 13693 3713 13699 3719
rect 13693 3667 13699 3673
rect 13718 3667 13746 3719
rect 13774 3713 13780 3719
rect 13774 3667 13780 3673
rect 13792 3667 13820 3719
rect 13855 3713 13861 3719
rect 13866 3713 13896 3719
rect 13936 3713 13940 3719
rect 13866 3673 13894 3713
rect 13855 3667 13861 3673
rect 13866 3667 13896 3673
rect 13936 3667 13940 3673
rect 13943 3667 13968 3719
rect 13972 3713 13978 3719
rect 13972 3667 13978 3673
rect 14017 3667 14042 3719
rect 14053 3713 14059 3719
rect 14053 3667 14059 3673
rect 14091 3667 14116 3719
rect 14134 3713 14140 3719
rect 14134 3667 14140 3673
rect 14165 3667 14190 3719
rect 14215 3713 14221 3719
rect 14215 3667 14221 3673
rect 14239 3667 14260 3719
rect 33770 3713 33772 3719
rect 33770 3667 33772 3673
rect 33775 3667 33800 3719
rect 33816 3713 33822 3719
rect 33816 3667 33822 3673
rect 33846 3667 33874 3719
rect 33897 3713 33903 3719
rect 33897 3667 33903 3673
rect 33920 3667 33948 3719
rect 33978 3713 33984 3719
rect 33978 3667 33984 3673
rect 33994 3667 34022 3719
rect 34059 3713 34065 3719
rect 34068 3713 34100 3719
rect 34140 3713 34142 3719
rect 34068 3673 34096 3713
rect 34059 3667 34065 3673
rect 34068 3667 34100 3673
rect 34140 3667 34142 3673
rect 34145 3667 34170 3719
rect 34175 3713 34181 3719
rect 34175 3667 34181 3673
rect 34219 3667 34244 3719
rect 34256 3713 34262 3719
rect 34256 3667 34262 3673
rect 34293 3667 34318 3719
rect 34338 3713 34344 3719
rect 34338 3667 34344 3673
rect 34367 3667 34392 3719
rect 34419 3713 34425 3719
rect 34441 3713 34471 3719
rect 34500 3713 34506 3719
rect 34441 3673 34466 3713
rect 34419 3667 34425 3673
rect 34441 3667 34471 3673
rect 34500 3667 34506 3673
rect 34515 3667 34540 3719
rect 34546 3713 34552 3719
rect 34581 3713 34586 3719
rect 34546 3667 34552 3673
rect 34581 3667 34586 3673
rect 34589 3667 34614 3719
rect 34627 3713 34633 3719
rect 34627 3667 34633 3673
rect 34660 3667 34661 3719
rect 34663 3667 34688 3719
rect 34708 3713 34714 3719
rect 34708 3667 34714 3673
rect 34734 3667 34762 3719
rect 34789 3713 34795 3719
rect 34789 3667 34795 3673
rect 34808 3667 34836 3719
rect 34870 3713 34876 3719
rect 34882 3713 34912 3719
rect 34952 3713 34956 3719
rect 34882 3673 34910 3713
rect 34870 3667 34876 3673
rect 34882 3667 34912 3673
rect 34952 3667 34956 3673
rect 34959 3667 34984 3719
rect 34987 3713 34993 3719
rect 34987 3667 34993 3673
rect 13024 3661 13083 3667
rect 13131 3661 13137 3667
rect 13154 3661 13160 3667
rect 13212 3661 13218 3667
rect 13235 3661 13241 3667
rect 13293 3661 13299 3667
rect 13316 3661 13322 3667
rect 13374 3661 13380 3667
rect 13398 3661 13404 3667
rect 13456 3661 13462 3667
rect 13479 3661 13485 3667
rect 13537 3661 13543 3667
rect 13560 3661 13566 3667
rect 13616 3661 13624 3667
rect 13641 3661 13646 3667
rect 13024 3621 13050 3661
rect 13052 3621 13083 3661
rect 13024 3615 13083 3621
rect 13131 3621 13154 3643
rect 13131 3615 13160 3621
rect 13212 3615 13228 3643
rect 13235 3615 13241 3621
rect 13293 3615 13302 3643
rect 13374 3621 13376 3643
rect 13316 3615 13322 3621
rect 13374 3615 13380 3621
rect 13397 3615 13404 3643
rect 13456 3615 13462 3621
rect 13471 3615 13485 3643
rect 13537 3615 13543 3621
rect 13545 3615 13566 3643
rect 13616 3621 13618 3661
rect 13644 3643 13646 3661
rect 13619 3621 13646 3643
rect 13616 3615 13646 3621
rect 13690 3661 13705 3667
rect 13718 3661 13786 3667
rect 13792 3661 13897 3667
rect 13943 3661 13946 3667
rect 13966 3661 13972 3667
rect 14024 3661 14030 3667
rect 14047 3661 14053 3667
rect 14105 3661 14111 3667
rect 14128 3661 14134 3667
rect 14186 3661 14192 3667
rect 14209 3661 14215 3667
rect 33818 3661 33828 3667
rect 33845 3661 33909 3667
rect 33920 3661 33990 3667
rect 33994 3661 34099 3667
rect 34146 3661 34152 3667
rect 34169 3661 34175 3667
rect 34227 3661 34233 3667
rect 34250 3661 34256 3667
rect 34308 3661 34314 3667
rect 34332 3661 34338 3667
rect 34390 3661 34396 3667
rect 34413 3661 34419 3667
rect 34471 3661 34477 3667
rect 34494 3661 34500 3667
rect 34552 3661 34558 3667
rect 34575 3661 34581 3667
rect 34632 3661 34639 3667
rect 34657 3661 34661 3667
rect 13690 3621 13699 3661
rect 13718 3621 13780 3661
rect 13792 3621 13861 3661
rect 13866 3621 13897 3661
rect 13690 3615 13705 3621
rect 13718 3615 13786 3621
rect 13792 3615 13897 3621
rect 13943 3621 13968 3643
rect 13943 3615 13972 3621
rect 14024 3615 14042 3643
rect 14047 3615 14053 3621
rect 14105 3615 14116 3643
rect 14186 3621 14190 3643
rect 14211 3621 14215 3643
rect 14128 3615 14134 3621
rect 14186 3615 14192 3621
rect 14209 3615 14215 3621
rect 33818 3621 33822 3661
rect 33846 3621 33903 3661
rect 33920 3621 33984 3661
rect 33994 3621 34065 3661
rect 34068 3621 34099 3661
rect 33818 3615 33828 3621
rect 33845 3615 33909 3621
rect 33920 3615 33990 3621
rect 33994 3615 34099 3621
rect 34146 3621 34170 3643
rect 34146 3615 34175 3621
rect 34227 3615 34244 3643
rect 34250 3615 34256 3621
rect 34308 3615 34318 3643
rect 34390 3621 34392 3643
rect 34332 3615 34338 3621
rect 34390 3615 34396 3621
rect 34413 3615 34419 3643
rect 34471 3615 34477 3621
rect 34487 3615 34500 3643
rect 34552 3615 34558 3621
rect 34561 3615 34581 3643
rect 34632 3621 34633 3661
rect 34660 3643 34661 3661
rect 34635 3621 34661 3643
rect 34632 3615 34661 3621
rect 34706 3661 34720 3667
rect 34734 3661 34801 3667
rect 34808 3661 34913 3667
rect 34959 3661 34962 3667
rect 34981 3661 34987 3667
rect 34706 3621 34714 3661
rect 34734 3621 34795 3661
rect 34808 3621 34876 3661
rect 34882 3621 34913 3661
rect 34706 3615 34720 3621
rect 34734 3615 34801 3621
rect 34808 3615 34913 3621
rect 34959 3621 34984 3643
rect 34959 3615 34987 3621
rect 13000 3610 13006 3615
rect 12907 3604 12932 3610
rect 12981 3604 13006 3610
rect 13044 3609 13050 3615
rect 13052 3609 13085 3615
rect 13125 3609 13126 3615
rect 13052 3604 13080 3609
rect 13129 3604 13154 3615
rect 13160 3609 13166 3615
rect 13203 3604 13228 3615
rect 13241 3609 13247 3615
rect 13277 3604 13302 3615
rect 13322 3609 13328 3615
rect 13351 3604 13376 3615
rect 13404 3609 13410 3615
rect 13425 3609 13456 3615
rect 13485 3609 13491 3615
rect 13425 3604 13450 3609
rect 13499 3604 13524 3615
rect 13531 3609 13537 3615
rect 13566 3609 13570 3615
rect 13573 3604 13598 3615
rect 13612 3609 13618 3615
rect 13644 3604 13646 3615
rect 13647 3604 13672 3615
rect 13693 3609 13699 3615
rect 13718 3604 13746 3615
rect 13774 3609 13780 3615
rect 13792 3604 13820 3615
rect 13855 3609 13861 3615
rect 13866 3609 13896 3615
rect 13936 3609 13940 3615
rect 13866 3604 13894 3609
rect 13943 3604 13968 3615
rect 13972 3609 13978 3615
rect 14017 3604 14042 3615
rect 14053 3609 14059 3615
rect 14091 3604 14116 3615
rect 14134 3609 14140 3615
rect 14165 3604 14190 3615
rect 14215 3609 14221 3615
rect 14239 3604 14260 3615
rect 33770 3609 33772 3615
rect 33775 3604 33800 3615
rect 33816 3609 33822 3615
rect 33846 3604 33874 3615
rect 33897 3609 33903 3615
rect 33920 3604 33948 3615
rect 33978 3609 33984 3615
rect 33994 3604 34022 3615
rect 34059 3609 34065 3615
rect 34068 3609 34100 3615
rect 34140 3609 34142 3615
rect 34068 3604 34096 3609
rect 34145 3604 34170 3615
rect 34175 3609 34181 3615
rect 34219 3604 34244 3615
rect 34256 3609 34262 3615
rect 34293 3604 34318 3615
rect 34338 3609 34344 3615
rect 34367 3604 34392 3615
rect 34419 3609 34425 3615
rect 34441 3609 34471 3615
rect 34500 3609 34506 3615
rect 34441 3604 34466 3609
rect 34515 3604 34540 3615
rect 34546 3609 34552 3615
rect 34581 3609 34586 3615
rect 34589 3604 34614 3615
rect 34627 3609 34633 3615
rect 34660 3604 34661 3615
rect 34663 3604 34688 3615
rect 34708 3609 34714 3615
rect 34734 3604 34762 3615
rect 34789 3609 34795 3615
rect 34808 3604 34836 3615
rect 34870 3609 34876 3615
rect 34882 3609 34912 3615
rect 34952 3609 34956 3615
rect 34882 3604 34910 3609
rect 34959 3604 34984 3615
rect 34987 3609 34993 3615
<< error_s >>
rect 35000 3615 35030 3634
rect 35028 3604 35030 3615
<< metal1 >>
rect 3270 17968 7575 18001
rect 3270 17852 3294 17968
rect 7570 17852 7575 17968
rect 3270 17819 7575 17852
rect 2275 17185 6745 17205
rect 2269 17170 6751 17185
rect 2269 16990 2276 17170
rect 6744 16990 6751 17170
rect 2269 16975 6751 16990
rect 6515 14295 6745 16975
rect 7405 15230 7575 17819
rect 7405 15060 8390 15230
rect 6515 14065 7695 14295
rect 7465 6285 7695 14065
rect 7465 6055 9310 6285
rect 9080 4975 9310 6055
rect 9080 4970 9558 4975
rect 9080 4967 9560 4970
rect 9080 4723 9312 4967
rect 9556 4723 9560 4967
rect 9080 4720 9560 4723
rect 9310 4715 9558 4720
rect 37180 3600 38650 3900
<< via1 >>
rect 3294 17852 7570 17968
rect 2276 16990 6744 17170
rect 9312 4723 9556 4967
<< metal2 >>
rect -3150 19580 -2820 19680
rect -1650 16075 -1560 18571
rect -4300 15965 -1560 16075
rect -4300 15315 -4190 15965
rect -1140 15470 -1050 18581
rect 1300 17115 1410 18621
rect 3300 18000 3410 18621
rect 3270 17995 3650 18000
rect 3270 17968 7581 17995
rect 3270 17852 3294 17968
rect 7570 17852 7581 17968
rect 3270 17825 7581 17852
rect 3270 17820 3650 17825
rect 2275 17170 6745 17191
rect 2275 17115 2276 17170
rect 1300 17005 2276 17115
rect 2275 16990 2276 17005
rect 6744 16990 6745 17170
rect 2275 16969 6745 16990
rect -6725 14780 -6405 14890
rect -6815 12910 -6445 13000
rect -6885 9910 -6415 10000
rect 7150 8781 9060 9029
rect -6785 6910 -6460 7000
rect 7150 4598 7398 8781
rect 9304 4967 9564 4969
rect 9304 4723 9312 4967
rect 9556 4723 9564 4967
rect 9304 4721 9564 4723
rect 5990 4480 7398 4598
rect 5984 4232 7398 4480
<< metal3 >>
rect -1380 20090 -1180 20620
rect -870 20146 -670 20610
rect 150 19916 270 20280
rect 2220 19916 2340 20380
rect -1900 16385 -1810 18570
rect -4745 16295 -1810 16385
<< metal4 >>
rect -6705 14980 -6435 15090
rect 36260 12000 39290 12860
rect -4030 3675 -3920 3940
rect -3330 3840 -3110 4560
rect -330 3940 -110 4700
rect 2670 3690 2890 4690
<< metal5 >>
rect -6700 14270 -4950 14590
use bias#0  bias_0
timestamp 1654643737
transform 1 0 -3740 0 1 20716
box 790 -2236 7180 -220
use opamp_wrapper  opamp_wrapper_0
timestamp 1654749028
transform 1 0 10500 0 1 5170
box -2280 -1640 26995 13665
use pixel_array#0  pixel_array_0
timestamp 1654643737
transform 1 0 -3550 0 1 11430
box -3000 -7600 9740 5000
<< labels >>
rlabel metal1 s 38350 3600 38650 3900 4 GND
port 1 nsew
rlabel metal3 s 230 20230 230 20230 4 OUT_IB
port 2 nsew
rlabel metal3 s 2220 20260 2340 20380 4 AMP_Ib
port 3 nsew
rlabel metal3 s -870 20410 -670 20610 4 NB2
port 4 nsew
rlabel metal3 s -1380 20420 -1180 20620 4 NB1
port 5 nsew
rlabel metal2 s -3150 19580 -2820 19680 4 SF_IB
port 6 nsew
rlabel metal4 s 38430 12000 39290 12860 4 AOUT
port 7 nsew
rlabel metal4 s -6705 14980 -6595 15090 4 VBIAS
port 8 nsew
rlabel metal2 s -6725 14780 -6615 14890 4 VREF
port 9 nsew
rlabel metal4 s -4030 3675 -3920 3785 4 CSA_VREF
port 10 nsew
rlabel metal4 s -3330 3840 -3110 4060 4 COL_SEL0
port 11 nsew
rlabel metal4 s -330 3940 -110 4160 4 COL_SEL1
port 12 nsew
rlabel metal4 s 2670 3690 2890 3910 4 COL_SEL2
port 13 nsew
rlabel metal2 s -6785 6910 -6695 7000 4 ROW_SEL2
port 14 nsew
rlabel metal2 s -6885 9910 -6795 10000 4 ROW_SEL1
port 15 nsew
rlabel metal2 s -6815 12910 -6725 13000 4 ROW_SEL0
port 16 nsew
rlabel metal5 s -6700 14270 -6380 14590 4 GRING
port 17 nsew
<< end >>
