magic
tech sky130A
timestamp 1654641414
<< nmoslvt >>
rect 270 -3400 1070 -3200
rect 1770 -3400 2570 -3200
rect 3270 -3400 4070 -3200
<< ndiff >>
rect 270 -3160 1070 -3150
rect 270 -3190 280 -3160
rect 1060 -3190 1070 -3160
rect 270 -3200 1070 -3190
rect 1770 -3160 2570 -3150
rect 1770 -3190 1780 -3160
rect 2560 -3190 2570 -3160
rect 1770 -3200 2570 -3190
rect 3270 -3160 4070 -3150
rect 3270 -3190 3280 -3160
rect 4060 -3190 4070 -3160
rect 3270 -3200 4070 -3190
rect 270 -3415 1070 -3400
rect 270 -3435 280 -3415
rect 1060 -3435 1070 -3415
rect 270 -3440 1070 -3435
rect 1770 -3415 2570 -3400
rect 1770 -3435 1780 -3415
rect 2560 -3435 2570 -3415
rect 1770 -3440 2570 -3435
rect 3270 -3415 4070 -3400
rect 3270 -3435 3280 -3415
rect 4060 -3435 4070 -3415
rect 3270 -3440 4070 -3435
<< ndiffc >>
rect 280 -3190 1060 -3160
rect 1780 -3190 2560 -3160
rect 3280 -3190 4060 -3160
rect 280 -3435 1060 -3415
rect 1780 -3435 2560 -3415
rect 3280 -3435 4060 -3415
<< poly >>
rect 255 -3245 270 -3200
rect 110 -3250 270 -3245
rect 110 -3350 120 -3250
rect 210 -3350 270 -3250
rect 110 -3355 270 -3350
rect 255 -3400 270 -3355
rect 1070 -3400 1085 -3200
rect 1755 -3245 1770 -3200
rect 1610 -3250 1770 -3245
rect 1610 -3350 1620 -3250
rect 1710 -3350 1770 -3250
rect 1610 -3355 1770 -3350
rect 1755 -3400 1770 -3355
rect 2570 -3400 2585 -3200
rect 3255 -3245 3270 -3200
rect 3110 -3250 3270 -3245
rect 3110 -3350 3120 -3250
rect 3210 -3350 3270 -3250
rect 3110 -3355 3270 -3350
rect 3255 -3400 3270 -3355
rect 4070 -3400 4085 -3200
<< polycont >>
rect 120 -3350 210 -3250
rect 1620 -3350 1710 -3250
rect 3120 -3350 3210 -3250
<< locali >>
rect 270 -3145 280 -3115
rect 1060 -3145 1070 -3115
rect 270 -3160 1070 -3145
rect 270 -3190 280 -3160
rect 1060 -3190 1070 -3160
rect 1770 -3145 1780 -3115
rect 2560 -3145 2570 -3115
rect 1770 -3160 2570 -3145
rect 1770 -3190 1780 -3160
rect 2560 -3190 2570 -3160
rect 3270 -3145 3280 -3115
rect 4060 -3145 4070 -3115
rect 3270 -3160 4070 -3145
rect 3270 -3190 3280 -3160
rect 4060 -3190 4070 -3160
rect 110 -3250 220 -3245
rect 110 -3350 120 -3250
rect 210 -3350 220 -3250
rect 110 -3355 220 -3350
rect 1610 -3250 1720 -3245
rect 1610 -3350 1620 -3250
rect 1710 -3350 1720 -3250
rect 1610 -3355 1720 -3350
rect 3110 -3250 3220 -3245
rect 3110 -3350 3120 -3250
rect 3210 -3350 3220 -3250
rect 3110 -3355 3220 -3350
rect 270 -3415 1070 -3400
rect 270 -3435 280 -3415
rect 1060 -3435 1070 -3415
rect 270 -3460 1070 -3435
rect 270 -3490 280 -3460
rect 1060 -3490 1070 -3460
rect 270 -3500 1070 -3490
rect 1770 -3415 2570 -3400
rect 1770 -3435 1780 -3415
rect 2560 -3435 2570 -3415
rect 1770 -3460 2570 -3435
rect 1770 -3490 1780 -3460
rect 2560 -3490 2570 -3460
rect 1770 -3500 2570 -3490
rect 3270 -3415 4070 -3400
rect 3270 -3435 3280 -3415
rect 4060 -3435 4070 -3415
rect 3270 -3460 4070 -3435
rect 3270 -3490 3280 -3460
rect 4060 -3490 4070 -3460
rect 3270 -3500 4070 -3490
<< viali >>
rect 280 -3145 1060 -3115
rect 1780 -3145 2560 -3115
rect 3280 -3145 4060 -3115
rect 120 -3350 210 -3250
rect 1620 -3350 1710 -3250
rect 3120 -3350 3210 -3250
rect 280 -3490 1060 -3460
rect 1780 -3490 2560 -3460
rect 3280 -3490 4060 -3460
<< metal1 >>
rect -885 1725 4000 1730
rect -450 1680 25 1725
rect 70 1680 1525 1725
rect 1570 1680 3025 1725
rect 3070 1680 4000 1725
rect -885 1675 4000 1680
rect -1000 1485 -900 1495
rect -1000 1440 20 1485
rect -1000 1410 0 1440
rect -1000 -15 -900 1410
rect -800 780 0 785
rect -800 745 -790 780
rect -590 745 -270 780
rect -130 745 0 780
rect -800 740 0 745
rect 4700 90 4800 1515
rect 4500 15 4800 90
rect -1000 -60 20 -15
rect -1000 -90 0 -60
rect -1000 -1515 -900 -90
rect -800 -720 0 -715
rect -800 -755 -790 -720
rect -590 -755 -270 -720
rect -130 -755 0 -720
rect -800 -760 0 -755
rect 4700 -1410 4800 15
rect 4500 -1485 4800 -1410
rect -1000 -1560 20 -1515
rect -1000 -1590 0 -1560
rect -1000 -3000 -900 -1590
rect -800 -2220 0 -2215
rect -800 -2255 -790 -2220
rect -590 -2255 -270 -2220
rect -130 -2255 0 -2220
rect -800 -2260 0 -2255
rect 4700 -2910 4800 -1485
rect 1430 -2955 1500 -2915
rect 4500 -2985 4800 -2910
rect 270 -3100 280 -3065
rect 1060 -3100 1070 -3065
rect 270 -3115 1070 -3100
rect 270 -3145 280 -3115
rect 1060 -3145 1070 -3115
rect 270 -3150 1070 -3145
rect 1770 -3100 1780 -3065
rect 2560 -3100 2570 -3065
rect 1770 -3115 2570 -3100
rect 1770 -3145 1780 -3115
rect 2560 -3145 2570 -3115
rect 1770 -3150 2570 -3145
rect 3270 -3100 3280 -3065
rect 4060 -3100 4070 -3065
rect 3270 -3115 4070 -3100
rect 3270 -3145 3280 -3115
rect 4060 -3145 4070 -3115
rect 3270 -3150 4070 -3145
rect 110 -3250 220 -3245
rect 110 -3350 120 -3250
rect 210 -3350 220 -3250
rect 110 -3355 220 -3350
rect 1610 -3250 1720 -3245
rect 1610 -3350 1620 -3250
rect 1710 -3350 1720 -3250
rect 1610 -3355 1720 -3350
rect 3110 -3250 3220 -3245
rect 3110 -3350 3120 -3250
rect 3210 -3350 3220 -3250
rect 3110 -3355 3220 -3350
rect 270 -3460 4870 -3450
rect 270 -3540 280 -3460
rect 270 -3550 4870 -3540
<< via1 >>
rect -885 1680 -450 1725
rect 25 1680 70 1725
rect 1525 1680 1570 1725
rect 3025 1680 3070 1725
rect -790 745 -590 780
rect -270 745 -130 780
rect -790 -755 -590 -720
rect -270 -755 -130 -720
rect -790 -2255 -590 -2220
rect -270 -2255 -130 -2220
rect 280 -3100 1060 -3065
rect 1780 -3100 2560 -3065
rect 3280 -3100 4060 -3065
rect 120 -3350 210 -3250
rect 1620 -3350 1710 -3250
rect 3120 -3350 3210 -3250
rect 280 -3490 1060 -3460
rect 1060 -3490 1780 -3460
rect 1780 -3490 2560 -3460
rect 2560 -3490 3280 -3460
rect 3280 -3490 4060 -3460
rect 4060 -3490 4870 -3460
rect 280 -3540 4870 -3490
<< metal2 >>
rect 0 2020 4500 2075
rect -1500 1725 -445 1730
rect -1500 1680 -885 1725
rect -450 1680 -445 1725
rect -1500 1675 -445 1680
rect -1500 780 -500 785
rect -1500 745 -790 780
rect -590 745 -500 780
rect -1500 740 -500 745
rect -375 115 -320 2000
rect 240 1825 295 1830
rect 30 1730 65 1800
rect 240 1780 245 1825
rect 290 1780 295 1825
rect 240 1775 295 1780
rect 20 1725 75 1730
rect 20 1680 25 1725
rect 70 1680 75 1725
rect 20 1675 75 1680
rect 30 1500 65 1675
rect 250 1500 285 1775
rect 510 1500 545 2020
rect 1740 1825 1795 1830
rect 1530 1730 1565 1800
rect 1740 1780 1745 1825
rect 1790 1780 1795 1825
rect 1740 1775 1795 1780
rect 1520 1725 1575 1730
rect 1520 1680 1525 1725
rect 1570 1680 1575 1725
rect 1520 1675 1575 1680
rect 1530 1500 1565 1675
rect 1750 1500 1785 1775
rect 2010 1500 2045 2020
rect 3240 1825 3295 1830
rect 3030 1730 3065 1800
rect 3240 1780 3245 1825
rect 3290 1780 3295 1825
rect 3240 1775 3295 1780
rect 3020 1725 3075 1730
rect 3020 1680 3025 1725
rect 3070 1680 3075 1725
rect 3020 1675 3075 1680
rect 3030 1500 3065 1675
rect 3250 1500 3285 1775
rect 3510 1500 3545 2020
rect -280 780 -130 785
rect -280 745 -270 780
rect -280 740 -130 745
rect -375 80 -370 115
rect -325 80 -320 115
rect -1500 -720 -500 -715
rect -1500 -755 -790 -720
rect -590 -755 -500 -720
rect -1500 -760 -500 -755
rect -375 -1385 -320 80
rect -280 -720 -130 -715
rect -280 -755 -270 -720
rect -280 -760 -130 -755
rect -375 -1420 -370 -1385
rect -325 -1420 -320 -1385
rect -1500 -2220 -500 -2215
rect -1500 -2255 -790 -2220
rect -590 -2255 -500 -2220
rect -1500 -2260 -500 -2255
rect -375 -2885 -320 -1420
rect -280 -2220 -130 -2215
rect -280 -2255 -270 -2220
rect -280 -2260 -130 -2255
rect -375 -2920 -370 -2885
rect -325 -2920 -320 -2885
rect -375 -3000 -320 -2920
rect 270 -3040 1390 -3030
rect 270 -3100 280 -3040
rect 1380 -3090 1390 -3040
rect 1060 -3100 1390 -3090
rect 1770 -3040 2890 -3030
rect 1770 -3100 1780 -3040
rect 2880 -3090 2890 -3040
rect 2560 -3100 2890 -3090
rect 3270 -3040 4390 -3030
rect 3270 -3100 3280 -3040
rect 4380 -3090 4390 -3040
rect 4060 -3100 4390 -3090
rect 110 -3250 220 -3245
rect 110 -3350 120 -3250
rect 210 -3350 220 -3250
rect 110 -3355 220 -3350
rect 1610 -3250 1720 -3245
rect 1610 -3350 1620 -3250
rect 1710 -3350 1720 -3250
rect 1610 -3355 1720 -3350
rect 3110 -3250 3220 -3245
rect 3110 -3350 3120 -3250
rect 3210 -3350 3220 -3250
rect 3110 -3355 3220 -3350
rect 270 -3460 4870 -3450
rect 270 -3540 280 -3460
rect 270 -3550 4870 -3540
<< via2 >>
rect 245 1780 290 1825
rect 1745 1780 1790 1825
rect 3245 1780 3290 1825
rect -270 745 -130 780
rect -370 80 -325 115
rect -270 -755 -130 -720
rect -370 -1420 -325 -1385
rect -270 -2255 -130 -2220
rect -370 -2920 -325 -2885
rect 280 -3065 1380 -3040
rect 280 -3090 1060 -3065
rect 1060 -3090 1380 -3065
rect 1780 -3065 2880 -3040
rect 1780 -3090 2560 -3065
rect 2560 -3090 2880 -3065
rect 3280 -3065 4380 -3040
rect 3280 -3090 4060 -3065
rect 4060 -3090 4380 -3065
rect 120 -3350 210 -3250
rect 1620 -3350 1710 -3250
rect 3120 -3350 3210 -3250
<< metal3 >>
rect -600 1420 -555 2500
rect 240 1825 295 1830
rect 240 1780 245 1825
rect 290 1780 295 1825
rect 240 1775 295 1780
rect 1740 1825 1795 1830
rect 1740 1780 1745 1825
rect 1790 1780 1795 1825
rect 1740 1775 1795 1780
rect 3240 1825 3295 1830
rect 3240 1780 3245 1825
rect 3290 1780 3295 1825
rect 3240 1775 3295 1780
rect -600 1375 100 1420
rect -600 -80 -555 1375
rect -240 1275 -185 1280
rect -280 1270 260 1275
rect -280 1235 -235 1270
rect -190 1235 260 1270
rect -280 1230 260 1235
rect -240 1225 -185 1230
rect -280 780 220 785
rect -280 745 -270 780
rect -130 745 220 780
rect -280 740 220 745
rect -380 115 20 125
rect -380 80 -370 115
rect -325 80 20 115
rect -375 70 -320 80
rect -600 -125 100 -80
rect -600 -1580 -555 -125
rect -240 -225 -185 -220
rect -280 -230 260 -225
rect -280 -265 -235 -230
rect -190 -265 260 -230
rect -280 -270 260 -265
rect -240 -275 -185 -270
rect -280 -720 220 -715
rect -280 -755 -270 -720
rect -130 -755 220 -720
rect -280 -760 220 -755
rect -380 -1385 20 -1375
rect -380 -1420 -370 -1385
rect -325 -1420 20 -1385
rect -375 -1430 -320 -1420
rect -600 -1625 100 -1580
rect -600 -2000 -555 -1625
rect -240 -1725 -185 -1720
rect -280 -1730 260 -1725
rect -280 -1765 -235 -1730
rect -190 -1765 260 -1730
rect -280 -1770 260 -1765
rect -240 -1775 -185 -1770
rect -280 -2220 220 -2215
rect -280 -2255 -270 -2220
rect -130 -2255 220 -2220
rect -280 -2260 220 -2255
rect -380 -2885 20 -2875
rect -380 -2920 -370 -2885
rect -325 -2920 20 -2885
rect -375 -2930 -320 -2920
rect 270 -3040 1390 -3030
rect 270 -3090 280 -3040
rect 1380 -3090 1390 -3040
rect 270 -3100 1390 -3090
rect 1770 -3040 2890 -3030
rect 1770 -3090 1780 -3040
rect 2880 -3090 2890 -3040
rect 1770 -3100 2890 -3090
rect 3270 -3040 4390 -3030
rect 3270 -3090 3280 -3040
rect 4380 -3090 4390 -3040
rect 3270 -3100 4390 -3090
rect 110 -3250 220 -3245
rect 110 -3350 120 -3250
rect 210 -3350 220 -3250
rect 110 -3355 220 -3350
rect 1610 -3250 1720 -3245
rect 1610 -3350 1620 -3250
rect 1710 -3350 1720 -3250
rect 1610 -3355 1720 -3350
rect 3110 -3250 3220 -3245
rect 3110 -3350 3120 -3250
rect 3210 -3350 3220 -3250
rect 3110 -3355 3220 -3350
<< via3 >>
rect 245 1780 290 1825
rect 1745 1780 1790 1825
rect 3245 1780 3290 1825
rect -235 1235 -190 1270
rect -235 -265 -190 -230
rect -235 -1765 -190 -1730
rect 280 -3090 1380 -3040
rect 1780 -3090 2880 -3040
rect 3280 -3090 4380 -3040
rect 120 -3350 210 -3250
rect 1620 -3350 1710 -3250
rect 3120 -3350 3210 -3250
<< metal4 >>
rect -1500 1825 4100 1830
rect -1500 1780 245 1825
rect 290 1780 1745 1825
rect 1790 1780 3245 1825
rect 3290 1780 4100 1825
rect -1500 1775 4100 1780
rect -240 1270 -185 1300
rect -240 1235 -235 1270
rect -190 1235 -185 1270
rect -240 -230 -185 1235
rect -240 -265 -235 -230
rect -190 -265 -185 -230
rect -240 -1730 -185 -265
rect -240 -1765 -235 -1730
rect -190 -1765 -185 -1730
rect -240 -3800 -185 -1765
rect 1315 -3030 1390 -3000
rect 2815 -3030 2890 -3000
rect 4315 -3030 4390 -3000
rect 270 -3040 1390 -3030
rect 270 -3090 280 -3040
rect 1380 -3090 1390 -3040
rect 270 -3100 1390 -3090
rect 1770 -3040 2890 -3030
rect 1770 -3090 1780 -3040
rect 2880 -3090 2890 -3040
rect 1770 -3100 2890 -3090
rect 3270 -3040 4390 -3030
rect 3270 -3090 3280 -3040
rect 4380 -3090 4390 -3040
rect 3270 -3100 4390 -3090
rect 110 -3250 220 -3245
rect 110 -3350 120 -3250
rect 210 -3350 220 -3250
rect 110 -3550 220 -3350
rect 1610 -3250 1720 -3245
rect 1610 -3350 1620 -3250
rect 1710 -3350 1720 -3250
rect 1610 -3550 1720 -3350
rect 3110 -3250 3220 -3245
rect 3110 -3350 3120 -3250
rect 3210 -3350 3220 -3250
rect 3110 -3550 3220 -3350
<< metal5 >>
rect -1000 1420 0 1580
rect 520 520 620 620
rect 2020 520 2120 620
rect 3520 520 3620 620
rect 520 -980 620 -880
rect 2020 -980 2120 -880
rect 3520 -980 3620 -880
rect 520 -2480 620 -2380
rect 2020 -2480 2120 -2380
rect 3520 -2480 3620 -2380
use pixel  pixel_2 ~/CMOS/TopmetalSe/magic
timestamp 1654624193
transform 1 0 1100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_0
timestamp 1654624193
transform 1 0 -1900 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_1
timestamp 1654624193
transform 1 0 -400 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_5
timestamp 1654624193
transform 1 0 1100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_8
timestamp 1654624193
transform 1 0 1100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_3
timestamp 1654624193
transform 1 0 -1900 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_4
timestamp 1654624193
transform 1 0 -400 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_6
timestamp 1654624193
transform 1 0 -1900 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_7
timestamp 1654624193
transform 1 0 -400 0 1 -1650
box 1820 -1430 3480 230
<< labels >>
rlabel metal2 250 1500 285 1800 1 VBIAS
port 202 n
rlabel metal2 30 1500 65 1800 1 VREF
port 203 n
rlabel metal2 510 1500 545 1800 1 NB2
port 204 n
rlabel metal1 -280 1440 20 1485 1 VDD
port 205 n
rlabel metal3 -280 1375 20 1420 1 SF_IB
port 206 n
rlabel metal3 -280 1230 20 1275 1 CSA_VREF
port 207 n
rlabel metal3 -280 80 20 125 1 NB1
port 208 n
rlabel metal3 -280 740 20 785 1 ROW_SEL0
port 209 n
rlabel metal2 1750 1500 1785 1800 1 VBIAS
rlabel metal2 1530 1500 1565 1800 1 VREF
rlabel metal2 2010 1500 2045 1800 1 NB2
rlabel metal2 3250 1500 3285 1800 1 VBIAS
rlabel metal2 3030 1500 3065 1800 1 VREF
rlabel metal2 3510 1500 3545 1800 1 NB2
rlabel metal1 4500 15 4800 60 1 GND
port 212 n
rlabel metal1 -280 -60 20 -15 1 VDD
rlabel metal3 -280 -125 20 -80 1 SF_IB
rlabel metal3 -280 -270 20 -225 1 CSA_VREF
rlabel metal3 -280 -1420 20 -1375 1 NB1
rlabel metal3 -280 -760 20 -715 1 ROW_SEL1
port 214 n
rlabel metal1 4500 -1485 4800 -1440 1 GND
rlabel metal1 -280 -1560 20 -1515 1 VDD
rlabel metal3 -280 -1625 20 -1580 1 SF_IB
rlabel metal3 -280 -1770 20 -1725 1 CSA_VREF
rlabel metal3 -280 -2920 20 -2875 1 NB1
rlabel metal3 -280 -2260 20 -2215 1 ROW_SEL2
port 220 n
rlabel metal1 4500 -2985 4800 -2940 1 GND
rlabel metal4 -500 1775 -500 1775 1 VBIAS
port 202 n
rlabel metal1 -500 1675 -500 1675 3 VREF
port 203 e
rlabel metal2 -1500 740 -1500 740 3 ROW_SEL0
port 209 e
rlabel metal2 -1500 -760 -1500 -760 3 ROW_SEL1
port 214 e
rlabel metal2 -1500 -2260 -1500 -2260 3 ROW_SEL2
port 220 e
rlabel metal5 520 520 620 620 1 PIX0_IN
port 244 n
rlabel metal4 -1500 1775 -1500 1830 1 VBIAS
port 202 n
rlabel metal2 -1500 1675 -1500 1725 3 VREF
port 203 e
rlabel metal2 0 2020 0 2020 1 NB2
port 204 n
rlabel metal1 -1000 0 -1000 0 1 VDD
port 205 n
rlabel space -580 2875 -580 2875 5 SF_IB
port 206 s
rlabel metal2 -370 1780 -370 1780 1 NB1
port 208 n
rlabel metal2 -1500 740 -1500 785 3 ROW_SEL0
port 209 e
rlabel metal5 -1000 1420 -1000 1420 1 GRING
port 245 n
rlabel metal5 2020 520 2120 620 1 PIX1_IN
port 246 n
rlabel metal5 3520 520 3620 620 1 PIX2_IN
port 247 n
rlabel metal1 4700 15 4700 15 1 GND
port 212 n
rlabel metal5 520 -980 620 -880 1 PIX3_IN
port 248 n
rlabel metal2 -1500 -760 -1500 -715 3 ROW_SEL1
port 214 e
rlabel metal5 2020 -980 2120 -880 1 PIX4_IN
port 249 n
rlabel metal5 3520 -980 3620 -880 1 PIX5_IN
port 250 n
rlabel metal5 520 -2480 620 -2380 1 PIX6_IN
port 251 n
rlabel metal4 1315 -3100 1390 -3000 1 PIX_OUT0
port 252 n
rlabel metal4 110 -3550 220 -3350 1 COL_SEL0
port 253 n
rlabel metal4 -240 -3800 -240 -3800 1 CSA_VREF
port 207 n
rlabel metal2 -1500 -2260 -1500 -2215 3 ROW_SEL2
port 220 e
rlabel metal5 2020 -2480 2120 -2380 1 PIX7_IN
port 254 n
rlabel metal4 2815 -3100 2890 -3000 1 PIX_OUT1
port 255 n
rlabel metal4 1610 -3550 1720 -3350 1 COL_SEL1
port 256 n
rlabel metal5 3520 -2480 3620 -2380 1 PIX8_IN
port 257 n
rlabel metal4 4315 -3100 4390 -3000 1 PIX_OUT2
port 258 n
rlabel metal2 4470 -3550 4470 -3550 1 ARRAY_OUT
port 259 n
rlabel metal4 3110 -3550 3220 -3350 1 COL_SEL2
port 260 n
<< end >>
