magic
tech sky130A
magscale 1 2
timestamp 1654646295
<< error_p >>
rect 6863 -221 6897 0
rect 6981 -221 7015 0
rect 7099 -221 7133 0
rect 7217 -221 7251 0
rect 7335 -221 7369 0
rect 7453 -221 7487 0
rect 7571 -221 7605 0
rect 7689 -221 7723 0
rect 7807 -221 7841 0
rect 20160 297 20173 1173
rect 20287 297 20321 1173
rect 20435 297 20469 1173
rect 20583 297 20617 1173
rect 20731 297 20765 1173
rect 20879 297 20913 1173
rect 21027 297 21061 1173
rect 21175 297 21209 1173
rect 21323 297 21357 1173
rect 21471 297 21505 1173
rect 21619 297 21653 1173
rect 21915 297 21949 1173
rect 20201 213 20259 247
rect 20349 213 20407 247
rect 20497 213 20555 247
rect 20645 213 20703 247
rect 20793 213 20851 247
rect 20941 213 20999 247
rect 21089 213 21147 247
rect 21237 213 21295 247
rect 21385 213 21443 247
rect 21533 213 21591 247
rect 21681 213 21739 247
rect 21829 213 21887 247
rect 20201 105 20259 139
rect 20349 105 20407 139
rect 20497 105 20555 139
rect 20645 105 20703 139
rect 20793 105 20851 139
rect 20941 105 20999 139
rect 21089 105 21147 139
rect 21237 105 21295 139
rect 21385 105 21443 139
rect 21533 105 21591 139
rect 21681 105 21739 139
rect 21829 105 21887 139
rect 7925 -221 7959 0
rect 10815 -821 10849 0
rect 10963 -821 10997 0
rect 11111 -821 11145 0
rect 11259 -821 11293 0
rect 11407 -821 11441 0
rect 11555 -821 11589 0
rect 11703 -821 11737 0
rect 11851 -821 11885 0
rect 11999 -821 12033 0
rect 12147 -821 12181 0
rect 12295 -821 12329 0
rect 12443 -821 12477 0
rect 12591 -821 12625 0
rect 12739 -821 12773 0
rect 12887 -821 12921 0
rect 13035 -821 13069 0
rect 13183 -821 13217 0
rect 13331 -821 13365 0
rect 13479 -821 13513 0
rect 13627 -821 13661 0
rect 13775 -821 13809 0
rect 13923 -821 13957 0
rect 14071 -821 14105 0
rect 14219 -821 14253 0
rect 14367 -821 14401 0
rect 14515 -821 14549 0
rect 14663 -821 14697 0
rect 14811 -821 14845 0
rect 14959 -821 14993 0
rect 15107 -821 15141 0
rect 15255 -821 15289 0
rect 15403 -821 15437 0
rect 15551 -821 15585 0
rect 15699 -821 15733 0
rect 15847 -821 15881 0
rect 15995 -821 16029 0
rect 16143 -821 16177 0
rect 16291 -821 16325 0
rect 16439 -821 16473 0
rect 16587 -821 16621 0
rect 16735 -821 16769 0
rect 16883 -821 16917 0
rect 17031 -821 17065 0
rect 17179 -821 17213 0
rect 17327 -821 17361 0
rect 17475 -821 17509 0
rect 17623 -821 17657 0
rect 17771 -821 17805 0
rect 17919 -821 17953 0
rect 18067 -821 18101 0
rect 18215 -821 18249 0
rect 18363 -821 18397 0
rect 18511 -821 18545 0
rect 18659 -821 18693 0
rect 18807 -821 18841 0
rect 18955 -821 18989 0
rect 19103 -821 19137 0
rect 19251 -821 19285 0
rect 19399 -821 19433 0
rect 19547 -821 19581 0
rect 19695 -821 19729 0
rect 19843 -821 19877 0
rect 19991 -821 20025 0
rect 20160 0 20173 55
rect 20139 -821 20173 0
rect 20287 -821 20321 55
rect 20435 -821 20469 55
rect 20583 -821 20617 55
rect 20731 -821 20765 55
rect 20879 -821 20913 55
rect 21027 -821 21061 55
rect 21175 -821 21209 55
rect 21323 -821 21357 55
rect 21471 -821 21505 55
rect 21619 -821 21653 55
<< error_s >>
rect 5679 10487 5713 11063
rect 11017 10486 11051 11062
rect 11135 10486 11169 11062
rect 11253 10486 11287 11062
rect 11371 10486 11405 11062
rect 11489 10486 11523 11062
rect 11607 10486 11641 11062
rect 11725 10486 11759 11062
rect 11843 10486 11877 11062
rect 11961 10486 11995 11062
rect 12079 10486 12113 11062
rect 12197 10486 12231 11062
rect 12315 10486 12349 11062
rect 12433 10486 12467 11062
rect 12551 10486 12585 11062
rect 12669 10486 12703 11062
rect 12787 10486 12821 11062
rect 12905 10486 12939 11062
rect 13023 10486 13057 11062
rect 13141 10486 13175 11062
rect 13259 10486 13293 11062
rect 13377 10486 13411 11062
rect 13495 10486 13529 11062
rect 13613 10486 13647 11062
rect 13731 10486 13765 11062
rect 15140 10486 15174 11062
rect 15258 10486 15292 11062
rect 15376 10486 15410 11062
rect 15494 10486 15528 11062
rect 15612 10486 15646 11062
rect 15730 10486 15764 11062
rect 15848 10486 15882 11062
rect 15966 10486 16000 11062
rect 16084 10486 16118 11062
rect 16202 10486 16236 11062
rect 16320 10486 16354 11062
rect 16438 10486 16472 11062
rect 16556 10486 16590 11062
rect 16674 10486 16708 11062
rect 16792 10486 16826 11062
rect 16910 10486 16944 11062
rect 17028 10486 17062 11062
rect 17146 10486 17180 11062
rect 17264 10486 17298 11062
rect 17382 10486 17416 11062
rect 17500 10486 17534 11062
rect 17618 10486 17652 11062
rect 17736 10486 17770 11062
rect 17854 10486 17888 11062
rect 19263 10486 19297 11062
rect 19381 10486 19415 11062
rect 19499 10486 19533 11062
rect 19617 10486 19651 11062
rect 19735 10486 19769 11062
rect 19853 10486 19887 11062
rect 19971 10486 20005 11062
rect 20089 10486 20123 11062
rect 20207 10486 20241 11062
rect 20325 10486 20359 11062
rect 20443 10486 20477 11062
rect 20561 10486 20595 11062
rect 20679 10486 20713 11062
rect 20797 10486 20831 11062
rect 20915 10486 20949 11062
rect 21033 10486 21067 11062
rect 21151 10486 21185 11062
rect 21269 10486 21303 11062
rect 21387 10486 21421 11062
rect 21505 10486 21539 11062
rect 21623 10486 21657 11062
rect 21741 10486 21775 11062
rect 21859 10486 21893 11062
rect 21977 10486 22011 11062
rect 3073 9727 9043 9761
rect 2977 8055 3011 9665
rect 3091 8990 3125 9566
rect 3209 8990 3243 9566
rect 3327 8990 3361 9566
rect 3445 8990 3479 9566
rect 3563 8990 3597 9566
rect 3681 8990 3715 9566
rect 3799 8990 3833 9566
rect 3917 8990 3951 9566
rect 4035 8990 4069 9566
rect 4153 8990 4187 9566
rect 4271 8990 4305 9566
rect 4389 8990 4423 9566
rect 4507 8990 4541 9566
rect 4625 8990 4659 9566
rect 4743 8990 4777 9566
rect 4861 8990 4895 9566
rect 4979 8990 5013 9566
rect 5097 8990 5131 9566
rect 5215 8990 5249 9566
rect 5333 8990 5367 9566
rect 5451 8990 5485 9566
rect 5569 8990 5603 9566
rect 5687 8990 5721 9566
rect 5805 8990 5839 9566
rect 5923 8990 5957 9566
rect 6041 8990 6075 9566
rect 6159 8990 6193 9566
rect 6277 8990 6311 9566
rect 6395 8990 6429 9566
rect 6513 8990 6547 9566
rect 6631 8990 6665 9566
rect 6749 8990 6783 9566
rect 6867 8990 6901 9566
rect 6985 8990 7019 9566
rect 7103 8990 7137 9566
rect 7221 8990 7255 9566
rect 7339 8990 7373 9566
rect 7457 8990 7491 9566
rect 7575 8990 7609 9566
rect 7693 8990 7727 9566
rect 7811 8990 7845 9566
rect 7929 8990 7963 9566
rect 8047 8990 8081 9566
rect 8165 8990 8199 9566
rect 8283 8990 8317 9566
rect 8401 8990 8435 9566
rect 8519 8990 8553 9566
rect 8637 8990 8671 9566
rect 8755 8990 8789 9566
rect 8873 8990 8907 9566
rect 8991 8990 9025 9566
rect 3091 8154 3125 8730
rect 3209 8154 3243 8730
rect 3327 8154 3361 8730
rect 3445 8154 3479 8730
rect 3563 8154 3597 8730
rect 3681 8154 3715 8730
rect 3799 8154 3833 8730
rect 3917 8154 3951 8730
rect 4035 8154 4069 8730
rect 4153 8154 4187 8730
rect 4271 8154 4305 8730
rect 4389 8154 4423 8730
rect 4507 8154 4541 8730
rect 4625 8154 4659 8730
rect 4743 8154 4777 8730
rect 4861 8154 4895 8730
rect 4979 8154 5013 8730
rect 5097 8154 5131 8730
rect 5215 8154 5249 8730
rect 5333 8154 5367 8730
rect 5451 8154 5485 8730
rect 5569 8154 5603 8730
rect 5687 8154 5721 8730
rect 5805 8154 5839 8730
rect 5923 8154 5957 8730
rect 6041 8154 6075 8730
rect 6159 8154 6193 8730
rect 6277 8154 6311 8730
rect 6395 8154 6429 8730
rect 6513 8154 6547 8730
rect 6631 8154 6665 8730
rect 6749 8154 6783 8730
rect 6867 8154 6901 8730
rect 6985 8154 7019 8730
rect 7103 8154 7137 8730
rect 7221 8154 7255 8730
rect 7339 8154 7373 8730
rect 7457 8154 7491 8730
rect 7575 8154 7609 8730
rect 7693 8154 7727 8730
rect 7811 8154 7845 8730
rect 7929 8154 7963 8730
rect 8047 8154 8081 8730
rect 8165 8154 8199 8730
rect 8283 8154 8317 8730
rect 8401 8154 8435 8730
rect 8519 8154 8553 8730
rect 8637 8154 8671 8730
rect 8755 8154 8789 8730
rect 8873 8154 8907 8730
rect 8991 8154 9025 8730
rect 9105 8055 9139 9665
rect 10781 9650 10815 10226
rect 10899 9650 10933 10226
rect 11017 9650 11051 10226
rect 11135 9650 11169 10226
rect 11253 9650 11287 10226
rect 11371 9650 11405 10226
rect 11489 9650 11523 10226
rect 11607 9650 11641 10226
rect 11725 9650 11759 10226
rect 11843 9650 11877 10226
rect 11961 9650 11995 10226
rect 12079 9650 12113 10226
rect 12197 9650 12231 10226
rect 12315 9650 12349 10226
rect 12433 9650 12467 10226
rect 12551 9650 12585 10226
rect 12669 9650 12703 10226
rect 12787 9650 12821 10226
rect 12905 9650 12939 10226
rect 13023 9650 13057 10226
rect 13141 9650 13175 10226
rect 13259 9650 13293 10226
rect 13377 9650 13411 10226
rect 13495 9650 13529 10226
rect 13613 9650 13647 10226
rect 13731 9650 13765 10226
rect 14904 9650 14938 10226
rect 15022 9650 15056 10226
rect 15140 9650 15174 10226
rect 15258 9650 15292 10226
rect 15376 9650 15410 10226
rect 15494 9650 15528 10226
rect 15612 9650 15646 10226
rect 15730 9650 15764 10226
rect 15848 9650 15882 10226
rect 15966 9650 16000 10226
rect 16084 9650 16118 10226
rect 16202 9650 16236 10226
rect 16320 9650 16354 10226
rect 16438 9650 16472 10226
rect 16556 9650 16590 10226
rect 16674 9650 16708 10226
rect 16792 9650 16826 10226
rect 16910 9650 16944 10226
rect 17028 9650 17062 10226
rect 17146 9650 17180 10226
rect 17264 9650 17298 10226
rect 17382 9650 17416 10226
rect 17500 9650 17534 10226
rect 17618 9650 17652 10226
rect 17736 9650 17770 10226
rect 17854 9650 17888 10226
rect 19027 9650 19061 10226
rect 19145 9650 19179 10226
rect 19263 9650 19297 10226
rect 19381 9650 19415 10226
rect 19499 9650 19533 10226
rect 19617 9650 19651 10226
rect 19735 9650 19769 10226
rect 19853 9650 19887 10226
rect 19971 9650 20005 10226
rect 20089 9650 20123 10226
rect 20207 9650 20241 10226
rect 20325 9650 20359 10226
rect 20443 9650 20477 10226
rect 20561 9650 20595 10226
rect 20679 9650 20713 10226
rect 20797 9650 20831 10226
rect 20915 9650 20949 10226
rect 21033 9650 21067 10226
rect 21151 9650 21185 10226
rect 21269 9650 21303 10226
rect 21387 9650 21421 10226
rect 21505 9650 21539 10226
rect 21623 9650 21657 10226
rect 21741 9650 21775 10226
rect 21859 9650 21893 10226
rect 21977 9650 22011 10226
rect 3073 7959 9043 7993
rect 3073 7677 9043 7711
rect 2977 6005 3011 7615
rect 3091 6940 3125 7516
rect 3209 6940 3243 7516
rect 3327 6940 3361 7516
rect 3445 6940 3479 7516
rect 3563 6940 3597 7516
rect 3681 6940 3715 7516
rect 3799 6940 3833 7516
rect 3917 6940 3951 7516
rect 4035 6940 4069 7516
rect 4153 6940 4187 7516
rect 4271 6940 4305 7516
rect 4389 6940 4423 7516
rect 4507 6940 4541 7516
rect 4625 6940 4659 7516
rect 4743 6940 4777 7516
rect 4861 6940 4895 7516
rect 4979 6940 5013 7516
rect 5097 6940 5131 7516
rect 5215 6940 5249 7516
rect 5333 6940 5367 7516
rect 5451 6940 5485 7516
rect 5569 6940 5603 7516
rect 5687 6940 5721 7516
rect 5805 6940 5839 7516
rect 5923 6940 5957 7516
rect 6041 6940 6075 7516
rect 6159 6940 6193 7516
rect 6277 6940 6311 7516
rect 6395 6940 6429 7516
rect 6513 6940 6547 7516
rect 6631 6940 6665 7516
rect 6749 6940 6783 7516
rect 6867 6940 6901 7516
rect 6985 6940 7019 7516
rect 7103 6940 7137 7516
rect 7221 6940 7255 7516
rect 7339 6940 7373 7516
rect 7457 6940 7491 7516
rect 7575 6940 7609 7516
rect 7693 6940 7727 7516
rect 7811 6940 7845 7516
rect 7929 6940 7963 7516
rect 8047 6940 8081 7516
rect 8165 6940 8199 7516
rect 8283 6940 8317 7516
rect 8401 6940 8435 7516
rect 8519 6940 8553 7516
rect 8637 6940 8671 7516
rect 8755 6940 8789 7516
rect 8873 6940 8907 7516
rect 8991 6940 9025 7516
rect 3091 6104 3125 6680
rect 3209 6104 3243 6680
rect 3327 6104 3361 6680
rect 3445 6104 3479 6680
rect 3563 6104 3597 6680
rect 3681 6104 3715 6680
rect 3799 6104 3833 6680
rect 3917 6104 3951 6680
rect 4035 6104 4069 6680
rect 4153 6104 4187 6680
rect 4271 6104 4305 6680
rect 4389 6104 4423 6680
rect 4507 6104 4541 6680
rect 4625 6104 4659 6680
rect 4743 6104 4777 6680
rect 4861 6104 4895 6680
rect 4979 6104 5013 6680
rect 5097 6104 5131 6680
rect 5215 6104 5249 6680
rect 5333 6104 5367 6680
rect 5451 6104 5485 6680
rect 5569 6104 5603 6680
rect 5687 6104 5721 6680
rect 5805 6104 5839 6680
rect 5923 6104 5957 6680
rect 6041 6104 6075 6680
rect 6159 6104 6193 6680
rect 6277 6104 6311 6680
rect 6395 6104 6429 6680
rect 6513 6104 6547 6680
rect 6631 6104 6665 6680
rect 6749 6104 6783 6680
rect 6867 6104 6901 6680
rect 6985 6104 7019 6680
rect 7103 6104 7137 6680
rect 7221 6104 7255 6680
rect 7339 6104 7373 6680
rect 7457 6104 7491 6680
rect 7575 6104 7609 6680
rect 7693 6104 7727 6680
rect 7811 6104 7845 6680
rect 7929 6104 7963 6680
rect 8047 6104 8081 6680
rect 8165 6104 8199 6680
rect 8283 6104 8317 6680
rect 8401 6104 8435 6680
rect 8519 6104 8553 6680
rect 8637 6104 8671 6680
rect 8755 6104 8789 6680
rect 8873 6104 8907 6680
rect 8991 6104 9025 6680
rect 9105 6005 9139 7615
rect 3073 5909 9043 5943
rect 3073 5627 9043 5661
rect 2977 3955 3011 5565
rect 3091 4890 3125 5466
rect 3209 4890 3243 5466
rect 3327 4890 3361 5466
rect 3445 4890 3479 5466
rect 3563 4890 3597 5466
rect 3681 4890 3715 5466
rect 3799 4890 3833 5466
rect 3917 4890 3951 5466
rect 4035 4890 4069 5466
rect 4153 4890 4187 5466
rect 4271 4890 4305 5466
rect 4389 4890 4423 5466
rect 4507 4890 4541 5466
rect 4625 4890 4659 5466
rect 4743 4890 4777 5466
rect 4861 4890 4895 5466
rect 4979 4890 5013 5466
rect 5097 4890 5131 5466
rect 5215 4890 5249 5466
rect 5333 4890 5367 5466
rect 5451 4890 5485 5466
rect 5569 4890 5603 5466
rect 5687 4890 5721 5466
rect 5805 4890 5839 5466
rect 5923 4890 5957 5466
rect 6041 4890 6075 5466
rect 6159 4890 6193 5466
rect 6277 4890 6311 5466
rect 6395 4890 6429 5466
rect 6513 4890 6547 5466
rect 6631 4890 6665 5466
rect 6749 4890 6783 5466
rect 6867 4890 6901 5466
rect 6985 4890 7019 5466
rect 7103 4890 7137 5466
rect 7221 4890 7255 5466
rect 7339 4890 7373 5466
rect 7457 4890 7491 5466
rect 7575 4890 7609 5466
rect 7693 4890 7727 5466
rect 7811 4890 7845 5466
rect 7929 4890 7963 5466
rect 8047 4890 8081 5466
rect 8165 4890 8199 5466
rect 8283 4890 8317 5466
rect 8401 4890 8435 5466
rect 8519 4890 8553 5466
rect 8637 4890 8671 5466
rect 8755 4890 8789 5466
rect 8873 4890 8907 5466
rect 8991 4890 9025 5466
rect 3091 4054 3125 4630
rect 3209 4054 3243 4630
rect 3327 4054 3361 4630
rect 3445 4054 3479 4630
rect 3563 4054 3597 4630
rect 3681 4054 3715 4630
rect 3799 4054 3833 4630
rect 3917 4054 3951 4630
rect 4035 4054 4069 4630
rect 4153 4054 4187 4630
rect 4271 4054 4305 4630
rect 4389 4054 4423 4630
rect 4507 4054 4541 4630
rect 4625 4054 4659 4630
rect 4743 4054 4777 4630
rect 4861 4054 4895 4630
rect 4979 4054 5013 4630
rect 5097 4054 5131 4630
rect 5215 4054 5249 4630
rect 5333 4054 5367 4630
rect 5451 4054 5485 4630
rect 5569 4054 5603 4630
rect 5687 4054 5721 4630
rect 5805 4054 5839 4630
rect 5923 4054 5957 4630
rect 6041 4054 6075 4630
rect 6159 4054 6193 4630
rect 6277 4054 6311 4630
rect 6395 4054 6429 4630
rect 6513 4054 6547 4630
rect 6631 4054 6665 4630
rect 6749 4054 6783 4630
rect 6867 4054 6901 4630
rect 6985 4054 7019 4630
rect 7103 4054 7137 4630
rect 7221 4054 7255 4630
rect 7339 4054 7373 4630
rect 7457 4054 7491 4630
rect 7575 4054 7609 4630
rect 7693 4054 7727 4630
rect 7811 4054 7845 4630
rect 7929 4054 7963 4630
rect 8047 4054 8081 4630
rect 8165 4054 8199 4630
rect 8283 4054 8317 4630
rect 8401 4054 8435 4630
rect 8519 4054 8553 4630
rect 8637 4054 8671 4630
rect 8755 4054 8789 4630
rect 8873 4054 8907 4630
rect 8991 4054 9025 4630
rect 9105 3955 9139 5565
rect 3073 3859 9043 3893
rect 3327 2840 3361 3416
rect 3445 2840 3479 3416
rect 3563 2840 3597 3416
rect 3681 2840 3715 3416
rect 3799 2840 3833 3416
rect 3917 2840 3951 3416
rect 4035 2840 4069 3416
rect 4153 2840 4187 3416
rect 4271 2840 4305 3416
rect 4389 2840 4423 3416
rect 4507 2840 4541 3416
rect 4625 2840 4659 3416
rect 4743 2840 4777 3416
rect 4861 2840 4895 3416
rect 4979 2840 5013 3416
rect 5097 2840 5131 3416
rect 5215 2840 5249 3416
rect 5333 2840 5367 3416
rect 5451 2840 5485 3416
rect 5569 2840 5603 3416
rect 5687 2840 5721 3416
rect 5805 2840 5839 3416
rect 5923 2840 5957 3416
rect 6041 2840 6075 3416
rect 6159 2840 6193 3416
rect 6277 2840 6311 3416
rect 6395 2840 6429 3416
rect 6513 2840 6547 3416
rect 6631 2840 6665 3416
rect 6749 2840 6783 3416
rect 6867 2840 6901 3416
rect 6985 2840 7019 3416
rect 7103 2840 7137 3416
rect 7221 2840 7255 3416
rect 7339 2840 7373 3416
rect 7457 2840 7491 3416
rect 7575 2840 7609 3416
rect 7693 2840 7727 3416
rect 7811 2840 7845 3416
rect 7929 2840 7963 3416
rect 8047 2840 8081 3416
rect 8165 2840 8199 3416
rect 8283 2840 8317 3416
rect 8401 2840 8435 3416
rect 8519 2840 8553 3416
rect 8637 2840 8671 3416
rect 8755 2840 8789 3416
rect 8873 2840 8907 3416
rect 8991 2840 9025 3416
rect 3091 2004 3125 2580
rect 3209 2004 3243 2580
rect 3327 2004 3361 2580
rect 3445 2004 3479 2580
rect 3563 2004 3597 2580
rect 3681 2004 3715 2580
rect 3799 2004 3833 2580
rect 3917 2004 3951 2580
rect 4035 2004 4069 2580
rect 4153 2004 4187 2580
rect 4271 2004 4305 2580
rect 4389 2004 4423 2580
rect 4507 2004 4541 2580
rect 4625 2004 4659 2580
rect 4743 2004 4777 2580
rect 4861 2004 4895 2580
rect 4979 2004 5013 2580
rect 5097 2004 5131 2580
rect 5215 2004 5249 2580
rect 5333 2004 5367 2580
rect 5451 2004 5485 2580
rect 5569 2004 5603 2580
rect 5687 2004 5721 2580
rect 5805 2004 5839 2580
rect 5923 2004 5957 2580
rect 6041 2004 6075 2580
rect 6159 2004 6193 2580
rect 6277 2004 6311 2580
rect 6395 2004 6429 2580
rect 6513 2004 6547 2580
rect 6631 2004 6665 2580
rect 6749 2004 6783 2580
rect 6867 2004 6901 2580
rect 6985 2004 7019 2580
rect 7103 2004 7137 2580
rect 7221 2004 7255 2580
rect 7339 2004 7373 2580
rect 7457 2004 7491 2580
rect 7575 2004 7609 2580
rect 7693 2004 7727 2580
rect 7811 2004 7845 2580
rect 7929 2004 7963 2580
rect 8047 2004 8081 2580
rect 8165 2004 8199 2580
rect 8283 2004 8317 2580
rect 8401 2004 8435 2580
rect 8519 2004 8553 2580
rect 8637 2004 8671 2580
rect 8755 2004 8789 2580
rect 8873 2004 8907 2580
rect 8991 2004 9025 2580
rect 4393 597 4427 1173
rect 4511 597 4545 1173
rect 4629 597 4663 1173
rect 4747 597 4781 1173
rect 4865 597 4899 1173
rect 4983 597 5017 1173
rect 5101 597 5135 1173
rect 5219 597 5253 1173
rect 5337 597 5371 1173
rect 5455 597 5489 1173
rect 5573 597 5607 1173
rect 5691 597 5725 1173
rect 5809 597 5843 1173
rect 5927 597 5961 1173
rect 6155 597 6189 1173
rect 6273 597 6307 1173
rect 6391 597 6425 1173
rect 6509 597 6543 1173
rect 6627 597 6661 1173
rect 6745 597 6779 1173
rect 6863 597 6897 1173
rect 6981 597 7015 1173
rect 7099 597 7133 1173
rect 7217 597 7251 1173
rect 7335 597 7369 1173
rect 7453 597 7487 1173
rect 7571 597 7605 1173
rect 7689 597 7723 1173
rect 7807 597 7841 1173
rect 7925 597 7959 1173
rect 9018 795 9052 1101
rect 9132 885 9166 1011
rect 9220 885 9254 1011
rect 9334 795 9368 1101
rect 9448 885 9482 1011
rect 9536 885 9570 1011
rect 9650 795 9684 1101
rect 9764 885 9798 1011
rect 9852 885 9886 1011
rect 9966 795 10000 1101
rect 10080 885 10114 1011
rect 10168 885 10202 1011
rect 10282 795 10316 1101
rect 10396 885 10430 1011
rect 10484 885 10518 1011
rect 10598 795 10632 1101
rect 4157 0 4191 355
rect 4275 0 4309 355
rect 4393 0 4427 355
rect 4511 0 4545 355
rect 4629 0 4663 355
rect 4747 0 4781 355
rect 4865 0 4899 355
rect 4983 0 5017 355
rect 5101 0 5135 355
rect 5219 0 5253 355
rect 5337 0 5371 355
rect 5455 0 5489 355
rect 5573 0 5607 355
rect 5691 0 5725 355
rect 5809 0 5843 355
rect 5927 0 5961 355
rect 6155 0 6189 355
rect 6273 0 6307 355
rect 6391 0 6425 355
rect 6509 0 6543 355
rect 6627 0 6661 355
rect 6745 0 6779 355
rect 6863 0 6897 355
rect 6981 0 7015 355
rect 7099 0 7133 355
rect 7217 0 7251 355
rect 7335 0 7369 355
rect 7453 0 7487 355
rect 7571 0 7605 355
rect 7689 0 7723 355
rect 7807 0 7841 355
rect 7925 0 7959 355
rect 10815 297 10849 1173
rect 10963 297 10997 1173
rect 11111 297 11145 1173
rect 11259 297 11293 1173
rect 11407 297 11441 1173
rect 11555 297 11589 1173
rect 11703 297 11737 1173
rect 11851 297 11885 1173
rect 11999 297 12033 1173
rect 12147 297 12181 1173
rect 12295 297 12329 1173
rect 12443 297 12477 1173
rect 12591 297 12625 1173
rect 12739 297 12773 1173
rect 12887 297 12921 1173
rect 13035 297 13069 1173
rect 13183 297 13217 1173
rect 13331 297 13365 1173
rect 13479 297 13513 1173
rect 13627 297 13661 1173
rect 13775 297 13809 1173
rect 13923 297 13957 1173
rect 14071 297 14105 1173
rect 14219 297 14253 1173
rect 14367 297 14401 1173
rect 14515 297 14549 1173
rect 14663 297 14697 1173
rect 14811 297 14845 1173
rect 14959 297 14993 1173
rect 15107 297 15141 1173
rect 15255 297 15289 1173
rect 15403 297 15437 1173
rect 15551 297 15585 1173
rect 15699 297 15733 1173
rect 15847 297 15881 1173
rect 15995 297 16029 1173
rect 16143 297 16177 1173
rect 16291 297 16325 1173
rect 16439 297 16473 1173
rect 16587 297 16621 1173
rect 16735 297 16769 1173
rect 16883 297 16917 1173
rect 17031 297 17065 1173
rect 17179 297 17213 1173
rect 17327 297 17361 1173
rect 17475 297 17509 1173
rect 17623 297 17657 1173
rect 17771 297 17805 1173
rect 17919 297 17953 1173
rect 18067 297 18101 1173
rect 18215 297 18249 1173
rect 18363 297 18397 1173
rect 18511 297 18545 1173
rect 18659 297 18693 1173
rect 18807 297 18841 1173
rect 18955 297 18989 1173
rect 19103 297 19137 1173
rect 19251 297 19285 1173
rect 19399 297 19433 1173
rect 19547 297 19581 1173
rect 19695 297 19729 1173
rect 19843 297 19877 1173
rect 19991 297 20025 1173
rect 20139 297 20160 1173
rect 11025 213 11083 247
rect 11173 213 11231 247
rect 11321 213 11379 247
rect 11469 213 11527 247
rect 11617 213 11675 247
rect 11765 213 11823 247
rect 11913 213 11971 247
rect 12061 213 12119 247
rect 12209 213 12267 247
rect 12357 213 12415 247
rect 12505 213 12563 247
rect 12653 213 12711 247
rect 12801 213 12859 247
rect 12949 213 13007 247
rect 13097 213 13155 247
rect 13245 213 13303 247
rect 13393 213 13451 247
rect 13541 213 13599 247
rect 13689 213 13747 247
rect 13837 213 13895 247
rect 13985 213 14043 247
rect 14133 213 14191 247
rect 14281 213 14339 247
rect 14429 213 14487 247
rect 14577 213 14635 247
rect 14725 213 14783 247
rect 14873 213 14931 247
rect 15021 213 15079 247
rect 15169 213 15227 247
rect 15317 213 15375 247
rect 15465 213 15523 247
rect 15613 213 15671 247
rect 15761 213 15819 247
rect 15909 213 15967 247
rect 16057 213 16115 247
rect 16205 213 16263 247
rect 16353 213 16411 247
rect 16501 213 16559 247
rect 16649 213 16707 247
rect 16797 213 16855 247
rect 16945 213 17003 247
rect 17093 213 17151 247
rect 17241 213 17299 247
rect 17389 213 17447 247
rect 17537 213 17595 247
rect 17685 213 17743 247
rect 17833 213 17891 247
rect 17981 213 18039 247
rect 18129 213 18187 247
rect 18277 213 18335 247
rect 18425 213 18483 247
rect 18573 213 18631 247
rect 18721 213 18779 247
rect 18869 213 18927 247
rect 19017 213 19075 247
rect 19165 213 19223 247
rect 19313 213 19371 247
rect 19461 213 19519 247
rect 19609 213 19667 247
rect 19757 213 19815 247
rect 19905 213 19963 247
rect 20053 213 20111 247
rect 11025 105 11083 139
rect 11173 105 11231 139
rect 11321 105 11379 139
rect 11469 105 11527 139
rect 11617 105 11675 139
rect 11765 105 11823 139
rect 11913 105 11971 139
rect 12061 105 12119 139
rect 12209 105 12267 139
rect 12357 105 12415 139
rect 12505 105 12563 139
rect 12653 105 12711 139
rect 12801 105 12859 139
rect 12949 105 13007 139
rect 13097 105 13155 139
rect 13245 105 13303 139
rect 13393 105 13451 139
rect 13541 105 13599 139
rect 13689 105 13747 139
rect 13837 105 13895 139
rect 13985 105 14043 139
rect 14133 105 14191 139
rect 14281 105 14339 139
rect 14429 105 14487 139
rect 14577 105 14635 139
rect 14725 105 14783 139
rect 14873 105 14931 139
rect 15021 105 15079 139
rect 15169 105 15227 139
rect 15317 105 15375 139
rect 15465 105 15523 139
rect 15613 105 15671 139
rect 15761 105 15819 139
rect 15909 105 15967 139
rect 16057 105 16115 139
rect 16205 105 16263 139
rect 16353 105 16411 139
rect 16501 105 16559 139
rect 16649 105 16707 139
rect 16797 105 16855 139
rect 16945 105 17003 139
rect 17093 105 17151 139
rect 17241 105 17299 139
rect 17389 105 17447 139
rect 17537 105 17595 139
rect 17685 105 17743 139
rect 17833 105 17891 139
rect 17981 105 18039 139
rect 18129 105 18187 139
rect 18277 105 18335 139
rect 18425 105 18483 139
rect 18573 105 18631 139
rect 18721 105 18779 139
rect 18869 105 18927 139
rect 19017 105 19075 139
rect 19165 105 19223 139
rect 19313 105 19371 139
rect 19461 105 19519 139
rect 19609 105 19667 139
rect 19757 105 19815 139
rect 19905 105 19963 139
rect 20053 105 20111 139
rect 10815 0 10849 55
rect 10963 0 10997 55
rect 11111 0 11145 55
rect 11259 0 11293 55
rect 11407 0 11441 55
rect 11555 0 11589 55
rect 11703 0 11737 55
rect 11851 0 11885 55
rect 11999 0 12033 55
rect 12147 0 12181 55
rect 12295 0 12329 55
rect 12443 0 12477 55
rect 12591 0 12625 55
rect 12739 0 12773 55
rect 12887 0 12921 55
rect 13035 0 13069 55
rect 13183 0 13217 55
rect 13331 0 13365 55
rect 13479 0 13513 55
rect 13627 0 13661 55
rect 13775 0 13809 55
rect 13923 0 13957 55
rect 14071 0 14105 55
rect 14219 0 14253 55
rect 14367 0 14401 55
rect 14515 0 14549 55
rect 14663 0 14697 55
rect 14811 0 14845 55
rect 14959 0 14993 55
rect 15107 0 15141 55
rect 15255 0 15289 55
rect 15403 0 15437 55
rect 15551 0 15585 55
rect 15699 0 15733 55
rect 15847 0 15881 55
rect 15995 0 16029 55
rect 16143 0 16177 55
rect 16291 0 16325 55
rect 16439 0 16473 55
rect 16587 0 16621 55
rect 16735 0 16769 55
rect 16883 0 16917 55
rect 17031 0 17065 55
rect 17179 0 17213 55
rect 17327 0 17361 55
rect 17475 0 17509 55
rect 17623 0 17657 55
rect 17771 0 17805 55
rect 17919 0 17953 55
rect 18067 0 18101 55
rect 18215 0 18249 55
rect 18363 0 18397 55
rect 18511 0 18545 55
rect 18659 0 18693 55
rect 18807 0 18841 55
rect 18955 0 18989 55
rect 19103 0 19137 55
rect 19251 0 19285 55
rect 19399 0 19433 55
rect 19547 0 19581 55
rect 19695 0 19729 55
rect 19843 0 19877 55
rect 19991 0 20025 55
rect 20139 0 20160 55
<< error_ps >>
rect 4157 -221 4191 0
rect 4275 -221 4309 0
rect 4393 -221 4427 0
rect 4511 -221 4545 0
rect 4629 -221 4663 0
rect 4747 -221 4781 0
rect 4865 -221 4899 0
rect 4983 -221 5017 0
rect 5101 -221 5135 0
rect 5219 -221 5253 0
rect 5337 -221 5371 0
rect 5455 -221 5489 0
rect 5573 -221 5607 0
rect 5691 -221 5725 0
rect 5809 -221 5843 0
rect 5927 -221 5961 0
rect 6155 -221 6189 0
rect 6273 -221 6307 0
rect 6391 -221 6425 0
rect 6509 -221 6543 0
rect 6627 -221 6661 0
rect 6745 -221 6779 0
<< pwell >>
rect -976 9244 676 10696
rect 254 -1586 1906 -94
<< nmoslvt >>
rect -950 9870 650 10270
rect 280 -850 1880 -450
<< ndiff >>
rect -950 10608 650 10670
rect -950 10302 -915 10608
rect 615 10302 650 10608
rect -950 10270 650 10302
rect -950 9815 650 9870
rect -950 9645 -915 9815
rect 615 9645 650 9815
rect -950 9610 650 9645
rect 280 -161 1880 -120
rect 280 -399 315 -161
rect 1845 -399 1880 -161
rect 280 -450 1880 -399
rect 280 -880 1880 -850
rect 280 -1050 315 -880
rect 1845 -1050 1880 -880
rect 280 -1080 1880 -1050
<< ndiffc >>
rect -915 10302 615 10608
rect -915 9645 615 9815
rect 315 -399 1845 -161
rect 315 -1050 1845 -880
<< psubdiff >>
rect -950 9559 650 9610
rect -950 9321 -915 9559
rect 615 9321 650 9559
rect -950 9270 650 9321
rect 280 -1116 1880 -1080
rect 280 -1354 315 -1116
rect 1845 -1354 1880 -1116
rect 280 -1560 1880 -1354
<< psubdiffcont >>
rect -915 9321 615 9559
rect 315 -1354 1845 -1116
<< poly >>
rect -980 10080 -950 10270
rect -1370 10060 -950 10080
rect -1370 9890 -1325 10060
rect -1155 9890 -950 10060
rect -1370 9870 -950 9890
rect 650 9870 680 10270
rect -110 -240 100 -230
rect -110 -410 -66 -240
rect 36 -410 100 -240
rect -110 -450 100 -410
rect -110 -500 280 -450
rect 250 -850 280 -500
rect 1880 -850 1910 -450
<< polycont >>
rect -1325 9890 -1155 10060
rect -66 -410 36 -240
<< locali >>
rect -950 10616 650 10650
rect -950 10294 -923 10616
rect 623 10294 650 10616
rect -950 10270 650 10294
rect -1690 10028 -1325 10060
rect -1155 10028 -1020 10060
rect -1690 9922 -1660 10028
rect -1050 9922 -1020 10028
rect -1690 9890 -1325 9922
rect -1155 9890 -1020 9922
rect -950 9815 650 9850
rect -950 9768 -915 9815
rect 615 9768 650 9815
rect -950 9302 -923 9768
rect 623 9302 650 9768
rect -950 9270 650 9302
rect 280 53 1880 60
rect -400 -272 -66 -240
rect -400 -378 -375 -272
rect -125 -378 -66 -272
rect -400 -410 -66 -378
rect 36 -410 100 -240
rect 280 -413 307 53
rect 1853 -413 1880 53
rect 280 -430 1880 -413
rect 280 -880 1880 -870
rect 280 -1050 315 -880
rect 1845 -1050 1880 -880
rect 280 -1116 1880 -1050
rect 280 -1326 315 -1116
rect 1845 -1326 1880 -1116
rect 280 -1504 307 -1326
rect 1853 -1504 1880 -1326
rect 280 -1550 1880 -1504
<< viali >>
rect -923 10608 623 10616
rect -923 10302 -915 10608
rect -915 10302 615 10608
rect 615 10302 623 10608
rect -923 10294 623 10302
rect -1660 9922 -1325 10028
rect -1325 9922 -1155 10028
rect -1155 9922 -1050 10028
rect -923 9645 -915 9768
rect -915 9645 615 9768
rect 615 9645 623 9768
rect -923 9559 623 9645
rect -923 9321 -915 9559
rect -915 9321 615 9559
rect 615 9321 623 9559
rect -923 9302 623 9321
rect -375 -378 -125 -272
rect 307 -161 1853 53
rect 307 -399 315 -161
rect 315 -399 1845 -161
rect 1845 -399 1853 -161
rect 307 -413 1853 -399
rect 307 -1354 315 -1326
rect 315 -1354 1845 -1326
rect 1845 -1354 1853 -1326
rect 307 -1504 1853 -1354
<< metal1 >>
rect 23020 11280 26995 11570
rect -950 10616 650 10630
rect -950 10294 -923 10616
rect 623 10294 650 10616
rect -950 10270 650 10294
rect -2210 10040 -1020 10060
rect -2210 9910 -2200 10040
rect -1030 9910 -1020 10040
rect -2210 9890 -1020 9910
rect -960 9768 650 9850
rect -960 9302 -923 9768
rect 623 9302 650 9768
rect -960 9220 650 9302
rect 280 53 1880 180
rect -500 -272 100 -240
rect -500 -388 -486 -272
rect -114 -388 100 -272
rect -500 -410 100 -388
rect 280 -413 307 53
rect 1853 -413 1880 53
rect 280 -430 1880 -413
rect -950 -1298 2500 -1280
rect -950 -1542 -914 -1298
rect 2274 -1542 2500 -1298
rect -950 -1560 2500 -1542
rect 24530 -1570 26980 -1270
<< via1 >>
rect -912 10301 612 10609
rect -2200 10028 -1030 10040
rect -2200 9922 -1660 10028
rect -1660 9922 -1050 10028
rect -1050 9922 -1030 10028
rect -2200 9910 -1030 9922
rect -912 9317 612 9753
rect -486 -378 -375 -272
rect -375 -378 -125 -272
rect -125 -378 -114 -272
rect -486 -388 -114 -378
rect 318 -398 1842 38
rect -914 -1326 2274 -1298
rect -914 -1504 307 -1326
rect 307 -1504 1853 -1326
rect 1853 -1504 2274 -1326
rect -914 -1542 2274 -1504
<< metal2 >>
rect -950 10609 650 10630
rect -950 10301 -912 10609
rect 612 10301 650 10609
rect -950 10270 650 10301
rect -950 10269 529 10270
rect -2280 10040 -1020 10060
rect -2280 9910 -2200 10040
rect -1030 9910 -1020 10040
rect -2280 9890 -1020 9910
rect -960 9763 650 9850
rect -960 9753 -898 9763
rect 598 9753 650 9763
rect -960 9317 -912 9753
rect 612 9317 650 9753
rect -960 9307 -898 9317
rect 598 9307 650 9317
rect -960 9220 650 9307
rect 1300 8348 2520 8450
rect 1300 7732 1357 8348
rect 2453 7732 2520 8348
rect 1300 7620 2520 7732
rect 280 3859 1890 3870
rect -1688 3611 2174 3859
rect 280 38 1890 3611
rect -1925 -260 -100 -240
rect -1925 -390 -1910 -260
rect -1200 -272 -100 -260
rect -1200 -388 -486 -272
rect -114 -388 -100 -272
rect -1200 -390 -100 -388
rect -1925 -410 -100 -390
rect 280 -398 318 38
rect 1842 -398 1890 38
rect 280 -430 1890 -398
rect -950 -1298 2490 -1280
rect -950 -1542 -914 -1298
rect 2274 -1542 2490 -1298
rect -950 -1560 2490 -1542
<< via2 >>
rect -898 9753 598 9763
rect -898 9317 598 9753
rect -898 9307 598 9317
rect 1357 7732 2453 8348
rect -1910 -390 -1200 -260
rect -908 -1528 2268 -1312
<< metal3 >>
rect -960 9763 650 9850
rect -960 9307 -898 9763
rect 598 9307 650 9763
rect -960 9220 650 9307
rect -2280 -260 -1180 -240
rect -2280 -390 -1910 -260
rect -1200 -390 -1180 -260
rect -2280 -410 -1180 -390
rect -950 -1280 -265 9220
rect 1300 8352 2520 8450
rect 1300 7728 1353 8352
rect 2457 7728 2520 8352
rect 1300 7620 2520 7728
rect -950 -1312 2490 -1280
rect -950 -1528 -908 -1312
rect 2268 -1528 2490 -1312
rect -950 -1560 2490 -1528
<< via3 >>
rect 1353 8348 2457 8352
rect 1353 7732 1357 8348
rect 1357 7732 2453 8348
rect 2453 7732 2457 8348
rect 1353 7728 2457 7732
<< metal4 >>
rect -2205 12835 26620 13665
rect -2205 8455 -1375 12835
rect -2205 8352 2515 8455
rect -2205 7728 1353 8352
rect 2457 7728 2515 8352
rect -2205 7625 2515 7728
rect 25795 7690 26620 12835
rect 24850 6830 26620 7690
use opamp_diego  opamp_diego_0 ~/CMOS/TopmetalSe/magic
timestamp 1654646295
transform 1 0 -1719 0 1 8388
box 2069 -9997 26971 3199
<< labels >>
rlabel metal1 s 26840 11440 26840 11440 4 VDD
port 1 nsew
rlabel metal4 s 26418 7258 26418 7258 4 AOUT
port 2 nsew
rlabel metal2 s -1078 -314 -1078 -314 4 OUT_IB
port 3 nsew
rlabel metal2 s -1576 3762 -1576 3762 4 ARRAY_OUT
port 5 nsew
rlabel metal1 s 26870 -1360 26870 -1360 4 GND
port 6 nsew
<< end >>
