magic
tech sky130A
magscale 1 2
timestamp 1654749028
<< error_s >>
rect 3033 11271 3041 11293
rect 3293 11271 3395 11280
rect 3765 11271 3867 11292
rect 4473 11271 4575 11277
rect 5291 11271 5393 11292
rect 5527 11271 5629 11277
rect 5999 11271 6101 11280
rect 6471 11271 6573 11289
rect 7289 11271 7391 11292
rect 7525 11271 7627 11277
rect 7997 11271 8099 11280
rect 8469 11271 8571 11289
rect 3061 11249 3069 11271
rect 3057 11204 3069 11249
rect 3321 11243 3367 11252
rect 3793 11243 3839 11264
rect 4501 11243 4547 11249
rect 5319 11243 5365 11264
rect 5555 11243 5601 11249
rect 6027 11243 6073 11252
rect 6499 11243 6545 11261
rect 7317 11243 7363 11264
rect 7553 11243 7599 11249
rect 8025 11243 8071 11252
rect 8497 11243 8543 11261
rect 16879 11223 16913 11257
rect 22112 11231 22139 11269
rect 22140 11259 22167 11269
rect 3085 11176 3089 11221
rect 22128 11203 22139 11231
rect 3889 11075 3979 11091
rect 3889 11063 3911 11075
rect 3917 11063 3951 11075
rect 3917 11055 3939 11063
rect 3957 11055 3979 11075
rect 4125 11075 4215 11091
rect 4125 11063 4147 11075
rect 4153 11063 4187 11075
rect 4153 11055 4175 11063
rect 4193 11055 4215 11075
rect 4361 11075 4451 11091
rect 4361 11063 4383 11075
rect 4389 11063 4423 11075
rect 4389 11055 4411 11063
rect 4429 11055 4451 11075
rect 4597 11075 4687 11091
rect 4597 11063 4619 11075
rect 4625 11063 4659 11075
rect 4625 11055 4647 11063
rect 4665 11055 4687 11075
rect 4833 11075 4923 11091
rect 4833 11063 4855 11075
rect 4861 11063 4895 11075
rect 4861 11055 4883 11063
rect 4901 11055 4923 11075
rect 6123 11075 6213 11091
rect 6123 11063 6145 11075
rect 6151 11063 6185 11075
rect 6151 11055 6173 11063
rect 6191 11055 6213 11075
rect 6595 11075 6685 11091
rect 6595 11063 6617 11075
rect 6623 11063 6657 11075
rect 6623 11055 6645 11063
rect 6663 11055 6685 11075
rect 7177 11075 7267 11091
rect 7177 11063 7199 11075
rect 7205 11063 7239 11075
rect 7205 11055 7227 11063
rect 7245 11055 7267 11075
rect 7649 11075 7739 11091
rect 7649 11063 7671 11075
rect 7677 11063 7711 11075
rect 7677 11055 7699 11063
rect 7717 11055 7739 11075
rect 8121 11075 8211 11091
rect 8121 11063 8143 11075
rect 8149 11063 8183 11075
rect 8149 11055 8171 11063
rect 8189 11055 8211 11075
rect 8593 11075 8683 11091
rect 8593 11063 8615 11075
rect 8621 11063 8655 11075
rect 8621 11055 8643 11063
rect 8661 11055 8683 11075
rect 11253 11062 11269 11078
rect 11271 11062 11287 11078
rect 11371 11062 11387 11078
rect 11389 11062 11405 11078
rect 11489 11062 11505 11078
rect 11507 11062 11523 11078
rect 11607 11062 11623 11078
rect 11625 11062 11641 11078
rect 11725 11062 11741 11078
rect 11743 11062 11759 11078
rect 11843 11062 11859 11078
rect 11861 11062 11877 11078
rect 11961 11062 11977 11078
rect 11979 11062 11995 11078
rect 12079 11062 12095 11078
rect 12097 11062 12113 11078
rect 12197 11062 12213 11078
rect 12215 11062 12231 11078
rect 12315 11062 12331 11078
rect 12333 11062 12349 11078
rect 12433 11062 12449 11078
rect 12451 11062 12467 11078
rect 12551 11062 12567 11078
rect 12569 11062 12585 11078
rect 12669 11062 12685 11078
rect 12687 11062 12703 11078
rect 12787 11062 12803 11078
rect 12805 11062 12821 11078
rect 12905 11062 12921 11078
rect 12923 11062 12939 11078
rect 13023 11062 13039 11078
rect 13041 11062 13057 11078
rect 13141 11062 13157 11078
rect 13159 11062 13175 11078
rect 13259 11062 13275 11078
rect 13277 11062 13293 11078
rect 13377 11062 13393 11078
rect 13395 11062 13411 11078
rect 13495 11062 13511 11078
rect 13513 11062 13529 11078
rect 13613 11062 13629 11078
rect 13631 11062 13647 11078
rect 13731 11062 13747 11078
rect 13749 11062 13765 11078
rect 15376 11062 15392 11078
rect 15394 11062 15410 11078
rect 15494 11062 15510 11078
rect 15512 11062 15528 11078
rect 15612 11062 15628 11078
rect 15630 11062 15646 11078
rect 15730 11062 15746 11078
rect 15748 11062 15764 11078
rect 15848 11062 15864 11078
rect 15866 11062 15882 11078
rect 15966 11062 15982 11078
rect 15984 11062 16000 11078
rect 16084 11062 16100 11078
rect 16102 11062 16118 11078
rect 16202 11062 16218 11078
rect 16220 11062 16236 11078
rect 16320 11062 16336 11078
rect 16338 11062 16354 11078
rect 16438 11062 16454 11078
rect 16456 11062 16472 11078
rect 16556 11062 16572 11078
rect 16574 11062 16590 11078
rect 16674 11062 16690 11078
rect 16692 11062 16708 11078
rect 16792 11062 16808 11078
rect 16810 11062 16826 11078
rect 16910 11062 16926 11078
rect 16928 11062 16944 11078
rect 17028 11062 17044 11078
rect 17046 11062 17062 11078
rect 17146 11062 17162 11078
rect 17164 11062 17180 11078
rect 17264 11062 17280 11078
rect 17282 11062 17298 11078
rect 17382 11062 17398 11078
rect 17400 11062 17416 11078
rect 17500 11062 17516 11078
rect 17518 11062 17534 11078
rect 17618 11062 17634 11078
rect 17636 11062 17652 11078
rect 17736 11062 17752 11078
rect 17754 11062 17770 11078
rect 17854 11062 17870 11078
rect 17872 11062 17888 11078
rect 19499 11062 19515 11078
rect 19517 11062 19533 11078
rect 19617 11062 19633 11078
rect 19635 11062 19651 11078
rect 19735 11062 19751 11078
rect 19753 11062 19769 11078
rect 19853 11062 19869 11078
rect 19871 11062 19887 11078
rect 19971 11062 19987 11078
rect 19989 11062 20005 11078
rect 20089 11062 20105 11078
rect 20107 11062 20123 11078
rect 20207 11062 20223 11078
rect 20225 11062 20241 11078
rect 20325 11062 20341 11078
rect 20343 11062 20359 11078
rect 20443 11062 20459 11078
rect 20461 11062 20477 11078
rect 20561 11062 20577 11078
rect 20579 11062 20595 11078
rect 20679 11062 20695 11078
rect 20697 11062 20713 11078
rect 20797 11062 20813 11078
rect 20815 11062 20831 11078
rect 20915 11062 20931 11078
rect 20933 11062 20949 11078
rect 21033 11062 21049 11078
rect 21051 11062 21067 11078
rect 21151 11062 21167 11078
rect 21169 11062 21185 11078
rect 21269 11062 21285 11078
rect 21287 11062 21303 11078
rect 21387 11062 21403 11078
rect 21405 11062 21421 11078
rect 21505 11062 21521 11078
rect 21523 11062 21539 11078
rect 21623 11062 21639 11078
rect 21641 11062 21657 11078
rect 21741 11062 21757 11078
rect 21759 11062 21775 11078
rect 21859 11062 21875 11078
rect 21877 11062 21893 11078
rect 21977 11062 21993 11078
rect 21995 11062 22011 11078
rect 3917 11035 3951 11055
rect 4153 11035 4187 11055
rect 4389 11035 4423 11055
rect 4625 11035 4659 11055
rect 4861 11035 4895 11055
rect 6151 11035 6185 11055
rect 6623 11035 6657 11055
rect 7205 11035 7239 11055
rect 7677 11035 7711 11055
rect 8149 11035 8183 11055
rect 8621 11035 8655 11055
rect 11237 11054 11303 11062
rect 11237 11046 11261 11054
rect 3889 10495 3898 10523
rect 3917 10475 3951 10515
rect 3970 10495 3979 10523
rect 4125 10495 4134 10523
rect 3957 10487 3979 10495
rect 4153 10475 4187 10515
rect 4206 10495 4215 10523
rect 4361 10495 4370 10523
rect 4193 10487 4215 10495
rect 4389 10475 4423 10515
rect 4442 10495 4451 10523
rect 4597 10495 4606 10523
rect 4429 10487 4451 10495
rect 4625 10475 4659 10515
rect 4678 10495 4687 10523
rect 4833 10495 4842 10523
rect 4665 10487 4687 10495
rect 4861 10475 4895 10515
rect 4914 10495 4923 10523
rect 6123 10495 6132 10523
rect 4901 10487 4923 10495
rect 6151 10475 6185 10515
rect 6204 10495 6213 10523
rect 6595 10495 6604 10523
rect 6191 10487 6213 10495
rect 6623 10475 6657 10515
rect 6676 10495 6685 10523
rect 7177 10495 7186 10523
rect 6663 10487 6685 10495
rect 7205 10475 7239 10515
rect 7258 10495 7267 10523
rect 7649 10495 7658 10523
rect 7245 10487 7267 10495
rect 7677 10475 7711 10515
rect 7730 10495 7739 10523
rect 8121 10495 8130 10523
rect 7717 10487 7739 10495
rect 8149 10475 8183 10515
rect 8202 10495 8211 10523
rect 8593 10495 8602 10523
rect 8189 10487 8211 10495
rect 8621 10475 8655 10515
rect 8674 10495 8683 10523
rect 11253 10502 11261 11046
rect 8661 10487 8683 10495
rect 11237 10494 11261 10502
rect 11279 11046 11303 11054
rect 11355 11054 11421 11062
rect 11355 11046 11379 11054
rect 11279 10502 11287 11046
rect 11371 10502 11379 11046
rect 11279 10494 11303 10502
rect 11237 10486 11303 10494
rect 11355 10494 11379 10502
rect 11397 11046 11421 11054
rect 11473 11054 11539 11062
rect 11473 11046 11497 11054
rect 11397 10502 11405 11046
rect 11489 10502 11497 11046
rect 11397 10494 11421 10502
rect 11355 10486 11421 10494
rect 11473 10494 11497 10502
rect 11515 11046 11539 11054
rect 11591 11054 11657 11062
rect 11591 11046 11615 11054
rect 11515 10502 11523 11046
rect 11607 10502 11615 11046
rect 11515 10494 11539 10502
rect 11473 10486 11539 10494
rect 11591 10494 11615 10502
rect 11633 11046 11657 11054
rect 11709 11054 11775 11062
rect 11709 11046 11733 11054
rect 11633 10502 11641 11046
rect 11725 10502 11733 11046
rect 11633 10494 11657 10502
rect 11591 10486 11657 10494
rect 11709 10494 11733 10502
rect 11751 11046 11775 11054
rect 11827 11054 11893 11062
rect 11827 11046 11851 11054
rect 11751 10502 11759 11046
rect 11843 10502 11851 11046
rect 11751 10494 11775 10502
rect 11709 10486 11775 10494
rect 11827 10494 11851 10502
rect 11869 11046 11893 11054
rect 11945 11054 12011 11062
rect 11945 11046 11969 11054
rect 11869 10502 11877 11046
rect 11961 10502 11969 11046
rect 11869 10494 11893 10502
rect 11827 10486 11893 10494
rect 11945 10494 11969 10502
rect 11987 11046 12011 11054
rect 12063 11054 12129 11062
rect 12063 11046 12087 11054
rect 11987 10502 11995 11046
rect 12079 10502 12087 11046
rect 11987 10494 12011 10502
rect 11945 10486 12011 10494
rect 12063 10494 12087 10502
rect 12105 11046 12129 11054
rect 12181 11054 12247 11062
rect 12181 11046 12205 11054
rect 12105 10502 12113 11046
rect 12197 10502 12205 11046
rect 12105 10494 12129 10502
rect 12063 10486 12129 10494
rect 12181 10494 12205 10502
rect 12223 11046 12247 11054
rect 12299 11054 12365 11062
rect 12299 11046 12323 11054
rect 12223 10502 12231 11046
rect 12315 10502 12323 11046
rect 12223 10494 12247 10502
rect 12181 10486 12247 10494
rect 12299 10494 12323 10502
rect 12341 11046 12365 11054
rect 12417 11054 12483 11062
rect 12417 11046 12441 11054
rect 12341 10502 12349 11046
rect 12433 10502 12441 11046
rect 12341 10494 12365 10502
rect 12299 10486 12365 10494
rect 12417 10494 12441 10502
rect 12459 11046 12483 11054
rect 12535 11054 12601 11062
rect 12535 11046 12559 11054
rect 12459 10502 12467 11046
rect 12551 10502 12559 11046
rect 12459 10494 12483 10502
rect 12417 10486 12483 10494
rect 12535 10494 12559 10502
rect 12577 11046 12601 11054
rect 12653 11054 12719 11062
rect 12653 11046 12677 11054
rect 12577 10502 12585 11046
rect 12669 10502 12677 11046
rect 12577 10494 12601 10502
rect 12535 10486 12601 10494
rect 12653 10494 12677 10502
rect 12695 11046 12719 11054
rect 12771 11054 12837 11062
rect 12771 11046 12795 11054
rect 12695 10502 12703 11046
rect 12787 10502 12795 11046
rect 12695 10494 12719 10502
rect 12653 10486 12719 10494
rect 12771 10494 12795 10502
rect 12813 11046 12837 11054
rect 12889 11054 12955 11062
rect 12889 11046 12913 11054
rect 12813 10502 12821 11046
rect 12905 10502 12913 11046
rect 12813 10494 12837 10502
rect 12771 10486 12837 10494
rect 12889 10494 12913 10502
rect 12931 11046 12955 11054
rect 13007 11054 13073 11062
rect 13007 11046 13031 11054
rect 12931 10502 12939 11046
rect 13023 10502 13031 11046
rect 12931 10494 12955 10502
rect 12889 10486 12955 10494
rect 13007 10494 13031 10502
rect 13049 11046 13073 11054
rect 13125 11054 13191 11062
rect 13125 11046 13149 11054
rect 13049 10502 13057 11046
rect 13141 10502 13149 11046
rect 13049 10494 13073 10502
rect 13007 10486 13073 10494
rect 13125 10494 13149 10502
rect 13167 11046 13191 11054
rect 13243 11054 13309 11062
rect 13243 11046 13267 11054
rect 13167 10502 13175 11046
rect 13259 10502 13267 11046
rect 13167 10494 13191 10502
rect 13125 10486 13191 10494
rect 13243 10494 13267 10502
rect 13285 11046 13309 11054
rect 13361 11054 13427 11062
rect 13361 11046 13385 11054
rect 13285 10502 13293 11046
rect 13377 10502 13385 11046
rect 13285 10494 13309 10502
rect 13243 10486 13309 10494
rect 13361 10494 13385 10502
rect 13403 11046 13427 11054
rect 13479 11054 13545 11062
rect 13479 11046 13503 11054
rect 13403 10502 13411 11046
rect 13495 10502 13503 11046
rect 13403 10494 13427 10502
rect 13361 10486 13427 10494
rect 13479 10494 13503 10502
rect 13521 11046 13545 11054
rect 13597 11054 13663 11062
rect 13597 11046 13621 11054
rect 13521 10502 13529 11046
rect 13613 10502 13621 11046
rect 13521 10494 13545 10502
rect 13479 10486 13545 10494
rect 13597 10494 13621 10502
rect 13639 11046 13663 11054
rect 13715 11054 13781 11062
rect 13715 11046 13739 11054
rect 13639 10502 13647 11046
rect 13731 10502 13739 11046
rect 13639 10494 13663 10502
rect 13597 10486 13663 10494
rect 13715 10494 13739 10502
rect 13757 11046 13781 11054
rect 15360 11054 15426 11062
rect 15360 11046 15384 11054
rect 13757 10502 13765 11046
rect 15376 10502 15384 11046
rect 13757 10494 13781 10502
rect 13715 10486 13781 10494
rect 15360 10494 15384 10502
rect 15402 11046 15426 11054
rect 15478 11054 15544 11062
rect 15478 11046 15502 11054
rect 15402 10502 15410 11046
rect 15494 10502 15502 11046
rect 15402 10494 15426 10502
rect 15360 10486 15426 10494
rect 15478 10494 15502 10502
rect 15520 11046 15544 11054
rect 15596 11054 15662 11062
rect 15596 11046 15620 11054
rect 15520 10502 15528 11046
rect 15612 10502 15620 11046
rect 15520 10494 15544 10502
rect 15478 10486 15544 10494
rect 15596 10494 15620 10502
rect 15638 11046 15662 11054
rect 15714 11054 15780 11062
rect 15714 11046 15738 11054
rect 15638 10502 15646 11046
rect 15730 10502 15738 11046
rect 15638 10494 15662 10502
rect 15596 10486 15662 10494
rect 15714 10494 15738 10502
rect 15756 11046 15780 11054
rect 15832 11054 15898 11062
rect 15832 11046 15856 11054
rect 15756 10502 15764 11046
rect 15848 10502 15856 11046
rect 15756 10494 15780 10502
rect 15714 10486 15780 10494
rect 15832 10494 15856 10502
rect 15874 11046 15898 11054
rect 15950 11054 16016 11062
rect 15950 11046 15974 11054
rect 15874 10502 15882 11046
rect 15966 10502 15974 11046
rect 15874 10494 15898 10502
rect 15832 10486 15898 10494
rect 15950 10494 15974 10502
rect 15992 11046 16016 11054
rect 16068 11054 16134 11062
rect 16068 11046 16092 11054
rect 15992 10502 16000 11046
rect 16084 10502 16092 11046
rect 15992 10494 16016 10502
rect 15950 10486 16016 10494
rect 16068 10494 16092 10502
rect 16110 11046 16134 11054
rect 16186 11054 16252 11062
rect 16186 11046 16210 11054
rect 16110 10502 16118 11046
rect 16202 10502 16210 11046
rect 16110 10494 16134 10502
rect 16068 10486 16134 10494
rect 16186 10494 16210 10502
rect 16228 11046 16252 11054
rect 16304 11054 16370 11062
rect 16304 11046 16328 11054
rect 16228 10502 16236 11046
rect 16320 10502 16328 11046
rect 16228 10494 16252 10502
rect 16186 10486 16252 10494
rect 16304 10494 16328 10502
rect 16346 11046 16370 11054
rect 16422 11054 16488 11062
rect 16422 11046 16446 11054
rect 16346 10502 16354 11046
rect 16438 10502 16446 11046
rect 16346 10494 16370 10502
rect 16304 10486 16370 10494
rect 16422 10494 16446 10502
rect 16464 11046 16488 11054
rect 16540 11054 16606 11062
rect 16540 11046 16564 11054
rect 16464 10502 16472 11046
rect 16556 10502 16564 11046
rect 16464 10494 16488 10502
rect 16422 10486 16488 10494
rect 16540 10494 16564 10502
rect 16582 11046 16606 11054
rect 16658 11054 16724 11062
rect 16658 11046 16682 11054
rect 16582 10502 16590 11046
rect 16674 10502 16682 11046
rect 16582 10494 16606 10502
rect 16540 10486 16606 10494
rect 16658 10494 16682 10502
rect 16700 11046 16724 11054
rect 16776 11054 16842 11062
rect 16776 11046 16800 11054
rect 16700 10502 16708 11046
rect 16792 10502 16800 11046
rect 16700 10494 16724 10502
rect 16658 10486 16724 10494
rect 16776 10494 16800 10502
rect 16818 11046 16842 11054
rect 16894 11054 16960 11062
rect 16894 11046 16918 11054
rect 16818 10502 16826 11046
rect 16910 10502 16918 11046
rect 16818 10494 16842 10502
rect 16776 10486 16842 10494
rect 16894 10494 16918 10502
rect 16936 11046 16960 11054
rect 17012 11054 17078 11062
rect 17012 11046 17036 11054
rect 16936 10502 16944 11046
rect 17028 10502 17036 11046
rect 16936 10494 16960 10502
rect 16894 10486 16960 10494
rect 17012 10494 17036 10502
rect 17054 11046 17078 11054
rect 17130 11054 17196 11062
rect 17130 11046 17154 11054
rect 17054 10502 17062 11046
rect 17146 10502 17154 11046
rect 17054 10494 17078 10502
rect 17012 10486 17078 10494
rect 17130 10494 17154 10502
rect 17172 11046 17196 11054
rect 17248 11054 17314 11062
rect 17248 11046 17272 11054
rect 17172 10502 17180 11046
rect 17264 10502 17272 11046
rect 17172 10494 17196 10502
rect 17130 10486 17196 10494
rect 17248 10494 17272 10502
rect 17290 11046 17314 11054
rect 17366 11054 17432 11062
rect 17366 11046 17390 11054
rect 17290 10502 17298 11046
rect 17382 10502 17390 11046
rect 17290 10494 17314 10502
rect 17248 10486 17314 10494
rect 17366 10494 17390 10502
rect 17408 11046 17432 11054
rect 17484 11054 17550 11062
rect 17484 11046 17508 11054
rect 17408 10502 17416 11046
rect 17500 10502 17508 11046
rect 17408 10494 17432 10502
rect 17366 10486 17432 10494
rect 17484 10494 17508 10502
rect 17526 11046 17550 11054
rect 17602 11054 17668 11062
rect 17602 11046 17626 11054
rect 17526 10502 17534 11046
rect 17618 10502 17626 11046
rect 17526 10494 17550 10502
rect 17484 10486 17550 10494
rect 17602 10494 17626 10502
rect 17644 11046 17668 11054
rect 17720 11054 17786 11062
rect 17720 11046 17744 11054
rect 17644 10502 17652 11046
rect 17736 10502 17744 11046
rect 17644 10494 17668 10502
rect 17602 10486 17668 10494
rect 17720 10494 17744 10502
rect 17762 11046 17786 11054
rect 17838 11054 17904 11062
rect 17838 11046 17862 11054
rect 17762 10502 17770 11046
rect 17854 10502 17862 11046
rect 17762 10494 17786 10502
rect 17720 10486 17786 10494
rect 17838 10494 17862 10502
rect 17880 11046 17904 11054
rect 19483 11054 19549 11062
rect 19483 11046 19507 11054
rect 17880 10502 17888 11046
rect 19499 10502 19507 11046
rect 17880 10494 17904 10502
rect 17838 10486 17904 10494
rect 19483 10494 19507 10502
rect 19525 11046 19549 11054
rect 19601 11054 19667 11062
rect 19601 11046 19625 11054
rect 19525 10502 19533 11046
rect 19617 10502 19625 11046
rect 19525 10494 19549 10502
rect 19483 10486 19549 10494
rect 19601 10494 19625 10502
rect 19643 11046 19667 11054
rect 19719 11054 19785 11062
rect 19719 11046 19743 11054
rect 19643 10502 19651 11046
rect 19735 10502 19743 11046
rect 19643 10494 19667 10502
rect 19601 10486 19667 10494
rect 19719 10494 19743 10502
rect 19761 11046 19785 11054
rect 19837 11054 19903 11062
rect 19837 11046 19861 11054
rect 19761 10502 19769 11046
rect 19853 10502 19861 11046
rect 19761 10494 19785 10502
rect 19719 10486 19785 10494
rect 19837 10494 19861 10502
rect 19879 11046 19903 11054
rect 19955 11054 20021 11062
rect 19955 11046 19979 11054
rect 19879 10502 19887 11046
rect 19971 10502 19979 11046
rect 19879 10494 19903 10502
rect 19837 10486 19903 10494
rect 19955 10494 19979 10502
rect 19997 11046 20021 11054
rect 20073 11054 20139 11062
rect 20073 11046 20097 11054
rect 19997 10502 20005 11046
rect 20089 10502 20097 11046
rect 19997 10494 20021 10502
rect 19955 10486 20021 10494
rect 20073 10494 20097 10502
rect 20115 11046 20139 11054
rect 20191 11054 20257 11062
rect 20191 11046 20215 11054
rect 20115 10502 20123 11046
rect 20207 10502 20215 11046
rect 20115 10494 20139 10502
rect 20073 10486 20139 10494
rect 20191 10494 20215 10502
rect 20233 11046 20257 11054
rect 20309 11054 20375 11062
rect 20309 11046 20333 11054
rect 20233 10502 20241 11046
rect 20325 10502 20333 11046
rect 20233 10494 20257 10502
rect 20191 10486 20257 10494
rect 20309 10494 20333 10502
rect 20351 11046 20375 11054
rect 20427 11054 20493 11062
rect 20427 11046 20451 11054
rect 20351 10502 20359 11046
rect 20443 10502 20451 11046
rect 20351 10494 20375 10502
rect 20309 10486 20375 10494
rect 20427 10494 20451 10502
rect 20469 11046 20493 11054
rect 20545 11054 20611 11062
rect 20545 11046 20569 11054
rect 20469 10502 20477 11046
rect 20561 10502 20569 11046
rect 20469 10494 20493 10502
rect 20427 10486 20493 10494
rect 20545 10494 20569 10502
rect 20587 11046 20611 11054
rect 20663 11054 20729 11062
rect 20663 11046 20687 11054
rect 20587 10502 20595 11046
rect 20679 10502 20687 11046
rect 20587 10494 20611 10502
rect 20545 10486 20611 10494
rect 20663 10494 20687 10502
rect 20705 11046 20729 11054
rect 20781 11054 20847 11062
rect 20781 11046 20805 11054
rect 20705 10502 20713 11046
rect 20797 10502 20805 11046
rect 20705 10494 20729 10502
rect 20663 10486 20729 10494
rect 20781 10494 20805 10502
rect 20823 11046 20847 11054
rect 20899 11054 20965 11062
rect 20899 11046 20923 11054
rect 20823 10502 20831 11046
rect 20915 10502 20923 11046
rect 20823 10494 20847 10502
rect 20781 10486 20847 10494
rect 20899 10494 20923 10502
rect 20941 11046 20965 11054
rect 21017 11054 21083 11062
rect 21017 11046 21041 11054
rect 20941 10502 20949 11046
rect 21033 10502 21041 11046
rect 20941 10494 20965 10502
rect 20899 10486 20965 10494
rect 21017 10494 21041 10502
rect 21059 11046 21083 11054
rect 21135 11054 21201 11062
rect 21135 11046 21159 11054
rect 21059 10502 21067 11046
rect 21151 10502 21159 11046
rect 21059 10494 21083 10502
rect 21017 10486 21083 10494
rect 21135 10494 21159 10502
rect 21177 11046 21201 11054
rect 21253 11054 21319 11062
rect 21253 11046 21277 11054
rect 21177 10502 21185 11046
rect 21269 10502 21277 11046
rect 21177 10494 21201 10502
rect 21135 10486 21201 10494
rect 21253 10494 21277 10502
rect 21295 11046 21319 11054
rect 21371 11054 21437 11062
rect 21371 11046 21395 11054
rect 21295 10502 21303 11046
rect 21387 10502 21395 11046
rect 21295 10494 21319 10502
rect 21253 10486 21319 10494
rect 21371 10494 21395 10502
rect 21413 11046 21437 11054
rect 21489 11054 21555 11062
rect 21489 11046 21513 11054
rect 21413 10502 21421 11046
rect 21505 10502 21513 11046
rect 21413 10494 21437 10502
rect 21371 10486 21437 10494
rect 21489 10494 21513 10502
rect 21531 11046 21555 11054
rect 21607 11054 21673 11062
rect 21607 11046 21631 11054
rect 21531 10502 21539 11046
rect 21623 10502 21631 11046
rect 21531 10494 21555 10502
rect 21489 10486 21555 10494
rect 21607 10494 21631 10502
rect 21649 11046 21673 11054
rect 21725 11054 21791 11062
rect 21725 11046 21749 11054
rect 21649 10502 21657 11046
rect 21741 10502 21749 11046
rect 21649 10494 21673 10502
rect 21607 10486 21673 10494
rect 21725 10494 21749 10502
rect 21767 11046 21791 11054
rect 21843 11054 21909 11062
rect 21843 11046 21867 11054
rect 21767 10502 21775 11046
rect 21859 10502 21867 11046
rect 21767 10494 21791 10502
rect 21725 10486 21791 10494
rect 21843 10494 21867 10502
rect 21885 11046 21909 11054
rect 21961 11054 22027 11062
rect 21961 11046 21985 11054
rect 21885 10502 21893 11046
rect 21977 10502 21985 11046
rect 21885 10494 21909 10502
rect 21843 10486 21909 10494
rect 21961 10494 21985 10502
rect 22003 11046 22027 11054
rect 22003 10502 22011 11046
rect 22003 10494 22027 10502
rect 21961 10486 22027 10494
rect 11253 10470 11269 10486
rect 11271 10470 11287 10486
rect 11371 10470 11387 10486
rect 11389 10470 11405 10486
rect 11489 10470 11505 10486
rect 11507 10470 11523 10486
rect 11607 10470 11623 10486
rect 11625 10470 11641 10486
rect 11725 10470 11741 10486
rect 11743 10470 11759 10486
rect 11843 10470 11859 10486
rect 11861 10470 11877 10486
rect 11961 10470 11977 10486
rect 11979 10470 11995 10486
rect 12079 10470 12095 10486
rect 12097 10470 12113 10486
rect 12197 10470 12213 10486
rect 12215 10470 12231 10486
rect 12315 10470 12331 10486
rect 12333 10470 12349 10486
rect 12433 10470 12449 10486
rect 12451 10470 12467 10486
rect 12551 10470 12567 10486
rect 12569 10470 12585 10486
rect 12669 10470 12685 10486
rect 12687 10470 12703 10486
rect 12787 10470 12803 10486
rect 12805 10470 12821 10486
rect 12905 10470 12921 10486
rect 12923 10470 12939 10486
rect 13023 10470 13039 10486
rect 13041 10470 13057 10486
rect 13141 10470 13157 10486
rect 13159 10470 13175 10486
rect 13259 10470 13275 10486
rect 13277 10470 13293 10486
rect 13377 10470 13393 10486
rect 13395 10470 13411 10486
rect 13495 10470 13511 10486
rect 13513 10470 13529 10486
rect 13613 10470 13629 10486
rect 13631 10470 13647 10486
rect 13731 10470 13747 10486
rect 13749 10470 13765 10486
rect 15376 10470 15392 10486
rect 15394 10470 15410 10486
rect 15494 10470 15510 10486
rect 15512 10470 15528 10486
rect 15612 10470 15628 10486
rect 15630 10470 15646 10486
rect 15730 10470 15746 10486
rect 15748 10470 15764 10486
rect 15848 10470 15864 10486
rect 15866 10470 15882 10486
rect 15966 10470 15982 10486
rect 15984 10470 16000 10486
rect 16084 10470 16100 10486
rect 16102 10470 16118 10486
rect 16202 10470 16218 10486
rect 16220 10470 16236 10486
rect 16320 10470 16336 10486
rect 16338 10470 16354 10486
rect 16438 10470 16454 10486
rect 16456 10470 16472 10486
rect 16556 10470 16572 10486
rect 16574 10470 16590 10486
rect 16674 10470 16690 10486
rect 16692 10470 16708 10486
rect 16792 10470 16808 10486
rect 16810 10470 16826 10486
rect 16910 10470 16926 10486
rect 16928 10470 16944 10486
rect 17028 10470 17044 10486
rect 17046 10470 17062 10486
rect 17146 10470 17162 10486
rect 17164 10470 17180 10486
rect 17264 10470 17280 10486
rect 17282 10470 17298 10486
rect 17382 10470 17398 10486
rect 17400 10470 17416 10486
rect 17500 10470 17516 10486
rect 17518 10470 17534 10486
rect 17618 10470 17634 10486
rect 17636 10470 17652 10486
rect 17736 10470 17752 10486
rect 17754 10470 17770 10486
rect 17854 10470 17870 10486
rect 17872 10470 17888 10486
rect 19499 10470 19515 10486
rect 19517 10470 19533 10486
rect 19617 10470 19633 10486
rect 19635 10470 19651 10486
rect 19735 10470 19751 10486
rect 19753 10470 19769 10486
rect 19853 10470 19869 10486
rect 19871 10470 19887 10486
rect 19971 10470 19987 10486
rect 19989 10470 20005 10486
rect 20089 10470 20105 10486
rect 20107 10470 20123 10486
rect 20207 10470 20223 10486
rect 20225 10470 20241 10486
rect 20325 10470 20341 10486
rect 20343 10470 20359 10486
rect 20443 10470 20459 10486
rect 20461 10470 20477 10486
rect 20561 10470 20577 10486
rect 20579 10470 20595 10486
rect 20679 10470 20695 10486
rect 20697 10470 20713 10486
rect 20797 10470 20813 10486
rect 20815 10470 20831 10486
rect 20915 10470 20931 10486
rect 20933 10470 20949 10486
rect 21033 10470 21049 10486
rect 21051 10470 21067 10486
rect 21151 10470 21167 10486
rect 21169 10470 21185 10486
rect 21269 10470 21285 10486
rect 21287 10470 21303 10486
rect 21387 10470 21403 10486
rect 21405 10470 21421 10486
rect 21505 10470 21521 10486
rect 21523 10470 21539 10486
rect 21623 10470 21639 10486
rect 21641 10470 21657 10486
rect 21741 10470 21757 10486
rect 21759 10470 21775 10486
rect 21859 10470 21875 10486
rect 21877 10470 21893 10486
rect 21977 10470 21993 10486
rect 21995 10470 22011 10486
rect 3150 10394 3184 10428
rect 3268 10394 3302 10428
rect 3386 10394 3420 10428
rect 3504 10394 3538 10428
rect 3622 10394 3656 10428
rect 3740 10394 3774 10428
rect 3858 10394 3892 10428
rect 3976 10394 4010 10428
rect 4094 10394 4128 10428
rect 4212 10394 4246 10428
rect 4330 10394 4364 10428
rect 4448 10394 4482 10428
rect 4566 10394 4600 10428
rect 4684 10394 4718 10428
rect 4802 10394 4836 10428
rect 5384 10394 5418 10428
rect 5502 10394 5536 10428
rect 5620 10394 5654 10428
rect 5738 10394 5772 10428
rect 5856 10394 5890 10428
rect 5974 10394 6008 10428
rect 10958 10427 10974 10443
rect 10976 10427 10992 10443
rect 15081 10427 15097 10443
rect 15099 10427 15115 10443
rect 19204 10427 19220 10443
rect 19222 10427 19238 10443
rect 10942 10423 10992 10427
rect 10942 10411 10958 10423
rect 11004 10411 11008 10427
rect 15065 10423 15115 10427
rect 15065 10411 15081 10423
rect 15127 10411 15131 10427
rect 19188 10423 19238 10427
rect 19188 10411 19204 10423
rect 19250 10411 19254 10427
rect 10946 10409 10958 10411
rect 15069 10409 15081 10411
rect 19192 10409 19204 10411
rect 10942 10393 10958 10409
rect 11004 10393 11008 10409
rect 15065 10393 15081 10409
rect 15127 10393 15131 10409
rect 19188 10393 19204 10409
rect 19250 10393 19254 10409
rect 10958 10377 10974 10393
rect 10976 10377 10992 10393
rect 15081 10377 15097 10393
rect 15099 10377 15115 10393
rect 19204 10377 19220 10393
rect 19222 10377 19238 10393
rect 10958 10319 10974 10335
rect 10976 10319 10992 10335
rect 15081 10319 15097 10335
rect 15099 10319 15115 10335
rect 19204 10319 19220 10335
rect 19222 10319 19238 10335
rect 10942 10303 10958 10319
rect 11004 10303 11008 10319
rect 15065 10303 15081 10319
rect 15127 10303 15131 10319
rect 19188 10303 19204 10319
rect 19250 10303 19254 10319
rect 10946 10301 10958 10303
rect 15069 10301 15081 10303
rect 19192 10301 19204 10303
rect 10942 10289 10958 10301
rect 10942 10285 10992 10289
rect 11004 10285 11008 10301
rect 15065 10289 15081 10301
rect 15065 10285 15115 10289
rect 15127 10285 15131 10301
rect 19188 10289 19204 10301
rect 19188 10285 19238 10289
rect 19250 10285 19254 10301
rect 10958 10269 10974 10285
rect 10976 10269 10992 10285
rect 15081 10269 15097 10285
rect 15099 10269 15115 10285
rect 19204 10269 19220 10285
rect 19222 10269 19238 10285
rect 11253 10226 11269 10242
rect 11271 10226 11287 10242
rect 11371 10226 11387 10242
rect 11389 10226 11405 10242
rect 11489 10226 11505 10242
rect 11507 10226 11523 10242
rect 11607 10226 11623 10242
rect 11625 10226 11641 10242
rect 11725 10226 11741 10242
rect 11743 10226 11759 10242
rect 11843 10226 11859 10242
rect 11861 10226 11877 10242
rect 11961 10226 11977 10242
rect 11979 10226 11995 10242
rect 12079 10226 12095 10242
rect 12097 10226 12113 10242
rect 12197 10226 12213 10242
rect 12215 10226 12231 10242
rect 12315 10226 12331 10242
rect 12333 10226 12349 10242
rect 12433 10226 12449 10242
rect 12451 10226 12467 10242
rect 12551 10226 12567 10242
rect 12569 10226 12585 10242
rect 12669 10226 12685 10242
rect 12687 10226 12703 10242
rect 12787 10226 12803 10242
rect 12805 10226 12821 10242
rect 12905 10226 12921 10242
rect 12923 10226 12939 10242
rect 13023 10226 13039 10242
rect 13041 10226 13057 10242
rect 13141 10226 13157 10242
rect 13159 10226 13175 10242
rect 13259 10226 13275 10242
rect 13277 10226 13293 10242
rect 13377 10226 13393 10242
rect 13395 10226 13411 10242
rect 13495 10226 13511 10242
rect 13513 10226 13529 10242
rect 13613 10226 13629 10242
rect 13631 10226 13647 10242
rect 13731 10226 13747 10242
rect 13749 10226 13765 10242
rect 15376 10226 15392 10242
rect 15394 10226 15410 10242
rect 15494 10226 15510 10242
rect 15512 10226 15528 10242
rect 15612 10226 15628 10242
rect 15630 10226 15646 10242
rect 15730 10226 15746 10242
rect 15748 10226 15764 10242
rect 15848 10226 15864 10242
rect 15866 10226 15882 10242
rect 15966 10226 15982 10242
rect 15984 10226 16000 10242
rect 16084 10226 16100 10242
rect 16102 10226 16118 10242
rect 16202 10226 16218 10242
rect 16220 10226 16236 10242
rect 16320 10226 16336 10242
rect 16338 10226 16354 10242
rect 16438 10226 16454 10242
rect 16456 10226 16472 10242
rect 16556 10226 16572 10242
rect 16574 10226 16590 10242
rect 16674 10226 16690 10242
rect 16692 10226 16708 10242
rect 16792 10226 16808 10242
rect 16810 10226 16826 10242
rect 16910 10226 16926 10242
rect 16928 10226 16944 10242
rect 17028 10226 17044 10242
rect 17046 10226 17062 10242
rect 17146 10226 17162 10242
rect 17164 10226 17180 10242
rect 17264 10226 17280 10242
rect 17282 10226 17298 10242
rect 17382 10226 17398 10242
rect 17400 10226 17416 10242
rect 17500 10226 17516 10242
rect 17518 10226 17534 10242
rect 17618 10226 17634 10242
rect 17636 10226 17652 10242
rect 17736 10226 17752 10242
rect 17754 10226 17770 10242
rect 17854 10226 17870 10242
rect 17872 10226 17888 10242
rect 19499 10226 19515 10242
rect 19517 10226 19533 10242
rect 19617 10226 19633 10242
rect 19635 10226 19651 10242
rect 19735 10226 19751 10242
rect 19753 10226 19769 10242
rect 19853 10226 19869 10242
rect 19871 10226 19887 10242
rect 19971 10226 19987 10242
rect 19989 10226 20005 10242
rect 20089 10226 20105 10242
rect 20107 10226 20123 10242
rect 20207 10226 20223 10242
rect 20225 10226 20241 10242
rect 20325 10226 20341 10242
rect 20343 10226 20359 10242
rect 20443 10226 20459 10242
rect 20461 10226 20477 10242
rect 20561 10226 20577 10242
rect 20579 10226 20595 10242
rect 20679 10226 20695 10242
rect 20697 10226 20713 10242
rect 20797 10226 20813 10242
rect 20815 10226 20831 10242
rect 20915 10226 20931 10242
rect 20933 10226 20949 10242
rect 21033 10226 21049 10242
rect 21051 10226 21067 10242
rect 21151 10226 21167 10242
rect 21169 10226 21185 10242
rect 21269 10226 21285 10242
rect 21287 10226 21303 10242
rect 21387 10226 21403 10242
rect 21405 10226 21421 10242
rect 21505 10226 21521 10242
rect 21523 10226 21539 10242
rect 21623 10226 21639 10242
rect 21641 10226 21657 10242
rect 21741 10226 21757 10242
rect 21759 10226 21775 10242
rect 21859 10226 21875 10242
rect 21877 10226 21893 10242
rect 21977 10226 21993 10242
rect 21995 10226 22011 10242
rect 11237 10218 11303 10226
rect 11237 10210 11261 10218
rect 2887 1950 2892 10158
rect 2915 1950 2920 10158
rect 2975 9679 2979 9986
rect 3003 9851 3007 9958
rect 3054 9883 3075 9958
rect 3082 9957 3088 9963
rect 3128 9957 3134 9963
rect 3318 9957 3324 9963
rect 3364 9957 3370 9963
rect 3554 9957 3560 9963
rect 3600 9957 3606 9963
rect 3790 9957 3796 9963
rect 3836 9957 3842 9963
rect 4026 9957 4032 9963
rect 4072 9957 4078 9963
rect 4262 9957 4268 9963
rect 4308 9957 4314 9963
rect 4498 9957 4504 9963
rect 4544 9957 4550 9963
rect 4734 9957 4740 9963
rect 4780 9957 4786 9963
rect 4970 9957 4976 9963
rect 5016 9957 5022 9963
rect 5206 9957 5212 9963
rect 5252 9957 5258 9963
rect 5442 9957 5448 9963
rect 5488 9957 5494 9963
rect 5678 9957 5684 9963
rect 5724 9957 5730 9963
rect 5914 9957 5920 9963
rect 5960 9957 5966 9963
rect 6150 9957 6156 9963
rect 6196 9957 6202 9963
rect 6386 9957 6392 9963
rect 6432 9957 6438 9963
rect 6622 9957 6628 9963
rect 6668 9957 6674 9963
rect 6858 9957 6864 9963
rect 6904 9957 6910 9963
rect 7094 9957 7100 9963
rect 7140 9957 7146 9963
rect 7330 9957 7336 9963
rect 7376 9957 7382 9963
rect 7566 9957 7572 9963
rect 7612 9957 7618 9963
rect 7802 9957 7808 9963
rect 7848 9957 7854 9963
rect 8038 9957 8044 9963
rect 8084 9957 8090 9963
rect 8274 9957 8280 9963
rect 8320 9957 8326 9963
rect 8510 9957 8516 9963
rect 8556 9957 8562 9963
rect 8746 9957 8752 9963
rect 8792 9957 8798 9963
rect 8982 9957 8988 9963
rect 9028 9957 9034 9963
rect 3076 9951 3103 9957
rect 3134 9951 3140 9957
rect 3312 9951 3318 9957
rect 3370 9951 3376 9957
rect 3548 9951 3554 9957
rect 3606 9951 3612 9957
rect 3784 9951 3790 9957
rect 3842 9951 3848 9957
rect 4020 9951 4026 9957
rect 4078 9951 4084 9957
rect 4256 9951 4262 9957
rect 4314 9951 4320 9957
rect 4492 9951 4498 9957
rect 4550 9951 4556 9957
rect 4728 9951 4734 9957
rect 4786 9951 4792 9957
rect 4964 9951 4970 9957
rect 5022 9951 5028 9957
rect 5200 9951 5206 9957
rect 5258 9951 5264 9957
rect 5436 9951 5442 9957
rect 5494 9951 5500 9957
rect 5672 9951 5678 9957
rect 5730 9951 5736 9957
rect 5908 9951 5914 9957
rect 5966 9951 5972 9957
rect 6144 9951 6150 9957
rect 6202 9951 6208 9957
rect 6380 9951 6386 9957
rect 6438 9951 6444 9957
rect 6616 9951 6622 9957
rect 6674 9951 6680 9957
rect 6852 9951 6858 9957
rect 6910 9951 6916 9957
rect 7088 9951 7094 9957
rect 7146 9951 7152 9957
rect 7324 9951 7330 9957
rect 7382 9951 7388 9957
rect 7560 9951 7566 9957
rect 7618 9951 7624 9957
rect 7796 9951 7802 9957
rect 7854 9951 7860 9957
rect 8032 9951 8038 9957
rect 8090 9951 8096 9957
rect 8268 9951 8274 9957
rect 8326 9951 8332 9957
rect 8504 9951 8510 9957
rect 8562 9951 8568 9957
rect 8740 9951 8746 9957
rect 8798 9951 8804 9957
rect 8976 9951 8982 9957
rect 9034 9951 9040 9957
rect 3082 9883 3103 9951
rect 2991 9849 3033 9851
rect 3003 9707 3007 9849
rect 3312 9707 3318 9713
rect 3370 9707 3376 9713
rect 3548 9707 3554 9713
rect 3606 9707 3612 9713
rect 3784 9707 3790 9713
rect 3842 9707 3848 9713
rect 4020 9707 4026 9713
rect 4078 9707 4084 9713
rect 4256 9707 4262 9713
rect 4314 9707 4320 9713
rect 4492 9707 4498 9713
rect 4550 9707 4556 9713
rect 4728 9707 4734 9713
rect 4786 9707 4792 9713
rect 4964 9707 4970 9713
rect 5022 9707 5028 9713
rect 5200 9707 5206 9713
rect 5258 9707 5264 9713
rect 5436 9707 5442 9713
rect 5494 9707 5500 9713
rect 5672 9707 5678 9713
rect 5730 9707 5736 9713
rect 5908 9707 5914 9713
rect 5966 9707 5972 9713
rect 6144 9707 6150 9713
rect 6202 9707 6208 9713
rect 6380 9707 6386 9713
rect 6438 9707 6444 9713
rect 6616 9707 6622 9713
rect 6674 9707 6680 9713
rect 6852 9707 6858 9713
rect 6910 9707 6916 9713
rect 7088 9707 7094 9713
rect 7146 9707 7152 9713
rect 7324 9707 7330 9713
rect 7382 9707 7388 9713
rect 7560 9707 7566 9713
rect 7618 9707 7624 9713
rect 7796 9707 7802 9713
rect 7854 9707 7860 9713
rect 8032 9707 8038 9713
rect 8090 9707 8096 9713
rect 8268 9707 8274 9713
rect 8326 9707 8332 9713
rect 8504 9707 8510 9713
rect 8562 9707 8568 9713
rect 8740 9707 8746 9713
rect 8798 9707 8804 9713
rect 8976 9707 8982 9713
rect 9034 9707 9040 9713
rect 3318 9701 3324 9707
rect 3364 9701 3370 9707
rect 3554 9701 3560 9707
rect 3600 9701 3606 9707
rect 3790 9701 3796 9707
rect 3836 9701 3842 9707
rect 4026 9701 4032 9707
rect 4072 9701 4078 9707
rect 4262 9701 4268 9707
rect 4308 9701 4314 9707
rect 4498 9701 4504 9707
rect 4544 9701 4550 9707
rect 4734 9701 4740 9707
rect 4780 9701 4786 9707
rect 4970 9701 4976 9707
rect 5016 9701 5022 9707
rect 5206 9701 5212 9707
rect 5252 9701 5258 9707
rect 5442 9701 5448 9707
rect 5488 9701 5494 9707
rect 5678 9701 5684 9707
rect 5724 9701 5730 9707
rect 5914 9701 5920 9707
rect 5960 9701 5966 9707
rect 6150 9701 6156 9707
rect 6196 9701 6202 9707
rect 6386 9701 6392 9707
rect 6432 9701 6438 9707
rect 6622 9701 6628 9707
rect 6668 9701 6674 9707
rect 6858 9701 6864 9707
rect 6904 9701 6910 9707
rect 7094 9701 7100 9707
rect 7140 9701 7146 9707
rect 7330 9701 7336 9707
rect 7376 9701 7382 9707
rect 7566 9701 7572 9707
rect 7612 9701 7618 9707
rect 7802 9701 7808 9707
rect 7848 9701 7854 9707
rect 8038 9701 8044 9707
rect 8084 9701 8090 9707
rect 8274 9701 8280 9707
rect 8320 9701 8326 9707
rect 8510 9701 8516 9707
rect 8556 9701 8562 9707
rect 8746 9701 8752 9707
rect 8792 9701 8798 9707
rect 8982 9701 8988 9707
rect 9028 9701 9034 9707
rect 11253 9666 11261 10210
rect 11237 9658 11261 9666
rect 11279 10210 11303 10218
rect 11355 10218 11421 10226
rect 11355 10210 11379 10218
rect 11279 9666 11287 10210
rect 11371 9666 11379 10210
rect 11279 9658 11303 9666
rect 11237 9650 11303 9658
rect 11355 9658 11379 9666
rect 11397 10210 11421 10218
rect 11473 10218 11539 10226
rect 11473 10210 11497 10218
rect 11397 9666 11405 10210
rect 11489 9666 11497 10210
rect 11397 9658 11421 9666
rect 11355 9650 11421 9658
rect 11473 9658 11497 9666
rect 11515 10210 11539 10218
rect 11591 10218 11657 10226
rect 11591 10210 11615 10218
rect 11515 9666 11523 10210
rect 11607 9666 11615 10210
rect 11515 9658 11539 9666
rect 11473 9650 11539 9658
rect 11591 9658 11615 9666
rect 11633 10210 11657 10218
rect 11709 10218 11775 10226
rect 11709 10210 11733 10218
rect 11633 9666 11641 10210
rect 11725 9666 11733 10210
rect 11633 9658 11657 9666
rect 11591 9650 11657 9658
rect 11709 9658 11733 9666
rect 11751 10210 11775 10218
rect 11827 10218 11893 10226
rect 11827 10210 11851 10218
rect 11751 9666 11759 10210
rect 11843 9666 11851 10210
rect 11751 9658 11775 9666
rect 11709 9650 11775 9658
rect 11827 9658 11851 9666
rect 11869 10210 11893 10218
rect 11945 10218 12011 10226
rect 11945 10210 11969 10218
rect 11869 9666 11877 10210
rect 11961 9666 11969 10210
rect 11869 9658 11893 9666
rect 11827 9650 11893 9658
rect 11945 9658 11969 9666
rect 11987 10210 12011 10218
rect 12063 10218 12129 10226
rect 12063 10210 12087 10218
rect 11987 9666 11995 10210
rect 12079 9666 12087 10210
rect 11987 9658 12011 9666
rect 11945 9650 12011 9658
rect 12063 9658 12087 9666
rect 12105 10210 12129 10218
rect 12181 10218 12247 10226
rect 12181 10210 12205 10218
rect 12105 9666 12113 10210
rect 12197 9666 12205 10210
rect 12105 9658 12129 9666
rect 12063 9650 12129 9658
rect 12181 9658 12205 9666
rect 12223 10210 12247 10218
rect 12299 10218 12365 10226
rect 12299 10210 12323 10218
rect 12223 9666 12231 10210
rect 12315 9666 12323 10210
rect 12223 9658 12247 9666
rect 12181 9650 12247 9658
rect 12299 9658 12323 9666
rect 12341 10210 12365 10218
rect 12417 10218 12483 10226
rect 12417 10210 12441 10218
rect 12341 9666 12349 10210
rect 12433 9666 12441 10210
rect 12341 9658 12365 9666
rect 12299 9650 12365 9658
rect 12417 9658 12441 9666
rect 12459 10210 12483 10218
rect 12535 10218 12601 10226
rect 12535 10210 12559 10218
rect 12459 9666 12467 10210
rect 12551 9666 12559 10210
rect 12459 9658 12483 9666
rect 12417 9650 12483 9658
rect 12535 9658 12559 9666
rect 12577 10210 12601 10218
rect 12653 10218 12719 10226
rect 12653 10210 12677 10218
rect 12577 9666 12585 10210
rect 12669 9666 12677 10210
rect 12577 9658 12601 9666
rect 12535 9650 12601 9658
rect 12653 9658 12677 9666
rect 12695 10210 12719 10218
rect 12771 10218 12837 10226
rect 12771 10210 12795 10218
rect 12695 9666 12703 10210
rect 12787 9666 12795 10210
rect 12695 9658 12719 9666
rect 12653 9650 12719 9658
rect 12771 9658 12795 9666
rect 12813 10210 12837 10218
rect 12889 10218 12955 10226
rect 12889 10210 12913 10218
rect 12813 9666 12821 10210
rect 12905 9666 12913 10210
rect 12813 9658 12837 9666
rect 12771 9650 12837 9658
rect 12889 9658 12913 9666
rect 12931 10210 12955 10218
rect 13007 10218 13073 10226
rect 13007 10210 13031 10218
rect 12931 9666 12939 10210
rect 13023 9666 13031 10210
rect 12931 9658 12955 9666
rect 12889 9650 12955 9658
rect 13007 9658 13031 9666
rect 13049 10210 13073 10218
rect 13125 10218 13191 10226
rect 13125 10210 13149 10218
rect 13049 9666 13057 10210
rect 13141 9666 13149 10210
rect 13049 9658 13073 9666
rect 13007 9650 13073 9658
rect 13125 9658 13149 9666
rect 13167 10210 13191 10218
rect 13243 10218 13309 10226
rect 13243 10210 13267 10218
rect 13167 9666 13175 10210
rect 13259 9666 13267 10210
rect 13167 9658 13191 9666
rect 13125 9650 13191 9658
rect 13243 9658 13267 9666
rect 13285 10210 13309 10218
rect 13361 10218 13427 10226
rect 13361 10210 13385 10218
rect 13285 9666 13293 10210
rect 13377 9666 13385 10210
rect 13285 9658 13309 9666
rect 13243 9650 13309 9658
rect 13361 9658 13385 9666
rect 13403 10210 13427 10218
rect 13479 10218 13545 10226
rect 13479 10210 13503 10218
rect 13403 9666 13411 10210
rect 13495 9666 13503 10210
rect 13403 9658 13427 9666
rect 13361 9650 13427 9658
rect 13479 9658 13503 9666
rect 13521 10210 13545 10218
rect 13597 10218 13663 10226
rect 13597 10210 13621 10218
rect 13521 9666 13529 10210
rect 13613 9666 13621 10210
rect 13521 9658 13545 9666
rect 13479 9650 13545 9658
rect 13597 9658 13621 9666
rect 13639 10210 13663 10218
rect 13715 10218 13781 10226
rect 13715 10210 13739 10218
rect 13639 9666 13647 10210
rect 13731 9666 13739 10210
rect 13639 9658 13663 9666
rect 13597 9650 13663 9658
rect 13715 9658 13739 9666
rect 13757 10210 13781 10218
rect 15360 10218 15426 10226
rect 15360 10210 15384 10218
rect 13757 9666 13765 10210
rect 15376 9666 15384 10210
rect 13757 9658 13781 9666
rect 13715 9650 13781 9658
rect 15360 9658 15384 9666
rect 15402 10210 15426 10218
rect 15478 10218 15544 10226
rect 15478 10210 15502 10218
rect 15402 9666 15410 10210
rect 15494 9666 15502 10210
rect 15402 9658 15426 9666
rect 15360 9650 15426 9658
rect 15478 9658 15502 9666
rect 15520 10210 15544 10218
rect 15596 10218 15662 10226
rect 15596 10210 15620 10218
rect 15520 9666 15528 10210
rect 15612 9666 15620 10210
rect 15520 9658 15544 9666
rect 15478 9650 15544 9658
rect 15596 9658 15620 9666
rect 15638 10210 15662 10218
rect 15714 10218 15780 10226
rect 15714 10210 15738 10218
rect 15638 9666 15646 10210
rect 15730 9666 15738 10210
rect 15638 9658 15662 9666
rect 15596 9650 15662 9658
rect 15714 9658 15738 9666
rect 15756 10210 15780 10218
rect 15832 10218 15898 10226
rect 15832 10210 15856 10218
rect 15756 9666 15764 10210
rect 15848 9666 15856 10210
rect 15756 9658 15780 9666
rect 15714 9650 15780 9658
rect 15832 9658 15856 9666
rect 15874 10210 15898 10218
rect 15950 10218 16016 10226
rect 15950 10210 15974 10218
rect 15874 9666 15882 10210
rect 15966 9666 15974 10210
rect 15874 9658 15898 9666
rect 15832 9650 15898 9658
rect 15950 9658 15974 9666
rect 15992 10210 16016 10218
rect 16068 10218 16134 10226
rect 16068 10210 16092 10218
rect 15992 9666 16000 10210
rect 16084 9666 16092 10210
rect 15992 9658 16016 9666
rect 15950 9650 16016 9658
rect 16068 9658 16092 9666
rect 16110 10210 16134 10218
rect 16186 10218 16252 10226
rect 16186 10210 16210 10218
rect 16110 9666 16118 10210
rect 16202 9666 16210 10210
rect 16110 9658 16134 9666
rect 16068 9650 16134 9658
rect 16186 9658 16210 9666
rect 16228 10210 16252 10218
rect 16304 10218 16370 10226
rect 16304 10210 16328 10218
rect 16228 9666 16236 10210
rect 16320 9666 16328 10210
rect 16228 9658 16252 9666
rect 16186 9650 16252 9658
rect 16304 9658 16328 9666
rect 16346 10210 16370 10218
rect 16422 10218 16488 10226
rect 16422 10210 16446 10218
rect 16346 9666 16354 10210
rect 16438 9666 16446 10210
rect 16346 9658 16370 9666
rect 16304 9650 16370 9658
rect 16422 9658 16446 9666
rect 16464 10210 16488 10218
rect 16540 10218 16606 10226
rect 16540 10210 16564 10218
rect 16464 9666 16472 10210
rect 16556 9666 16564 10210
rect 16464 9658 16488 9666
rect 16422 9650 16488 9658
rect 16540 9658 16564 9666
rect 16582 10210 16606 10218
rect 16658 10218 16724 10226
rect 16658 10210 16682 10218
rect 16582 9666 16590 10210
rect 16674 9666 16682 10210
rect 16582 9658 16606 9666
rect 16540 9650 16606 9658
rect 16658 9658 16682 9666
rect 16700 10210 16724 10218
rect 16776 10218 16842 10226
rect 16776 10210 16800 10218
rect 16700 9666 16708 10210
rect 16792 9666 16800 10210
rect 16700 9658 16724 9666
rect 16658 9650 16724 9658
rect 16776 9658 16800 9666
rect 16818 10210 16842 10218
rect 16894 10218 16960 10226
rect 16894 10210 16918 10218
rect 16818 9666 16826 10210
rect 16910 9666 16918 10210
rect 16818 9658 16842 9666
rect 16776 9650 16842 9658
rect 16894 9658 16918 9666
rect 16936 10210 16960 10218
rect 17012 10218 17078 10226
rect 17012 10210 17036 10218
rect 16936 9666 16944 10210
rect 17028 9666 17036 10210
rect 16936 9658 16960 9666
rect 16894 9650 16960 9658
rect 17012 9658 17036 9666
rect 17054 10210 17078 10218
rect 17130 10218 17196 10226
rect 17130 10210 17154 10218
rect 17054 9666 17062 10210
rect 17146 9666 17154 10210
rect 17054 9658 17078 9666
rect 17012 9650 17078 9658
rect 17130 9658 17154 9666
rect 17172 10210 17196 10218
rect 17248 10218 17314 10226
rect 17248 10210 17272 10218
rect 17172 9666 17180 10210
rect 17264 9666 17272 10210
rect 17172 9658 17196 9666
rect 17130 9650 17196 9658
rect 17248 9658 17272 9666
rect 17290 10210 17314 10218
rect 17366 10218 17432 10226
rect 17366 10210 17390 10218
rect 17290 9666 17298 10210
rect 17382 9666 17390 10210
rect 17290 9658 17314 9666
rect 17248 9650 17314 9658
rect 17366 9658 17390 9666
rect 17408 10210 17432 10218
rect 17484 10218 17550 10226
rect 17484 10210 17508 10218
rect 17408 9666 17416 10210
rect 17500 9666 17508 10210
rect 17408 9658 17432 9666
rect 17366 9650 17432 9658
rect 17484 9658 17508 9666
rect 17526 10210 17550 10218
rect 17602 10218 17668 10226
rect 17602 10210 17626 10218
rect 17526 9666 17534 10210
rect 17618 9666 17626 10210
rect 17526 9658 17550 9666
rect 17484 9650 17550 9658
rect 17602 9658 17626 9666
rect 17644 10210 17668 10218
rect 17720 10218 17786 10226
rect 17720 10210 17744 10218
rect 17644 9666 17652 10210
rect 17736 9666 17744 10210
rect 17644 9658 17668 9666
rect 17602 9650 17668 9658
rect 17720 9658 17744 9666
rect 17762 10210 17786 10218
rect 17838 10218 17904 10226
rect 17838 10210 17862 10218
rect 17762 9666 17770 10210
rect 17854 9666 17862 10210
rect 17762 9658 17786 9666
rect 17720 9650 17786 9658
rect 17838 9658 17862 9666
rect 17880 10210 17904 10218
rect 19483 10218 19549 10226
rect 19483 10210 19507 10218
rect 17880 9666 17888 10210
rect 19499 9666 19507 10210
rect 17880 9658 17904 9666
rect 17838 9650 17904 9658
rect 19483 9658 19507 9666
rect 19525 10210 19549 10218
rect 19601 10218 19667 10226
rect 19601 10210 19625 10218
rect 19525 9666 19533 10210
rect 19617 9666 19625 10210
rect 19525 9658 19549 9666
rect 19483 9650 19549 9658
rect 19601 9658 19625 9666
rect 19643 10210 19667 10218
rect 19719 10218 19785 10226
rect 19719 10210 19743 10218
rect 19643 9666 19651 10210
rect 19735 9666 19743 10210
rect 19643 9658 19667 9666
rect 19601 9650 19667 9658
rect 19719 9658 19743 9666
rect 19761 10210 19785 10218
rect 19837 10218 19903 10226
rect 19837 10210 19861 10218
rect 19761 9666 19769 10210
rect 19853 9666 19861 10210
rect 19761 9658 19785 9666
rect 19719 9650 19785 9658
rect 19837 9658 19861 9666
rect 19879 10210 19903 10218
rect 19955 10218 20021 10226
rect 19955 10210 19979 10218
rect 19879 9666 19887 10210
rect 19971 9666 19979 10210
rect 19879 9658 19903 9666
rect 19837 9650 19903 9658
rect 19955 9658 19979 9666
rect 19997 10210 20021 10218
rect 20073 10218 20139 10226
rect 20073 10210 20097 10218
rect 19997 9666 20005 10210
rect 20089 9666 20097 10210
rect 19997 9658 20021 9666
rect 19955 9650 20021 9658
rect 20073 9658 20097 9666
rect 20115 10210 20139 10218
rect 20191 10218 20257 10226
rect 20191 10210 20215 10218
rect 20115 9666 20123 10210
rect 20207 9666 20215 10210
rect 20115 9658 20139 9666
rect 20073 9650 20139 9658
rect 20191 9658 20215 9666
rect 20233 10210 20257 10218
rect 20309 10218 20375 10226
rect 20309 10210 20333 10218
rect 20233 9666 20241 10210
rect 20325 9666 20333 10210
rect 20233 9658 20257 9666
rect 20191 9650 20257 9658
rect 20309 9658 20333 9666
rect 20351 10210 20375 10218
rect 20427 10218 20493 10226
rect 20427 10210 20451 10218
rect 20351 9666 20359 10210
rect 20443 9666 20451 10210
rect 20351 9658 20375 9666
rect 20309 9650 20375 9658
rect 20427 9658 20451 9666
rect 20469 10210 20493 10218
rect 20545 10218 20611 10226
rect 20545 10210 20569 10218
rect 20469 9666 20477 10210
rect 20561 9666 20569 10210
rect 20469 9658 20493 9666
rect 20427 9650 20493 9658
rect 20545 9658 20569 9666
rect 20587 10210 20611 10218
rect 20663 10218 20729 10226
rect 20663 10210 20687 10218
rect 20587 9666 20595 10210
rect 20679 9666 20687 10210
rect 20587 9658 20611 9666
rect 20545 9650 20611 9658
rect 20663 9658 20687 9666
rect 20705 10210 20729 10218
rect 20781 10218 20847 10226
rect 20781 10210 20805 10218
rect 20705 9666 20713 10210
rect 20797 9666 20805 10210
rect 20705 9658 20729 9666
rect 20663 9650 20729 9658
rect 20781 9658 20805 9666
rect 20823 10210 20847 10218
rect 20899 10218 20965 10226
rect 20899 10210 20923 10218
rect 20823 9666 20831 10210
rect 20915 9666 20923 10210
rect 20823 9658 20847 9666
rect 20781 9650 20847 9658
rect 20899 9658 20923 9666
rect 20941 10210 20965 10218
rect 21017 10218 21083 10226
rect 21017 10210 21041 10218
rect 20941 9666 20949 10210
rect 21033 9666 21041 10210
rect 20941 9658 20965 9666
rect 20899 9650 20965 9658
rect 21017 9658 21041 9666
rect 21059 10210 21083 10218
rect 21135 10218 21201 10226
rect 21135 10210 21159 10218
rect 21059 9666 21067 10210
rect 21151 9666 21159 10210
rect 21059 9658 21083 9666
rect 21017 9650 21083 9658
rect 21135 9658 21159 9666
rect 21177 10210 21201 10218
rect 21253 10218 21319 10226
rect 21253 10210 21277 10218
rect 21177 9666 21185 10210
rect 21269 9666 21277 10210
rect 21177 9658 21201 9666
rect 21135 9650 21201 9658
rect 21253 9658 21277 9666
rect 21295 10210 21319 10218
rect 21371 10218 21437 10226
rect 21371 10210 21395 10218
rect 21295 9666 21303 10210
rect 21387 9666 21395 10210
rect 21295 9658 21319 9666
rect 21253 9650 21319 9658
rect 21371 9658 21395 9666
rect 21413 10210 21437 10218
rect 21489 10218 21555 10226
rect 21489 10210 21513 10218
rect 21413 9666 21421 10210
rect 21505 9666 21513 10210
rect 21413 9658 21437 9666
rect 21371 9650 21437 9658
rect 21489 9658 21513 9666
rect 21531 10210 21555 10218
rect 21607 10218 21673 10226
rect 21607 10210 21631 10218
rect 21531 9666 21539 10210
rect 21623 9666 21631 10210
rect 21531 9658 21555 9666
rect 21489 9650 21555 9658
rect 21607 9658 21631 9666
rect 21649 10210 21673 10218
rect 21725 10218 21791 10226
rect 21725 10210 21749 10218
rect 21649 9666 21657 10210
rect 21741 9666 21749 10210
rect 21649 9658 21673 9666
rect 21607 9650 21673 9658
rect 21725 9658 21749 9666
rect 21767 10210 21791 10218
rect 21843 10218 21909 10226
rect 21843 10210 21867 10218
rect 21767 9666 21775 10210
rect 21859 9666 21867 10210
rect 21767 9658 21791 9666
rect 21725 9650 21791 9658
rect 21843 9658 21867 9666
rect 21885 10210 21909 10218
rect 21961 10218 22027 10226
rect 21961 10210 21985 10218
rect 21885 9666 21893 10210
rect 21977 9666 21985 10210
rect 21885 9658 21909 9666
rect 21843 9650 21909 9658
rect 21961 9658 21985 9666
rect 22003 10210 22027 10218
rect 22003 9666 22011 10210
rect 22003 9658 22027 9666
rect 21961 9650 22027 9658
rect 11253 9634 11269 9650
rect 11271 9634 11287 9650
rect 11371 9634 11387 9650
rect 11389 9634 11405 9650
rect 11489 9634 11505 9650
rect 11507 9634 11523 9650
rect 11607 9634 11623 9650
rect 11625 9634 11641 9650
rect 11725 9634 11741 9650
rect 11743 9634 11759 9650
rect 11843 9634 11859 9650
rect 11861 9634 11877 9650
rect 11961 9634 11977 9650
rect 11979 9634 11995 9650
rect 12079 9634 12095 9650
rect 12097 9634 12113 9650
rect 12197 9634 12213 9650
rect 12215 9634 12231 9650
rect 12315 9634 12331 9650
rect 12333 9634 12349 9650
rect 12433 9634 12449 9650
rect 12451 9634 12467 9650
rect 12551 9634 12567 9650
rect 12569 9634 12585 9650
rect 12669 9634 12685 9650
rect 12687 9634 12703 9650
rect 12787 9634 12803 9650
rect 12805 9634 12821 9650
rect 12905 9634 12921 9650
rect 12923 9634 12939 9650
rect 13023 9634 13039 9650
rect 13041 9634 13057 9650
rect 13141 9634 13157 9650
rect 13159 9634 13175 9650
rect 13259 9634 13275 9650
rect 13277 9634 13293 9650
rect 13377 9634 13393 9650
rect 13395 9634 13411 9650
rect 13495 9634 13511 9650
rect 13513 9634 13529 9650
rect 13613 9634 13629 9650
rect 13631 9634 13647 9650
rect 13731 9634 13747 9650
rect 13749 9634 13765 9650
rect 15376 9634 15392 9650
rect 15394 9634 15410 9650
rect 15494 9634 15510 9650
rect 15512 9634 15528 9650
rect 15612 9634 15628 9650
rect 15630 9634 15646 9650
rect 15730 9634 15746 9650
rect 15748 9634 15764 9650
rect 15848 9634 15864 9650
rect 15866 9634 15882 9650
rect 15966 9634 15982 9650
rect 15984 9634 16000 9650
rect 16084 9634 16100 9650
rect 16102 9634 16118 9650
rect 16202 9634 16218 9650
rect 16220 9634 16236 9650
rect 16320 9634 16336 9650
rect 16338 9634 16354 9650
rect 16438 9634 16454 9650
rect 16456 9634 16472 9650
rect 16556 9634 16572 9650
rect 16574 9634 16590 9650
rect 16674 9634 16690 9650
rect 16692 9634 16708 9650
rect 16792 9634 16808 9650
rect 16810 9634 16826 9650
rect 16910 9634 16926 9650
rect 16928 9634 16944 9650
rect 17028 9634 17044 9650
rect 17046 9634 17062 9650
rect 17146 9634 17162 9650
rect 17164 9634 17180 9650
rect 17264 9634 17280 9650
rect 17282 9634 17298 9650
rect 17382 9634 17398 9650
rect 17400 9634 17416 9650
rect 17500 9634 17516 9650
rect 17518 9634 17534 9650
rect 17618 9634 17634 9650
rect 17636 9634 17652 9650
rect 17736 9634 17752 9650
rect 17754 9634 17770 9650
rect 17854 9634 17870 9650
rect 17872 9634 17888 9650
rect 19499 9634 19515 9650
rect 19517 9634 19533 9650
rect 19617 9634 19633 9650
rect 19635 9634 19651 9650
rect 19735 9634 19751 9650
rect 19753 9634 19769 9650
rect 19853 9634 19869 9650
rect 19871 9634 19887 9650
rect 19971 9634 19987 9650
rect 19989 9634 20005 9650
rect 20089 9634 20105 9650
rect 20107 9634 20123 9650
rect 20207 9634 20223 9650
rect 20225 9634 20241 9650
rect 20325 9634 20341 9650
rect 20343 9634 20359 9650
rect 20443 9634 20459 9650
rect 20461 9634 20477 9650
rect 20561 9634 20577 9650
rect 20579 9634 20595 9650
rect 20679 9634 20695 9650
rect 20697 9634 20713 9650
rect 20797 9634 20813 9650
rect 20815 9634 20831 9650
rect 20915 9634 20931 9650
rect 20933 9634 20949 9650
rect 21033 9634 21049 9650
rect 21051 9634 21067 9650
rect 21151 9634 21167 9650
rect 21169 9634 21185 9650
rect 21269 9634 21285 9650
rect 21287 9634 21303 9650
rect 21387 9634 21403 9650
rect 21405 9634 21421 9650
rect 21505 9634 21521 9650
rect 21523 9634 21539 9650
rect 21623 9634 21639 9650
rect 21641 9634 21657 9650
rect 21741 9634 21757 9650
rect 21759 9634 21775 9650
rect 21859 9634 21875 9650
rect 21877 9634 21893 9650
rect 21977 9634 21993 9650
rect 21995 9634 22011 9650
rect 10760 9455 10794 9489
rect 16193 9147 16252 9310
rect 16253 9087 16312 9250
rect 16598 9060 16637 9250
rect 16658 9120 16697 9310
rect 20359 9144 20375 9342
rect 20419 9084 20435 9282
rect 2990 7905 3030 7909
rect 3563 7510 3597 7516
rect 3563 7502 3569 7510
rect 3591 7502 3597 7510
rect 3799 7510 3833 7516
rect 3799 7502 3805 7510
rect 3827 7502 3833 7510
rect 4035 7510 4069 7516
rect 4035 7502 4041 7510
rect 4063 7502 4069 7510
rect 4271 7510 4305 7516
rect 4271 7502 4277 7510
rect 4299 7502 4305 7510
rect 4507 7510 4541 7516
rect 4507 7502 4513 7510
rect 4535 7502 4541 7510
rect 4743 7510 4777 7516
rect 4743 7502 4749 7510
rect 4771 7502 4777 7510
rect 4979 7510 5013 7516
rect 4979 7502 4985 7510
rect 5007 7502 5013 7510
rect 5215 7510 5249 7516
rect 5215 7502 5221 7510
rect 5243 7502 5249 7510
rect 5451 7510 5485 7516
rect 5451 7502 5457 7510
rect 5479 7502 5485 7510
rect 5687 7510 5721 7516
rect 5687 7502 5693 7510
rect 5715 7502 5721 7510
rect 5923 7510 5957 7516
rect 5923 7502 5929 7510
rect 5951 7502 5957 7510
rect 6159 7510 6193 7516
rect 6159 7502 6165 7510
rect 6187 7502 6193 7510
rect 6395 7510 6429 7516
rect 6395 7502 6401 7510
rect 6423 7502 6429 7510
rect 6631 7510 6665 7516
rect 6631 7502 6637 7510
rect 6659 7502 6665 7510
rect 6867 7510 6901 7516
rect 6867 7502 6873 7510
rect 6895 7502 6901 7510
rect 7103 7510 7137 7516
rect 7103 7502 7109 7510
rect 7131 7502 7137 7510
rect 7339 7510 7373 7516
rect 7339 7502 7345 7510
rect 7367 7502 7373 7510
rect 7575 7510 7609 7516
rect 7575 7502 7581 7510
rect 7603 7502 7609 7510
rect 7811 7510 7845 7516
rect 7811 7502 7817 7510
rect 7839 7502 7845 7510
rect 8047 7510 8081 7516
rect 8047 7502 8053 7510
rect 8075 7502 8081 7510
rect 8283 7510 8317 7516
rect 8283 7502 8289 7510
rect 8311 7502 8317 7510
rect 8519 7510 8553 7516
rect 8519 7502 8525 7510
rect 8547 7502 8553 7510
rect 8755 7510 8789 7516
rect 8755 7502 8761 7510
rect 8783 7502 8789 7510
rect 8991 7510 9025 7516
rect 8991 7502 8997 7510
rect 9019 7502 9025 7510
rect 2984 5855 3024 5858
rect 2992 5767 3029 5771
rect 2990 3805 3029 3831
rect 2988 3717 3034 3721
rect 4035 3416 4051 3432
rect 4053 3416 4069 3432
rect 4153 3416 4169 3432
rect 4171 3416 4187 3432
rect 4271 3416 4287 3432
rect 4289 3416 4305 3432
rect 4389 3416 4405 3432
rect 4407 3416 4423 3432
rect 7339 3416 7355 3432
rect 7357 3416 7373 3432
rect 7457 3416 7473 3432
rect 7475 3416 7491 3432
rect 7575 3416 7591 3432
rect 7593 3416 7609 3432
rect 7693 3416 7709 3432
rect 7711 3416 7727 3432
rect 7811 3416 7827 3432
rect 7829 3416 7845 3432
rect 7929 3416 7945 3432
rect 7947 3416 7963 3432
rect 8047 3416 8063 3432
rect 8065 3416 8081 3432
rect 8165 3416 8181 3432
rect 8183 3416 8199 3432
rect 8283 3416 8299 3432
rect 8301 3416 8317 3432
rect 8401 3416 8417 3432
rect 8419 3416 8435 3432
rect 8519 3416 8535 3432
rect 8537 3416 8553 3432
rect 8637 3416 8653 3432
rect 8655 3416 8671 3432
rect 4019 3408 4085 3416
rect 4019 3400 4043 3408
rect 4035 2856 4043 3400
rect 4019 2848 4043 2856
rect 4061 3400 4085 3408
rect 4137 3408 4203 3416
rect 4137 3400 4161 3408
rect 4061 2856 4069 3400
rect 4153 2856 4161 3400
rect 4061 2848 4085 2856
rect 4019 2840 4085 2848
rect 4137 2848 4161 2856
rect 4179 3400 4203 3408
rect 4255 3408 4321 3416
rect 4255 3400 4279 3408
rect 4179 2856 4187 3400
rect 4271 2856 4279 3400
rect 4179 2848 4203 2856
rect 4137 2840 4203 2848
rect 4255 2848 4279 2856
rect 4297 3400 4321 3408
rect 4373 3408 4439 3416
rect 4373 3400 4397 3408
rect 4297 2856 4305 3400
rect 4389 2856 4397 3400
rect 4297 2848 4321 2856
rect 4255 2840 4321 2848
rect 4373 2848 4397 2856
rect 4415 3400 4439 3408
rect 7323 3408 7389 3416
rect 7323 3400 7347 3408
rect 4415 2856 4423 3400
rect 7339 2856 7347 3400
rect 4415 2848 4439 2856
rect 4373 2840 4439 2848
rect 7323 2848 7347 2856
rect 7365 3400 7389 3408
rect 7441 3408 7507 3416
rect 7441 3400 7465 3408
rect 7365 2856 7373 3400
rect 7457 2856 7465 3400
rect 7365 2848 7389 2856
rect 7323 2840 7389 2848
rect 7441 2848 7465 2856
rect 7483 3400 7507 3408
rect 7559 3408 7625 3416
rect 7559 3400 7583 3408
rect 7483 2856 7491 3400
rect 7575 2856 7583 3400
rect 7483 2848 7507 2856
rect 7441 2840 7507 2848
rect 7559 2848 7583 2856
rect 7601 3400 7625 3408
rect 7677 3408 7743 3416
rect 7677 3400 7701 3408
rect 7601 2856 7609 3400
rect 7693 2856 7701 3400
rect 7601 2848 7625 2856
rect 7559 2840 7625 2848
rect 7677 2848 7701 2856
rect 7719 3400 7743 3408
rect 7795 3408 7861 3416
rect 7795 3400 7819 3408
rect 7719 2856 7727 3400
rect 7811 2856 7819 3400
rect 7719 2848 7743 2856
rect 7677 2840 7743 2848
rect 7795 2848 7819 2856
rect 7837 3400 7861 3408
rect 7913 3408 7979 3416
rect 7913 3400 7937 3408
rect 7837 2856 7845 3400
rect 7929 2856 7937 3400
rect 7837 2848 7861 2856
rect 7795 2840 7861 2848
rect 7913 2848 7937 2856
rect 7955 3400 7979 3408
rect 8031 3408 8097 3416
rect 8031 3400 8055 3408
rect 7955 2856 7963 3400
rect 8047 2856 8055 3400
rect 7955 2848 7979 2856
rect 7913 2840 7979 2848
rect 8031 2848 8055 2856
rect 8073 3400 8097 3408
rect 8149 3408 8215 3416
rect 8149 3400 8173 3408
rect 8073 2856 8081 3400
rect 8165 2856 8173 3400
rect 8073 2848 8097 2856
rect 8031 2840 8097 2848
rect 8149 2848 8173 2856
rect 8191 3400 8215 3408
rect 8267 3408 8333 3416
rect 8267 3400 8291 3408
rect 8191 2856 8199 3400
rect 8283 2856 8291 3400
rect 8191 2848 8215 2856
rect 8149 2840 8215 2848
rect 8267 2848 8291 2856
rect 8309 3400 8333 3408
rect 8385 3408 8451 3416
rect 8385 3400 8409 3408
rect 8309 2856 8317 3400
rect 8401 2856 8409 3400
rect 8309 2848 8333 2856
rect 8267 2840 8333 2848
rect 8385 2848 8409 2856
rect 8427 3400 8451 3408
rect 8503 3408 8569 3416
rect 8503 3400 8527 3408
rect 8427 2856 8435 3400
rect 8519 2856 8527 3400
rect 8427 2848 8451 2856
rect 8385 2840 8451 2848
rect 8503 2848 8527 2856
rect 8545 3400 8569 3408
rect 8621 3408 8687 3416
rect 8621 3400 8645 3408
rect 8545 2856 8553 3400
rect 8637 2856 8645 3400
rect 8545 2848 8569 2856
rect 8503 2840 8569 2848
rect 8621 2848 8645 2856
rect 8663 3400 8687 3408
rect 8663 2856 8671 3400
rect 8663 2848 8687 2856
rect 8621 2840 8687 2848
rect 4035 2824 4051 2840
rect 4053 2824 4069 2840
rect 4153 2824 4169 2840
rect 4171 2824 4187 2840
rect 4271 2824 4287 2840
rect 4289 2824 4305 2840
rect 4389 2824 4405 2840
rect 4407 2824 4423 2840
rect 7339 2824 7355 2840
rect 7357 2824 7373 2840
rect 7457 2824 7473 2840
rect 7475 2824 7491 2840
rect 7575 2824 7591 2840
rect 7593 2824 7609 2840
rect 7693 2824 7709 2840
rect 7711 2824 7727 2840
rect 7811 2824 7827 2840
rect 7829 2824 7845 2840
rect 7929 2824 7945 2840
rect 7947 2824 7963 2840
rect 8047 2824 8063 2840
rect 8065 2824 8081 2840
rect 8165 2824 8181 2840
rect 8183 2824 8199 2840
rect 8283 2824 8299 2840
rect 8301 2824 8317 2840
rect 8401 2824 8417 2840
rect 8419 2824 8435 2840
rect 8519 2824 8535 2840
rect 8537 2824 8553 2840
rect 8637 2824 8653 2840
rect 8655 2824 8671 2840
rect 4035 2580 4051 2596
rect 4053 2580 4069 2596
rect 4153 2580 4169 2596
rect 4171 2580 4187 2596
rect 4271 2580 4287 2596
rect 4289 2580 4305 2596
rect 4389 2580 4405 2596
rect 4407 2580 4423 2596
rect 7339 2580 7355 2596
rect 7357 2580 7373 2596
rect 7457 2580 7473 2596
rect 7475 2580 7491 2596
rect 7575 2580 7591 2596
rect 7593 2580 7609 2596
rect 7693 2580 7709 2596
rect 7711 2580 7727 2596
rect 7811 2580 7827 2596
rect 7829 2580 7845 2596
rect 7929 2580 7945 2596
rect 7947 2580 7963 2596
rect 8047 2580 8063 2596
rect 8065 2580 8081 2596
rect 8165 2580 8181 2596
rect 8183 2580 8199 2596
rect 8283 2580 8299 2596
rect 8301 2580 8317 2596
rect 8401 2580 8417 2596
rect 8419 2580 8435 2596
rect 8519 2580 8535 2596
rect 8537 2580 8553 2596
rect 8637 2580 8653 2596
rect 8655 2580 8671 2596
rect 4019 2572 4085 2580
rect 4019 2564 4043 2572
rect 4035 2020 4043 2564
rect 4019 2012 4043 2020
rect 4061 2564 4085 2572
rect 4137 2572 4203 2580
rect 4137 2564 4161 2572
rect 4061 2020 4069 2564
rect 4153 2020 4161 2564
rect 4061 2012 4085 2020
rect 4019 2004 4085 2012
rect 4137 2012 4161 2020
rect 4179 2564 4203 2572
rect 4255 2572 4321 2580
rect 4255 2564 4279 2572
rect 4179 2020 4187 2564
rect 4271 2020 4279 2564
rect 4179 2012 4203 2020
rect 4137 2004 4203 2012
rect 4255 2012 4279 2020
rect 4297 2564 4321 2572
rect 4373 2572 4439 2580
rect 4373 2564 4397 2572
rect 4297 2020 4305 2564
rect 4389 2020 4397 2564
rect 4297 2012 4321 2020
rect 4255 2004 4321 2012
rect 4373 2012 4397 2020
rect 4415 2564 4439 2572
rect 7323 2572 7389 2580
rect 7323 2564 7347 2572
rect 4415 2020 4423 2564
rect 7339 2020 7347 2564
rect 4415 2012 4439 2020
rect 4373 2004 4439 2012
rect 7323 2012 7347 2020
rect 7365 2564 7389 2572
rect 7441 2572 7507 2580
rect 7441 2564 7465 2572
rect 7365 2020 7373 2564
rect 7457 2020 7465 2564
rect 7365 2012 7389 2020
rect 7323 2004 7389 2012
rect 7441 2012 7465 2020
rect 7483 2564 7507 2572
rect 7559 2572 7625 2580
rect 7559 2564 7583 2572
rect 7483 2020 7491 2564
rect 7575 2020 7583 2564
rect 7483 2012 7507 2020
rect 7441 2004 7507 2012
rect 7559 2012 7583 2020
rect 7601 2564 7625 2572
rect 7677 2572 7743 2580
rect 7677 2564 7701 2572
rect 7601 2020 7609 2564
rect 7693 2020 7701 2564
rect 7601 2012 7625 2020
rect 7559 2004 7625 2012
rect 7677 2012 7701 2020
rect 7719 2564 7743 2572
rect 7795 2572 7861 2580
rect 7795 2564 7819 2572
rect 7719 2020 7727 2564
rect 7811 2020 7819 2564
rect 7719 2012 7743 2020
rect 7677 2004 7743 2012
rect 7795 2012 7819 2020
rect 7837 2564 7861 2572
rect 7913 2572 7979 2580
rect 7913 2564 7937 2572
rect 7837 2020 7845 2564
rect 7929 2020 7937 2564
rect 7837 2012 7861 2020
rect 7795 2004 7861 2012
rect 7913 2012 7937 2020
rect 7955 2564 7979 2572
rect 8031 2572 8097 2580
rect 8031 2564 8055 2572
rect 7955 2020 7963 2564
rect 8047 2020 8055 2564
rect 7955 2012 7979 2020
rect 7913 2004 7979 2012
rect 8031 2012 8055 2020
rect 8073 2564 8097 2572
rect 8149 2572 8215 2580
rect 8149 2564 8173 2572
rect 8073 2020 8081 2564
rect 8165 2020 8173 2564
rect 8073 2012 8097 2020
rect 8031 2004 8097 2012
rect 8149 2012 8173 2020
rect 8191 2564 8215 2572
rect 8267 2572 8333 2580
rect 8267 2564 8291 2572
rect 8191 2020 8199 2564
rect 8283 2020 8291 2564
rect 8191 2012 8215 2020
rect 8149 2004 8215 2012
rect 8267 2012 8291 2020
rect 8309 2564 8333 2572
rect 8385 2572 8451 2580
rect 8385 2564 8409 2572
rect 8309 2020 8317 2564
rect 8401 2020 8409 2564
rect 8309 2012 8333 2020
rect 8267 2004 8333 2012
rect 8385 2012 8409 2020
rect 8427 2564 8451 2572
rect 8503 2572 8569 2580
rect 8503 2564 8527 2572
rect 8427 2020 8435 2564
rect 8519 2020 8527 2564
rect 8427 2012 8451 2020
rect 8385 2004 8451 2012
rect 8503 2012 8527 2020
rect 8545 2564 8569 2572
rect 8621 2572 8687 2580
rect 8621 2564 8645 2572
rect 8545 2020 8553 2564
rect 8637 2020 8645 2564
rect 8545 2012 8569 2020
rect 8503 2004 8569 2012
rect 8621 2012 8645 2020
rect 8663 2564 8687 2572
rect 8663 2020 8671 2564
rect 8663 2012 8687 2020
rect 8621 2004 8687 2012
rect 4035 1988 4051 2004
rect 4053 1988 4069 2004
rect 4153 1988 4169 2004
rect 4171 1988 4187 2004
rect 4271 1988 4287 2004
rect 4289 1988 4305 2004
rect 4389 1988 4405 2004
rect 4407 1988 4423 2004
rect 7339 1988 7355 2004
rect 7357 1988 7373 2004
rect 7457 1988 7473 2004
rect 7475 1988 7491 2004
rect 7575 1988 7591 2004
rect 7593 1988 7609 2004
rect 7693 1988 7709 2004
rect 7711 1988 7727 2004
rect 7811 1988 7827 2004
rect 7829 1988 7845 2004
rect 7929 1988 7945 2004
rect 7947 1988 7963 2004
rect 8047 1988 8063 2004
rect 8065 1988 8081 2004
rect 8165 1988 8181 2004
rect 8183 1988 8199 2004
rect 8283 1988 8299 2004
rect 8301 1988 8317 2004
rect 8401 1988 8417 2004
rect 8419 1988 8435 2004
rect 8519 1988 8535 2004
rect 8537 1988 8553 2004
rect 8637 1988 8653 2004
rect 8655 1988 8671 2004
rect 2919 1878 2937 1932
rect 2947 1878 2965 1932
rect 2956 1850 2965 1878
rect 3318 1863 3324 1869
rect 3364 1863 3370 1869
rect 3554 1863 3560 1869
rect 3600 1863 3606 1869
rect 3790 1863 3796 1869
rect 3836 1863 3842 1869
rect 4026 1863 4032 1869
rect 4072 1863 4078 1869
rect 4262 1863 4268 1869
rect 4308 1863 4314 1869
rect 4498 1863 4504 1869
rect 4544 1863 4550 1869
rect 4734 1863 4740 1869
rect 4780 1863 4786 1869
rect 4970 1863 4976 1869
rect 5016 1863 5022 1869
rect 5206 1863 5212 1869
rect 5252 1863 5258 1869
rect 5442 1863 5448 1869
rect 5488 1863 5494 1869
rect 5678 1863 5684 1869
rect 5724 1863 5730 1869
rect 5914 1863 5920 1869
rect 5960 1863 5966 1869
rect 6150 1863 6156 1869
rect 6196 1863 6202 1869
rect 6386 1863 6392 1869
rect 6432 1863 6438 1869
rect 6622 1863 6628 1869
rect 6668 1863 6674 1869
rect 6858 1863 6864 1869
rect 6904 1863 6910 1869
rect 7094 1863 7100 1869
rect 7140 1863 7146 1869
rect 7330 1863 7336 1869
rect 7376 1863 7382 1869
rect 7566 1863 7572 1869
rect 7612 1863 7618 1869
rect 7802 1863 7808 1869
rect 7848 1863 7854 1869
rect 8038 1863 8044 1869
rect 8084 1863 8090 1869
rect 8274 1863 8280 1869
rect 8320 1863 8326 1869
rect 8510 1863 8516 1869
rect 8556 1863 8562 1869
rect 8746 1863 8752 1869
rect 8792 1863 8798 1869
rect 8982 1863 8988 1869
rect 9028 1863 9034 1869
rect 3312 1857 3318 1863
rect 3370 1857 3376 1863
rect 3548 1857 3554 1863
rect 3606 1857 3612 1863
rect 3784 1857 3790 1863
rect 3842 1857 3848 1863
rect 4020 1857 4026 1863
rect 4078 1857 4084 1863
rect 4256 1857 4262 1863
rect 4314 1857 4320 1863
rect 4492 1857 4498 1863
rect 4550 1857 4556 1863
rect 4728 1857 4734 1863
rect 4786 1857 4792 1863
rect 4964 1857 4970 1863
rect 5022 1857 5028 1863
rect 5200 1857 5206 1863
rect 5258 1857 5264 1863
rect 5436 1857 5442 1863
rect 5494 1857 5500 1863
rect 5672 1857 5678 1863
rect 5730 1857 5736 1863
rect 5908 1857 5914 1863
rect 5966 1857 5972 1863
rect 6144 1857 6150 1863
rect 6202 1857 6208 1863
rect 6380 1857 6386 1863
rect 6438 1857 6444 1863
rect 6616 1857 6622 1863
rect 6674 1857 6680 1863
rect 6852 1857 6858 1863
rect 6910 1857 6916 1863
rect 7088 1857 7094 1863
rect 7146 1857 7152 1863
rect 7324 1857 7330 1863
rect 7382 1857 7388 1863
rect 7560 1857 7566 1863
rect 7618 1857 7624 1863
rect 7796 1857 7802 1863
rect 7854 1857 7860 1863
rect 8032 1857 8038 1863
rect 8090 1857 8096 1863
rect 8268 1857 8274 1863
rect 8326 1857 8332 1863
rect 8504 1857 8510 1863
rect 8562 1857 8568 1863
rect 8740 1857 8746 1863
rect 8798 1857 8804 1863
rect 8976 1857 8982 1863
rect 9034 1857 9040 1863
rect 3313 1778 9103 1791
rect 3277 1742 9067 1755
rect 15714 1645 15738 1731
rect 16050 1647 16076 1731
rect 3312 1613 3318 1619
rect 3370 1613 3376 1619
rect 3548 1613 3554 1619
rect 3606 1613 3612 1619
rect 3784 1613 3790 1619
rect 3842 1613 3848 1619
rect 4020 1613 4026 1619
rect 4078 1613 4084 1619
rect 4256 1613 4262 1619
rect 4314 1613 4320 1619
rect 4492 1613 4498 1619
rect 4550 1613 4556 1619
rect 4728 1613 4734 1619
rect 4786 1613 4792 1619
rect 4964 1613 4970 1619
rect 5022 1613 5028 1619
rect 5200 1613 5206 1619
rect 5258 1613 5264 1619
rect 5436 1613 5442 1619
rect 5494 1613 5500 1619
rect 5672 1613 5678 1619
rect 5730 1613 5736 1619
rect 5908 1613 5914 1619
rect 5966 1613 5972 1619
rect 6144 1613 6150 1619
rect 6202 1613 6208 1619
rect 6380 1613 6386 1619
rect 6438 1613 6444 1619
rect 6616 1613 6622 1619
rect 6674 1613 6680 1619
rect 6852 1613 6858 1619
rect 6910 1613 6916 1619
rect 7088 1613 7094 1619
rect 7146 1613 7152 1619
rect 7324 1613 7330 1619
rect 7382 1613 7388 1619
rect 7560 1613 7566 1619
rect 7618 1613 7624 1619
rect 7796 1613 7802 1619
rect 7854 1613 7860 1619
rect 8032 1613 8038 1619
rect 8090 1613 8096 1619
rect 8268 1613 8274 1619
rect 8326 1613 8332 1619
rect 8504 1613 8510 1619
rect 8562 1613 8568 1619
rect 8740 1613 8746 1619
rect 8798 1613 8804 1619
rect 8976 1613 8982 1619
rect 9034 1613 9040 1619
rect 3318 1607 3324 1613
rect 3364 1607 3370 1613
rect 3554 1607 3560 1613
rect 3600 1607 3606 1613
rect 3790 1607 3796 1613
rect 3836 1607 3842 1613
rect 4026 1607 4032 1613
rect 4072 1607 4078 1613
rect 4262 1607 4268 1613
rect 4308 1607 4314 1613
rect 4498 1607 4504 1613
rect 4544 1607 4550 1613
rect 4734 1607 4740 1613
rect 4780 1607 4786 1613
rect 4970 1607 4976 1613
rect 5016 1607 5022 1613
rect 5206 1607 5212 1613
rect 5252 1607 5258 1613
rect 5442 1607 5448 1613
rect 5488 1607 5494 1613
rect 5678 1607 5684 1613
rect 5724 1607 5730 1613
rect 5914 1607 5920 1613
rect 5960 1607 5966 1613
rect 6150 1607 6156 1613
rect 6196 1607 6202 1613
rect 6386 1607 6392 1613
rect 6432 1607 6438 1613
rect 6622 1607 6628 1613
rect 6668 1607 6674 1613
rect 6858 1607 6864 1613
rect 6904 1607 6910 1613
rect 7094 1607 7100 1613
rect 7140 1607 7146 1613
rect 7330 1607 7336 1613
rect 7376 1607 7382 1613
rect 7566 1607 7572 1613
rect 7612 1607 7618 1613
rect 7802 1607 7808 1613
rect 7848 1607 7854 1613
rect 8038 1607 8044 1613
rect 8084 1607 8090 1613
rect 8274 1607 8280 1613
rect 8320 1607 8326 1613
rect 8510 1607 8516 1613
rect 8556 1607 8562 1613
rect 8746 1607 8752 1613
rect 8792 1607 8798 1613
rect 8982 1607 8988 1613
rect 9028 1607 9034 1613
rect 4629 1173 4645 1189
rect 4647 1173 4663 1189
rect 4747 1173 4763 1189
rect 4765 1173 4781 1189
rect 4865 1173 4881 1189
rect 4883 1173 4899 1189
rect 4983 1173 4999 1189
rect 5001 1173 5017 1189
rect 6155 1173 6171 1189
rect 6173 1173 6189 1189
rect 6273 1173 6289 1189
rect 6291 1173 6307 1189
rect 6391 1173 6407 1189
rect 6409 1173 6425 1189
rect 6509 1173 6525 1189
rect 6527 1173 6543 1189
rect 6627 1173 6643 1189
rect 6645 1173 6661 1189
rect 6745 1173 6761 1189
rect 6763 1173 6779 1189
rect 6863 1173 6879 1189
rect 6881 1173 6897 1189
rect 6981 1173 6997 1189
rect 6999 1173 7015 1189
rect 7099 1173 7115 1189
rect 7117 1173 7133 1189
rect 7217 1173 7233 1189
rect 7235 1173 7251 1189
rect 7335 1173 7351 1189
rect 7353 1173 7369 1189
rect 7453 1173 7469 1189
rect 7471 1173 7487 1189
rect 7571 1173 7587 1189
rect 7589 1173 7605 1189
rect 7689 1173 7705 1189
rect 7707 1173 7723 1189
rect 7807 1173 7823 1189
rect 7825 1173 7841 1189
rect 7925 1173 7941 1189
rect 7943 1173 7959 1189
rect 4613 1165 4679 1173
rect 4613 1157 4637 1165
rect 4629 613 4637 1157
rect 4613 605 4637 613
rect 4655 1157 4679 1165
rect 4731 1165 4797 1173
rect 4731 1157 4755 1165
rect 4655 613 4663 1157
rect 4747 613 4755 1157
rect 4655 605 4679 613
rect 4613 597 4679 605
rect 4731 605 4755 613
rect 4773 1157 4797 1165
rect 4849 1165 4915 1173
rect 4849 1157 4873 1165
rect 4773 613 4781 1157
rect 4865 613 4873 1157
rect 4773 605 4797 613
rect 4731 597 4797 605
rect 4849 605 4873 613
rect 4891 1157 4915 1165
rect 4967 1165 5033 1173
rect 4967 1157 4991 1165
rect 4891 613 4899 1157
rect 4983 613 4991 1157
rect 4891 605 4915 613
rect 4849 597 4915 605
rect 4967 605 4991 613
rect 5009 1157 5033 1165
rect 6139 1165 6205 1173
rect 6139 1157 6163 1165
rect 5009 613 5017 1157
rect 6155 613 6163 1157
rect 5009 605 5033 613
rect 4967 597 5033 605
rect 6139 605 6163 613
rect 6181 1157 6205 1165
rect 6257 1165 6323 1173
rect 6257 1157 6281 1165
rect 6181 613 6189 1157
rect 6273 613 6281 1157
rect 6181 605 6205 613
rect 6139 597 6205 605
rect 6257 605 6281 613
rect 6299 1157 6323 1165
rect 6375 1165 6441 1173
rect 6375 1157 6399 1165
rect 6299 613 6307 1157
rect 6391 613 6399 1157
rect 6299 605 6323 613
rect 6257 597 6323 605
rect 6375 605 6399 613
rect 6417 1157 6441 1165
rect 6493 1165 6559 1173
rect 6493 1157 6517 1165
rect 6417 613 6425 1157
rect 6509 613 6517 1157
rect 6417 605 6441 613
rect 6375 597 6441 605
rect 6493 605 6517 613
rect 6535 1157 6559 1165
rect 6611 1165 6677 1173
rect 6611 1157 6635 1165
rect 6535 613 6543 1157
rect 6627 613 6635 1157
rect 6535 605 6559 613
rect 6493 597 6559 605
rect 6611 605 6635 613
rect 6653 1157 6677 1165
rect 6729 1165 6795 1173
rect 6729 1157 6753 1165
rect 6653 613 6661 1157
rect 6745 613 6753 1157
rect 6653 605 6677 613
rect 6611 597 6677 605
rect 6729 605 6753 613
rect 6771 1157 6795 1165
rect 6847 1165 6913 1173
rect 6847 1157 6871 1165
rect 6771 613 6779 1157
rect 6863 613 6871 1157
rect 6771 605 6795 613
rect 6729 597 6795 605
rect 6847 605 6871 613
rect 6889 1157 6913 1165
rect 6965 1165 7031 1173
rect 6965 1157 6989 1165
rect 6889 613 6897 1157
rect 6981 613 6989 1157
rect 6889 605 6913 613
rect 6847 597 6913 605
rect 6965 605 6989 613
rect 7007 1157 7031 1165
rect 7083 1165 7149 1173
rect 7083 1157 7107 1165
rect 7007 613 7015 1157
rect 7099 613 7107 1157
rect 7007 605 7031 613
rect 6965 597 7031 605
rect 7083 605 7107 613
rect 7125 1157 7149 1165
rect 7201 1165 7267 1173
rect 7201 1157 7225 1165
rect 7125 613 7133 1157
rect 7217 613 7225 1157
rect 7125 605 7149 613
rect 7083 597 7149 605
rect 7201 605 7225 613
rect 7243 1157 7267 1165
rect 7319 1165 7385 1173
rect 7319 1157 7343 1165
rect 7243 613 7251 1157
rect 7335 613 7343 1157
rect 7243 605 7267 613
rect 7201 597 7267 605
rect 7319 605 7343 613
rect 7361 1157 7385 1165
rect 7437 1165 7503 1173
rect 7437 1157 7461 1165
rect 7361 613 7369 1157
rect 7453 613 7461 1157
rect 7361 605 7385 613
rect 7319 597 7385 605
rect 7437 605 7461 613
rect 7479 1157 7503 1165
rect 7555 1165 7621 1173
rect 7555 1157 7579 1165
rect 7479 613 7487 1157
rect 7571 613 7579 1157
rect 7479 605 7503 613
rect 7437 597 7503 605
rect 7555 605 7579 613
rect 7597 1157 7621 1165
rect 7673 1165 7739 1173
rect 7673 1157 7697 1165
rect 7597 613 7605 1157
rect 7689 613 7697 1157
rect 7597 605 7621 613
rect 7555 597 7621 605
rect 7673 605 7697 613
rect 7715 1157 7739 1165
rect 7791 1165 7857 1173
rect 7791 1157 7815 1165
rect 7715 613 7723 1157
rect 7807 613 7815 1157
rect 7715 605 7739 613
rect 7673 597 7739 605
rect 7791 605 7815 613
rect 7833 1157 7857 1165
rect 7909 1165 7975 1173
rect 7909 1157 7933 1165
rect 7833 613 7841 1157
rect 7925 613 7933 1157
rect 7833 605 7857 613
rect 7791 597 7857 605
rect 7909 605 7933 613
rect 7951 1157 7975 1165
rect 8702 1163 8736 1197
rect 11999 1173 12015 1189
rect 12017 1173 12033 1189
rect 12147 1173 12163 1189
rect 12165 1173 12181 1189
rect 12295 1173 12311 1189
rect 12313 1173 12329 1189
rect 12443 1173 12459 1189
rect 12461 1173 12477 1189
rect 12591 1173 12607 1189
rect 12609 1173 12625 1189
rect 12739 1173 12755 1189
rect 12757 1173 12773 1189
rect 12887 1173 12903 1189
rect 12905 1173 12921 1189
rect 13035 1173 13051 1189
rect 13053 1173 13069 1189
rect 13183 1173 13199 1189
rect 13201 1173 13217 1189
rect 13331 1173 13347 1189
rect 13349 1173 13365 1189
rect 13479 1173 13495 1189
rect 13497 1173 13513 1189
rect 13627 1173 13643 1189
rect 13645 1173 13661 1189
rect 13775 1173 13791 1189
rect 13793 1173 13809 1189
rect 13923 1173 13939 1189
rect 13941 1173 13957 1189
rect 14071 1173 14087 1189
rect 14089 1173 14105 1189
rect 14219 1173 14235 1189
rect 14237 1173 14253 1189
rect 14367 1173 14383 1189
rect 14385 1173 14401 1189
rect 14515 1173 14531 1189
rect 14533 1173 14549 1189
rect 14663 1173 14679 1189
rect 14681 1173 14697 1189
rect 14811 1173 14827 1189
rect 14829 1173 14845 1189
rect 14959 1173 14975 1189
rect 14977 1173 14993 1189
rect 15107 1173 15123 1189
rect 15125 1173 15141 1189
rect 15255 1173 15271 1189
rect 15273 1173 15289 1189
rect 15403 1173 15419 1189
rect 15421 1173 15437 1189
rect 15551 1173 15567 1189
rect 15569 1173 15585 1189
rect 15699 1173 15715 1189
rect 15717 1173 15733 1189
rect 15847 1173 15863 1189
rect 15865 1173 15881 1189
rect 15995 1173 16011 1189
rect 16013 1173 16029 1189
rect 16143 1173 16159 1189
rect 16161 1173 16177 1189
rect 16291 1173 16307 1189
rect 16309 1173 16325 1189
rect 16439 1173 16455 1189
rect 16457 1173 16473 1189
rect 16587 1173 16603 1189
rect 16605 1173 16621 1189
rect 16735 1173 16751 1189
rect 16753 1173 16769 1189
rect 16883 1173 16899 1189
rect 16901 1173 16917 1189
rect 17031 1173 17047 1189
rect 17049 1173 17065 1189
rect 17179 1173 17195 1189
rect 17197 1173 17213 1189
rect 17327 1173 17343 1189
rect 17345 1173 17361 1189
rect 17475 1173 17491 1189
rect 17493 1173 17509 1189
rect 17623 1173 17639 1189
rect 17641 1173 17657 1189
rect 17771 1173 17787 1189
rect 17789 1173 17805 1189
rect 17919 1173 17935 1189
rect 17937 1173 17953 1189
rect 18067 1173 18083 1189
rect 18085 1173 18101 1189
rect 18215 1173 18231 1189
rect 18233 1173 18249 1189
rect 18363 1173 18379 1189
rect 18381 1173 18397 1189
rect 18511 1173 18527 1189
rect 18529 1173 18545 1189
rect 18659 1173 18675 1189
rect 18677 1173 18693 1189
rect 18807 1173 18823 1189
rect 18825 1173 18841 1189
rect 18955 1173 18971 1189
rect 18973 1173 18989 1189
rect 19103 1173 19119 1189
rect 19121 1173 19137 1189
rect 19251 1173 19267 1189
rect 19269 1173 19285 1189
rect 19399 1173 19415 1189
rect 19417 1173 19433 1189
rect 19547 1173 19563 1189
rect 19565 1173 19581 1189
rect 19695 1173 19711 1189
rect 19713 1173 19729 1189
rect 19843 1173 19859 1189
rect 19861 1173 19877 1189
rect 19991 1173 20007 1189
rect 20009 1173 20025 1189
rect 20139 1173 20155 1189
rect 20157 1173 20160 1189
rect 11983 1165 12049 1173
rect 11983 1157 12007 1165
rect 7951 613 7959 1157
rect 8702 1129 8736 1154
rect 9208 873 9232 1023
rect 9524 873 9548 1023
rect 9840 873 9864 1023
rect 10156 873 10180 1023
rect 10472 873 10496 1023
rect 8702 748 8736 787
rect 9018 773 9052 787
rect 8994 739 9052 773
rect 9334 739 9368 787
rect 9650 739 9684 787
rect 9966 739 10000 787
rect 10282 739 10316 787
rect 10598 739 10632 787
rect 9028 733 9052 739
rect 8775 699 8809 733
rect 8848 699 8882 733
rect 8921 699 8955 733
rect 9067 699 9101 733
rect 9140 699 9174 733
rect 9213 699 9247 733
rect 9286 699 9320 733
rect 9359 699 9393 733
rect 9432 699 9466 733
rect 9505 699 9539 733
rect 9578 699 9612 733
rect 9651 699 9685 733
rect 9724 699 9758 733
rect 9797 699 9831 733
rect 9870 699 9904 733
rect 9943 699 9977 733
rect 10016 699 10050 733
rect 10089 699 10123 733
rect 10162 699 10196 733
rect 10235 699 10269 733
rect 10308 699 10342 733
rect 10381 699 10415 733
rect 10454 699 10488 733
rect 10527 699 10561 733
rect 10600 699 10634 733
rect 7951 605 7975 613
rect 7909 597 7975 605
rect 4629 581 4645 597
rect 4647 581 4663 597
rect 4747 581 4763 597
rect 4765 581 4781 597
rect 4865 581 4881 597
rect 4883 581 4899 597
rect 4983 581 4999 597
rect 5001 581 5017 597
rect 6155 581 6171 597
rect 6173 581 6189 597
rect 6273 581 6289 597
rect 6291 581 6307 597
rect 6391 581 6407 597
rect 6409 581 6425 597
rect 6509 581 6525 597
rect 6527 581 6543 597
rect 6627 581 6643 597
rect 6645 581 6661 597
rect 6745 581 6761 597
rect 6763 581 6779 597
rect 6863 581 6879 597
rect 6881 581 6897 597
rect 6981 581 6997 597
rect 6999 581 7015 597
rect 7099 581 7115 597
rect 7117 581 7133 597
rect 7217 581 7233 597
rect 7235 581 7251 597
rect 7335 581 7351 597
rect 7353 581 7369 597
rect 7453 581 7469 597
rect 7471 581 7487 597
rect 7571 581 7587 597
rect 7589 581 7605 597
rect 7689 581 7705 597
rect 7707 581 7723 597
rect 7807 581 7823 597
rect 7825 581 7841 597
rect 7925 581 7941 597
rect 7943 581 7959 597
rect 6184 563 6278 577
rect 6184 547 6198 563
rect 6214 547 6248 555
rect 6214 513 6228 547
rect 6248 513 6256 547
rect 6264 513 6278 563
rect 6302 563 6396 577
rect 6302 547 6316 563
rect 6332 547 6366 555
rect 6332 513 6346 547
rect 6366 513 6374 547
rect 6382 513 6396 563
rect 6420 563 6514 577
rect 6420 547 6434 563
rect 6450 547 6484 555
rect 6450 513 6464 547
rect 6484 513 6492 547
rect 6500 513 6514 563
rect 6538 563 6632 577
rect 6538 547 6552 563
rect 6568 547 6602 555
rect 6568 513 6582 547
rect 6602 513 6610 547
rect 6618 513 6632 563
rect 6656 563 6750 577
rect 6656 547 6670 563
rect 6686 547 6720 555
rect 6686 513 6700 547
rect 6720 513 6728 547
rect 6736 513 6750 563
rect 6774 563 6868 577
rect 6774 547 6788 563
rect 6804 547 6838 555
rect 6804 513 6818 547
rect 6838 513 6846 547
rect 6854 513 6868 563
rect 6892 563 6986 577
rect 6892 547 6906 563
rect 6922 547 6956 555
rect 6922 513 6936 547
rect 6956 513 6964 547
rect 6972 513 6986 563
rect 7010 563 7104 577
rect 7010 547 7024 563
rect 7040 547 7074 555
rect 7040 513 7054 547
rect 7074 513 7082 547
rect 7090 513 7104 563
rect 7128 563 7222 577
rect 7128 547 7142 563
rect 7158 547 7192 555
rect 7158 513 7172 547
rect 7192 513 7200 547
rect 7208 513 7222 563
rect 7246 563 7340 577
rect 7246 547 7260 563
rect 7276 547 7310 555
rect 7276 513 7290 547
rect 7310 513 7318 547
rect 7326 513 7340 563
rect 7364 563 7458 577
rect 7364 547 7378 563
rect 7394 547 7428 555
rect 7394 513 7408 547
rect 7428 513 7436 547
rect 7444 513 7458 563
rect 7482 563 7576 577
rect 7482 547 7496 563
rect 7512 547 7546 555
rect 7512 513 7526 547
rect 7546 513 7554 547
rect 7562 513 7576 563
rect 7600 563 7694 577
rect 7600 547 7614 563
rect 7630 547 7664 555
rect 7630 513 7644 547
rect 7664 513 7672 547
rect 7680 513 7694 563
rect 7718 563 7812 577
rect 7718 547 7732 563
rect 7748 547 7782 555
rect 7748 513 7762 547
rect 7782 513 7790 547
rect 7798 513 7812 563
rect 7836 563 7930 577
rect 7836 547 7850 563
rect 7866 547 7900 555
rect 7866 513 7880 547
rect 7900 513 7908 547
rect 7916 513 7930 563
rect 6184 439 6198 469
rect 6214 439 6248 447
rect 6214 419 6228 439
rect 6248 419 6256 439
rect 6214 405 6256 419
rect 6264 405 6278 469
rect 6302 439 6316 469
rect 6332 439 6366 447
rect 6332 419 6346 439
rect 6366 419 6374 439
rect 6332 405 6374 419
rect 6382 405 6396 469
rect 6420 439 6434 469
rect 6450 439 6484 447
rect 6450 419 6464 439
rect 6484 419 6492 439
rect 6450 405 6492 419
rect 6500 405 6514 469
rect 6538 439 6552 469
rect 6568 439 6602 447
rect 6568 419 6582 439
rect 6602 419 6610 439
rect 6568 405 6610 419
rect 6618 405 6632 469
rect 6656 439 6670 469
rect 6686 439 6720 447
rect 6686 419 6700 439
rect 6720 419 6728 439
rect 6686 405 6728 419
rect 6736 405 6750 469
rect 6774 439 6788 469
rect 6804 439 6838 447
rect 6804 419 6818 439
rect 6838 419 6846 439
rect 6804 405 6846 419
rect 6854 405 6868 469
rect 6892 439 6906 469
rect 6922 439 6956 447
rect 6922 419 6936 439
rect 6956 419 6964 439
rect 6922 405 6964 419
rect 6972 405 6986 469
rect 7010 439 7024 469
rect 7040 439 7074 447
rect 7040 419 7054 439
rect 7074 419 7082 439
rect 7040 405 7082 419
rect 7090 405 7104 469
rect 7128 439 7142 469
rect 7158 439 7192 447
rect 7158 419 7172 439
rect 7192 419 7200 439
rect 7158 405 7200 419
rect 7208 405 7222 469
rect 7246 439 7260 469
rect 7276 439 7310 447
rect 7276 419 7290 439
rect 7310 419 7318 439
rect 7276 405 7318 419
rect 7326 405 7340 469
rect 7364 439 7378 469
rect 7394 439 7428 447
rect 7394 419 7408 439
rect 7428 419 7436 439
rect 7394 405 7436 419
rect 7444 405 7458 469
rect 7482 439 7496 469
rect 7512 439 7546 447
rect 7512 419 7526 439
rect 7546 419 7554 439
rect 7512 405 7554 419
rect 7562 405 7576 469
rect 7600 439 7614 469
rect 7630 439 7664 447
rect 7630 419 7644 439
rect 7664 419 7672 439
rect 7630 405 7672 419
rect 7680 405 7694 469
rect 7718 439 7732 469
rect 7748 439 7782 447
rect 7748 419 7762 439
rect 7782 419 7790 439
rect 7748 405 7790 419
rect 7798 405 7812 469
rect 7836 439 7850 469
rect 7866 439 7900 447
rect 7866 419 7880 439
rect 7900 419 7908 439
rect 7866 405 7908 419
rect 7916 405 7930 469
rect 4629 355 4645 371
rect 4647 355 4663 371
rect 4747 355 4763 371
rect 4765 355 4781 371
rect 4865 355 4881 371
rect 4883 355 4899 371
rect 4983 355 4999 371
rect 5001 355 5017 371
rect 6155 355 6171 371
rect 6173 355 6189 371
rect 6273 355 6289 371
rect 6291 355 6307 371
rect 6391 355 6407 371
rect 6409 355 6425 371
rect 6509 355 6525 371
rect 6527 355 6543 371
rect 6627 355 6643 371
rect 6645 355 6661 371
rect 6745 355 6761 371
rect 6763 355 6779 371
rect 6863 355 6879 371
rect 6881 355 6897 371
rect 6981 355 6997 371
rect 6999 355 7015 371
rect 7099 355 7115 371
rect 7117 355 7133 371
rect 7217 355 7233 371
rect 7235 355 7251 371
rect 7335 355 7351 371
rect 7353 355 7369 371
rect 7453 355 7469 371
rect 7471 355 7487 371
rect 7571 355 7587 371
rect 7589 355 7605 371
rect 7689 355 7705 371
rect 7707 355 7723 371
rect 7807 355 7823 371
rect 7825 355 7841 371
rect 7925 355 7941 371
rect 7943 355 7959 371
rect 4613 347 4679 355
rect 4613 339 4637 347
rect 4629 0 4637 339
rect 4655 339 4679 347
rect 4731 347 4797 355
rect 4731 339 4755 347
rect 4655 0 4663 339
rect 4747 0 4755 339
rect 4773 339 4797 347
rect 4849 347 4915 355
rect 4849 339 4873 347
rect 4773 0 4781 339
rect 4865 0 4873 339
rect 4891 339 4915 347
rect 4967 347 5033 355
rect 4967 339 4991 347
rect 4891 0 4899 339
rect 4983 0 4991 339
rect 5009 339 5033 347
rect 6139 347 6205 355
rect 6139 339 6163 347
rect 5009 0 5017 339
rect 6155 0 6163 339
rect 6181 339 6205 347
rect 6257 347 6323 355
rect 6257 339 6281 347
rect 6181 0 6189 339
rect 6273 0 6281 339
rect 6299 339 6323 347
rect 6375 347 6441 355
rect 6375 339 6399 347
rect 6299 0 6307 339
rect 6391 0 6399 339
rect 6417 339 6441 347
rect 6493 347 6559 355
rect 6493 339 6517 347
rect 6417 0 6425 339
rect 6509 0 6517 339
rect 6535 339 6559 347
rect 6611 347 6677 355
rect 6611 339 6635 347
rect 6535 0 6543 339
rect 6627 0 6635 339
rect 6653 339 6677 347
rect 6729 347 6795 355
rect 6729 339 6753 347
rect 6653 0 6661 339
rect 6745 0 6753 339
rect 6771 339 6795 347
rect 6847 347 6913 355
rect 6847 339 6871 347
rect 6771 0 6779 339
rect 6863 0 6871 339
rect 6889 339 6913 347
rect 6965 347 7031 355
rect 6965 339 6989 347
rect 6889 0 6897 339
rect 6981 0 6989 339
rect 7007 339 7031 347
rect 7083 347 7149 355
rect 7083 339 7107 347
rect 7007 0 7015 339
rect 7099 0 7107 339
rect 7125 339 7149 347
rect 7201 347 7267 355
rect 7201 339 7225 347
rect 7125 0 7133 339
rect 7217 0 7225 339
rect 7243 339 7267 347
rect 7319 347 7385 355
rect 7319 339 7343 347
rect 7243 0 7251 339
rect 7335 0 7343 339
rect 7361 339 7385 347
rect 7437 347 7503 355
rect 7437 339 7461 347
rect 7361 0 7369 339
rect 7453 0 7461 339
rect 7479 339 7503 347
rect 7555 347 7621 355
rect 7555 339 7579 347
rect 7479 0 7487 339
rect 7571 0 7579 339
rect 7597 339 7621 347
rect 7673 347 7739 355
rect 7673 339 7697 347
rect 7597 0 7605 339
rect 7689 0 7697 339
rect 7715 339 7739 347
rect 7791 347 7857 355
rect 7791 339 7815 347
rect 7715 0 7723 339
rect 7807 0 7815 339
rect 7833 339 7857 347
rect 7909 347 7975 355
rect 7909 339 7933 347
rect 7833 0 7841 339
rect 7925 0 7933 339
rect 7951 339 7975 347
rect 7951 0 7959 339
rect 11999 313 12007 1157
rect 11983 305 12007 313
rect 12025 1157 12049 1165
rect 12131 1165 12197 1173
rect 12131 1157 12155 1165
rect 12025 313 12033 1157
rect 12147 313 12155 1157
rect 12025 305 12049 313
rect 11983 297 12049 305
rect 12131 305 12155 313
rect 12173 1157 12197 1165
rect 12279 1165 12345 1173
rect 12279 1157 12303 1165
rect 12173 313 12181 1157
rect 12295 313 12303 1157
rect 12173 305 12197 313
rect 12131 297 12197 305
rect 12279 305 12303 313
rect 12321 1157 12345 1165
rect 12427 1165 12493 1173
rect 12427 1157 12451 1165
rect 12321 313 12329 1157
rect 12443 313 12451 1157
rect 12321 305 12345 313
rect 12279 297 12345 305
rect 12427 305 12451 313
rect 12469 1157 12493 1165
rect 12575 1165 12641 1173
rect 12575 1157 12599 1165
rect 12469 313 12477 1157
rect 12591 313 12599 1157
rect 12469 305 12493 313
rect 12427 297 12493 305
rect 12575 305 12599 313
rect 12617 1157 12641 1165
rect 12723 1165 12789 1173
rect 12723 1157 12747 1165
rect 12617 313 12625 1157
rect 12739 313 12747 1157
rect 12617 305 12641 313
rect 12575 297 12641 305
rect 12723 305 12747 313
rect 12765 1157 12789 1165
rect 12871 1165 12937 1173
rect 12871 1157 12895 1165
rect 12765 313 12773 1157
rect 12887 313 12895 1157
rect 12765 305 12789 313
rect 12723 297 12789 305
rect 12871 305 12895 313
rect 12913 1157 12937 1165
rect 13019 1165 13085 1173
rect 13019 1157 13043 1165
rect 12913 313 12921 1157
rect 13035 313 13043 1157
rect 12913 305 12937 313
rect 12871 297 12937 305
rect 13019 305 13043 313
rect 13061 1157 13085 1165
rect 13167 1165 13233 1173
rect 13167 1157 13191 1165
rect 13061 313 13069 1157
rect 13183 313 13191 1157
rect 13061 305 13085 313
rect 13019 297 13085 305
rect 13167 305 13191 313
rect 13209 1157 13233 1165
rect 13315 1165 13381 1173
rect 13315 1157 13339 1165
rect 13209 313 13217 1157
rect 13331 313 13339 1157
rect 13209 305 13233 313
rect 13167 297 13233 305
rect 13315 305 13339 313
rect 13357 1157 13381 1165
rect 13463 1165 13529 1173
rect 13463 1157 13487 1165
rect 13357 313 13365 1157
rect 13479 313 13487 1157
rect 13357 305 13381 313
rect 13315 297 13381 305
rect 13463 305 13487 313
rect 13505 1157 13529 1165
rect 13611 1165 13677 1173
rect 13611 1157 13635 1165
rect 13505 313 13513 1157
rect 13627 313 13635 1157
rect 13505 305 13529 313
rect 13463 297 13529 305
rect 13611 305 13635 313
rect 13653 1157 13677 1165
rect 13759 1165 13825 1173
rect 13759 1157 13783 1165
rect 13653 313 13661 1157
rect 13775 313 13783 1157
rect 13653 305 13677 313
rect 13611 297 13677 305
rect 13759 305 13783 313
rect 13801 1157 13825 1165
rect 13907 1165 13973 1173
rect 13907 1157 13931 1165
rect 13801 313 13809 1157
rect 13923 313 13931 1157
rect 13801 305 13825 313
rect 13759 297 13825 305
rect 13907 305 13931 313
rect 13949 1157 13973 1165
rect 14055 1165 14121 1173
rect 14055 1157 14079 1165
rect 13949 313 13957 1157
rect 14071 313 14079 1157
rect 13949 305 13973 313
rect 13907 297 13973 305
rect 14055 305 14079 313
rect 14097 1157 14121 1165
rect 14203 1165 14269 1173
rect 14203 1157 14227 1165
rect 14097 313 14105 1157
rect 14219 313 14227 1157
rect 14097 305 14121 313
rect 14055 297 14121 305
rect 14203 305 14227 313
rect 14245 1157 14269 1165
rect 14351 1165 14417 1173
rect 14351 1157 14375 1165
rect 14245 313 14253 1157
rect 14367 313 14375 1157
rect 14245 305 14269 313
rect 14203 297 14269 305
rect 14351 305 14375 313
rect 14393 1157 14417 1165
rect 14499 1165 14565 1173
rect 14499 1157 14523 1165
rect 14393 313 14401 1157
rect 14515 313 14523 1157
rect 14393 305 14417 313
rect 14351 297 14417 305
rect 14499 305 14523 313
rect 14541 1157 14565 1165
rect 14647 1165 14713 1173
rect 14647 1157 14671 1165
rect 14541 313 14549 1157
rect 14663 313 14671 1157
rect 14541 305 14565 313
rect 14499 297 14565 305
rect 14647 305 14671 313
rect 14689 1157 14713 1165
rect 14795 1165 14861 1173
rect 14795 1157 14819 1165
rect 14689 313 14697 1157
rect 14811 313 14819 1157
rect 14689 305 14713 313
rect 14647 297 14713 305
rect 14795 305 14819 313
rect 14837 1157 14861 1165
rect 14943 1165 15009 1173
rect 14943 1157 14967 1165
rect 14837 313 14845 1157
rect 14959 313 14967 1157
rect 14837 305 14861 313
rect 14795 297 14861 305
rect 14943 305 14967 313
rect 14985 1157 15009 1165
rect 15091 1165 15157 1173
rect 15091 1157 15115 1165
rect 14985 313 14993 1157
rect 15107 313 15115 1157
rect 14985 305 15009 313
rect 14943 297 15009 305
rect 15091 305 15115 313
rect 15133 1157 15157 1165
rect 15239 1165 15305 1173
rect 15239 1157 15263 1165
rect 15133 313 15141 1157
rect 15255 313 15263 1157
rect 15133 305 15157 313
rect 15091 297 15157 305
rect 15239 305 15263 313
rect 15281 1157 15305 1165
rect 15387 1165 15453 1173
rect 15387 1157 15411 1165
rect 15281 313 15289 1157
rect 15403 313 15411 1157
rect 15281 305 15305 313
rect 15239 297 15305 305
rect 15387 305 15411 313
rect 15429 1157 15453 1165
rect 15535 1165 15601 1173
rect 15535 1157 15559 1165
rect 15429 313 15437 1157
rect 15551 313 15559 1157
rect 15429 305 15453 313
rect 15387 297 15453 305
rect 15535 305 15559 313
rect 15577 1157 15601 1165
rect 15683 1165 15749 1173
rect 15683 1157 15707 1165
rect 15577 313 15585 1157
rect 15699 313 15707 1157
rect 15577 305 15601 313
rect 15535 297 15601 305
rect 15683 305 15707 313
rect 15725 1157 15749 1165
rect 15831 1165 15897 1173
rect 15831 1157 15855 1165
rect 15725 313 15733 1157
rect 15847 313 15855 1157
rect 15725 305 15749 313
rect 15683 297 15749 305
rect 15831 305 15855 313
rect 15873 1157 15897 1165
rect 15979 1165 16045 1173
rect 15979 1157 16003 1165
rect 15873 313 15881 1157
rect 15995 313 16003 1157
rect 15873 305 15897 313
rect 15831 297 15897 305
rect 15979 305 16003 313
rect 16021 1157 16045 1165
rect 16127 1165 16193 1173
rect 16127 1157 16151 1165
rect 16021 313 16029 1157
rect 16143 313 16151 1157
rect 16021 305 16045 313
rect 15979 297 16045 305
rect 16127 305 16151 313
rect 16169 1157 16193 1165
rect 16275 1165 16341 1173
rect 16275 1157 16299 1165
rect 16169 313 16177 1157
rect 16291 313 16299 1157
rect 16169 305 16193 313
rect 16127 297 16193 305
rect 16275 305 16299 313
rect 16317 1157 16341 1165
rect 16423 1165 16489 1173
rect 16423 1157 16447 1165
rect 16317 313 16325 1157
rect 16439 313 16447 1157
rect 16317 305 16341 313
rect 16275 297 16341 305
rect 16423 305 16447 313
rect 16465 1157 16489 1165
rect 16571 1165 16637 1173
rect 16571 1157 16595 1165
rect 16465 313 16473 1157
rect 16587 313 16595 1157
rect 16465 305 16489 313
rect 16423 297 16489 305
rect 16571 305 16595 313
rect 16613 1157 16637 1165
rect 16719 1165 16785 1173
rect 16719 1157 16743 1165
rect 16613 313 16621 1157
rect 16735 313 16743 1157
rect 16613 305 16637 313
rect 16571 297 16637 305
rect 16719 305 16743 313
rect 16761 1157 16785 1165
rect 16867 1165 16933 1173
rect 16867 1157 16891 1165
rect 16761 313 16769 1157
rect 16883 313 16891 1157
rect 16761 305 16785 313
rect 16719 297 16785 305
rect 16867 305 16891 313
rect 16909 1157 16933 1165
rect 17015 1165 17081 1173
rect 17015 1157 17039 1165
rect 16909 313 16917 1157
rect 17031 313 17039 1157
rect 16909 305 16933 313
rect 16867 297 16933 305
rect 17015 305 17039 313
rect 17057 1157 17081 1165
rect 17163 1165 17229 1173
rect 17163 1157 17187 1165
rect 17057 313 17065 1157
rect 17179 313 17187 1157
rect 17057 305 17081 313
rect 17015 297 17081 305
rect 17163 305 17187 313
rect 17205 1157 17229 1165
rect 17311 1165 17377 1173
rect 17311 1157 17335 1165
rect 17205 313 17213 1157
rect 17327 313 17335 1157
rect 17205 305 17229 313
rect 17163 297 17229 305
rect 17311 305 17335 313
rect 17353 1157 17377 1165
rect 17459 1165 17525 1173
rect 17459 1157 17483 1165
rect 17353 313 17361 1157
rect 17475 313 17483 1157
rect 17353 305 17377 313
rect 17311 297 17377 305
rect 17459 305 17483 313
rect 17501 1157 17525 1165
rect 17607 1165 17673 1173
rect 17607 1157 17631 1165
rect 17501 313 17509 1157
rect 17623 313 17631 1157
rect 17501 305 17525 313
rect 17459 297 17525 305
rect 17607 305 17631 313
rect 17649 1157 17673 1165
rect 17755 1165 17821 1173
rect 17755 1157 17779 1165
rect 17649 313 17657 1157
rect 17771 313 17779 1157
rect 17649 305 17673 313
rect 17607 297 17673 305
rect 17755 305 17779 313
rect 17797 1157 17821 1165
rect 17903 1165 17969 1173
rect 17903 1157 17927 1165
rect 17797 313 17805 1157
rect 17919 313 17927 1157
rect 17797 305 17821 313
rect 17755 297 17821 305
rect 17903 305 17927 313
rect 17945 1157 17969 1165
rect 18051 1165 18117 1173
rect 18051 1157 18075 1165
rect 17945 313 17953 1157
rect 18067 313 18075 1157
rect 17945 305 17969 313
rect 17903 297 17969 305
rect 18051 305 18075 313
rect 18093 1157 18117 1165
rect 18199 1165 18265 1173
rect 18199 1157 18223 1165
rect 18093 313 18101 1157
rect 18215 313 18223 1157
rect 18093 305 18117 313
rect 18051 297 18117 305
rect 18199 305 18223 313
rect 18241 1157 18265 1165
rect 18347 1165 18413 1173
rect 18347 1157 18371 1165
rect 18241 313 18249 1157
rect 18363 313 18371 1157
rect 18241 305 18265 313
rect 18199 297 18265 305
rect 18347 305 18371 313
rect 18389 1157 18413 1165
rect 18495 1165 18561 1173
rect 18495 1157 18519 1165
rect 18389 313 18397 1157
rect 18511 313 18519 1157
rect 18389 305 18413 313
rect 18347 297 18413 305
rect 18495 305 18519 313
rect 18537 1157 18561 1165
rect 18643 1165 18709 1173
rect 18643 1157 18667 1165
rect 18537 313 18545 1157
rect 18659 313 18667 1157
rect 18537 305 18561 313
rect 18495 297 18561 305
rect 18643 305 18667 313
rect 18685 1157 18709 1165
rect 18791 1165 18857 1173
rect 18791 1157 18815 1165
rect 18685 313 18693 1157
rect 18807 313 18815 1157
rect 18685 305 18709 313
rect 18643 297 18709 305
rect 18791 305 18815 313
rect 18833 1157 18857 1165
rect 18939 1165 19005 1173
rect 18939 1157 18963 1165
rect 18833 313 18841 1157
rect 18955 313 18963 1157
rect 18833 305 18857 313
rect 18791 297 18857 305
rect 18939 305 18963 313
rect 18981 1157 19005 1165
rect 19087 1165 19153 1173
rect 19087 1157 19111 1165
rect 18981 313 18989 1157
rect 19103 313 19111 1157
rect 18981 305 19005 313
rect 18939 297 19005 305
rect 19087 305 19111 313
rect 19129 1157 19153 1165
rect 19235 1165 19301 1173
rect 19235 1157 19259 1165
rect 19129 313 19137 1157
rect 19251 313 19259 1157
rect 19129 305 19153 313
rect 19087 297 19153 305
rect 19235 305 19259 313
rect 19277 1157 19301 1165
rect 19383 1165 19449 1173
rect 19383 1157 19407 1165
rect 19277 313 19285 1157
rect 19399 313 19407 1157
rect 19277 305 19301 313
rect 19235 297 19301 305
rect 19383 305 19407 313
rect 19425 1157 19449 1165
rect 19531 1165 19597 1173
rect 19531 1157 19555 1165
rect 19425 313 19433 1157
rect 19547 313 19555 1157
rect 19425 305 19449 313
rect 19383 297 19449 305
rect 19531 305 19555 313
rect 19573 1157 19597 1165
rect 19679 1165 19745 1173
rect 19679 1157 19703 1165
rect 19573 313 19581 1157
rect 19695 313 19703 1157
rect 19573 305 19597 313
rect 19531 297 19597 305
rect 19679 305 19703 313
rect 19721 1157 19745 1165
rect 19827 1165 19893 1173
rect 19827 1157 19851 1165
rect 19721 313 19729 1157
rect 19843 313 19851 1157
rect 19721 305 19745 313
rect 19679 297 19745 305
rect 19827 305 19851 313
rect 19869 1157 19893 1165
rect 19975 1165 20041 1173
rect 19975 1157 19999 1165
rect 19869 313 19877 1157
rect 19991 313 19999 1157
rect 19869 305 19893 313
rect 19827 297 19893 305
rect 19975 305 19999 313
rect 20017 1157 20041 1165
rect 20123 1165 20160 1173
rect 20123 1157 20147 1165
rect 20017 313 20025 1157
rect 20139 313 20147 1157
rect 20017 305 20041 313
rect 19975 297 20041 305
rect 20123 305 20147 313
rect 20123 297 20160 305
rect 11999 281 12015 297
rect 12017 281 12033 297
rect 12147 281 12163 297
rect 12165 281 12181 297
rect 12295 281 12311 297
rect 12313 281 12329 297
rect 12443 281 12459 297
rect 12461 281 12477 297
rect 12591 281 12607 297
rect 12609 281 12625 297
rect 12739 281 12755 297
rect 12757 281 12773 297
rect 12887 281 12903 297
rect 12905 281 12921 297
rect 13035 281 13051 297
rect 13053 281 13069 297
rect 13183 281 13199 297
rect 13201 281 13217 297
rect 13331 281 13347 297
rect 13349 281 13365 297
rect 13479 281 13495 297
rect 13497 281 13513 297
rect 13627 281 13643 297
rect 13645 281 13661 297
rect 13775 281 13791 297
rect 13793 281 13809 297
rect 13923 281 13939 297
rect 13941 281 13957 297
rect 14071 281 14087 297
rect 14089 281 14105 297
rect 14219 281 14235 297
rect 14237 281 14253 297
rect 14367 281 14383 297
rect 14385 281 14401 297
rect 14515 281 14531 297
rect 14533 281 14549 297
rect 14663 281 14679 297
rect 14681 281 14697 297
rect 14811 281 14827 297
rect 14829 281 14845 297
rect 14959 281 14975 297
rect 14977 281 14993 297
rect 15107 281 15123 297
rect 15125 281 15141 297
rect 15255 281 15271 297
rect 15273 281 15289 297
rect 15403 281 15419 297
rect 15421 281 15437 297
rect 15551 281 15567 297
rect 15569 281 15585 297
rect 15699 281 15715 297
rect 15717 281 15733 297
rect 15847 281 15863 297
rect 15865 281 15881 297
rect 15995 281 16011 297
rect 16013 281 16029 297
rect 16143 281 16159 297
rect 16161 281 16177 297
rect 16291 281 16307 297
rect 16309 281 16325 297
rect 16439 281 16455 297
rect 16457 281 16473 297
rect 16587 281 16603 297
rect 16605 281 16621 297
rect 16735 281 16751 297
rect 16753 281 16769 297
rect 16883 281 16899 297
rect 16901 281 16917 297
rect 17031 281 17047 297
rect 17049 281 17065 297
rect 17179 281 17195 297
rect 17197 281 17213 297
rect 17327 281 17343 297
rect 17345 281 17361 297
rect 17475 281 17491 297
rect 17493 281 17509 297
rect 17623 281 17639 297
rect 17641 281 17657 297
rect 17771 281 17787 297
rect 17789 281 17805 297
rect 17919 281 17935 297
rect 17937 281 17953 297
rect 18067 281 18083 297
rect 18085 281 18101 297
rect 18215 281 18231 297
rect 18233 281 18249 297
rect 18363 281 18379 297
rect 18381 281 18397 297
rect 18511 281 18527 297
rect 18529 281 18545 297
rect 18659 281 18675 297
rect 18677 281 18693 297
rect 18807 281 18823 297
rect 18825 281 18841 297
rect 18955 281 18971 297
rect 18973 281 18989 297
rect 19103 281 19119 297
rect 19121 281 19137 297
rect 19251 281 19267 297
rect 19269 281 19285 297
rect 19399 281 19415 297
rect 19417 281 19433 297
rect 19547 281 19563 297
rect 19565 281 19581 297
rect 19695 281 19711 297
rect 19713 281 19729 297
rect 19843 281 19859 297
rect 19861 281 19877 297
rect 19991 281 20007 297
rect 20009 281 20025 297
rect 20139 281 20155 297
rect 20157 281 20160 297
rect 12919 263 13037 277
rect 12919 247 12933 263
rect 12949 247 13007 255
rect 12949 213 12963 247
rect 13023 213 13037 263
rect 13067 263 13185 277
rect 13067 247 13081 263
rect 13097 247 13155 255
rect 13097 213 13111 247
rect 13171 213 13185 263
rect 13215 263 13333 277
rect 13215 247 13229 263
rect 13245 247 13303 255
rect 13245 213 13259 247
rect 13319 213 13333 263
rect 13363 263 13481 277
rect 13363 247 13377 263
rect 13393 247 13451 255
rect 13393 213 13407 247
rect 13467 213 13481 263
rect 13511 263 13629 277
rect 13511 247 13525 263
rect 13541 247 13599 255
rect 13541 213 13555 247
rect 13615 213 13629 263
rect 13659 263 13777 277
rect 13659 247 13673 263
rect 13689 247 13747 255
rect 13689 213 13703 247
rect 13763 213 13777 263
rect 16767 263 16885 277
rect 16767 247 16781 263
rect 16797 247 16855 255
rect 16797 213 16811 247
rect 16871 213 16885 263
rect 16915 263 17033 277
rect 16915 247 16929 263
rect 16945 247 17003 255
rect 16945 213 16959 247
rect 17019 213 17033 263
rect 17063 263 17181 277
rect 17063 247 17077 263
rect 17093 247 17151 255
rect 17093 213 17107 247
rect 17167 213 17181 263
rect 17211 263 17329 277
rect 17211 247 17225 263
rect 17241 247 17299 255
rect 17241 213 17255 247
rect 17315 213 17329 263
rect 17359 263 17477 277
rect 17359 247 17373 263
rect 17389 247 17447 255
rect 17389 213 17403 247
rect 17463 213 17477 263
rect 18099 263 18217 277
rect 18099 247 18113 263
rect 18129 247 18187 255
rect 18129 213 18143 247
rect 18203 213 18217 263
rect 18247 263 18365 277
rect 18247 247 18261 263
rect 18277 247 18335 255
rect 18277 213 18291 247
rect 18351 213 18365 263
rect 18395 263 18513 277
rect 18395 247 18409 263
rect 18425 247 18483 255
rect 18425 213 18439 247
rect 18499 213 18513 263
rect 18543 263 18661 277
rect 18543 247 18557 263
rect 18573 247 18631 255
rect 18573 213 18587 247
rect 18647 213 18661 263
rect 18691 263 18809 277
rect 18691 247 18705 263
rect 18721 247 18779 255
rect 18721 213 18735 247
rect 18795 213 18809 263
rect 18839 263 18957 277
rect 18839 247 18853 263
rect 18869 247 18927 255
rect 18869 213 18883 247
rect 18943 213 18957 263
rect 18987 263 19105 277
rect 18987 247 19001 263
rect 19017 247 19075 255
rect 19017 213 19031 247
rect 19091 213 19105 263
rect 19135 263 19253 277
rect 19135 247 19149 263
rect 19165 247 19223 255
rect 19165 213 19179 247
rect 19239 213 19253 263
rect 19283 263 19401 277
rect 19283 247 19297 263
rect 19313 247 19371 255
rect 19313 213 19327 247
rect 19387 213 19401 263
rect 19431 263 19549 277
rect 19431 247 19445 263
rect 19461 247 19519 255
rect 19461 213 19475 247
rect 19535 213 19549 263
rect 19579 263 19697 277
rect 19579 247 19593 263
rect 19609 247 19667 255
rect 19609 213 19623 247
rect 19683 213 19697 263
rect 19727 263 19845 277
rect 19727 247 19741 263
rect 19757 247 19815 255
rect 19757 213 19771 247
rect 19831 213 19845 263
rect 19875 263 19993 277
rect 19875 247 19889 263
rect 19905 247 19963 255
rect 19905 213 19919 247
rect 19979 213 19993 263
rect 20023 263 20141 277
rect 20023 247 20037 263
rect 20053 247 20111 255
rect 20053 213 20067 247
rect 20127 213 20141 263
rect 12919 139 12933 169
rect 12949 139 13007 147
rect 12949 119 12963 139
rect 12949 105 13007 119
rect 13023 105 13037 169
rect 13067 139 13081 169
rect 13097 139 13155 147
rect 13097 119 13111 139
rect 13097 105 13155 119
rect 13171 105 13185 169
rect 13215 139 13229 169
rect 13245 139 13303 147
rect 13245 119 13259 139
rect 13245 105 13303 119
rect 13319 105 13333 169
rect 13363 139 13377 169
rect 13393 139 13451 147
rect 13393 119 13407 139
rect 13393 105 13451 119
rect 13467 105 13481 169
rect 13511 139 13525 169
rect 13541 139 13599 147
rect 13541 119 13555 139
rect 13541 105 13599 119
rect 13615 105 13629 169
rect 13659 139 13673 169
rect 13689 139 13747 147
rect 13689 119 13703 139
rect 13689 105 13747 119
rect 13763 105 13777 169
rect 16767 139 16781 169
rect 16797 139 16855 147
rect 16797 119 16811 139
rect 16797 105 16855 119
rect 16871 105 16885 169
rect 16915 139 16929 169
rect 16945 139 17003 147
rect 16945 119 16959 139
rect 16945 105 17003 119
rect 17019 105 17033 169
rect 17063 139 17077 169
rect 17093 139 17151 147
rect 17093 119 17107 139
rect 17093 105 17151 119
rect 17167 105 17181 169
rect 17211 139 17225 169
rect 17241 139 17299 147
rect 17241 119 17255 139
rect 17241 105 17299 119
rect 17315 105 17329 169
rect 17359 139 17373 169
rect 17389 139 17447 147
rect 17389 119 17403 139
rect 17389 105 17447 119
rect 17463 105 17477 169
rect 18099 139 18113 169
rect 18129 139 18187 147
rect 18129 119 18143 139
rect 18129 105 18187 119
rect 18203 105 18217 169
rect 18247 139 18261 169
rect 18277 139 18335 147
rect 18277 119 18291 139
rect 18277 105 18335 119
rect 18351 105 18365 169
rect 18395 139 18409 169
rect 18425 139 18483 147
rect 18425 119 18439 139
rect 18425 105 18483 119
rect 18499 105 18513 169
rect 18543 139 18557 169
rect 18573 139 18631 147
rect 18573 119 18587 139
rect 18573 105 18631 119
rect 18647 105 18661 169
rect 18691 139 18705 169
rect 18721 139 18779 147
rect 18721 119 18735 139
rect 18721 105 18779 119
rect 18795 105 18809 169
rect 18839 139 18853 169
rect 18869 139 18927 147
rect 18869 119 18883 139
rect 18869 105 18927 119
rect 18943 105 18957 169
rect 18987 139 19001 169
rect 19017 139 19075 147
rect 19017 119 19031 139
rect 19017 105 19075 119
rect 19091 105 19105 169
rect 19135 139 19149 169
rect 19165 139 19223 147
rect 19165 119 19179 139
rect 19165 105 19223 119
rect 19239 105 19253 169
rect 19283 139 19297 169
rect 19313 139 19371 147
rect 19313 119 19327 139
rect 19313 105 19371 119
rect 19387 105 19401 169
rect 19431 139 19445 169
rect 19461 139 19519 147
rect 19461 119 19475 139
rect 19461 105 19519 119
rect 19535 105 19549 169
rect 19579 139 19593 169
rect 19609 139 19667 147
rect 19609 119 19623 139
rect 19609 105 19667 119
rect 19683 105 19697 169
rect 19727 139 19741 169
rect 19757 139 19815 147
rect 19757 119 19771 139
rect 19757 105 19815 119
rect 19831 105 19845 169
rect 19875 139 19889 169
rect 19905 139 19963 147
rect 19905 119 19919 139
rect 19905 105 19963 119
rect 19979 105 19993 169
rect 20023 139 20037 169
rect 20053 139 20111 147
rect 20053 119 20067 139
rect 20053 105 20111 119
rect 20127 105 20141 169
rect 19695 55 19711 71
rect 19713 55 19729 71
rect 19843 55 19859 71
rect 19861 55 19877 71
rect 19991 55 20007 71
rect 20009 55 20025 71
rect 20139 55 20155 71
rect 20157 55 20160 71
rect 19679 47 19745 55
rect 19679 39 19703 47
rect 19695 0 19703 39
rect 19721 39 19745 47
rect 19827 47 19893 55
rect 19827 39 19851 47
rect 19721 0 19729 39
rect 19843 0 19851 39
rect 19869 39 19893 47
rect 19975 47 20041 55
rect 19975 39 19999 47
rect 19869 0 19877 39
rect 19991 0 19999 39
rect 20017 39 20041 47
rect 20123 47 20160 55
rect 20123 39 20147 47
rect 20017 0 20025 39
rect 20139 0 20147 39
rect 2337 -467 2361 -462
rect 2395 -467 2433 -462
rect 2467 -467 2515 -462
rect 2549 -467 2587 -462
rect 2621 -467 2669 -462
rect 2703 -467 2741 -462
rect 2775 -467 2823 -462
rect 2857 -467 2895 -462
rect 2929 -467 2977 -462
rect 3011 -467 3049 -462
rect 3083 -467 3131 -462
rect 3165 -467 3203 -462
rect 3237 -467 3285 -462
rect 3319 -467 3357 -462
rect 3391 -467 3439 -462
rect 3473 -467 3511 -462
rect 3545 -467 3593 -462
rect 3627 -467 3665 -462
rect 3699 -467 3747 -462
rect 2337 -483 2377 -467
rect 2379 -483 2449 -467
rect 2451 -483 2531 -467
rect 2533 -483 2603 -467
rect 2605 -483 2685 -467
rect 2687 -483 2757 -467
rect 2759 -483 2839 -467
rect 2841 -483 2911 -467
rect 2913 -483 2993 -467
rect 2995 -483 3065 -467
rect 3067 -483 3147 -467
rect 3149 -483 3219 -467
rect 3221 -483 3301 -467
rect 3303 -483 3373 -467
rect 3375 -483 3455 -467
rect 3457 -483 3527 -467
rect 3529 -483 3609 -467
rect 3611 -483 3681 -467
rect 3683 -483 3760 -467
rect 2337 -488 3760 -483
rect 2345 -490 2411 -488
rect 2417 -490 2483 -488
rect 2499 -490 2565 -488
rect 2571 -490 2637 -488
rect 2653 -490 2719 -488
rect 2725 -490 2791 -488
rect 2807 -490 2873 -488
rect 2879 -490 2945 -488
rect 2961 -490 3027 -488
rect 3033 -490 3099 -488
rect 3115 -490 3181 -488
rect 3187 -490 3253 -488
rect 3269 -490 3335 -488
rect 3341 -490 3407 -488
rect 3423 -490 3489 -488
rect 3495 -490 3561 -488
rect 3577 -490 3643 -488
rect 3649 -490 3715 -488
rect 3731 -490 3760 -488
rect 2337 -516 3760 -490
rect 2345 -517 2411 -516
rect 2417 -517 2483 -516
rect 2499 -517 2565 -516
rect 2571 -517 2637 -516
rect 2653 -517 2719 -516
rect 2725 -517 2791 -516
rect 2807 -517 2873 -516
rect 2879 -517 2945 -516
rect 2961 -517 3027 -516
rect 3033 -517 3099 -516
rect 3115 -517 3181 -516
rect 3187 -517 3253 -516
rect 3269 -517 3335 -516
rect 3341 -517 3407 -516
rect 3423 -517 3489 -516
rect 3495 -517 3561 -516
rect 3577 -517 3643 -516
rect 3649 -517 3715 -516
rect 3731 -517 3760 -516
rect 2361 -533 2377 -517
rect 2379 -533 2395 -517
rect 2433 -533 2449 -517
rect 2451 -533 2467 -517
rect 2515 -533 2531 -517
rect 2533 -533 2549 -517
rect 2587 -533 2603 -517
rect 2605 -533 2621 -517
rect 2669 -533 2685 -517
rect 2687 -533 2703 -517
rect 2741 -533 2757 -517
rect 2759 -533 2775 -517
rect 2823 -533 2839 -517
rect 2841 -533 2857 -517
rect 2895 -533 2911 -517
rect 2913 -533 2929 -517
rect 2977 -533 2993 -517
rect 2995 -533 3011 -517
rect 3049 -533 3065 -517
rect 3067 -533 3083 -517
rect 3131 -533 3147 -517
rect 3149 -533 3165 -517
rect 3203 -533 3219 -517
rect 3221 -533 3237 -517
rect 3285 -533 3301 -517
rect 3303 -533 3319 -517
rect 3357 -533 3373 -517
rect 3375 -533 3391 -517
rect 3439 -533 3455 -517
rect 3457 -533 3473 -517
rect 3511 -533 3527 -517
rect 3529 -533 3545 -517
rect 3593 -533 3609 -517
rect 3611 -533 3627 -517
rect 3665 -533 3681 -517
rect 3683 -533 3699 -517
rect 3747 -533 3760 -517
rect 2361 -557 2377 -541
rect 2379 -557 2395 -541
rect 2433 -557 2449 -541
rect 2451 -557 2467 -541
rect 2515 -557 2531 -541
rect 2533 -557 2549 -541
rect 2587 -557 2603 -541
rect 2605 -557 2621 -541
rect 2669 -557 2685 -541
rect 2687 -557 2703 -541
rect 2741 -557 2757 -541
rect 2759 -557 2775 -541
rect 2823 -557 2839 -541
rect 2841 -557 2857 -541
rect 2895 -557 2911 -541
rect 2913 -557 2929 -541
rect 2977 -557 2993 -541
rect 2995 -557 3011 -541
rect 3049 -557 3065 -541
rect 3067 -557 3083 -541
rect 3131 -557 3147 -541
rect 3149 -557 3165 -541
rect 3203 -557 3219 -541
rect 3221 -557 3237 -541
rect 3285 -557 3301 -541
rect 3303 -557 3319 -541
rect 3357 -557 3373 -541
rect 3375 -557 3391 -541
rect 3439 -557 3455 -541
rect 3457 -557 3473 -541
rect 3511 -557 3527 -541
rect 3529 -557 3545 -541
rect 3593 -557 3609 -541
rect 3611 -557 3627 -541
rect 3665 -557 3681 -541
rect 3683 -557 3699 -541
rect 3747 -557 3760 -541
rect 2345 -573 2411 -557
rect 2417 -573 2483 -557
rect 2499 -573 2565 -557
rect 2571 -573 2637 -557
rect 2653 -573 2719 -557
rect 2725 -573 2791 -557
rect 2807 -573 2873 -557
rect 2879 -573 2945 -557
rect 2961 -573 3027 -557
rect 3033 -573 3099 -557
rect 3115 -573 3181 -557
rect 3187 -573 3253 -557
rect 3269 -573 3335 -557
rect 3341 -573 3407 -557
rect 3423 -573 3489 -557
rect 3495 -573 3561 -557
rect 3577 -573 3643 -557
rect 3649 -573 3715 -557
rect 3731 -573 3760 -557
rect 2361 -575 2395 -573
rect 2433 -575 2467 -573
rect 2515 -575 2549 -573
rect 2587 -575 2621 -573
rect 2669 -575 2703 -573
rect 2741 -575 2775 -573
rect 2823 -575 2857 -573
rect 2895 -575 2929 -573
rect 2977 -575 3011 -573
rect 3049 -575 3083 -573
rect 3131 -575 3165 -573
rect 3203 -575 3237 -573
rect 3285 -575 3319 -573
rect 3357 -575 3391 -573
rect 3439 -575 3473 -573
rect 3511 -575 3545 -573
rect 3593 -575 3627 -573
rect 3665 -575 3699 -573
rect 3747 -575 3760 -573
rect 2345 -591 2411 -575
rect 2417 -591 2483 -575
rect 2499 -591 2565 -575
rect 2571 -591 2637 -575
rect 2653 -591 2719 -575
rect 2725 -591 2791 -575
rect 2807 -591 2873 -575
rect 2879 -591 2945 -575
rect 2961 -591 3027 -575
rect 3033 -591 3099 -575
rect 3115 -591 3181 -575
rect 3187 -591 3253 -575
rect 3269 -591 3335 -575
rect 3341 -591 3407 -575
rect 3423 -591 3489 -575
rect 3495 -591 3561 -575
rect 3577 -591 3643 -575
rect 3649 -591 3715 -575
rect 3731 -591 3760 -575
rect 2361 -607 2377 -591
rect 2379 -607 2395 -591
rect 2433 -607 2449 -591
rect 2451 -607 2467 -591
rect 2515 -607 2531 -591
rect 2533 -607 2549 -591
rect 2587 -607 2603 -591
rect 2605 -607 2621 -591
rect 2669 -607 2685 -591
rect 2687 -607 2703 -591
rect 2741 -607 2757 -591
rect 2759 -607 2775 -591
rect 2823 -607 2839 -591
rect 2841 -607 2857 -591
rect 2895 -607 2911 -591
rect 2913 -607 2929 -591
rect 2977 -607 2993 -591
rect 2995 -607 3011 -591
rect 3049 -607 3065 -591
rect 3067 -607 3083 -591
rect 3131 -607 3147 -591
rect 3149 -607 3165 -591
rect 3203 -607 3219 -591
rect 3221 -607 3237 -591
rect 3285 -607 3301 -591
rect 3303 -607 3319 -591
rect 3357 -607 3373 -591
rect 3375 -607 3391 -591
rect 3439 -607 3455 -591
rect 3457 -607 3473 -591
rect 3511 -607 3527 -591
rect 3529 -607 3545 -591
rect 3593 -607 3609 -591
rect 3611 -607 3627 -591
rect 3665 -607 3681 -591
rect 3683 -607 3699 -591
rect 3747 -607 3760 -591
rect 2361 -631 2377 -615
rect 2379 -631 2395 -615
rect 2433 -631 2449 -615
rect 2451 -631 2467 -615
rect 2515 -631 2531 -615
rect 2533 -631 2549 -615
rect 2587 -631 2603 -615
rect 2605 -631 2621 -615
rect 2669 -631 2685 -615
rect 2687 -631 2703 -615
rect 2741 -631 2757 -615
rect 2759 -631 2775 -615
rect 2823 -631 2839 -615
rect 2841 -631 2857 -615
rect 2895 -631 2911 -615
rect 2913 -631 2929 -615
rect 2977 -631 2993 -615
rect 2995 -631 3011 -615
rect 3049 -631 3065 -615
rect 3067 -631 3083 -615
rect 3131 -631 3147 -615
rect 3149 -631 3165 -615
rect 3203 -631 3219 -615
rect 3221 -631 3237 -615
rect 3285 -631 3301 -615
rect 3303 -631 3319 -615
rect 3357 -631 3373 -615
rect 3375 -631 3391 -615
rect 3439 -631 3455 -615
rect 3457 -631 3473 -615
rect 3511 -631 3527 -615
rect 3529 -631 3545 -615
rect 3593 -631 3609 -615
rect 3611 -631 3627 -615
rect 3665 -631 3681 -615
rect 3683 -631 3699 -615
rect 3747 -631 3760 -615
rect 2345 -647 2411 -631
rect 2417 -647 2483 -631
rect 2499 -647 2565 -631
rect 2571 -647 2637 -631
rect 2653 -647 2719 -631
rect 2725 -647 2791 -631
rect 2807 -647 2873 -631
rect 2879 -647 2945 -631
rect 2961 -647 3027 -631
rect 3033 -647 3099 -631
rect 3115 -647 3181 -631
rect 3187 -647 3253 -631
rect 3269 -647 3335 -631
rect 3341 -647 3407 -631
rect 3423 -647 3489 -631
rect 3495 -647 3561 -631
rect 3577 -647 3643 -631
rect 3649 -647 3715 -631
rect 3731 -647 3760 -631
rect 2361 -649 2395 -647
rect 2433 -649 2467 -647
rect 2515 -649 2549 -647
rect 2587 -649 2621 -647
rect 2669 -649 2703 -647
rect 2741 -649 2775 -647
rect 2823 -649 2857 -647
rect 2895 -649 2929 -647
rect 2977 -649 3011 -647
rect 3049 -649 3083 -647
rect 3131 -649 3165 -647
rect 3203 -649 3237 -647
rect 3285 -649 3319 -647
rect 3357 -649 3391 -647
rect 3439 -649 3473 -647
rect 3511 -649 3545 -647
rect 3593 -649 3627 -647
rect 3665 -649 3699 -647
rect 3747 -649 3760 -647
rect 2345 -665 2411 -649
rect 2417 -665 2483 -649
rect 2499 -665 2565 -649
rect 2571 -665 2637 -649
rect 2653 -665 2719 -649
rect 2725 -665 2791 -649
rect 2807 -665 2873 -649
rect 2879 -665 2945 -649
rect 2961 -665 3027 -649
rect 3033 -665 3099 -649
rect 3115 -665 3181 -649
rect 3187 -665 3253 -649
rect 3269 -665 3335 -649
rect 3341 -665 3407 -649
rect 3423 -665 3489 -649
rect 3495 -665 3561 -649
rect 3577 -665 3643 -649
rect 3649 -665 3715 -649
rect 3731 -665 3760 -649
rect 2361 -681 2377 -665
rect 2379 -681 2395 -665
rect 2433 -681 2449 -665
rect 2451 -681 2467 -665
rect 2515 -681 2531 -665
rect 2533 -681 2549 -665
rect 2587 -681 2603 -665
rect 2605 -681 2621 -665
rect 2669 -681 2685 -665
rect 2687 -681 2703 -665
rect 2741 -681 2757 -665
rect 2759 -681 2775 -665
rect 2823 -681 2839 -665
rect 2841 -681 2857 -665
rect 2895 -681 2911 -665
rect 2913 -681 2929 -665
rect 2977 -681 2993 -665
rect 2995 -681 3011 -665
rect 3049 -681 3065 -665
rect 3067 -681 3083 -665
rect 3131 -681 3147 -665
rect 3149 -681 3165 -665
rect 3203 -681 3219 -665
rect 3221 -681 3237 -665
rect 3285 -681 3301 -665
rect 3303 -681 3319 -665
rect 3357 -681 3373 -665
rect 3375 -681 3391 -665
rect 3439 -681 3455 -665
rect 3457 -681 3473 -665
rect 3511 -681 3527 -665
rect 3529 -681 3545 -665
rect 3593 -681 3609 -665
rect 3611 -681 3627 -665
rect 3665 -681 3681 -665
rect 3683 -681 3699 -665
rect 3747 -681 3760 -665
rect 2361 -705 2377 -689
rect 2379 -705 2395 -689
rect 2433 -705 2449 -689
rect 2451 -705 2467 -689
rect 2515 -705 2531 -689
rect 2533 -705 2549 -689
rect 2587 -705 2603 -689
rect 2605 -705 2621 -689
rect 2669 -705 2685 -689
rect 2687 -705 2703 -689
rect 2741 -705 2757 -689
rect 2759 -705 2775 -689
rect 2823 -705 2839 -689
rect 2841 -705 2857 -689
rect 2895 -705 2911 -689
rect 2913 -705 2929 -689
rect 2977 -705 2993 -689
rect 2995 -705 3011 -689
rect 3049 -705 3065 -689
rect 3067 -705 3083 -689
rect 3131 -705 3147 -689
rect 3149 -705 3165 -689
rect 3203 -705 3219 -689
rect 3221 -705 3237 -689
rect 3285 -705 3301 -689
rect 3303 -705 3319 -689
rect 3357 -705 3373 -689
rect 3375 -705 3391 -689
rect 3439 -705 3455 -689
rect 3457 -705 3473 -689
rect 3511 -705 3527 -689
rect 3529 -705 3545 -689
rect 3593 -705 3609 -689
rect 3611 -705 3627 -689
rect 3665 -705 3681 -689
rect 3683 -705 3699 -689
rect 3747 -705 3760 -689
rect 2345 -721 2411 -705
rect 2417 -721 2483 -705
rect 2499 -721 2565 -705
rect 2571 -721 2637 -705
rect 2653 -721 2719 -705
rect 2725 -721 2791 -705
rect 2807 -721 2873 -705
rect 2879 -721 2945 -705
rect 2961 -721 3027 -705
rect 3033 -721 3099 -705
rect 3115 -721 3181 -705
rect 3187 -721 3253 -705
rect 3269 -721 3335 -705
rect 3341 -721 3407 -705
rect 3423 -721 3489 -705
rect 3495 -721 3561 -705
rect 3577 -721 3643 -705
rect 3649 -721 3715 -705
rect 3731 -721 3760 -705
rect 2361 -723 2395 -721
rect 2433 -723 2467 -721
rect 2515 -723 2549 -721
rect 2587 -723 2621 -721
rect 2669 -723 2703 -721
rect 2741 -723 2775 -721
rect 2823 -723 2857 -721
rect 2895 -723 2929 -721
rect 2977 -723 3011 -721
rect 3049 -723 3083 -721
rect 3131 -723 3165 -721
rect 3203 -723 3237 -721
rect 3285 -723 3319 -721
rect 3357 -723 3391 -721
rect 3439 -723 3473 -721
rect 3511 -723 3545 -721
rect 3593 -723 3627 -721
rect 3665 -723 3699 -721
rect 3747 -723 3760 -721
rect 2345 -739 2411 -723
rect 2417 -739 2483 -723
rect 2499 -739 2565 -723
rect 2571 -739 2637 -723
rect 2653 -739 2719 -723
rect 2725 -739 2791 -723
rect 2807 -739 2873 -723
rect 2879 -739 2945 -723
rect 2961 -739 3027 -723
rect 3033 -739 3099 -723
rect 3115 -739 3181 -723
rect 3187 -739 3253 -723
rect 3269 -739 3335 -723
rect 3341 -739 3407 -723
rect 3423 -739 3489 -723
rect 3495 -739 3561 -723
rect 3577 -739 3643 -723
rect 3649 -739 3715 -723
rect 3731 -739 3760 -723
rect 2361 -755 2377 -739
rect 2379 -755 2395 -739
rect 2433 -755 2449 -739
rect 2451 -755 2467 -739
rect 2515 -755 2531 -739
rect 2533 -755 2549 -739
rect 2587 -755 2603 -739
rect 2605 -755 2621 -739
rect 2669 -755 2685 -739
rect 2687 -755 2703 -739
rect 2741 -755 2757 -739
rect 2759 -755 2775 -739
rect 2823 -755 2839 -739
rect 2841 -755 2857 -739
rect 2895 -755 2911 -739
rect 2913 -755 2929 -739
rect 2977 -755 2993 -739
rect 2995 -755 3011 -739
rect 3049 -755 3065 -739
rect 3067 -755 3083 -739
rect 3131 -755 3147 -739
rect 3149 -755 3165 -739
rect 3203 -755 3219 -739
rect 3221 -755 3237 -739
rect 3285 -755 3301 -739
rect 3303 -755 3319 -739
rect 3357 -755 3373 -739
rect 3375 -755 3391 -739
rect 3439 -755 3455 -739
rect 3457 -755 3473 -739
rect 3511 -755 3527 -739
rect 3529 -755 3545 -739
rect 3593 -755 3609 -739
rect 3611 -755 3627 -739
rect 3665 -755 3681 -739
rect 3683 -755 3699 -739
rect 3747 -755 3760 -739
rect 2361 -779 2377 -763
rect 2379 -779 2395 -763
rect 2433 -779 2449 -763
rect 2451 -779 2467 -763
rect 2515 -779 2531 -763
rect 2533 -779 2549 -763
rect 2587 -779 2603 -763
rect 2605 -779 2621 -763
rect 2669 -779 2685 -763
rect 2687 -779 2703 -763
rect 2741 -779 2757 -763
rect 2759 -779 2775 -763
rect 2823 -779 2839 -763
rect 2841 -779 2857 -763
rect 2895 -779 2911 -763
rect 2913 -779 2929 -763
rect 2977 -779 2993 -763
rect 2995 -779 3011 -763
rect 3049 -779 3065 -763
rect 3067 -779 3083 -763
rect 3131 -779 3147 -763
rect 3149 -779 3165 -763
rect 3203 -779 3219 -763
rect 3221 -779 3237 -763
rect 3285 -779 3301 -763
rect 3303 -779 3319 -763
rect 3357 -779 3373 -763
rect 3375 -779 3391 -763
rect 3439 -779 3455 -763
rect 3457 -779 3473 -763
rect 3511 -779 3527 -763
rect 3529 -779 3545 -763
rect 3593 -779 3609 -763
rect 3611 -779 3627 -763
rect 3665 -779 3681 -763
rect 3683 -779 3699 -763
rect 3747 -779 3760 -763
rect 2345 -795 2411 -779
rect 2417 -795 2483 -779
rect 2499 -795 2565 -779
rect 2571 -795 2637 -779
rect 2653 -795 2719 -779
rect 2725 -795 2791 -779
rect 2807 -795 2873 -779
rect 2879 -795 2945 -779
rect 2961 -795 3027 -779
rect 3033 -795 3099 -779
rect 3115 -795 3181 -779
rect 3187 -795 3253 -779
rect 3269 -795 3335 -779
rect 3341 -795 3407 -779
rect 3423 -795 3489 -779
rect 3495 -795 3561 -779
rect 3577 -795 3643 -779
rect 3649 -795 3715 -779
rect 3731 -795 3760 -779
rect 2361 -797 2395 -795
rect 2433 -797 2467 -795
rect 2515 -797 2549 -795
rect 2587 -797 2621 -795
rect 2669 -797 2703 -795
rect 2741 -797 2775 -795
rect 2823 -797 2857 -795
rect 2895 -797 2929 -795
rect 2977 -797 3011 -795
rect 3049 -797 3083 -795
rect 3131 -797 3165 -795
rect 3203 -797 3237 -795
rect 3285 -797 3319 -795
rect 3357 -797 3391 -795
rect 3439 -797 3473 -795
rect 3511 -797 3545 -795
rect 3593 -797 3627 -795
rect 3665 -797 3699 -795
rect 3747 -797 3760 -795
rect 2345 -813 2411 -797
rect 2417 -813 2483 -797
rect 2499 -813 2565 -797
rect 2571 -813 2637 -797
rect 2653 -813 2719 -797
rect 2725 -813 2791 -797
rect 2807 -813 2873 -797
rect 2879 -813 2945 -797
rect 2961 -813 3027 -797
rect 3033 -813 3099 -797
rect 3115 -813 3181 -797
rect 3187 -813 3253 -797
rect 3269 -813 3335 -797
rect 3341 -813 3407 -797
rect 3423 -813 3489 -797
rect 3495 -813 3561 -797
rect 3577 -813 3643 -797
rect 3649 -813 3715 -797
rect 3731 -813 3760 -797
rect 2361 -829 2377 -813
rect 2379 -829 2395 -813
rect 2433 -829 2449 -813
rect 2451 -829 2467 -813
rect 2515 -829 2531 -813
rect 2533 -829 2549 -813
rect 2587 -829 2603 -813
rect 2605 -829 2621 -813
rect 2669 -829 2685 -813
rect 2687 -829 2703 -813
rect 2741 -829 2757 -813
rect 2759 -829 2775 -813
rect 2823 -829 2839 -813
rect 2841 -829 2857 -813
rect 2895 -829 2911 -813
rect 2913 -829 2929 -813
rect 2977 -829 2993 -813
rect 2995 -829 3011 -813
rect 3049 -829 3065 -813
rect 3067 -829 3083 -813
rect 3131 -829 3147 -813
rect 3149 -829 3165 -813
rect 3203 -829 3219 -813
rect 3221 -829 3237 -813
rect 3285 -829 3301 -813
rect 3303 -829 3319 -813
rect 3357 -829 3373 -813
rect 3375 -829 3391 -813
rect 3439 -829 3455 -813
rect 3457 -829 3473 -813
rect 3511 -829 3527 -813
rect 3529 -829 3545 -813
rect 3593 -829 3609 -813
rect 3611 -829 3627 -813
rect 3665 -829 3681 -813
rect 3683 -829 3699 -813
rect 3747 -829 3760 -813
rect 2361 -853 2377 -837
rect 2379 -853 2395 -837
rect 2433 -853 2449 -837
rect 2451 -853 2467 -837
rect 2515 -853 2531 -837
rect 2533 -853 2549 -837
rect 2587 -853 2603 -837
rect 2605 -853 2621 -837
rect 2669 -853 2685 -837
rect 2687 -853 2703 -837
rect 2741 -853 2757 -837
rect 2759 -853 2775 -837
rect 2823 -853 2839 -837
rect 2841 -853 2857 -837
rect 2895 -853 2911 -837
rect 2913 -853 2929 -837
rect 2977 -853 2993 -837
rect 2995 -853 3011 -837
rect 3049 -853 3065 -837
rect 3067 -853 3083 -837
rect 3131 -853 3147 -837
rect 3149 -853 3165 -837
rect 3203 -853 3219 -837
rect 3221 -853 3237 -837
rect 3285 -853 3301 -837
rect 3303 -853 3319 -837
rect 3357 -853 3373 -837
rect 3375 -853 3391 -837
rect 3439 -853 3455 -837
rect 3457 -853 3473 -837
rect 3511 -853 3527 -837
rect 3529 -853 3545 -837
rect 3593 -853 3609 -837
rect 3611 -853 3627 -837
rect 3665 -853 3681 -837
rect 3683 -853 3699 -837
rect 3747 -853 3760 -837
rect 2345 -869 2411 -853
rect 2417 -869 2483 -853
rect 2499 -869 2565 -853
rect 2571 -869 2637 -853
rect 2653 -869 2719 -853
rect 2725 -869 2791 -853
rect 2807 -869 2873 -853
rect 2879 -869 2945 -853
rect 2961 -869 3027 -853
rect 3033 -869 3099 -853
rect 3115 -869 3181 -853
rect 3187 -869 3253 -853
rect 3269 -869 3335 -853
rect 3341 -869 3407 -853
rect 3423 -869 3489 -853
rect 3495 -869 3561 -853
rect 3577 -869 3643 -853
rect 3649 -869 3715 -853
rect 3731 -869 3760 -853
rect 2361 -871 2395 -869
rect 2433 -871 2467 -869
rect 2515 -871 2549 -869
rect 2587 -871 2621 -869
rect 2669 -871 2703 -869
rect 2741 -871 2775 -869
rect 2823 -871 2857 -869
rect 2895 -871 2929 -869
rect 2977 -871 3011 -869
rect 3049 -871 3083 -869
rect 3131 -871 3165 -869
rect 3203 -871 3237 -869
rect 3285 -871 3319 -869
rect 3357 -871 3391 -869
rect 3439 -871 3473 -869
rect 3511 -871 3545 -869
rect 3593 -871 3627 -869
rect 3665 -871 3699 -869
rect 3747 -871 3760 -869
rect 2345 -887 2411 -871
rect 2417 -887 2483 -871
rect 2499 -887 2565 -871
rect 2571 -887 2637 -871
rect 2653 -887 2719 -871
rect 2725 -887 2791 -871
rect 2807 -887 2873 -871
rect 2879 -887 2945 -871
rect 2961 -887 3027 -871
rect 3033 -887 3099 -871
rect 3115 -887 3181 -871
rect 3187 -887 3253 -871
rect 3269 -887 3335 -871
rect 3341 -887 3407 -871
rect 3423 -887 3489 -871
rect 3495 -887 3561 -871
rect 3577 -887 3643 -871
rect 3649 -887 3715 -871
rect 3731 -887 3760 -871
rect 2361 -903 2377 -887
rect 2379 -903 2395 -887
rect 2433 -903 2449 -887
rect 2451 -903 2467 -887
rect 2515 -903 2531 -887
rect 2533 -903 2549 -887
rect 2587 -903 2603 -887
rect 2605 -903 2621 -887
rect 2669 -903 2685 -887
rect 2687 -903 2703 -887
rect 2741 -903 2757 -887
rect 2759 -903 2775 -887
rect 2823 -903 2839 -887
rect 2841 -903 2857 -887
rect 2895 -903 2911 -887
rect 2913 -903 2929 -887
rect 2977 -903 2993 -887
rect 2995 -903 3011 -887
rect 3049 -903 3065 -887
rect 3067 -903 3083 -887
rect 3131 -903 3147 -887
rect 3149 -903 3165 -887
rect 3203 -903 3219 -887
rect 3221 -903 3237 -887
rect 3285 -903 3301 -887
rect 3303 -903 3319 -887
rect 3357 -903 3373 -887
rect 3375 -903 3391 -887
rect 3439 -903 3455 -887
rect 3457 -903 3473 -887
rect 3511 -903 3527 -887
rect 3529 -903 3545 -887
rect 3593 -903 3609 -887
rect 3611 -903 3627 -887
rect 3665 -903 3681 -887
rect 3683 -903 3699 -887
rect 3747 -903 3760 -887
rect 2361 -927 2377 -911
rect 2379 -927 2395 -911
rect 2433 -927 2449 -911
rect 2451 -927 2467 -911
rect 2515 -927 2531 -911
rect 2533 -927 2549 -911
rect 2587 -927 2603 -911
rect 2605 -927 2621 -911
rect 2669 -927 2685 -911
rect 2687 -927 2703 -911
rect 2741 -927 2757 -911
rect 2759 -927 2775 -911
rect 2823 -927 2839 -911
rect 2841 -927 2857 -911
rect 2895 -927 2911 -911
rect 2913 -927 2929 -911
rect 2977 -927 2993 -911
rect 2995 -927 3011 -911
rect 3049 -927 3065 -911
rect 3067 -927 3083 -911
rect 3131 -927 3147 -911
rect 3149 -927 3165 -911
rect 3203 -927 3219 -911
rect 3221 -927 3237 -911
rect 3285 -927 3301 -911
rect 3303 -927 3319 -911
rect 3357 -927 3373 -911
rect 3375 -927 3391 -911
rect 3439 -927 3455 -911
rect 3457 -927 3473 -911
rect 3511 -927 3527 -911
rect 3529 -927 3545 -911
rect 3593 -927 3609 -911
rect 3611 -927 3627 -911
rect 3665 -927 3681 -911
rect 3683 -927 3699 -911
rect 3747 -927 3760 -911
rect 2345 -943 2411 -927
rect 2417 -943 2483 -927
rect 2499 -943 2565 -927
rect 2571 -943 2637 -927
rect 2653 -943 2719 -927
rect 2725 -943 2791 -927
rect 2807 -943 2873 -927
rect 2879 -943 2945 -927
rect 2961 -943 3027 -927
rect 3033 -943 3099 -927
rect 3115 -943 3181 -927
rect 3187 -943 3253 -927
rect 3269 -943 3335 -927
rect 3341 -943 3407 -927
rect 3423 -943 3489 -927
rect 3495 -943 3561 -927
rect 3577 -943 3643 -927
rect 3649 -943 3715 -927
rect 3731 -943 3760 -927
rect 2361 -945 2395 -943
rect 2433 -945 2467 -943
rect 2515 -945 2549 -943
rect 2587 -945 2621 -943
rect 2669 -945 2703 -943
rect 2741 -945 2775 -943
rect 2823 -945 2857 -943
rect 2895 -945 2929 -943
rect 2977 -945 3011 -943
rect 3049 -945 3083 -943
rect 3131 -945 3165 -943
rect 3203 -945 3237 -943
rect 3285 -945 3319 -943
rect 3357 -945 3391 -943
rect 3439 -945 3473 -943
rect 3511 -945 3545 -943
rect 3593 -945 3627 -943
rect 3665 -945 3699 -943
rect 3747 -945 3760 -943
rect 2345 -961 2411 -945
rect 2417 -961 2483 -945
rect 2499 -961 2565 -945
rect 2571 -961 2637 -945
rect 2653 -961 2719 -945
rect 2725 -961 2791 -945
rect 2807 -961 2873 -945
rect 2879 -961 2945 -945
rect 2961 -961 3027 -945
rect 3033 -961 3099 -945
rect 3115 -961 3181 -945
rect 3187 -961 3253 -945
rect 3269 -961 3335 -945
rect 3341 -961 3407 -945
rect 3423 -961 3489 -945
rect 3495 -961 3561 -945
rect 3577 -961 3643 -945
rect 3649 -961 3715 -945
rect 3731 -961 3760 -945
rect 2361 -977 2377 -961
rect 2379 -977 2395 -961
rect 2433 -977 2449 -961
rect 2451 -977 2467 -961
rect 2515 -977 2531 -961
rect 2533 -977 2549 -961
rect 2587 -977 2603 -961
rect 2605 -977 2621 -961
rect 2669 -977 2685 -961
rect 2687 -977 2703 -961
rect 2741 -977 2757 -961
rect 2759 -977 2775 -961
rect 2823 -977 2839 -961
rect 2841 -977 2857 -961
rect 2895 -977 2911 -961
rect 2913 -977 2929 -961
rect 2977 -977 2993 -961
rect 2995 -977 3011 -961
rect 3049 -977 3065 -961
rect 3067 -977 3083 -961
rect 3131 -977 3147 -961
rect 3149 -977 3165 -961
rect 3203 -977 3219 -961
rect 3221 -977 3237 -961
rect 3285 -977 3301 -961
rect 3303 -977 3319 -961
rect 3357 -977 3373 -961
rect 3375 -977 3391 -961
rect 3439 -977 3455 -961
rect 3457 -977 3473 -961
rect 3511 -977 3527 -961
rect 3529 -977 3545 -961
rect 3593 -977 3609 -961
rect 3611 -977 3627 -961
rect 3665 -977 3681 -961
rect 3683 -977 3699 -961
rect 3747 -977 3760 -961
rect 2361 -1001 2377 -985
rect 2379 -1001 2395 -985
rect 2433 -1001 2449 -985
rect 2451 -1001 2467 -985
rect 2515 -1001 2531 -985
rect 2533 -1001 2549 -985
rect 2587 -1001 2603 -985
rect 2605 -1001 2621 -985
rect 2669 -1001 2685 -985
rect 2687 -1001 2703 -985
rect 2741 -1001 2757 -985
rect 2759 -1001 2775 -985
rect 2823 -1001 2839 -985
rect 2841 -1001 2857 -985
rect 2895 -1001 2911 -985
rect 2913 -1001 2929 -985
rect 2977 -1001 2993 -985
rect 2995 -1001 3011 -985
rect 3049 -1001 3065 -985
rect 3067 -1001 3083 -985
rect 3131 -1001 3147 -985
rect 3149 -1001 3165 -985
rect 3203 -1001 3219 -985
rect 3221 -1001 3237 -985
rect 3285 -1001 3301 -985
rect 3303 -1001 3319 -985
rect 3357 -1001 3373 -985
rect 3375 -1001 3391 -985
rect 3439 -1001 3455 -985
rect 3457 -1001 3473 -985
rect 3511 -1001 3527 -985
rect 3529 -1001 3545 -985
rect 3593 -1001 3609 -985
rect 3611 -1001 3627 -985
rect 3665 -1001 3681 -985
rect 3683 -1001 3699 -985
rect 3747 -1001 3760 -985
rect 2345 -1017 2411 -1001
rect 2417 -1017 2483 -1001
rect 2499 -1017 2565 -1001
rect 2571 -1017 2637 -1001
rect 2653 -1017 2719 -1001
rect 2725 -1017 2791 -1001
rect 2807 -1017 2873 -1001
rect 2879 -1017 2945 -1001
rect 2961 -1017 3027 -1001
rect 3033 -1017 3099 -1001
rect 3115 -1017 3181 -1001
rect 3187 -1017 3253 -1001
rect 3269 -1017 3335 -1001
rect 3341 -1017 3407 -1001
rect 3423 -1017 3489 -1001
rect 3495 -1017 3561 -1001
rect 3577 -1017 3643 -1001
rect 3649 -1017 3715 -1001
rect 3731 -1017 3760 -1001
rect 2361 -1019 2395 -1017
rect 2433 -1019 2467 -1017
rect 2515 -1019 2549 -1017
rect 2587 -1019 2621 -1017
rect 2669 -1019 2703 -1017
rect 2741 -1019 2775 -1017
rect 2823 -1019 2857 -1017
rect 2895 -1019 2929 -1017
rect 2977 -1019 3011 -1017
rect 3049 -1019 3083 -1017
rect 3131 -1019 3165 -1017
rect 3203 -1019 3237 -1017
rect 3285 -1019 3319 -1017
rect 3357 -1019 3391 -1017
rect 3439 -1019 3473 -1017
rect 3511 -1019 3545 -1017
rect 3593 -1019 3627 -1017
rect 3665 -1019 3699 -1017
rect 3747 -1019 3760 -1017
rect 2345 -1035 2411 -1019
rect 2417 -1035 2483 -1019
rect 2499 -1035 2565 -1019
rect 2571 -1035 2637 -1019
rect 2653 -1035 2719 -1019
rect 2725 -1035 2791 -1019
rect 2807 -1035 2873 -1019
rect 2879 -1035 2945 -1019
rect 2961 -1035 3027 -1019
rect 3033 -1035 3099 -1019
rect 3115 -1035 3181 -1019
rect 3187 -1035 3253 -1019
rect 3269 -1035 3335 -1019
rect 3341 -1035 3407 -1019
rect 3423 -1035 3489 -1019
rect 3495 -1035 3561 -1019
rect 3577 -1035 3643 -1019
rect 3649 -1035 3715 -1019
rect 3731 -1035 3760 -1019
rect 2361 -1051 2377 -1035
rect 2379 -1051 2395 -1035
rect 2433 -1051 2449 -1035
rect 2451 -1051 2467 -1035
rect 2515 -1051 2531 -1035
rect 2533 -1051 2549 -1035
rect 2587 -1051 2603 -1035
rect 2605 -1051 2621 -1035
rect 2669 -1051 2685 -1035
rect 2687 -1051 2703 -1035
rect 2741 -1051 2757 -1035
rect 2759 -1051 2775 -1035
rect 2823 -1051 2839 -1035
rect 2841 -1051 2857 -1035
rect 2895 -1051 2911 -1035
rect 2913 -1051 2929 -1035
rect 2977 -1051 2993 -1035
rect 2995 -1051 3011 -1035
rect 3049 -1051 3065 -1035
rect 3067 -1051 3083 -1035
rect 3131 -1051 3147 -1035
rect 3149 -1051 3165 -1035
rect 3203 -1051 3219 -1035
rect 3221 -1051 3237 -1035
rect 3285 -1051 3301 -1035
rect 3303 -1051 3319 -1035
rect 3357 -1051 3373 -1035
rect 3375 -1051 3391 -1035
rect 3439 -1051 3455 -1035
rect 3457 -1051 3473 -1035
rect 3511 -1051 3527 -1035
rect 3529 -1051 3545 -1035
rect 3593 -1051 3609 -1035
rect 3611 -1051 3627 -1035
rect 3665 -1051 3681 -1035
rect 3683 -1051 3699 -1035
rect 3747 -1051 3760 -1035
rect 2407 -1280 2432 -1270
rect 2481 -1280 2506 -1270
rect 2552 -1289 2580 -1270
rect 2544 -1295 2550 -1289
rect 2552 -1295 2585 -1289
rect 2625 -1295 2626 -1289
rect 2629 -1295 2654 -1270
rect 2660 -1295 2666 -1289
rect 2703 -1295 2728 -1270
rect 2741 -1295 2747 -1289
rect 2777 -1295 2802 -1270
rect 2822 -1295 2828 -1289
rect 2851 -1295 2876 -1270
rect 2925 -1289 2950 -1270
rect 2904 -1295 2910 -1289
rect 2925 -1295 2956 -1289
rect 2985 -1295 2991 -1289
rect 2999 -1295 3024 -1270
rect 3031 -1295 3037 -1289
rect 3066 -1295 3070 -1289
rect 3073 -1295 3098 -1270
rect 3112 -1295 3118 -1289
rect 3144 -1295 3146 -1270
rect 3147 -1295 3172 -1270
rect 3193 -1295 3199 -1289
rect 3218 -1295 3246 -1270
rect 3274 -1295 3280 -1289
rect 3292 -1295 3320 -1270
rect 3366 -1289 3394 -1270
rect 3355 -1295 3361 -1289
rect 3366 -1295 3396 -1289
rect 3436 -1295 3440 -1289
rect 3443 -1295 3468 -1270
rect 3472 -1295 3478 -1289
rect 3517 -1295 3542 -1270
rect 3553 -1295 3559 -1289
rect 3591 -1295 3616 -1270
rect 3634 -1295 3640 -1289
rect 3665 -1295 3690 -1270
rect 3715 -1295 3721 -1289
rect 3739 -1295 3760 -1270
rect 23270 -1295 23272 -1289
rect 23275 -1295 23300 -1270
rect 23316 -1295 23322 -1289
rect 23346 -1295 23374 -1270
rect 23397 -1295 23403 -1289
rect 23420 -1295 23448 -1270
rect 23478 -1295 23484 -1289
rect 23494 -1295 23522 -1270
rect 23568 -1289 23596 -1270
rect 23559 -1295 23565 -1289
rect 23568 -1295 23600 -1289
rect 23640 -1295 23642 -1289
rect 23645 -1295 23670 -1270
rect 23675 -1295 23681 -1289
rect 23719 -1295 23744 -1270
rect 23756 -1295 23762 -1289
rect 23793 -1295 23818 -1270
rect 23838 -1295 23844 -1289
rect 23867 -1295 23892 -1270
rect 23941 -1289 23966 -1270
rect 23919 -1295 23925 -1289
rect 23941 -1295 23971 -1289
rect 24000 -1295 24006 -1289
rect 24015 -1295 24040 -1270
rect 24046 -1295 24052 -1289
rect 24081 -1295 24086 -1289
rect 24089 -1295 24114 -1270
rect 24127 -1295 24133 -1289
rect 24160 -1295 24161 -1270
rect 24163 -1295 24188 -1270
rect 24208 -1295 24214 -1289
rect 24234 -1295 24262 -1270
rect 24289 -1295 24295 -1289
rect 24308 -1295 24336 -1270
rect 24382 -1289 24410 -1270
rect 24370 -1295 24376 -1289
rect 24382 -1295 24412 -1289
rect 24452 -1295 24456 -1289
rect 24459 -1295 24484 -1270
rect 24487 -1295 24493 -1289
rect 2524 -1301 2583 -1295
rect 2631 -1301 2637 -1295
rect 2654 -1301 2660 -1295
rect 2712 -1301 2718 -1295
rect 2735 -1301 2741 -1295
rect 2793 -1301 2799 -1295
rect 2816 -1301 2822 -1295
rect 2874 -1301 2880 -1295
rect 2898 -1301 2904 -1295
rect 2956 -1301 2962 -1295
rect 2979 -1301 2985 -1295
rect 3037 -1301 3043 -1295
rect 3060 -1301 3066 -1295
rect 3116 -1301 3124 -1295
rect 3141 -1301 3146 -1295
rect 2524 -1341 2550 -1301
rect 2552 -1341 2583 -1301
rect 2524 -1347 2583 -1341
rect 2631 -1341 2654 -1319
rect 2631 -1347 2660 -1341
rect 2712 -1347 2728 -1319
rect 2735 -1347 2741 -1341
rect 2793 -1347 2802 -1319
rect 2874 -1341 2876 -1319
rect 2816 -1347 2822 -1341
rect 2874 -1347 2880 -1341
rect 2897 -1347 2904 -1319
rect 2956 -1347 2962 -1341
rect 2971 -1347 2985 -1319
rect 3037 -1347 3043 -1341
rect 3045 -1347 3066 -1319
rect 3116 -1341 3118 -1301
rect 3144 -1319 3146 -1301
rect 3119 -1341 3146 -1319
rect 3116 -1347 3146 -1341
rect 3190 -1301 3205 -1295
rect 3218 -1301 3286 -1295
rect 3292 -1301 3397 -1295
rect 3443 -1301 3446 -1295
rect 3466 -1301 3472 -1295
rect 3524 -1301 3530 -1295
rect 3547 -1301 3553 -1295
rect 3605 -1301 3611 -1295
rect 3628 -1301 3634 -1295
rect 3686 -1301 3692 -1295
rect 3709 -1301 3715 -1295
rect 23318 -1301 23328 -1295
rect 23345 -1301 23409 -1295
rect 23420 -1301 23490 -1295
rect 23494 -1301 23599 -1295
rect 23646 -1301 23652 -1295
rect 23669 -1301 23675 -1295
rect 23727 -1301 23733 -1295
rect 23750 -1301 23756 -1295
rect 23808 -1301 23814 -1295
rect 23832 -1301 23838 -1295
rect 23890 -1301 23896 -1295
rect 23913 -1301 23919 -1295
rect 23971 -1301 23977 -1295
rect 23994 -1301 24000 -1295
rect 24052 -1301 24058 -1295
rect 24075 -1301 24081 -1295
rect 24132 -1301 24139 -1295
rect 24157 -1301 24161 -1295
rect 3190 -1341 3199 -1301
rect 3218 -1341 3280 -1301
rect 3292 -1341 3361 -1301
rect 3366 -1341 3397 -1301
rect 3190 -1347 3205 -1341
rect 3218 -1347 3286 -1341
rect 3292 -1347 3397 -1341
rect 3443 -1341 3468 -1319
rect 3443 -1347 3472 -1341
rect 3524 -1347 3542 -1319
rect 3547 -1347 3553 -1341
rect 3605 -1347 3616 -1319
rect 3686 -1341 3690 -1319
rect 3711 -1341 3715 -1319
rect 3628 -1347 3634 -1341
rect 3686 -1347 3692 -1341
rect 3709 -1347 3715 -1341
rect 23318 -1341 23322 -1301
rect 23346 -1341 23403 -1301
rect 23420 -1341 23484 -1301
rect 23494 -1341 23565 -1301
rect 23568 -1341 23599 -1301
rect 23318 -1347 23328 -1341
rect 23345 -1347 23409 -1341
rect 23420 -1347 23490 -1341
rect 23494 -1347 23599 -1341
rect 23646 -1341 23670 -1319
rect 23646 -1347 23675 -1341
rect 23727 -1347 23744 -1319
rect 23750 -1347 23756 -1341
rect 23808 -1347 23818 -1319
rect 23890 -1341 23892 -1319
rect 23832 -1347 23838 -1341
rect 23890 -1347 23896 -1341
rect 23913 -1347 23919 -1319
rect 23971 -1347 23977 -1341
rect 23987 -1347 24000 -1319
rect 24052 -1347 24058 -1341
rect 24061 -1347 24081 -1319
rect 24132 -1341 24133 -1301
rect 24160 -1319 24161 -1301
rect 24135 -1341 24161 -1319
rect 24132 -1347 24161 -1341
rect 24206 -1301 24220 -1295
rect 24234 -1301 24301 -1295
rect 24308 -1301 24413 -1295
rect 24459 -1301 24462 -1295
rect 24481 -1301 24487 -1295
rect 24206 -1341 24214 -1301
rect 24234 -1341 24295 -1301
rect 24308 -1341 24376 -1301
rect 24382 -1341 24413 -1301
rect 24206 -1347 24220 -1341
rect 24234 -1347 24301 -1341
rect 24308 -1347 24413 -1341
rect 24459 -1341 24484 -1319
rect 24459 -1347 24487 -1341
rect 2544 -1353 2550 -1347
rect 2552 -1353 2585 -1347
rect 2625 -1353 2626 -1347
rect 2552 -1393 2580 -1353
rect 2544 -1399 2550 -1393
rect 2552 -1399 2585 -1393
rect 2625 -1399 2626 -1393
rect 2629 -1399 2654 -1347
rect 2660 -1353 2666 -1347
rect 2660 -1399 2666 -1393
rect 2703 -1399 2728 -1347
rect 2741 -1353 2747 -1347
rect 2741 -1399 2747 -1393
rect 2777 -1399 2802 -1347
rect 2822 -1353 2828 -1347
rect 2822 -1399 2828 -1393
rect 2851 -1399 2876 -1347
rect 2904 -1353 2910 -1347
rect 2925 -1353 2956 -1347
rect 2985 -1353 2991 -1347
rect 2925 -1393 2950 -1353
rect 2904 -1399 2910 -1393
rect 2925 -1399 2956 -1393
rect 2985 -1399 2991 -1393
rect 2999 -1399 3024 -1347
rect 3031 -1353 3037 -1347
rect 3066 -1353 3070 -1347
rect 3031 -1399 3037 -1393
rect 3066 -1399 3070 -1393
rect 3073 -1399 3098 -1347
rect 3112 -1353 3118 -1347
rect 3112 -1399 3118 -1393
rect 3144 -1399 3146 -1347
rect 3147 -1399 3172 -1347
rect 3193 -1353 3199 -1347
rect 3193 -1399 3199 -1393
rect 3218 -1399 3246 -1347
rect 3274 -1353 3280 -1347
rect 3274 -1399 3280 -1393
rect 3292 -1399 3320 -1347
rect 3355 -1353 3361 -1347
rect 3366 -1353 3396 -1347
rect 3436 -1353 3440 -1347
rect 3366 -1393 3394 -1353
rect 3355 -1399 3361 -1393
rect 3366 -1399 3396 -1393
rect 3436 -1399 3440 -1393
rect 3443 -1399 3468 -1347
rect 3472 -1353 3478 -1347
rect 3472 -1399 3478 -1393
rect 3517 -1399 3542 -1347
rect 3553 -1353 3559 -1347
rect 3553 -1399 3559 -1393
rect 3591 -1399 3616 -1347
rect 3634 -1353 3640 -1347
rect 3634 -1399 3640 -1393
rect 3665 -1399 3690 -1347
rect 3715 -1353 3721 -1347
rect 3715 -1399 3721 -1393
rect 3739 -1399 3760 -1347
rect 23270 -1353 23272 -1347
rect 23270 -1399 23272 -1393
rect 23275 -1399 23300 -1347
rect 23316 -1353 23322 -1347
rect 23316 -1399 23322 -1393
rect 23346 -1399 23374 -1347
rect 23397 -1353 23403 -1347
rect 23397 -1399 23403 -1393
rect 23420 -1399 23448 -1347
rect 23478 -1353 23484 -1347
rect 23478 -1399 23484 -1393
rect 23494 -1399 23522 -1347
rect 23559 -1353 23565 -1347
rect 23568 -1353 23600 -1347
rect 23640 -1353 23642 -1347
rect 23568 -1393 23596 -1353
rect 23559 -1399 23565 -1393
rect 23568 -1399 23600 -1393
rect 23640 -1399 23642 -1393
rect 23645 -1399 23670 -1347
rect 23675 -1353 23681 -1347
rect 23675 -1399 23681 -1393
rect 23719 -1399 23744 -1347
rect 23756 -1353 23762 -1347
rect 23756 -1399 23762 -1393
rect 23793 -1399 23818 -1347
rect 23838 -1353 23844 -1347
rect 23838 -1399 23844 -1393
rect 23867 -1399 23892 -1347
rect 23919 -1353 23925 -1347
rect 23941 -1353 23971 -1347
rect 24000 -1353 24006 -1347
rect 23941 -1393 23966 -1353
rect 23919 -1399 23925 -1393
rect 23941 -1399 23971 -1393
rect 24000 -1399 24006 -1393
rect 24015 -1399 24040 -1347
rect 24046 -1353 24052 -1347
rect 24081 -1353 24086 -1347
rect 24046 -1399 24052 -1393
rect 24081 -1399 24086 -1393
rect 24089 -1399 24114 -1347
rect 24127 -1353 24133 -1347
rect 24127 -1399 24133 -1393
rect 24160 -1399 24161 -1347
rect 24163 -1399 24188 -1347
rect 24208 -1353 24214 -1347
rect 24208 -1399 24214 -1393
rect 24234 -1399 24262 -1347
rect 24289 -1353 24295 -1347
rect 24289 -1399 24295 -1393
rect 24308 -1399 24336 -1347
rect 24370 -1353 24376 -1347
rect 24382 -1353 24412 -1347
rect 24452 -1353 24456 -1347
rect 24382 -1393 24410 -1353
rect 24370 -1399 24376 -1393
rect 24382 -1399 24412 -1393
rect 24452 -1399 24456 -1393
rect 24459 -1399 24484 -1347
rect 24487 -1353 24493 -1347
rect 24487 -1399 24493 -1393
rect 2524 -1405 2583 -1399
rect 2631 -1405 2637 -1399
rect 2654 -1405 2660 -1399
rect 2712 -1405 2718 -1399
rect 2735 -1405 2741 -1399
rect 2793 -1405 2799 -1399
rect 2816 -1405 2822 -1399
rect 2874 -1405 2880 -1399
rect 2898 -1405 2904 -1399
rect 2956 -1405 2962 -1399
rect 2979 -1405 2985 -1399
rect 3037 -1405 3043 -1399
rect 3060 -1405 3066 -1399
rect 3116 -1405 3124 -1399
rect 3141 -1405 3146 -1399
rect 2524 -1445 2550 -1405
rect 2552 -1445 2583 -1405
rect 2524 -1451 2583 -1445
rect 2631 -1445 2654 -1423
rect 2631 -1451 2660 -1445
rect 2712 -1451 2728 -1423
rect 2735 -1451 2741 -1445
rect 2793 -1451 2802 -1423
rect 2874 -1445 2876 -1423
rect 2816 -1451 2822 -1445
rect 2874 -1451 2880 -1445
rect 2897 -1451 2904 -1423
rect 2956 -1451 2962 -1445
rect 2971 -1451 2985 -1423
rect 3037 -1451 3043 -1445
rect 3045 -1451 3066 -1423
rect 3116 -1445 3118 -1405
rect 3144 -1423 3146 -1405
rect 3119 -1445 3146 -1423
rect 3116 -1451 3146 -1445
rect 3190 -1405 3205 -1399
rect 3218 -1405 3286 -1399
rect 3292 -1405 3397 -1399
rect 3443 -1405 3446 -1399
rect 3466 -1405 3472 -1399
rect 3524 -1405 3530 -1399
rect 3547 -1405 3553 -1399
rect 3605 -1405 3611 -1399
rect 3628 -1405 3634 -1399
rect 3686 -1405 3692 -1399
rect 3709 -1405 3715 -1399
rect 23318 -1405 23328 -1399
rect 23345 -1405 23409 -1399
rect 23420 -1405 23490 -1399
rect 23494 -1405 23599 -1399
rect 23646 -1405 23652 -1399
rect 23669 -1405 23675 -1399
rect 23727 -1405 23733 -1399
rect 23750 -1405 23756 -1399
rect 23808 -1405 23814 -1399
rect 23832 -1405 23838 -1399
rect 23890 -1405 23896 -1399
rect 23913 -1405 23919 -1399
rect 23971 -1405 23977 -1399
rect 23994 -1405 24000 -1399
rect 24052 -1405 24058 -1399
rect 24075 -1405 24081 -1399
rect 24132 -1405 24139 -1399
rect 24157 -1405 24161 -1399
rect 3190 -1445 3199 -1405
rect 3218 -1445 3280 -1405
rect 3292 -1445 3361 -1405
rect 3366 -1445 3397 -1405
rect 3190 -1451 3205 -1445
rect 3218 -1451 3286 -1445
rect 3292 -1451 3397 -1445
rect 3443 -1445 3468 -1423
rect 3443 -1451 3472 -1445
rect 3524 -1451 3542 -1423
rect 3547 -1451 3553 -1445
rect 3605 -1451 3616 -1423
rect 3686 -1445 3690 -1423
rect 3711 -1445 3715 -1423
rect 3628 -1451 3634 -1445
rect 3686 -1451 3692 -1445
rect 3709 -1451 3715 -1445
rect 23318 -1445 23322 -1405
rect 23346 -1445 23403 -1405
rect 23420 -1445 23484 -1405
rect 23494 -1445 23565 -1405
rect 23568 -1445 23599 -1405
rect 23318 -1451 23328 -1445
rect 23345 -1451 23409 -1445
rect 23420 -1451 23490 -1445
rect 23494 -1451 23599 -1445
rect 23646 -1445 23670 -1423
rect 23646 -1451 23675 -1445
rect 23727 -1451 23744 -1423
rect 23750 -1451 23756 -1445
rect 23808 -1451 23818 -1423
rect 23890 -1445 23892 -1423
rect 23832 -1451 23838 -1445
rect 23890 -1451 23896 -1445
rect 23913 -1451 23919 -1423
rect 23971 -1451 23977 -1445
rect 23987 -1451 24000 -1423
rect 24052 -1451 24058 -1445
rect 24061 -1451 24081 -1423
rect 24132 -1445 24133 -1405
rect 24160 -1423 24161 -1405
rect 24135 -1445 24161 -1423
rect 24132 -1451 24161 -1445
rect 24206 -1405 24220 -1399
rect 24234 -1405 24301 -1399
rect 24308 -1405 24413 -1399
rect 24459 -1405 24462 -1399
rect 24481 -1405 24487 -1399
rect 24206 -1445 24214 -1405
rect 24234 -1445 24295 -1405
rect 24308 -1445 24376 -1405
rect 24382 -1445 24413 -1405
rect 24206 -1451 24220 -1445
rect 24234 -1451 24301 -1445
rect 24308 -1451 24413 -1445
rect 24459 -1445 24484 -1423
rect 24459 -1451 24487 -1445
rect 2544 -1457 2550 -1451
rect 2552 -1457 2585 -1451
rect 2625 -1457 2626 -1451
rect 2552 -1497 2580 -1457
rect 2544 -1503 2550 -1497
rect 2552 -1503 2585 -1497
rect 2625 -1503 2626 -1497
rect 2629 -1503 2654 -1451
rect 2660 -1457 2666 -1451
rect 2660 -1503 2666 -1497
rect 2703 -1503 2728 -1451
rect 2741 -1457 2747 -1451
rect 2741 -1503 2747 -1497
rect 2777 -1503 2802 -1451
rect 2822 -1457 2828 -1451
rect 2822 -1503 2828 -1497
rect 2851 -1503 2876 -1451
rect 2904 -1457 2910 -1451
rect 2925 -1457 2956 -1451
rect 2985 -1457 2991 -1451
rect 2925 -1497 2950 -1457
rect 2904 -1503 2910 -1497
rect 2925 -1503 2956 -1497
rect 2985 -1503 2991 -1497
rect 2999 -1503 3024 -1451
rect 3031 -1457 3037 -1451
rect 3066 -1457 3070 -1451
rect 3031 -1503 3037 -1497
rect 3066 -1503 3070 -1497
rect 3073 -1503 3098 -1451
rect 3112 -1457 3118 -1451
rect 3112 -1503 3118 -1497
rect 3144 -1503 3146 -1451
rect 3147 -1503 3172 -1451
rect 3193 -1457 3199 -1451
rect 3193 -1503 3199 -1497
rect 3218 -1503 3246 -1451
rect 3274 -1457 3280 -1451
rect 3274 -1503 3280 -1497
rect 3292 -1503 3320 -1451
rect 3355 -1457 3361 -1451
rect 3366 -1457 3396 -1451
rect 3436 -1457 3440 -1451
rect 3366 -1497 3394 -1457
rect 3355 -1503 3361 -1497
rect 3366 -1503 3396 -1497
rect 3436 -1503 3440 -1497
rect 3443 -1503 3468 -1451
rect 3472 -1457 3478 -1451
rect 3472 -1503 3478 -1497
rect 3517 -1503 3542 -1451
rect 3553 -1457 3559 -1451
rect 3553 -1503 3559 -1497
rect 3591 -1503 3616 -1451
rect 3634 -1457 3640 -1451
rect 3634 -1503 3640 -1497
rect 3665 -1503 3690 -1451
rect 3715 -1457 3721 -1451
rect 3715 -1503 3721 -1497
rect 3739 -1503 3760 -1451
rect 23270 -1457 23272 -1451
rect 23270 -1503 23272 -1497
rect 23275 -1503 23300 -1451
rect 23316 -1457 23322 -1451
rect 23316 -1503 23322 -1497
rect 23346 -1503 23374 -1451
rect 23397 -1457 23403 -1451
rect 23397 -1503 23403 -1497
rect 23420 -1503 23448 -1451
rect 23478 -1457 23484 -1451
rect 23478 -1503 23484 -1497
rect 23494 -1503 23522 -1451
rect 23559 -1457 23565 -1451
rect 23568 -1457 23600 -1451
rect 23640 -1457 23642 -1451
rect 23568 -1497 23596 -1457
rect 23559 -1503 23565 -1497
rect 23568 -1503 23600 -1497
rect 23640 -1503 23642 -1497
rect 23645 -1503 23670 -1451
rect 23675 -1457 23681 -1451
rect 23675 -1503 23681 -1497
rect 23719 -1503 23744 -1451
rect 23756 -1457 23762 -1451
rect 23756 -1503 23762 -1497
rect 23793 -1503 23818 -1451
rect 23838 -1457 23844 -1451
rect 23838 -1503 23844 -1497
rect 23867 -1503 23892 -1451
rect 23919 -1457 23925 -1451
rect 23941 -1457 23971 -1451
rect 24000 -1457 24006 -1451
rect 23941 -1497 23966 -1457
rect 23919 -1503 23925 -1497
rect 23941 -1503 23971 -1497
rect 24000 -1503 24006 -1497
rect 24015 -1503 24040 -1451
rect 24046 -1457 24052 -1451
rect 24081 -1457 24086 -1451
rect 24046 -1503 24052 -1497
rect 24081 -1503 24086 -1497
rect 24089 -1503 24114 -1451
rect 24127 -1457 24133 -1451
rect 24127 -1503 24133 -1497
rect 24160 -1503 24161 -1451
rect 24163 -1503 24188 -1451
rect 24208 -1457 24214 -1451
rect 24208 -1503 24214 -1497
rect 24234 -1503 24262 -1451
rect 24289 -1457 24295 -1451
rect 24289 -1503 24295 -1497
rect 24308 -1503 24336 -1451
rect 24370 -1457 24376 -1451
rect 24382 -1457 24412 -1451
rect 24452 -1457 24456 -1451
rect 24382 -1497 24410 -1457
rect 24370 -1503 24376 -1497
rect 24382 -1503 24412 -1497
rect 24452 -1503 24456 -1497
rect 24459 -1503 24484 -1451
rect 24487 -1457 24493 -1451
rect 24487 -1503 24493 -1497
rect 2524 -1509 2583 -1503
rect 2631 -1509 2637 -1503
rect 2654 -1509 2660 -1503
rect 2712 -1509 2718 -1503
rect 2735 -1509 2741 -1503
rect 2793 -1509 2799 -1503
rect 2816 -1509 2822 -1503
rect 2874 -1509 2880 -1503
rect 2898 -1509 2904 -1503
rect 2956 -1509 2962 -1503
rect 2979 -1509 2985 -1503
rect 3037 -1509 3043 -1503
rect 3060 -1509 3066 -1503
rect 3116 -1509 3124 -1503
rect 3141 -1509 3146 -1503
rect 2524 -1549 2550 -1509
rect 2552 -1549 2583 -1509
rect 2524 -1555 2583 -1549
rect 2631 -1549 2654 -1527
rect 2631 -1555 2660 -1549
rect 2712 -1555 2728 -1527
rect 2735 -1555 2741 -1549
rect 2793 -1555 2802 -1527
rect 2874 -1549 2876 -1527
rect 2816 -1555 2822 -1549
rect 2874 -1555 2880 -1549
rect 2897 -1555 2904 -1527
rect 2956 -1555 2962 -1549
rect 2971 -1555 2985 -1527
rect 3037 -1555 3043 -1549
rect 3045 -1555 3066 -1527
rect 3116 -1549 3118 -1509
rect 3144 -1527 3146 -1509
rect 3119 -1549 3146 -1527
rect 3116 -1555 3146 -1549
rect 3190 -1509 3205 -1503
rect 3218 -1509 3286 -1503
rect 3292 -1509 3397 -1503
rect 3443 -1509 3446 -1503
rect 3466 -1509 3472 -1503
rect 3524 -1509 3530 -1503
rect 3547 -1509 3553 -1503
rect 3605 -1509 3611 -1503
rect 3628 -1509 3634 -1503
rect 3686 -1509 3692 -1503
rect 3709 -1509 3715 -1503
rect 23318 -1509 23328 -1503
rect 23345 -1509 23409 -1503
rect 23420 -1509 23490 -1503
rect 23494 -1509 23599 -1503
rect 23646 -1509 23652 -1503
rect 23669 -1509 23675 -1503
rect 23727 -1509 23733 -1503
rect 23750 -1509 23756 -1503
rect 23808 -1509 23814 -1503
rect 23832 -1509 23838 -1503
rect 23890 -1509 23896 -1503
rect 23913 -1509 23919 -1503
rect 23971 -1509 23977 -1503
rect 23994 -1509 24000 -1503
rect 24052 -1509 24058 -1503
rect 24075 -1509 24081 -1503
rect 24132 -1509 24139 -1503
rect 24157 -1509 24161 -1503
rect 3190 -1549 3199 -1509
rect 3218 -1549 3280 -1509
rect 3292 -1549 3361 -1509
rect 3366 -1549 3397 -1509
rect 3190 -1555 3205 -1549
rect 3218 -1555 3286 -1549
rect 3292 -1555 3397 -1549
rect 3443 -1549 3468 -1527
rect 3443 -1555 3472 -1549
rect 3524 -1555 3542 -1527
rect 3547 -1555 3553 -1549
rect 3605 -1555 3616 -1527
rect 3686 -1549 3690 -1527
rect 3711 -1549 3715 -1527
rect 3628 -1555 3634 -1549
rect 3686 -1555 3692 -1549
rect 3709 -1555 3715 -1549
rect 23318 -1549 23322 -1509
rect 23346 -1549 23403 -1509
rect 23420 -1549 23484 -1509
rect 23494 -1549 23565 -1509
rect 23568 -1549 23599 -1509
rect 23318 -1555 23328 -1549
rect 23345 -1555 23409 -1549
rect 23420 -1555 23490 -1549
rect 23494 -1555 23599 -1549
rect 23646 -1549 23670 -1527
rect 23646 -1555 23675 -1549
rect 23727 -1555 23744 -1527
rect 23750 -1555 23756 -1549
rect 23808 -1555 23818 -1527
rect 23890 -1549 23892 -1527
rect 23832 -1555 23838 -1549
rect 23890 -1555 23896 -1549
rect 23913 -1555 23919 -1527
rect 23971 -1555 23977 -1549
rect 23987 -1555 24000 -1527
rect 24052 -1555 24058 -1549
rect 24061 -1555 24081 -1527
rect 24132 -1549 24133 -1509
rect 24160 -1527 24161 -1509
rect 24135 -1549 24161 -1527
rect 24132 -1555 24161 -1549
rect 24206 -1509 24220 -1503
rect 24234 -1509 24301 -1503
rect 24308 -1509 24413 -1503
rect 24459 -1509 24462 -1503
rect 24481 -1509 24487 -1503
rect 24206 -1549 24214 -1509
rect 24234 -1549 24295 -1509
rect 24308 -1549 24376 -1509
rect 24382 -1549 24413 -1509
rect 24206 -1555 24220 -1549
rect 24234 -1555 24301 -1549
rect 24308 -1555 24413 -1549
rect 24459 -1549 24484 -1527
rect 24459 -1555 24487 -1549
rect 24500 -1555 24530 -1536
rect 2500 -1560 2506 -1555
rect 2407 -1566 2432 -1560
rect 2481 -1566 2506 -1560
rect 2544 -1561 2550 -1555
rect 2552 -1561 2585 -1555
rect 2625 -1561 2626 -1555
rect 2552 -1566 2580 -1561
rect 2629 -1566 2654 -1555
rect 2660 -1561 2666 -1555
rect 2703 -1566 2728 -1555
rect 2741 -1561 2747 -1555
rect 2777 -1566 2802 -1555
rect 2822 -1561 2828 -1555
rect 2851 -1566 2876 -1555
rect 2904 -1561 2910 -1555
rect 2925 -1561 2956 -1555
rect 2985 -1561 2991 -1555
rect 2925 -1566 2950 -1561
rect 2999 -1566 3024 -1555
rect 3031 -1561 3037 -1555
rect 3066 -1561 3070 -1555
rect 3073 -1566 3098 -1555
rect 3112 -1561 3118 -1555
rect 3144 -1566 3146 -1555
rect 3147 -1566 3172 -1555
rect 3193 -1561 3199 -1555
rect 3218 -1566 3246 -1555
rect 3274 -1561 3280 -1555
rect 3292 -1566 3320 -1555
rect 3355 -1561 3361 -1555
rect 3366 -1561 3396 -1555
rect 3436 -1561 3440 -1555
rect 3366 -1566 3394 -1561
rect 3443 -1566 3468 -1555
rect 3472 -1561 3478 -1555
rect 3517 -1566 3542 -1555
rect 3553 -1561 3559 -1555
rect 3591 -1566 3616 -1555
rect 3634 -1561 3640 -1555
rect 3665 -1566 3690 -1555
rect 3715 -1561 3721 -1555
rect 3739 -1566 3760 -1555
rect 23270 -1561 23272 -1555
rect 23275 -1566 23300 -1555
rect 23316 -1561 23322 -1555
rect 23346 -1566 23374 -1555
rect 23397 -1561 23403 -1555
rect 23420 -1566 23448 -1555
rect 23478 -1561 23484 -1555
rect 23494 -1566 23522 -1555
rect 23559 -1561 23565 -1555
rect 23568 -1561 23600 -1555
rect 23640 -1561 23642 -1555
rect 23568 -1566 23596 -1561
rect 23645 -1566 23670 -1555
rect 23675 -1561 23681 -1555
rect 23719 -1566 23744 -1555
rect 23756 -1561 23762 -1555
rect 23793 -1566 23818 -1555
rect 23838 -1561 23844 -1555
rect 23867 -1566 23892 -1555
rect 23919 -1561 23925 -1555
rect 23941 -1561 23971 -1555
rect 24000 -1561 24006 -1555
rect 23941 -1566 23966 -1561
rect 24015 -1566 24040 -1555
rect 24046 -1561 24052 -1555
rect 24081 -1561 24086 -1555
rect 24089 -1566 24114 -1555
rect 24127 -1561 24133 -1555
rect 24160 -1566 24161 -1555
rect 24163 -1566 24188 -1555
rect 24208 -1561 24214 -1555
rect 24234 -1566 24262 -1555
rect 24289 -1561 24295 -1555
rect 24308 -1566 24336 -1555
rect 24370 -1561 24376 -1555
rect 24382 -1561 24412 -1555
rect 24452 -1561 24456 -1555
rect 24382 -1566 24410 -1561
rect 24459 -1566 24484 -1555
rect 24487 -1561 24493 -1555
rect 24528 -1566 24530 -1555
<< pwell >>
rect -976 9244 676 10696
rect 254 -1586 1906 -94
<< nmoslvt >>
rect -950 9870 650 10270
rect 280 -850 1880 -450
<< ndiff >>
rect -950 10608 650 10670
rect -950 10302 -915 10608
rect 615 10302 650 10608
rect -950 10270 650 10302
rect -950 9815 650 9870
rect -950 9645 -915 9815
rect 615 9645 650 9815
rect -950 9610 650 9645
rect 280 -161 1880 -120
rect 280 -399 315 -161
rect 1845 -399 1880 -161
rect 280 -450 1880 -399
rect 280 -880 1880 -850
rect 280 -1050 315 -880
rect 1845 -1050 1880 -880
rect 280 -1080 1880 -1050
<< ndiffc >>
rect -915 10302 615 10608
rect -915 9645 615 9815
rect 315 -399 1845 -161
rect 315 -1050 1845 -880
<< psubdiff >>
rect -950 9559 650 9610
rect -950 9321 -915 9559
rect 615 9321 650 9559
rect -950 9270 650 9321
rect 280 -1116 1880 -1080
rect 280 -1354 315 -1116
rect 1845 -1354 1880 -1116
rect 280 -1560 1880 -1354
<< psubdiffcont >>
rect -915 9321 615 9559
rect 315 -1354 1845 -1116
<< poly >>
rect -980 10080 -950 10270
rect -1370 10060 -950 10080
rect -1370 9890 -1325 10060
rect -1155 9890 -950 10060
rect -1370 9870 -950 9890
rect 650 9870 680 10270
rect -110 -240 100 -230
rect -110 -410 -66 -240
rect 36 -410 100 -240
rect -110 -450 100 -410
rect -110 -500 280 -450
rect 250 -850 280 -500
rect 1880 -850 1910 -450
<< polycont >>
rect -1325 9890 -1155 10060
rect -66 -410 36 -240
<< locali >>
rect -950 10616 650 10650
rect -950 10294 -923 10616
rect 623 10294 650 10616
rect -950 10270 650 10294
rect -1690 10028 -1325 10060
rect -1155 10028 -1020 10060
rect -1690 9922 -1660 10028
rect -1050 9922 -1020 10028
rect -1690 9890 -1325 9922
rect -1155 9890 -1020 9922
rect -950 9815 650 9850
rect -950 9768 -915 9815
rect 615 9768 650 9815
rect -950 9302 -923 9768
rect 623 9302 650 9768
rect -950 9270 650 9302
rect 280 53 1880 60
rect -400 -272 -66 -240
rect -400 -378 -375 -272
rect -125 -378 -66 -272
rect -400 -410 -66 -378
rect 36 -410 100 -240
rect 280 -413 307 53
rect 1853 -413 1880 53
rect 280 -430 1880 -413
rect 280 -880 1880 -870
rect 280 -1050 315 -880
rect 1845 -1050 1880 -880
rect 280 -1116 1880 -1050
rect 280 -1326 315 -1116
rect 1845 -1326 1880 -1116
rect 280 -1504 307 -1326
rect 1853 -1504 1880 -1326
rect 280 -1550 1880 -1504
<< viali >>
rect -923 10608 623 10616
rect -923 10302 -915 10608
rect -915 10302 615 10608
rect 615 10302 623 10608
rect -923 10294 623 10302
rect -1660 9922 -1325 10028
rect -1325 9922 -1155 10028
rect -1155 9922 -1050 10028
rect -923 9645 -915 9768
rect -915 9645 615 9768
rect 615 9645 623 9768
rect -923 9559 623 9645
rect -923 9321 -915 9559
rect -915 9321 615 9559
rect 615 9321 623 9559
rect -923 9302 623 9321
rect -375 -378 -125 -272
rect 307 -161 1853 53
rect 307 -399 315 -161
rect 315 -399 1845 -161
rect 1845 -399 1853 -161
rect 307 -413 1853 -399
rect 307 -1354 315 -1326
rect 315 -1354 1845 -1326
rect 1845 -1354 1853 -1326
rect 307 -1504 1853 -1354
<< metal1 >>
rect 23020 11280 26995 11570
rect -950 10616 650 10630
rect -950 10294 -923 10616
rect 623 10294 650 10616
rect -950 10270 650 10294
rect -2210 10040 -1020 10060
rect -2210 9910 -2200 10040
rect -1030 9910 -1020 10040
rect -2210 9890 -1020 9910
rect -960 9768 650 9850
rect -960 9302 -923 9768
rect 623 9302 650 9768
rect -960 9220 650 9302
rect 280 53 1880 180
rect -500 -272 100 -240
rect -500 -388 -486 -272
rect -114 -388 100 -272
rect -500 -410 100 -388
rect 280 -413 307 53
rect 1853 -413 1880 53
rect 280 -430 1880 -413
rect -950 -1298 2500 -1280
rect -950 -1542 -914 -1298
rect 2274 -1542 2500 -1298
rect -950 -1560 2500 -1542
rect 24530 -1570 26980 -1270
<< via1 >>
rect -912 10301 612 10609
rect -2200 10028 -1030 10040
rect -2200 9922 -1660 10028
rect -1660 9922 -1050 10028
rect -1050 9922 -1030 10028
rect -2200 9910 -1030 9922
rect -912 9317 612 9753
rect -486 -378 -375 -272
rect -375 -378 -125 -272
rect -125 -378 -114 -272
rect -486 -388 -114 -378
rect 318 -398 1842 38
rect -914 -1326 2274 -1298
rect -914 -1504 307 -1326
rect 307 -1504 1853 -1326
rect 1853 -1504 2274 -1326
rect -914 -1542 2274 -1504
<< metal2 >>
rect -950 10609 650 10630
rect -950 10301 -912 10609
rect 612 10301 650 10609
rect -950 10270 650 10301
rect -950 10269 529 10270
rect -2280 10040 -1020 10060
rect -2280 9910 -2200 10040
rect -1030 9910 -1020 10040
rect -2280 9890 -1020 9910
rect -960 9763 650 9850
rect -960 9753 -898 9763
rect 598 9753 650 9763
rect -960 9317 -912 9753
rect 612 9317 650 9753
rect -960 9307 -898 9317
rect 598 9307 650 9317
rect -960 9220 650 9307
rect 1300 8348 2520 8450
rect 1300 7732 1357 8348
rect 2453 7732 2520 8348
rect 1300 7620 2520 7732
rect 280 3859 1890 3870
rect -1688 3611 2174 3859
rect 280 38 1890 3611
rect -1925 -260 -100 -240
rect -1925 -390 -1910 -260
rect -1200 -272 -100 -260
rect -1200 -388 -486 -272
rect -114 -388 -100 -272
rect -1200 -390 -100 -388
rect -1925 -410 -100 -390
rect 280 -398 318 38
rect 1842 -398 1890 38
rect 280 -430 1890 -398
rect -950 -1298 2490 -1280
rect -950 -1542 -914 -1298
rect 2274 -1542 2490 -1298
rect -950 -1560 2490 -1542
<< via2 >>
rect -898 9753 598 9763
rect -898 9317 598 9753
rect -898 9307 598 9317
rect 1357 7732 2453 8348
rect -1910 -390 -1200 -260
rect -908 -1528 2268 -1312
<< metal3 >>
rect -960 9763 650 9850
rect -960 9307 -898 9763
rect 598 9307 650 9763
rect -960 9220 650 9307
rect -2280 -260 -1180 -240
rect -2280 -390 -1910 -260
rect -1200 -390 -1180 -260
rect -2280 -410 -1180 -390
rect -950 -1280 -265 9220
rect 1300 8352 2520 8450
rect 1300 7728 1353 8352
rect 2457 7728 2520 8352
rect 1300 7620 2520 7728
rect -950 -1312 2490 -1280
rect -950 -1528 -908 -1312
rect 2268 -1528 2490 -1312
rect -950 -1560 2490 -1528
<< via3 >>
rect 1353 8348 2457 8352
rect 1353 7732 1357 8348
rect 1357 7732 2453 8348
rect 2453 7732 2457 8348
rect 1353 7728 2457 7732
<< metal4 >>
rect -2205 12835 26620 13665
rect -2205 8455 -1375 12835
rect -2205 8352 2515 8455
rect -2205 7728 1353 8352
rect 2457 7728 2515 8352
rect -2205 7625 2515 7728
rect 25795 7690 26620 12835
rect 24850 6830 26620 7690
use opamp_diego  opamp_diego_0
timestamp 1654624193
transform 1 0 -1719 0 1 8388
box 2069 -10028 26971 3199
<< labels >>
rlabel metal1 s 26840 11440 26840 11440 4 VDD
port 1 nsew
rlabel metal4 s 26418 7258 26418 7258 4 AOUT
port 2 nsew
rlabel metal2 s -1078 -314 -1078 -314 4 OUT_IB
port 3 nsew
rlabel metal2 s -1576 3762 -1576 3762 4 ARRAY_OUT
port 5 nsew
rlabel metal1 s 26870 -1360 26870 -1360 4 GND
port 6 nsew
<< end >>
