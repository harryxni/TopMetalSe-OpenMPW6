magic
tech sky130A
magscale 1 2
timestamp 1654643737
<< error_p >>
rect -855 -347 -797 -341
rect -737 -347 -679 -341
rect -619 -347 -561 -341
rect -501 -347 -443 -341
rect -383 -347 -325 -341
rect -265 -347 -207 -341
rect -147 -347 -89 -341
rect -29 -347 29 -341
rect 89 -347 147 -341
rect 207 -347 265 -341
rect 325 -347 383 -341
rect 443 -347 501 -341
rect 561 -347 619 -341
rect 679 -347 737 -341
rect 797 -347 855 -341
rect -855 -381 -843 -347
rect -737 -381 -725 -347
rect -619 -381 -607 -347
rect -501 -381 -489 -347
rect -383 -381 -371 -347
rect -265 -381 -253 -347
rect -147 -381 -135 -347
rect -29 -381 -17 -347
rect 89 -381 101 -347
rect 207 -381 219 -347
rect 325 -381 337 -347
rect 443 -381 455 -347
rect 561 -381 573 -347
rect 679 -381 691 -347
rect 797 -381 809 -347
rect -855 -387 -797 -381
rect -737 -387 -679 -381
rect -619 -387 -561 -381
rect -501 -387 -443 -381
rect -383 -387 -325 -381
rect -265 -387 -207 -381
rect -147 -387 -89 -381
rect -29 -387 29 -381
rect 89 -387 147 -381
rect 207 -387 265 -381
rect 325 -387 383 -381
rect 443 -387 501 -381
rect 561 -387 619 -381
rect 679 -387 737 -381
rect 797 -387 855 -381
<< nwell >>
rect -1052 -519 1052 519
<< pmos >>
rect -856 -300 -796 300
rect -738 -300 -678 300
rect -620 -300 -560 300
rect -502 -300 -442 300
rect -384 -300 -324 300
rect -266 -300 -206 300
rect -148 -300 -88 300
rect -30 -300 30 300
rect 88 -300 148 300
rect 206 -300 266 300
rect 324 -300 384 300
rect 442 -300 502 300
rect 560 -300 620 300
rect 678 -300 738 300
rect 796 -300 856 300
<< pdiff >>
rect -914 255 -856 300
rect -914 221 -902 255
rect -868 221 -856 255
rect -914 187 -856 221
rect -914 153 -902 187
rect -868 153 -856 187
rect -914 119 -856 153
rect -914 85 -902 119
rect -868 85 -856 119
rect -914 51 -856 85
rect -914 17 -902 51
rect -868 17 -856 51
rect -914 -17 -856 17
rect -914 -51 -902 -17
rect -868 -51 -856 -17
rect -914 -85 -856 -51
rect -914 -119 -902 -85
rect -868 -119 -856 -85
rect -914 -153 -856 -119
rect -914 -187 -902 -153
rect -868 -187 -856 -153
rect -914 -221 -856 -187
rect -914 -255 -902 -221
rect -868 -255 -856 -221
rect -914 -300 -856 -255
rect -796 255 -738 300
rect -796 221 -784 255
rect -750 221 -738 255
rect -796 187 -738 221
rect -796 153 -784 187
rect -750 153 -738 187
rect -796 119 -738 153
rect -796 85 -784 119
rect -750 85 -738 119
rect -796 51 -738 85
rect -796 17 -784 51
rect -750 17 -738 51
rect -796 -17 -738 17
rect -796 -51 -784 -17
rect -750 -51 -738 -17
rect -796 -85 -738 -51
rect -796 -119 -784 -85
rect -750 -119 -738 -85
rect -796 -153 -738 -119
rect -796 -187 -784 -153
rect -750 -187 -738 -153
rect -796 -221 -738 -187
rect -796 -255 -784 -221
rect -750 -255 -738 -221
rect -796 -300 -738 -255
rect -678 255 -620 300
rect -678 221 -666 255
rect -632 221 -620 255
rect -678 187 -620 221
rect -678 153 -666 187
rect -632 153 -620 187
rect -678 119 -620 153
rect -678 85 -666 119
rect -632 85 -620 119
rect -678 51 -620 85
rect -678 17 -666 51
rect -632 17 -620 51
rect -678 -17 -620 17
rect -678 -51 -666 -17
rect -632 -51 -620 -17
rect -678 -85 -620 -51
rect -678 -119 -666 -85
rect -632 -119 -620 -85
rect -678 -153 -620 -119
rect -678 -187 -666 -153
rect -632 -187 -620 -153
rect -678 -221 -620 -187
rect -678 -255 -666 -221
rect -632 -255 -620 -221
rect -678 -300 -620 -255
rect -560 255 -502 300
rect -560 221 -548 255
rect -514 221 -502 255
rect -560 187 -502 221
rect -560 153 -548 187
rect -514 153 -502 187
rect -560 119 -502 153
rect -560 85 -548 119
rect -514 85 -502 119
rect -560 51 -502 85
rect -560 17 -548 51
rect -514 17 -502 51
rect -560 -17 -502 17
rect -560 -51 -548 -17
rect -514 -51 -502 -17
rect -560 -85 -502 -51
rect -560 -119 -548 -85
rect -514 -119 -502 -85
rect -560 -153 -502 -119
rect -560 -187 -548 -153
rect -514 -187 -502 -153
rect -560 -221 -502 -187
rect -560 -255 -548 -221
rect -514 -255 -502 -221
rect -560 -300 -502 -255
rect -442 255 -384 300
rect -442 221 -430 255
rect -396 221 -384 255
rect -442 187 -384 221
rect -442 153 -430 187
rect -396 153 -384 187
rect -442 119 -384 153
rect -442 85 -430 119
rect -396 85 -384 119
rect -442 51 -384 85
rect -442 17 -430 51
rect -396 17 -384 51
rect -442 -17 -384 17
rect -442 -51 -430 -17
rect -396 -51 -384 -17
rect -442 -85 -384 -51
rect -442 -119 -430 -85
rect -396 -119 -384 -85
rect -442 -153 -384 -119
rect -442 -187 -430 -153
rect -396 -187 -384 -153
rect -442 -221 -384 -187
rect -442 -255 -430 -221
rect -396 -255 -384 -221
rect -442 -300 -384 -255
rect -324 255 -266 300
rect -324 221 -312 255
rect -278 221 -266 255
rect -324 187 -266 221
rect -324 153 -312 187
rect -278 153 -266 187
rect -324 119 -266 153
rect -324 85 -312 119
rect -278 85 -266 119
rect -324 51 -266 85
rect -324 17 -312 51
rect -278 17 -266 51
rect -324 -17 -266 17
rect -324 -51 -312 -17
rect -278 -51 -266 -17
rect -324 -85 -266 -51
rect -324 -119 -312 -85
rect -278 -119 -266 -85
rect -324 -153 -266 -119
rect -324 -187 -312 -153
rect -278 -187 -266 -153
rect -324 -221 -266 -187
rect -324 -255 -312 -221
rect -278 -255 -266 -221
rect -324 -300 -266 -255
rect -206 255 -148 300
rect -206 221 -194 255
rect -160 221 -148 255
rect -206 187 -148 221
rect -206 153 -194 187
rect -160 153 -148 187
rect -206 119 -148 153
rect -206 85 -194 119
rect -160 85 -148 119
rect -206 51 -148 85
rect -206 17 -194 51
rect -160 17 -148 51
rect -206 -17 -148 17
rect -206 -51 -194 -17
rect -160 -51 -148 -17
rect -206 -85 -148 -51
rect -206 -119 -194 -85
rect -160 -119 -148 -85
rect -206 -153 -148 -119
rect -206 -187 -194 -153
rect -160 -187 -148 -153
rect -206 -221 -148 -187
rect -206 -255 -194 -221
rect -160 -255 -148 -221
rect -206 -300 -148 -255
rect -88 255 -30 300
rect -88 221 -76 255
rect -42 221 -30 255
rect -88 187 -30 221
rect -88 153 -76 187
rect -42 153 -30 187
rect -88 119 -30 153
rect -88 85 -76 119
rect -42 85 -30 119
rect -88 51 -30 85
rect -88 17 -76 51
rect -42 17 -30 51
rect -88 -17 -30 17
rect -88 -51 -76 -17
rect -42 -51 -30 -17
rect -88 -85 -30 -51
rect -88 -119 -76 -85
rect -42 -119 -30 -85
rect -88 -153 -30 -119
rect -88 -187 -76 -153
rect -42 -187 -30 -153
rect -88 -221 -30 -187
rect -88 -255 -76 -221
rect -42 -255 -30 -221
rect -88 -300 -30 -255
rect 30 255 88 300
rect 30 221 42 255
rect 76 221 88 255
rect 30 187 88 221
rect 30 153 42 187
rect 76 153 88 187
rect 30 119 88 153
rect 30 85 42 119
rect 76 85 88 119
rect 30 51 88 85
rect 30 17 42 51
rect 76 17 88 51
rect 30 -17 88 17
rect 30 -51 42 -17
rect 76 -51 88 -17
rect 30 -85 88 -51
rect 30 -119 42 -85
rect 76 -119 88 -85
rect 30 -153 88 -119
rect 30 -187 42 -153
rect 76 -187 88 -153
rect 30 -221 88 -187
rect 30 -255 42 -221
rect 76 -255 88 -221
rect 30 -300 88 -255
rect 148 255 206 300
rect 148 221 160 255
rect 194 221 206 255
rect 148 187 206 221
rect 148 153 160 187
rect 194 153 206 187
rect 148 119 206 153
rect 148 85 160 119
rect 194 85 206 119
rect 148 51 206 85
rect 148 17 160 51
rect 194 17 206 51
rect 148 -17 206 17
rect 148 -51 160 -17
rect 194 -51 206 -17
rect 148 -85 206 -51
rect 148 -119 160 -85
rect 194 -119 206 -85
rect 148 -153 206 -119
rect 148 -187 160 -153
rect 194 -187 206 -153
rect 148 -221 206 -187
rect 148 -255 160 -221
rect 194 -255 206 -221
rect 148 -300 206 -255
rect 266 255 324 300
rect 266 221 278 255
rect 312 221 324 255
rect 266 187 324 221
rect 266 153 278 187
rect 312 153 324 187
rect 266 119 324 153
rect 266 85 278 119
rect 312 85 324 119
rect 266 51 324 85
rect 266 17 278 51
rect 312 17 324 51
rect 266 -17 324 17
rect 266 -51 278 -17
rect 312 -51 324 -17
rect 266 -85 324 -51
rect 266 -119 278 -85
rect 312 -119 324 -85
rect 266 -153 324 -119
rect 266 -187 278 -153
rect 312 -187 324 -153
rect 266 -221 324 -187
rect 266 -255 278 -221
rect 312 -255 324 -221
rect 266 -300 324 -255
rect 384 255 442 300
rect 384 221 396 255
rect 430 221 442 255
rect 384 187 442 221
rect 384 153 396 187
rect 430 153 442 187
rect 384 119 442 153
rect 384 85 396 119
rect 430 85 442 119
rect 384 51 442 85
rect 384 17 396 51
rect 430 17 442 51
rect 384 -17 442 17
rect 384 -51 396 -17
rect 430 -51 442 -17
rect 384 -85 442 -51
rect 384 -119 396 -85
rect 430 -119 442 -85
rect 384 -153 442 -119
rect 384 -187 396 -153
rect 430 -187 442 -153
rect 384 -221 442 -187
rect 384 -255 396 -221
rect 430 -255 442 -221
rect 384 -300 442 -255
rect 502 255 560 300
rect 502 221 514 255
rect 548 221 560 255
rect 502 187 560 221
rect 502 153 514 187
rect 548 153 560 187
rect 502 119 560 153
rect 502 85 514 119
rect 548 85 560 119
rect 502 51 560 85
rect 502 17 514 51
rect 548 17 560 51
rect 502 -17 560 17
rect 502 -51 514 -17
rect 548 -51 560 -17
rect 502 -85 560 -51
rect 502 -119 514 -85
rect 548 -119 560 -85
rect 502 -153 560 -119
rect 502 -187 514 -153
rect 548 -187 560 -153
rect 502 -221 560 -187
rect 502 -255 514 -221
rect 548 -255 560 -221
rect 502 -300 560 -255
rect 620 255 678 300
rect 620 221 632 255
rect 666 221 678 255
rect 620 187 678 221
rect 620 153 632 187
rect 666 153 678 187
rect 620 119 678 153
rect 620 85 632 119
rect 666 85 678 119
rect 620 51 678 85
rect 620 17 632 51
rect 666 17 678 51
rect 620 -17 678 17
rect 620 -51 632 -17
rect 666 -51 678 -17
rect 620 -85 678 -51
rect 620 -119 632 -85
rect 666 -119 678 -85
rect 620 -153 678 -119
rect 620 -187 632 -153
rect 666 -187 678 -153
rect 620 -221 678 -187
rect 620 -255 632 -221
rect 666 -255 678 -221
rect 620 -300 678 -255
rect 738 255 796 300
rect 738 221 750 255
rect 784 221 796 255
rect 738 187 796 221
rect 738 153 750 187
rect 784 153 796 187
rect 738 119 796 153
rect 738 85 750 119
rect 784 85 796 119
rect 738 51 796 85
rect 738 17 750 51
rect 784 17 796 51
rect 738 -17 796 17
rect 738 -51 750 -17
rect 784 -51 796 -17
rect 738 -85 796 -51
rect 738 -119 750 -85
rect 784 -119 796 -85
rect 738 -153 796 -119
rect 738 -187 750 -153
rect 784 -187 796 -153
rect 738 -221 796 -187
rect 738 -255 750 -221
rect 784 -255 796 -221
rect 738 -300 796 -255
rect 856 255 914 300
rect 856 221 868 255
rect 902 221 914 255
rect 856 187 914 221
rect 856 153 868 187
rect 902 153 914 187
rect 856 119 914 153
rect 856 85 868 119
rect 902 85 914 119
rect 856 51 914 85
rect 856 17 868 51
rect 902 17 914 51
rect 856 -17 914 17
rect 856 -51 868 -17
rect 902 -51 914 -17
rect 856 -85 914 -51
rect 856 -119 868 -85
rect 902 -119 914 -85
rect 856 -153 914 -119
rect 856 -187 868 -153
rect 902 -187 914 -153
rect 856 -221 914 -187
rect 856 -255 868 -221
rect 902 -255 914 -221
rect 856 -300 914 -255
<< pdiffc >>
rect -902 221 -868 255
rect -902 153 -868 187
rect -902 85 -868 119
rect -902 17 -868 51
rect -902 -51 -868 -17
rect -902 -119 -868 -85
rect -902 -187 -868 -153
rect -902 -255 -868 -221
rect -784 221 -750 255
rect -784 153 -750 187
rect -784 85 -750 119
rect -784 17 -750 51
rect -784 -51 -750 -17
rect -784 -119 -750 -85
rect -784 -187 -750 -153
rect -784 -255 -750 -221
rect -666 221 -632 255
rect -666 153 -632 187
rect -666 85 -632 119
rect -666 17 -632 51
rect -666 -51 -632 -17
rect -666 -119 -632 -85
rect -666 -187 -632 -153
rect -666 -255 -632 -221
rect -548 221 -514 255
rect -548 153 -514 187
rect -548 85 -514 119
rect -548 17 -514 51
rect -548 -51 -514 -17
rect -548 -119 -514 -85
rect -548 -187 -514 -153
rect -548 -255 -514 -221
rect -430 221 -396 255
rect -430 153 -396 187
rect -430 85 -396 119
rect -430 17 -396 51
rect -430 -51 -396 -17
rect -430 -119 -396 -85
rect -430 -187 -396 -153
rect -430 -255 -396 -221
rect -312 221 -278 255
rect -312 153 -278 187
rect -312 85 -278 119
rect -312 17 -278 51
rect -312 -51 -278 -17
rect -312 -119 -278 -85
rect -312 -187 -278 -153
rect -312 -255 -278 -221
rect -194 221 -160 255
rect -194 153 -160 187
rect -194 85 -160 119
rect -194 17 -160 51
rect -194 -51 -160 -17
rect -194 -119 -160 -85
rect -194 -187 -160 -153
rect -194 -255 -160 -221
rect -76 221 -42 255
rect -76 153 -42 187
rect -76 85 -42 119
rect -76 17 -42 51
rect -76 -51 -42 -17
rect -76 -119 -42 -85
rect -76 -187 -42 -153
rect -76 -255 -42 -221
rect 42 221 76 255
rect 42 153 76 187
rect 42 85 76 119
rect 42 17 76 51
rect 42 -51 76 -17
rect 42 -119 76 -85
rect 42 -187 76 -153
rect 42 -255 76 -221
rect 160 221 194 255
rect 160 153 194 187
rect 160 85 194 119
rect 160 17 194 51
rect 160 -51 194 -17
rect 160 -119 194 -85
rect 160 -187 194 -153
rect 160 -255 194 -221
rect 278 221 312 255
rect 278 153 312 187
rect 278 85 312 119
rect 278 17 312 51
rect 278 -51 312 -17
rect 278 -119 312 -85
rect 278 -187 312 -153
rect 278 -255 312 -221
rect 396 221 430 255
rect 396 153 430 187
rect 396 85 430 119
rect 396 17 430 51
rect 396 -51 430 -17
rect 396 -119 430 -85
rect 396 -187 430 -153
rect 396 -255 430 -221
rect 514 221 548 255
rect 514 153 548 187
rect 514 85 548 119
rect 514 17 548 51
rect 514 -51 548 -17
rect 514 -119 548 -85
rect 514 -187 548 -153
rect 514 -255 548 -221
rect 632 221 666 255
rect 632 153 666 187
rect 632 85 666 119
rect 632 17 666 51
rect 632 -51 666 -17
rect 632 -119 666 -85
rect 632 -187 666 -153
rect 632 -255 666 -221
rect 750 221 784 255
rect 750 153 784 187
rect 750 85 784 119
rect 750 17 784 51
rect 750 -51 784 -17
rect 750 -119 784 -85
rect 750 -187 784 -153
rect 750 -255 784 -221
rect 868 221 902 255
rect 868 153 902 187
rect 868 85 902 119
rect 868 17 902 51
rect 868 -51 902 -17
rect 868 -119 902 -85
rect 868 -187 902 -153
rect 868 -255 902 -221
<< nsubdiff >>
rect -1016 449 -901 483
rect -867 449 -833 483
rect -799 449 -765 483
rect -731 449 -697 483
rect -663 449 -629 483
rect -595 449 -561 483
rect -527 449 -493 483
rect -459 449 -425 483
rect -391 449 -357 483
rect -323 449 -289 483
rect -255 449 -221 483
rect -187 449 -153 483
rect -119 449 -85 483
rect -51 449 -17 483
rect 17 449 51 483
rect 85 449 119 483
rect 153 449 187 483
rect 221 449 255 483
rect 289 449 323 483
rect 357 449 391 483
rect 425 449 459 483
rect 493 449 527 483
rect 561 449 595 483
rect 629 449 663 483
rect 697 449 731 483
rect 765 449 799 483
rect 833 449 867 483
rect 901 449 1016 483
rect -1016 357 -982 449
rect 982 357 1016 449
rect -1016 289 -982 323
rect -1016 221 -982 255
rect -1016 153 -982 187
rect -1016 85 -982 119
rect -1016 17 -982 51
rect -1016 -51 -982 -17
rect -1016 -119 -982 -85
rect -1016 -187 -982 -153
rect -1016 -255 -982 -221
rect -1016 -323 -982 -289
rect 982 289 1016 323
rect 982 221 1016 255
rect 982 153 1016 187
rect 982 85 1016 119
rect 982 17 1016 51
rect 982 -51 1016 -17
rect 982 -119 1016 -85
rect 982 -187 1016 -153
rect 982 -255 1016 -221
rect 982 -323 1016 -289
rect -1016 -449 -982 -357
rect 982 -449 1016 -357
rect -1016 -483 -901 -449
rect -867 -483 -833 -449
rect -799 -483 -765 -449
rect -731 -483 -697 -449
rect -663 -483 -629 -449
rect -595 -483 -561 -449
rect -527 -483 -493 -449
rect -459 -483 -425 -449
rect -391 -483 -357 -449
rect -323 -483 -289 -449
rect -255 -483 -221 -449
rect -187 -483 -153 -449
rect -119 -483 -85 -449
rect -51 -483 -17 -449
rect 17 -483 51 -449
rect 85 -483 119 -449
rect 153 -483 187 -449
rect 221 -483 255 -449
rect 289 -483 323 -449
rect 357 -483 391 -449
rect 425 -483 459 -449
rect 493 -483 527 -449
rect 561 -483 595 -449
rect 629 -483 663 -449
rect 697 -483 731 -449
rect 765 -483 799 -449
rect 833 -483 867 -449
rect 901 -483 1016 -449
<< nsubdiffcont >>
rect -901 449 -867 483
rect -833 449 -799 483
rect -765 449 -731 483
rect -697 449 -663 483
rect -629 449 -595 483
rect -561 449 -527 483
rect -493 449 -459 483
rect -425 449 -391 483
rect -357 449 -323 483
rect -289 449 -255 483
rect -221 449 -187 483
rect -153 449 -119 483
rect -85 449 -51 483
rect -17 449 17 483
rect 51 449 85 483
rect 119 449 153 483
rect 187 449 221 483
rect 255 449 289 483
rect 323 449 357 483
rect 391 449 425 483
rect 459 449 493 483
rect 527 449 561 483
rect 595 449 629 483
rect 663 449 697 483
rect 731 449 765 483
rect 799 449 833 483
rect 867 449 901 483
rect -1016 323 -982 357
rect 982 323 1016 357
rect -1016 255 -982 289
rect -1016 187 -982 221
rect -1016 119 -982 153
rect -1016 51 -982 85
rect -1016 -17 -982 17
rect -1016 -85 -982 -51
rect -1016 -153 -982 -119
rect -1016 -221 -982 -187
rect -1016 -289 -982 -255
rect 982 255 1016 289
rect 982 187 1016 221
rect 982 119 1016 153
rect 982 51 1016 85
rect 982 -17 1016 17
rect 982 -85 1016 -51
rect 982 -153 1016 -119
rect 982 -221 1016 -187
rect 982 -289 1016 -255
rect -1016 -357 -982 -323
rect 982 -357 1016 -323
rect -901 -483 -867 -449
rect -833 -483 -799 -449
rect -765 -483 -731 -449
rect -697 -483 -663 -449
rect -629 -483 -595 -449
rect -561 -483 -527 -449
rect -493 -483 -459 -449
rect -425 -483 -391 -449
rect -357 -483 -323 -449
rect -289 -483 -255 -449
rect -221 -483 -187 -449
rect -153 -483 -119 -449
rect -85 -483 -51 -449
rect -17 -483 17 -449
rect 51 -483 85 -449
rect 119 -483 153 -449
rect 187 -483 221 -449
rect 255 -483 289 -449
rect 323 -483 357 -449
rect 391 -483 425 -449
rect 459 -483 493 -449
rect 527 -483 561 -449
rect 595 -483 629 -449
rect 663 -483 697 -449
rect 731 -483 765 -449
rect 799 -483 833 -449
rect 867 -483 901 -449
<< poly >>
rect -731 397 -682 399
rect -859 331 -793 397
rect -741 331 -675 397
rect -623 331 -557 397
rect -505 331 -439 397
rect -387 331 -321 397
rect -269 331 -203 397
rect -151 331 -85 397
rect -33 331 33 397
rect 85 331 151 397
rect 203 331 269 397
rect 321 331 387 397
rect 439 331 505 397
rect 557 331 623 397
rect 675 331 741 397
rect 793 331 859 397
rect -856 300 -796 331
rect -738 300 -678 331
rect -620 300 -560 331
rect -502 300 -442 331
rect -384 300 -324 331
rect -266 300 -206 331
rect -148 300 -88 331
rect -30 300 30 331
rect 88 300 148 331
rect 206 300 266 331
rect 324 300 384 331
rect 442 300 502 331
rect 560 300 620 331
rect 678 300 738 331
rect 796 300 856 331
rect -856 -331 -796 -300
rect -738 -331 -678 -300
rect -620 -331 -560 -300
rect -502 -331 -442 -300
rect -384 -331 -324 -300
rect -266 -331 -206 -300
rect -148 -331 -88 -300
rect -30 -331 30 -300
rect 88 -331 148 -300
rect 206 -331 266 -300
rect 324 -331 384 -300
rect 442 -331 502 -300
rect 560 -331 620 -300
rect 678 -331 738 -300
rect 796 -331 856 -300
rect -859 -347 -793 -331
rect -859 -381 -843 -347
rect -809 -381 -793 -347
rect -859 -397 -793 -381
rect -741 -347 -675 -331
rect -741 -381 -725 -347
rect -691 -381 -675 -347
rect -741 -397 -675 -381
rect -623 -347 -557 -331
rect -623 -381 -607 -347
rect -573 -381 -557 -347
rect -623 -397 -557 -381
rect -505 -347 -439 -331
rect -505 -381 -489 -347
rect -455 -381 -439 -347
rect -505 -397 -439 -381
rect -387 -347 -321 -331
rect -387 -381 -371 -347
rect -337 -381 -321 -347
rect -387 -397 -321 -381
rect -269 -347 -203 -331
rect -269 -381 -253 -347
rect -219 -381 -203 -347
rect -269 -397 -203 -381
rect -151 -347 -85 -331
rect -151 -381 -135 -347
rect -101 -381 -85 -347
rect -151 -397 -85 -381
rect -33 -347 33 -331
rect -33 -381 -17 -347
rect 17 -381 33 -347
rect -33 -397 33 -381
rect 85 -347 151 -331
rect 85 -381 101 -347
rect 135 -381 151 -347
rect 85 -397 151 -381
rect 203 -347 269 -331
rect 203 -381 219 -347
rect 253 -381 269 -347
rect 203 -397 269 -381
rect 321 -347 387 -331
rect 321 -381 337 -347
rect 371 -381 387 -347
rect 321 -397 387 -381
rect 439 -347 505 -331
rect 439 -381 455 -347
rect 489 -381 505 -347
rect 439 -397 505 -381
rect 557 -347 623 -331
rect 557 -381 573 -347
rect 607 -381 623 -347
rect 557 -397 623 -381
rect 675 -347 741 -331
rect 675 -381 691 -347
rect 725 -381 741 -347
rect 675 -397 741 -381
rect 793 -347 859 -331
rect 793 -381 809 -347
rect 843 -381 859 -347
rect 793 -397 859 -381
<< polycont >>
rect -843 -381 -809 -347
rect -725 -381 -691 -347
rect -607 -381 -573 -347
rect -489 -381 -455 -347
rect -371 -381 -337 -347
rect -253 -381 -219 -347
rect -135 -381 -101 -347
rect -17 -381 17 -347
rect 101 -381 135 -347
rect 219 -381 253 -347
rect 337 -381 371 -347
rect 455 -381 489 -347
rect 573 -381 607 -347
rect 691 -381 725 -347
rect 809 -381 843 -347
<< locali >>
rect -1016 449 -901 483
rect -867 449 -833 483
rect -799 449 -765 483
rect -731 449 -697 483
rect -663 449 -629 483
rect -595 449 -561 483
rect -527 449 -493 483
rect -459 449 -425 483
rect -391 449 -357 483
rect -323 449 -289 483
rect -255 449 -221 483
rect -187 449 -153 483
rect -119 449 -85 483
rect -51 449 -17 483
rect 17 449 51 483
rect 85 449 119 483
rect 153 449 187 483
rect 221 449 255 483
rect 289 449 323 483
rect 357 449 391 483
rect 425 449 459 483
rect 493 449 527 483
rect 561 449 595 483
rect 629 449 663 483
rect 697 449 731 483
rect 765 449 799 483
rect 833 449 867 483
rect 901 449 1016 483
rect -1016 357 -982 449
rect -1016 289 -982 323
rect 982 357 1016 449
rect -1016 221 -982 255
rect -1016 153 -982 187
rect -1016 85 -982 119
rect -1016 17 -982 51
rect -1016 -51 -982 -17
rect -1016 -119 -982 -85
rect -1016 -187 -982 -153
rect -1016 -255 -982 -221
rect -1016 -323 -982 -289
rect -902 269 -868 304
rect -902 197 -868 221
rect -902 125 -868 153
rect -902 53 -868 85
rect -902 -17 -868 17
rect -902 -85 -868 -53
rect -902 -153 -868 -125
rect -902 -221 -868 -197
rect -902 -304 -868 -269
rect -784 269 -750 304
rect -784 197 -750 221
rect -784 125 -750 153
rect -784 53 -750 85
rect -784 -17 -750 17
rect -784 -85 -750 -53
rect -784 -153 -750 -125
rect -784 -221 -750 -197
rect -784 -304 -750 -269
rect -666 269 -632 304
rect -666 197 -632 221
rect -666 125 -632 153
rect -666 53 -632 85
rect -666 -17 -632 17
rect -666 -85 -632 -53
rect -666 -153 -632 -125
rect -666 -221 -632 -197
rect -666 -304 -632 -269
rect -548 269 -514 304
rect -548 197 -514 221
rect -548 125 -514 153
rect -548 53 -514 85
rect -548 -17 -514 17
rect -548 -85 -514 -53
rect -548 -153 -514 -125
rect -548 -221 -514 -197
rect -548 -304 -514 -269
rect -430 269 -396 304
rect -430 197 -396 221
rect -430 125 -396 153
rect -430 53 -396 85
rect -430 -17 -396 17
rect -430 -85 -396 -53
rect -430 -153 -396 -125
rect -430 -221 -396 -197
rect -430 -304 -396 -269
rect -312 269 -278 304
rect -312 197 -278 221
rect -312 125 -278 153
rect -312 53 -278 85
rect -312 -17 -278 17
rect -312 -85 -278 -53
rect -312 -153 -278 -125
rect -312 -221 -278 -197
rect -312 -304 -278 -269
rect -194 269 -160 304
rect -194 197 -160 221
rect -194 125 -160 153
rect -194 53 -160 85
rect -194 -17 -160 17
rect -194 -85 -160 -53
rect -194 -153 -160 -125
rect -194 -221 -160 -197
rect -194 -304 -160 -269
rect -76 269 -42 304
rect -76 197 -42 221
rect -76 125 -42 153
rect -76 53 -42 85
rect -76 -17 -42 17
rect -76 -85 -42 -53
rect -76 -153 -42 -125
rect -76 -221 -42 -197
rect -76 -304 -42 -269
rect 42 269 76 304
rect 42 197 76 221
rect 42 125 76 153
rect 42 53 76 85
rect 42 -17 76 17
rect 42 -85 76 -53
rect 42 -153 76 -125
rect 42 -221 76 -197
rect 42 -304 76 -269
rect 160 269 194 304
rect 160 197 194 221
rect 160 125 194 153
rect 160 53 194 85
rect 160 -17 194 17
rect 160 -85 194 -53
rect 160 -153 194 -125
rect 160 -221 194 -197
rect 160 -304 194 -269
rect 278 269 312 304
rect 278 197 312 221
rect 278 125 312 153
rect 278 53 312 85
rect 278 -17 312 17
rect 278 -85 312 -53
rect 278 -153 312 -125
rect 278 -221 312 -197
rect 278 -304 312 -269
rect 396 269 430 304
rect 396 197 430 221
rect 396 125 430 153
rect 396 53 430 85
rect 396 -17 430 17
rect 396 -85 430 -53
rect 396 -153 430 -125
rect 396 -221 430 -197
rect 396 -304 430 -269
rect 514 269 548 304
rect 514 197 548 221
rect 514 125 548 153
rect 514 53 548 85
rect 514 -17 548 17
rect 514 -85 548 -53
rect 514 -153 548 -125
rect 514 -221 548 -197
rect 514 -304 548 -269
rect 632 269 666 304
rect 632 197 666 221
rect 632 125 666 153
rect 632 53 666 85
rect 632 -17 666 17
rect 632 -85 666 -53
rect 632 -153 666 -125
rect 632 -221 666 -197
rect 632 -304 666 -269
rect 750 269 784 304
rect 750 197 784 221
rect 750 125 784 153
rect 750 53 784 85
rect 750 -17 784 17
rect 750 -85 784 -53
rect 750 -153 784 -125
rect 750 -221 784 -197
rect 750 -304 784 -269
rect 868 269 902 304
rect 868 197 902 221
rect 868 125 902 153
rect 868 53 902 85
rect 868 -17 902 17
rect 868 -85 902 -53
rect 868 -153 902 -125
rect 868 -221 902 -197
rect 868 -304 902 -269
rect 982 289 1016 323
rect 982 221 1016 255
rect 982 153 1016 187
rect 982 85 1016 119
rect 982 17 1016 51
rect 982 -51 1016 -17
rect 982 -119 1016 -85
rect 982 -187 1016 -153
rect 982 -255 1016 -221
rect 982 -323 1016 -289
rect -1016 -449 -982 -357
rect -859 -381 -843 -347
rect -809 -381 -793 -347
rect -741 -381 -725 -347
rect -691 -381 -675 -347
rect -623 -381 -607 -347
rect -573 -381 -557 -347
rect -505 -381 -489 -347
rect -455 -381 -439 -347
rect -387 -381 -371 -347
rect -337 -381 -321 -347
rect -269 -381 -253 -347
rect -219 -381 -203 -347
rect -151 -381 -135 -347
rect -101 -381 -85 -347
rect -33 -381 -17 -347
rect 17 -381 33 -347
rect 85 -381 101 -347
rect 135 -381 151 -347
rect 203 -381 219 -347
rect 253 -381 269 -347
rect 321 -381 337 -347
rect 371 -381 387 -347
rect 439 -381 455 -347
rect 489 -381 505 -347
rect 557 -381 573 -347
rect 607 -381 623 -347
rect 675 -381 691 -347
rect 725 -381 741 -347
rect 793 -381 809 -347
rect 843 -381 859 -347
rect 982 -449 1016 -357
rect -1016 -483 -901 -449
rect -867 -483 -833 -449
rect -799 -483 -765 -449
rect -731 -483 -697 -449
rect -663 -483 -629 -449
rect -595 -483 -561 -449
rect -527 -483 -493 -449
rect -459 -483 -425 -449
rect -391 -483 -357 -449
rect -323 -483 -289 -449
rect -255 -483 -221 -449
rect -187 -483 -153 -449
rect -119 -483 -85 -449
rect -51 -483 -17 -449
rect 17 -483 51 -449
rect 85 -483 119 -449
rect 153 -483 187 -449
rect 221 -483 255 -449
rect 289 -483 323 -449
rect 357 -483 391 -449
rect 425 -483 459 -449
rect 493 -483 527 -449
rect 561 -483 595 -449
rect 629 -483 663 -449
rect 697 -483 731 -449
rect 765 -483 799 -449
rect 833 -483 867 -449
rect 901 -483 1016 -449
<< viali >>
rect -902 255 -868 269
rect -902 235 -868 255
rect -902 187 -868 197
rect -902 163 -868 187
rect -902 119 -868 125
rect -902 91 -868 119
rect -902 51 -868 53
rect -902 19 -868 51
rect -902 -51 -868 -19
rect -902 -53 -868 -51
rect -902 -119 -868 -91
rect -902 -125 -868 -119
rect -902 -187 -868 -163
rect -902 -197 -868 -187
rect -902 -255 -868 -235
rect -902 -269 -868 -255
rect -784 255 -750 269
rect -784 235 -750 255
rect -784 187 -750 197
rect -784 163 -750 187
rect -784 119 -750 125
rect -784 91 -750 119
rect -784 51 -750 53
rect -784 19 -750 51
rect -784 -51 -750 -19
rect -784 -53 -750 -51
rect -784 -119 -750 -91
rect -784 -125 -750 -119
rect -784 -187 -750 -163
rect -784 -197 -750 -187
rect -784 -255 -750 -235
rect -784 -269 -750 -255
rect -666 255 -632 269
rect -666 235 -632 255
rect -666 187 -632 197
rect -666 163 -632 187
rect -666 119 -632 125
rect -666 91 -632 119
rect -666 51 -632 53
rect -666 19 -632 51
rect -666 -51 -632 -19
rect -666 -53 -632 -51
rect -666 -119 -632 -91
rect -666 -125 -632 -119
rect -666 -187 -632 -163
rect -666 -197 -632 -187
rect -666 -255 -632 -235
rect -666 -269 -632 -255
rect -548 255 -514 269
rect -548 235 -514 255
rect -548 187 -514 197
rect -548 163 -514 187
rect -548 119 -514 125
rect -548 91 -514 119
rect -548 51 -514 53
rect -548 19 -514 51
rect -548 -51 -514 -19
rect -548 -53 -514 -51
rect -548 -119 -514 -91
rect -548 -125 -514 -119
rect -548 -187 -514 -163
rect -548 -197 -514 -187
rect -548 -255 -514 -235
rect -548 -269 -514 -255
rect -430 255 -396 269
rect -430 235 -396 255
rect -430 187 -396 197
rect -430 163 -396 187
rect -430 119 -396 125
rect -430 91 -396 119
rect -430 51 -396 53
rect -430 19 -396 51
rect -430 -51 -396 -19
rect -430 -53 -396 -51
rect -430 -119 -396 -91
rect -430 -125 -396 -119
rect -430 -187 -396 -163
rect -430 -197 -396 -187
rect -430 -255 -396 -235
rect -430 -269 -396 -255
rect -312 255 -278 269
rect -312 235 -278 255
rect -312 187 -278 197
rect -312 163 -278 187
rect -312 119 -278 125
rect -312 91 -278 119
rect -312 51 -278 53
rect -312 19 -278 51
rect -312 -51 -278 -19
rect -312 -53 -278 -51
rect -312 -119 -278 -91
rect -312 -125 -278 -119
rect -312 -187 -278 -163
rect -312 -197 -278 -187
rect -312 -255 -278 -235
rect -312 -269 -278 -255
rect -194 255 -160 269
rect -194 235 -160 255
rect -194 187 -160 197
rect -194 163 -160 187
rect -194 119 -160 125
rect -194 91 -160 119
rect -194 51 -160 53
rect -194 19 -160 51
rect -194 -51 -160 -19
rect -194 -53 -160 -51
rect -194 -119 -160 -91
rect -194 -125 -160 -119
rect -194 -187 -160 -163
rect -194 -197 -160 -187
rect -194 -255 -160 -235
rect -194 -269 -160 -255
rect -76 255 -42 269
rect -76 235 -42 255
rect -76 187 -42 197
rect -76 163 -42 187
rect -76 119 -42 125
rect -76 91 -42 119
rect -76 51 -42 53
rect -76 19 -42 51
rect -76 -51 -42 -19
rect -76 -53 -42 -51
rect -76 -119 -42 -91
rect -76 -125 -42 -119
rect -76 -187 -42 -163
rect -76 -197 -42 -187
rect -76 -255 -42 -235
rect -76 -269 -42 -255
rect 42 255 76 269
rect 42 235 76 255
rect 42 187 76 197
rect 42 163 76 187
rect 42 119 76 125
rect 42 91 76 119
rect 42 51 76 53
rect 42 19 76 51
rect 42 -51 76 -19
rect 42 -53 76 -51
rect 42 -119 76 -91
rect 42 -125 76 -119
rect 42 -187 76 -163
rect 42 -197 76 -187
rect 42 -255 76 -235
rect 42 -269 76 -255
rect 160 255 194 269
rect 160 235 194 255
rect 160 187 194 197
rect 160 163 194 187
rect 160 119 194 125
rect 160 91 194 119
rect 160 51 194 53
rect 160 19 194 51
rect 160 -51 194 -19
rect 160 -53 194 -51
rect 160 -119 194 -91
rect 160 -125 194 -119
rect 160 -187 194 -163
rect 160 -197 194 -187
rect 160 -255 194 -235
rect 160 -269 194 -255
rect 278 255 312 269
rect 278 235 312 255
rect 278 187 312 197
rect 278 163 312 187
rect 278 119 312 125
rect 278 91 312 119
rect 278 51 312 53
rect 278 19 312 51
rect 278 -51 312 -19
rect 278 -53 312 -51
rect 278 -119 312 -91
rect 278 -125 312 -119
rect 278 -187 312 -163
rect 278 -197 312 -187
rect 278 -255 312 -235
rect 278 -269 312 -255
rect 396 255 430 269
rect 396 235 430 255
rect 396 187 430 197
rect 396 163 430 187
rect 396 119 430 125
rect 396 91 430 119
rect 396 51 430 53
rect 396 19 430 51
rect 396 -51 430 -19
rect 396 -53 430 -51
rect 396 -119 430 -91
rect 396 -125 430 -119
rect 396 -187 430 -163
rect 396 -197 430 -187
rect 396 -255 430 -235
rect 396 -269 430 -255
rect 514 255 548 269
rect 514 235 548 255
rect 514 187 548 197
rect 514 163 548 187
rect 514 119 548 125
rect 514 91 548 119
rect 514 51 548 53
rect 514 19 548 51
rect 514 -51 548 -19
rect 514 -53 548 -51
rect 514 -119 548 -91
rect 514 -125 548 -119
rect 514 -187 548 -163
rect 514 -197 548 -187
rect 514 -255 548 -235
rect 514 -269 548 -255
rect 632 255 666 269
rect 632 235 666 255
rect 632 187 666 197
rect 632 163 666 187
rect 632 119 666 125
rect 632 91 666 119
rect 632 51 666 53
rect 632 19 666 51
rect 632 -51 666 -19
rect 632 -53 666 -51
rect 632 -119 666 -91
rect 632 -125 666 -119
rect 632 -187 666 -163
rect 632 -197 666 -187
rect 632 -255 666 -235
rect 632 -269 666 -255
rect 750 255 784 269
rect 750 235 784 255
rect 750 187 784 197
rect 750 163 784 187
rect 750 119 784 125
rect 750 91 784 119
rect 750 51 784 53
rect 750 19 784 51
rect 750 -51 784 -19
rect 750 -53 784 -51
rect 750 -119 784 -91
rect 750 -125 784 -119
rect 750 -187 784 -163
rect 750 -197 784 -187
rect 750 -255 784 -235
rect 750 -269 784 -255
rect 868 255 902 269
rect 868 235 902 255
rect 868 187 902 197
rect 868 163 902 187
rect 868 119 902 125
rect 868 91 902 119
rect 868 51 902 53
rect 868 19 902 51
rect 868 -51 902 -19
rect 868 -53 902 -51
rect 868 -119 902 -91
rect 868 -125 902 -119
rect 868 -187 902 -163
rect 868 -197 902 -187
rect 868 -255 902 -235
rect 868 -269 902 -255
rect -843 -381 -809 -347
rect -725 -381 -691 -347
rect -607 -381 -573 -347
rect -489 -381 -455 -347
rect -371 -381 -337 -347
rect -253 -381 -219 -347
rect -135 -381 -101 -347
rect -17 -381 17 -347
rect 101 -381 135 -347
rect 219 -381 253 -347
rect 337 -381 371 -347
rect 455 -381 489 -347
rect 573 -381 607 -347
rect 691 -381 725 -347
rect 809 -381 843 -347
<< metal1 >>
rect -908 269 -862 300
rect -908 235 -902 269
rect -868 235 -862 269
rect -908 197 -862 235
rect -908 163 -902 197
rect -868 163 -862 197
rect -908 125 -862 163
rect -908 91 -902 125
rect -868 91 -862 125
rect -908 53 -862 91
rect -908 19 -902 53
rect -868 19 -862 53
rect -908 -19 -862 19
rect -908 -53 -902 -19
rect -868 -53 -862 -19
rect -908 -91 -862 -53
rect -908 -125 -902 -91
rect -868 -125 -862 -91
rect -908 -163 -862 -125
rect -908 -197 -902 -163
rect -868 -197 -862 -163
rect -908 -235 -862 -197
rect -908 -269 -902 -235
rect -868 -269 -862 -235
rect -908 -300 -862 -269
rect -790 269 -744 300
rect -790 235 -784 269
rect -750 235 -744 269
rect -790 197 -744 235
rect -790 163 -784 197
rect -750 163 -744 197
rect -790 125 -744 163
rect -790 91 -784 125
rect -750 91 -744 125
rect -790 53 -744 91
rect -790 19 -784 53
rect -750 19 -744 53
rect -790 -19 -744 19
rect -790 -53 -784 -19
rect -750 -53 -744 -19
rect -790 -91 -744 -53
rect -790 -125 -784 -91
rect -750 -125 -744 -91
rect -790 -163 -744 -125
rect -790 -197 -784 -163
rect -750 -197 -744 -163
rect -790 -235 -744 -197
rect -790 -269 -784 -235
rect -750 -269 -744 -235
rect -790 -300 -744 -269
rect -672 269 -626 300
rect -672 235 -666 269
rect -632 235 -626 269
rect -672 197 -626 235
rect -672 163 -666 197
rect -632 163 -626 197
rect -672 125 -626 163
rect -672 91 -666 125
rect -632 91 -626 125
rect -672 53 -626 91
rect -672 19 -666 53
rect -632 19 -626 53
rect -672 -19 -626 19
rect -672 -53 -666 -19
rect -632 -53 -626 -19
rect -672 -91 -626 -53
rect -672 -125 -666 -91
rect -632 -125 -626 -91
rect -672 -163 -626 -125
rect -672 -197 -666 -163
rect -632 -197 -626 -163
rect -672 -235 -626 -197
rect -672 -269 -666 -235
rect -632 -269 -626 -235
rect -672 -300 -626 -269
rect -554 269 -508 300
rect -554 235 -548 269
rect -514 235 -508 269
rect -554 197 -508 235
rect -554 163 -548 197
rect -514 163 -508 197
rect -554 125 -508 163
rect -554 91 -548 125
rect -514 91 -508 125
rect -554 53 -508 91
rect -554 19 -548 53
rect -514 19 -508 53
rect -554 -19 -508 19
rect -554 -53 -548 -19
rect -514 -53 -508 -19
rect -554 -91 -508 -53
rect -554 -125 -548 -91
rect -514 -125 -508 -91
rect -554 -163 -508 -125
rect -554 -197 -548 -163
rect -514 -197 -508 -163
rect -554 -235 -508 -197
rect -554 -269 -548 -235
rect -514 -269 -508 -235
rect -554 -300 -508 -269
rect -436 269 -390 300
rect -436 235 -430 269
rect -396 235 -390 269
rect -436 197 -390 235
rect -436 163 -430 197
rect -396 163 -390 197
rect -436 125 -390 163
rect -436 91 -430 125
rect -396 91 -390 125
rect -436 53 -390 91
rect -436 19 -430 53
rect -396 19 -390 53
rect -436 -19 -390 19
rect -436 -53 -430 -19
rect -396 -53 -390 -19
rect -436 -91 -390 -53
rect -436 -125 -430 -91
rect -396 -125 -390 -91
rect -436 -163 -390 -125
rect -436 -197 -430 -163
rect -396 -197 -390 -163
rect -436 -235 -390 -197
rect -436 -269 -430 -235
rect -396 -269 -390 -235
rect -436 -300 -390 -269
rect -318 269 -272 300
rect -318 235 -312 269
rect -278 235 -272 269
rect -318 197 -272 235
rect -318 163 -312 197
rect -278 163 -272 197
rect -318 125 -272 163
rect -318 91 -312 125
rect -278 91 -272 125
rect -318 53 -272 91
rect -318 19 -312 53
rect -278 19 -272 53
rect -318 -19 -272 19
rect -318 -53 -312 -19
rect -278 -53 -272 -19
rect -318 -91 -272 -53
rect -318 -125 -312 -91
rect -278 -125 -272 -91
rect -318 -163 -272 -125
rect -318 -197 -312 -163
rect -278 -197 -272 -163
rect -318 -235 -272 -197
rect -318 -269 -312 -235
rect -278 -269 -272 -235
rect -318 -300 -272 -269
rect -200 269 -154 300
rect -200 235 -194 269
rect -160 235 -154 269
rect -200 197 -154 235
rect -200 163 -194 197
rect -160 163 -154 197
rect -200 125 -154 163
rect -200 91 -194 125
rect -160 91 -154 125
rect -200 53 -154 91
rect -200 19 -194 53
rect -160 19 -154 53
rect -200 -19 -154 19
rect -200 -53 -194 -19
rect -160 -53 -154 -19
rect -200 -91 -154 -53
rect -200 -125 -194 -91
rect -160 -125 -154 -91
rect -200 -163 -154 -125
rect -200 -197 -194 -163
rect -160 -197 -154 -163
rect -200 -235 -154 -197
rect -200 -269 -194 -235
rect -160 -269 -154 -235
rect -200 -300 -154 -269
rect -82 269 -36 300
rect -82 235 -76 269
rect -42 235 -36 269
rect -82 197 -36 235
rect -82 163 -76 197
rect -42 163 -36 197
rect -82 125 -36 163
rect -82 91 -76 125
rect -42 91 -36 125
rect -82 53 -36 91
rect -82 19 -76 53
rect -42 19 -36 53
rect -82 -19 -36 19
rect -82 -53 -76 -19
rect -42 -53 -36 -19
rect -82 -91 -36 -53
rect -82 -125 -76 -91
rect -42 -125 -36 -91
rect -82 -163 -36 -125
rect -82 -197 -76 -163
rect -42 -197 -36 -163
rect -82 -235 -36 -197
rect -82 -269 -76 -235
rect -42 -269 -36 -235
rect -82 -300 -36 -269
rect 36 269 82 300
rect 36 235 42 269
rect 76 235 82 269
rect 36 197 82 235
rect 36 163 42 197
rect 76 163 82 197
rect 36 125 82 163
rect 36 91 42 125
rect 76 91 82 125
rect 36 53 82 91
rect 36 19 42 53
rect 76 19 82 53
rect 36 -19 82 19
rect 36 -53 42 -19
rect 76 -53 82 -19
rect 36 -91 82 -53
rect 36 -125 42 -91
rect 76 -125 82 -91
rect 36 -163 82 -125
rect 36 -197 42 -163
rect 76 -197 82 -163
rect 36 -235 82 -197
rect 36 -269 42 -235
rect 76 -269 82 -235
rect 36 -300 82 -269
rect 154 269 200 300
rect 154 235 160 269
rect 194 235 200 269
rect 154 197 200 235
rect 154 163 160 197
rect 194 163 200 197
rect 154 125 200 163
rect 154 91 160 125
rect 194 91 200 125
rect 154 53 200 91
rect 154 19 160 53
rect 194 19 200 53
rect 154 -19 200 19
rect 154 -53 160 -19
rect 194 -53 200 -19
rect 154 -91 200 -53
rect 154 -125 160 -91
rect 194 -125 200 -91
rect 154 -163 200 -125
rect 154 -197 160 -163
rect 194 -197 200 -163
rect 154 -235 200 -197
rect 154 -269 160 -235
rect 194 -269 200 -235
rect 154 -300 200 -269
rect 272 269 318 300
rect 272 235 278 269
rect 312 235 318 269
rect 272 197 318 235
rect 272 163 278 197
rect 312 163 318 197
rect 272 125 318 163
rect 272 91 278 125
rect 312 91 318 125
rect 272 53 318 91
rect 272 19 278 53
rect 312 19 318 53
rect 272 -19 318 19
rect 272 -53 278 -19
rect 312 -53 318 -19
rect 272 -91 318 -53
rect 272 -125 278 -91
rect 312 -125 318 -91
rect 272 -163 318 -125
rect 272 -197 278 -163
rect 312 -197 318 -163
rect 272 -235 318 -197
rect 272 -269 278 -235
rect 312 -269 318 -235
rect 272 -300 318 -269
rect 390 269 436 300
rect 390 235 396 269
rect 430 235 436 269
rect 390 197 436 235
rect 390 163 396 197
rect 430 163 436 197
rect 390 125 436 163
rect 390 91 396 125
rect 430 91 436 125
rect 390 53 436 91
rect 390 19 396 53
rect 430 19 436 53
rect 390 -19 436 19
rect 390 -53 396 -19
rect 430 -53 436 -19
rect 390 -91 436 -53
rect 390 -125 396 -91
rect 430 -125 436 -91
rect 390 -163 436 -125
rect 390 -197 396 -163
rect 430 -197 436 -163
rect 390 -235 436 -197
rect 390 -269 396 -235
rect 430 -269 436 -235
rect 390 -300 436 -269
rect 508 269 554 300
rect 508 235 514 269
rect 548 235 554 269
rect 508 197 554 235
rect 508 163 514 197
rect 548 163 554 197
rect 508 125 554 163
rect 508 91 514 125
rect 548 91 554 125
rect 508 53 554 91
rect 508 19 514 53
rect 548 19 554 53
rect 508 -19 554 19
rect 508 -53 514 -19
rect 548 -53 554 -19
rect 508 -91 554 -53
rect 508 -125 514 -91
rect 548 -125 554 -91
rect 508 -163 554 -125
rect 508 -197 514 -163
rect 548 -197 554 -163
rect 508 -235 554 -197
rect 508 -269 514 -235
rect 548 -269 554 -235
rect 508 -300 554 -269
rect 626 269 672 300
rect 626 235 632 269
rect 666 235 672 269
rect 626 197 672 235
rect 626 163 632 197
rect 666 163 672 197
rect 626 125 672 163
rect 626 91 632 125
rect 666 91 672 125
rect 626 53 672 91
rect 626 19 632 53
rect 666 19 672 53
rect 626 -19 672 19
rect 626 -53 632 -19
rect 666 -53 672 -19
rect 626 -91 672 -53
rect 626 -125 632 -91
rect 666 -125 672 -91
rect 626 -163 672 -125
rect 626 -197 632 -163
rect 666 -197 672 -163
rect 626 -235 672 -197
rect 626 -269 632 -235
rect 666 -269 672 -235
rect 626 -300 672 -269
rect 744 269 790 300
rect 744 235 750 269
rect 784 235 790 269
rect 744 197 790 235
rect 744 163 750 197
rect 784 163 790 197
rect 744 125 790 163
rect 744 91 750 125
rect 784 91 790 125
rect 744 53 790 91
rect 744 19 750 53
rect 784 19 790 53
rect 744 -19 790 19
rect 744 -53 750 -19
rect 784 -53 790 -19
rect 744 -91 790 -53
rect 744 -125 750 -91
rect 784 -125 790 -91
rect 744 -163 790 -125
rect 744 -197 750 -163
rect 784 -197 790 -163
rect 744 -235 790 -197
rect 744 -269 750 -235
rect 784 -269 790 -235
rect 744 -300 790 -269
rect 862 269 908 300
rect 862 235 868 269
rect 902 235 908 269
rect 862 197 908 235
rect 862 163 868 197
rect 902 163 908 197
rect 862 125 908 163
rect 862 91 868 125
rect 902 91 908 125
rect 862 53 908 91
rect 862 19 868 53
rect 902 19 908 53
rect 862 -19 908 19
rect 862 -53 868 -19
rect 902 -53 908 -19
rect 862 -91 908 -53
rect 862 -125 868 -91
rect 902 -125 908 -91
rect 862 -163 908 -125
rect 862 -197 868 -163
rect 902 -197 908 -163
rect 862 -235 908 -197
rect 862 -269 868 -235
rect 902 -269 908 -235
rect 862 -300 908 -269
rect -855 -347 -797 -341
rect -855 -381 -843 -347
rect -809 -381 -797 -347
rect -855 -387 -797 -381
rect -737 -347 -679 -341
rect -737 -381 -725 -347
rect -691 -381 -679 -347
rect -737 -387 -679 -381
rect -619 -347 -561 -341
rect -619 -381 -607 -347
rect -573 -381 -561 -347
rect -619 -387 -561 -381
rect -501 -347 -443 -341
rect -501 -381 -489 -347
rect -455 -381 -443 -347
rect -501 -387 -443 -381
rect -383 -347 -325 -341
rect -383 -381 -371 -347
rect -337 -381 -325 -347
rect -383 -387 -325 -381
rect -265 -347 -207 -341
rect -265 -381 -253 -347
rect -219 -381 -207 -347
rect -265 -387 -207 -381
rect -147 -347 -89 -341
rect -147 -381 -135 -347
rect -101 -381 -89 -347
rect -147 -387 -89 -381
rect -29 -347 29 -341
rect -29 -381 -17 -347
rect 17 -381 29 -347
rect -29 -387 29 -381
rect 89 -347 147 -341
rect 89 -381 101 -347
rect 135 -381 147 -347
rect 89 -387 147 -381
rect 207 -347 265 -341
rect 207 -381 219 -347
rect 253 -381 265 -347
rect 207 -387 265 -381
rect 325 -347 383 -341
rect 325 -381 337 -347
rect 371 -381 383 -347
rect 325 -387 383 -381
rect 443 -347 501 -341
rect 443 -381 455 -347
rect 489 -381 501 -347
rect 443 -387 501 -381
rect 561 -347 619 -341
rect 561 -381 573 -347
rect 607 -381 619 -347
rect 561 -387 619 -381
rect 679 -347 737 -341
rect 679 -381 691 -347
rect 725 -381 737 -347
rect 679 -387 737 -381
rect 797 -347 855 -341
rect 797 -381 809 -347
rect 843 -381 855 -347
rect 797 -387 855 -381
<< properties >>
string FIXED_BBOX -999 -466 999 466
<< end >>
