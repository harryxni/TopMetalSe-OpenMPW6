magic
tech sky130A
magscale 1 2
timestamp 1654753044
<< metal1 >>
rect 147045 6626 148460 7016
rect 154020 5336 155975 5706
rect 303400 1370 306810 1570
rect -730 1130 1200 1330
rect 303400 -1630 306810 -1430
rect -730 -1870 1200 -1670
rect 303400 -4630 306810 -4430
rect -730 -4870 1200 -4670
rect 303400 -7630 306810 -7430
rect -730 -7870 1200 -7670
rect 303400 -10630 306810 -10430
rect -730 -10870 1200 -10670
rect 303400 -13630 306810 -13430
rect -730 -13870 1200 -13670
rect 303400 -16630 306810 -16430
rect -730 -16870 1200 -16670
rect 303400 -19630 306810 -19430
rect -730 -19870 1200 -19670
rect 303400 -22630 306810 -22430
rect -730 -22870 1200 -22670
rect 303400 -25630 306810 -25430
rect -730 -25870 1200 -25670
rect 303400 -28630 306810 -28430
rect -730 -28870 1200 -28670
rect 303400 -31630 306810 -31430
rect -730 -31870 1200 -31670
rect 303400 -34630 306810 -34430
rect -730 -34870 1200 -34670
rect 303400 -37630 306810 -37430
rect -730 -37870 1200 -37670
rect 303400 -40630 306810 -40430
rect -730 -40870 1200 -40670
rect 303400 -43630 306810 -43430
rect -730 -43870 1200 -43670
rect 303400 -46630 306810 -46430
rect -730 -46870 1200 -46670
rect 303400 -49630 306810 -49430
rect -730 -49870 1200 -49670
rect 303400 -52630 306810 -52430
rect -730 -52870 1200 -52670
rect 303400 -55630 306810 -55430
rect -730 -55870 1200 -55670
rect 303400 -58630 306810 -58430
rect -730 -58870 1200 -58670
rect 303400 -61630 306810 -61430
rect -730 -61870 1200 -61670
rect 303400 -64630 306810 -64430
rect -730 -64870 1200 -64670
rect 303400 -67630 306810 -67430
rect -730 -67870 1200 -67670
rect 303400 -70630 306810 -70430
rect -730 -70870 1200 -70670
rect 303400 -73630 306810 -73430
rect -730 -73870 1200 -73670
rect 303400 -76630 306810 -76430
rect -730 -76870 1200 -76670
rect 303400 -79630 306810 -79430
rect -730 -79870 1200 -79670
rect 303400 -82630 306810 -82430
rect -730 -82870 1200 -82670
rect 303400 -85630 306810 -85430
rect -730 -85870 1200 -85670
rect 303400 -88630 306810 -88430
rect -730 -88870 1200 -88670
rect 303400 -91630 306810 -91430
rect -730 -91870 1200 -91670
rect 303400 -94630 306810 -94430
rect -730 -94870 1200 -94670
rect 303400 -97630 306810 -97430
rect -730 -97870 1200 -97670
rect 303400 -100630 306810 -100430
rect -730 -100870 1200 -100670
rect 303400 -103630 306810 -103430
rect -730 -103870 1200 -103670
rect 303400 -106630 306810 -106430
rect -730 -106870 1200 -106670
rect 303400 -109630 306810 -109430
rect -730 -109870 1200 -109670
rect 303400 -112630 306810 -112430
rect -730 -112870 1200 -112670
rect 303400 -115630 306810 -115430
rect -730 -115870 1200 -115670
rect 303400 -118630 306810 -118430
rect -730 -118870 1200 -118670
rect 303400 -121630 306810 -121430
rect -730 -121870 1200 -121670
rect 303400 -124630 306810 -124430
rect -730 -124870 1200 -124670
rect 303400 -127630 306810 -127430
rect -730 -127870 1200 -127670
rect 303400 -130630 306810 -130430
rect -730 -130870 1200 -130670
rect 303400 -133630 306810 -133430
rect -730 -133870 1200 -133670
rect 303400 -136630 306810 -136430
rect -730 -136870 1200 -136670
rect 303400 -139630 306810 -139430
rect -730 -139870 1200 -139670
rect 303400 -142630 306810 -142430
rect -730 -142870 1200 -142670
rect 303400 -145630 306810 -145430
rect -730 -145870 1200 -145670
rect 303400 -148630 306810 -148430
rect -730 -148870 1200 -148670
rect 303400 -151630 306810 -151430
rect -730 -151870 1200 -151670
rect 303400 -154630 306810 -154430
rect -730 -154870 1200 -154670
rect 303400 -157630 306810 -157430
rect -730 -157870 1200 -157670
rect 303400 -160630 306810 -160430
rect -730 -160870 1200 -160670
rect 303400 -163630 306810 -163430
rect -730 -163870 1200 -163670
rect 303400 -166630 306810 -166430
rect -730 -166870 1200 -166670
rect 303400 -169630 306810 -169430
rect -730 -169870 1200 -169670
rect 303400 -172630 306810 -172430
rect -730 -172870 1200 -172670
rect 303400 -175630 306810 -175430
rect -730 -175870 1200 -175670
rect 303400 -178630 306810 -178430
rect -730 -178870 1200 -178670
rect 303400 -181630 306810 -181430
rect -730 -181870 1200 -181670
rect 303400 -184630 306810 -184430
rect -730 -184870 1200 -184670
rect 303400 -187630 306810 -187430
rect -730 -187870 1200 -187670
rect 303400 -190630 306810 -190430
rect -730 -190870 1200 -190670
rect 303400 -193630 306810 -193430
rect -730 -193870 1200 -193670
rect 303400 -196630 306810 -196430
rect -730 -196870 1200 -196670
rect 303400 -199630 306810 -199430
rect -730 -199870 1200 -199670
rect 303400 -202630 306810 -202430
rect -730 -202870 1200 -202670
rect 303400 -205630 306810 -205430
rect -730 -205870 1200 -205670
rect 303400 -208630 306810 -208430
rect -730 -208870 1200 -208670
rect 303400 -211630 306810 -211430
rect -730 -211870 1200 -211670
rect 303400 -214630 306810 -214430
rect -730 -214870 1200 -214670
rect 303400 -217630 306810 -217430
rect -730 -217870 1200 -217670
rect 303400 -220630 306810 -220430
rect -730 -220870 1200 -220670
rect 303400 -223630 306810 -223430
rect -730 -223870 1200 -223670
rect 303400 -226630 306810 -226430
rect -730 -226870 1200 -226670
rect 303400 -229630 306810 -229430
rect -730 -229870 1200 -229670
rect 303400 -232630 306810 -232430
rect -730 -232870 1200 -232670
rect 303400 -235630 306810 -235430
rect -730 -235870 1200 -235670
rect 303400 -238630 306810 -238430
rect -730 -238870 1200 -238670
rect 303400 -241630 306810 -241430
rect -730 -241870 1200 -241670
rect 303400 -244630 306810 -244430
rect -730 -244870 1200 -244670
rect 303400 -247630 306810 -247430
rect -730 -247870 1200 -247670
rect 303400 -250630 306810 -250430
rect -730 -250870 1200 -250670
rect 303400 -253630 306810 -253430
rect -730 -253870 1200 -253670
rect 303400 -256630 306810 -256430
rect -730 -256870 1200 -256670
rect 303400 -259630 306810 -259430
rect -730 -259870 1200 -259670
rect 303400 -262630 306810 -262430
rect -730 -262870 1200 -262670
rect 303400 -265630 306810 -265430
rect -730 -265870 1200 -265670
rect 303400 -268630 306810 -268430
rect -730 -268870 1200 -268670
rect 303400 -271630 306810 -271430
rect -730 -271870 1200 -271670
rect 303400 -274630 306810 -274430
rect -730 -274870 1200 -274670
rect 303400 -277630 306810 -277430
rect -730 -277870 1200 -277670
rect 303400 -280630 306810 -280430
rect -730 -280870 1200 -280670
rect 303400 -283630 306810 -283430
rect -730 -283870 1200 -283670
rect 334985 -285211 335905 -284921
rect 303400 -286630 306810 -286430
rect -730 -286870 1200 -286670
rect 303400 -289630 306810 -289430
rect -730 -289870 1200 -289670
rect 303400 -292630 306810 -292430
rect -730 -292870 1200 -292670
rect 303400 -295630 306810 -295430
rect -730 -295870 1200 -295670
rect 334860 -298061 335870 -297761
rect 303400 -298630 306810 -298430
rect -730 -298870 1200 -298670
<< metal2 >>
rect 149300 3585 149390 5091
rect 2250 3475 149390 3585
rect 2250 2435 2360 3475
rect 147975 3465 149390 3475
rect 149810 2635 149900 5101
rect 152250 3670 152360 5141
rect 154250 4285 154360 5141
rect 305310 4285 305480 4300
rect 154250 4115 305480 4285
rect 152250 3496 152360 3505
rect -265 1950 125 2060
rect 305310 -285550 305480 4115
rect 305310 -285720 307605 -285550
rect 307435 -286430 307605 -285720
rect 307435 -286600 307860 -286430
rect 307435 -286605 307605 -286600
rect 304781 -292906 305029 -292880
rect 308336 -292906 308584 -292626
rect 304781 -293154 308584 -292906
rect 304781 -299300 305029 -293154
rect 303570 -299500 305030 -299300
<< via2 >>
rect 152250 3505 152360 3670
<< metal3 >>
rect 149050 3945 149140 5090
rect 1800 3855 149140 3945
rect 1800 3435 1890 3855
rect 149050 3850 149140 3855
rect 304505 3675 304675 3690
rect 152240 3670 304675 3675
rect 152240 3505 152250 3670
rect 152360 3505 304675 3670
rect 152245 3500 152365 3505
rect 304505 -296731 304675 3505
rect 304505 -296901 306255 -296731
<< metal4 >>
rect -265 2150 110 2260
rect 334040 -289661 336790 -288801
rect 2520 -300385 2630 -299885
use bias  bias_0
timestamp 1654639008
transform 1 0 147210 0 1 7236
box 790 -2236 7180 -220
use opamp_wrapper  opamp_wrapper_0
timestamp 1654750071
transform 1 0 310080 0 1 -296491
box -2280 -1640 26995 13665
use pixel_array100x100  pixel_array100x100_0
timestamp 1654753044
transform 1 0 3000 0 1 -1400
box -3000 -298600 300740 5750
<< labels >>
rlabel metal1 335570 -298061 335870 -297761 1 GND
port 1 n
rlabel metal1 335615 -285211 335905 -284921 1 VDD
port 2 n
rlabel metal4 335930 -289661 336790 -288801 1 AOUT
port 3 n
rlabel metal1 147045 6626 147435 7016 1 VDD
port 2 n
rlabel metal1 155605 5336 155975 5706 1 GND
port 1 n
rlabel metal4 -265 2150 -155 2260 1 VBIAS
port 4 n
rlabel metal2 -265 1950 -155 2060 1 VREF
port 5 n
rlabel metal4 2520 -300385 2630 -300275 1 CSA_VREF
port 6 n
<< end >>
