VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pixel_array#0
  CLASS BLOCK ;
  FOREIGN pixel_array#0 ;
  ORIGIN 15.000 38.000 ;
  SIZE 63.700 BY 63.000 ;
  PIN VBIAS
    ANTENNAGATEAREA 14.400000 ;
    PORT
      LAYER li1 ;
        RECT 2.850 10.750 3.100 11.200 ;
        RECT 17.850 10.750 18.100 11.200 ;
        RECT 32.850 10.750 33.100 11.200 ;
        RECT 2.700 10.250 3.100 10.750 ;
        RECT 17.700 10.250 18.100 10.750 ;
        RECT 32.700 10.250 33.100 10.750 ;
        RECT 2.850 -4.250 3.100 -3.800 ;
        RECT 17.850 -4.250 18.100 -3.800 ;
        RECT 32.850 -4.250 33.100 -3.800 ;
        RECT 2.700 -4.750 3.100 -4.250 ;
        RECT 17.700 -4.750 18.100 -4.250 ;
        RECT 32.700 -4.750 33.100 -4.250 ;
        RECT 2.850 -19.250 3.100 -18.800 ;
        RECT 17.850 -19.250 18.100 -18.800 ;
        RECT 32.850 -19.250 33.100 -18.800 ;
        RECT 2.700 -19.750 3.100 -19.250 ;
        RECT 17.700 -19.750 18.100 -19.250 ;
        RECT 32.700 -19.750 33.100 -19.250 ;
      LAYER mcon ;
        RECT 2.890 10.915 3.060 11.085 ;
        RECT 17.890 10.915 18.060 11.085 ;
        RECT 32.890 10.915 33.060 11.085 ;
        RECT 2.890 -4.085 3.060 -3.915 ;
        RECT 17.890 -4.085 18.060 -3.915 ;
        RECT 32.890 -4.085 33.060 -3.915 ;
        RECT 2.890 -19.085 3.060 -18.915 ;
        RECT 17.890 -19.085 18.060 -18.915 ;
        RECT 32.890 -19.085 33.060 -18.915 ;
      LAYER met1 ;
        RECT 2.400 11.200 3.150 11.550 ;
        RECT 17.400 11.200 18.150 11.550 ;
        RECT 32.400 11.200 33.150 11.550 ;
        RECT 2.800 10.750 3.150 11.200 ;
        RECT 17.800 10.750 18.150 11.200 ;
        RECT 32.800 10.750 33.150 11.200 ;
        RECT 2.850 10.450 3.100 10.750 ;
        RECT 17.850 10.450 18.100 10.750 ;
        RECT 32.850 10.450 33.100 10.750 ;
        RECT 2.400 -3.800 3.150 -3.450 ;
        RECT 17.400 -3.800 18.150 -3.450 ;
        RECT 32.400 -3.800 33.150 -3.450 ;
        RECT 2.800 -4.250 3.150 -3.800 ;
        RECT 17.800 -4.250 18.150 -3.800 ;
        RECT 32.800 -4.250 33.150 -3.800 ;
        RECT 2.850 -4.550 3.100 -4.250 ;
        RECT 17.850 -4.550 18.100 -4.250 ;
        RECT 32.850 -4.550 33.100 -4.250 ;
        RECT 2.400 -18.800 3.150 -18.450 ;
        RECT 17.400 -18.800 18.150 -18.450 ;
        RECT 32.400 -18.800 33.150 -18.450 ;
        RECT 2.800 -19.250 3.150 -18.800 ;
        RECT 17.800 -19.250 18.150 -18.800 ;
        RECT 32.800 -19.250 33.150 -18.800 ;
        RECT 2.850 -19.550 3.100 -19.250 ;
        RECT 17.850 -19.550 18.100 -19.250 ;
        RECT 32.850 -19.550 33.100 -19.250 ;
      LAYER via ;
        RECT 2.495 11.270 2.755 11.530 ;
        RECT 17.495 11.270 17.755 11.530 ;
        RECT 32.495 11.270 32.755 11.530 ;
        RECT 2.495 -3.730 2.755 -3.470 ;
        RECT 17.495 -3.730 17.755 -3.470 ;
        RECT 32.495 -3.730 32.755 -3.470 ;
        RECT 2.495 -18.730 2.755 -18.470 ;
        RECT 17.495 -18.730 17.755 -18.470 ;
        RECT 32.495 -18.730 32.755 -18.470 ;
      LAYER met2 ;
        RECT 2.400 17.750 2.950 18.300 ;
        RECT 17.400 17.750 17.950 18.300 ;
        RECT 32.400 17.750 32.950 18.300 ;
        RECT 2.500 11.550 2.850 17.750 ;
        RECT 17.500 11.550 17.850 17.750 ;
        RECT 32.500 11.550 32.850 17.750 ;
        RECT 2.400 11.200 2.900 11.550 ;
        RECT 17.400 11.200 17.900 11.550 ;
        RECT 32.400 11.200 32.900 11.550 ;
        RECT 2.500 -3.450 2.850 11.200 ;
        RECT 17.500 -3.450 17.850 11.200 ;
        RECT 32.500 -3.450 32.850 11.200 ;
        RECT 2.400 -3.800 2.900 -3.450 ;
        RECT 17.400 -3.800 17.900 -3.450 ;
        RECT 32.400 -3.800 32.900 -3.450 ;
        RECT 2.500 -18.450 2.850 -3.800 ;
        RECT 17.500 -18.450 17.850 -3.800 ;
        RECT 32.500 -18.450 32.850 -3.800 ;
        RECT 2.400 -18.800 2.900 -18.450 ;
        RECT 17.400 -18.800 17.900 -18.450 ;
        RECT 32.400 -18.800 32.900 -18.450 ;
        RECT 2.500 -30.000 2.850 -18.800 ;
        RECT 17.500 -30.000 17.850 -18.800 ;
        RECT 32.500 -30.000 32.850 -18.800 ;
      LAYER via2 ;
        RECT 2.535 17.885 2.815 18.165 ;
        RECT 17.535 17.885 17.815 18.165 ;
        RECT 32.535 17.885 32.815 18.165 ;
      LAYER met3 ;
        RECT 2.400 17.750 2.950 18.300 ;
        RECT 17.400 17.750 17.950 18.300 ;
        RECT 32.400 17.750 32.950 18.300 ;
      LAYER via3 ;
        RECT 2.515 17.865 2.835 18.185 ;
        RECT 17.515 17.865 17.835 18.185 ;
        RECT 32.515 17.865 32.835 18.185 ;
      LAYER met4 ;
        RECT -15.000 17.750 41.000 18.300 ;
    END
  END VBIAS
  PIN VREF
    ANTENNAGATEAREA 9.450000 ;
    PORT
      LAYER li1 ;
        RECT 0.250 2.000 0.700 2.750 ;
        RECT 15.250 2.000 15.700 2.750 ;
        RECT 30.250 2.000 30.700 2.750 ;
        RECT 0.250 -13.000 0.700 -12.250 ;
        RECT 15.250 -13.000 15.700 -12.250 ;
        RECT 30.250 -13.000 30.700 -12.250 ;
        RECT 0.250 -28.000 0.700 -27.250 ;
        RECT 15.250 -28.000 15.700 -27.250 ;
        RECT 30.250 -28.000 30.700 -27.250 ;
      LAYER mcon ;
        RECT 0.390 2.540 0.560 2.710 ;
        RECT 15.390 2.540 15.560 2.710 ;
        RECT 30.390 2.540 30.560 2.710 ;
        RECT 0.390 -12.460 0.560 -12.290 ;
        RECT 15.390 -12.460 15.560 -12.290 ;
        RECT 30.390 -12.460 30.560 -12.290 ;
        RECT 0.390 -27.460 0.560 -27.290 ;
        RECT 15.390 -27.460 15.560 -27.290 ;
        RECT 30.390 -27.460 30.560 -27.290 ;
      LAYER met1 ;
        RECT -8.850 16.750 40.000 17.300 ;
        RECT 0.250 2.450 0.700 3.200 ;
        RECT 15.250 2.450 15.700 3.200 ;
        RECT 30.250 2.450 30.700 3.200 ;
        RECT 0.250 -12.550 0.700 -11.800 ;
        RECT 15.250 -12.550 15.700 -11.800 ;
        RECT 30.250 -12.550 30.700 -11.800 ;
        RECT 0.250 -27.550 0.700 -26.800 ;
        RECT 15.250 -27.550 15.700 -26.800 ;
        RECT 30.250 -27.550 30.700 -26.800 ;
      LAYER via ;
        RECT -8.725 16.895 -8.465 17.155 ;
        RECT -8.405 16.895 -8.145 17.155 ;
        RECT -8.085 16.895 -7.825 17.155 ;
        RECT -7.765 16.895 -7.505 17.155 ;
        RECT -7.445 16.895 -7.185 17.155 ;
        RECT -7.125 16.895 -6.865 17.155 ;
        RECT -6.805 16.895 -6.545 17.155 ;
        RECT -6.485 16.895 -6.225 17.155 ;
        RECT -6.165 16.895 -5.905 17.155 ;
        RECT -5.845 16.895 -5.585 17.155 ;
        RECT -5.525 16.895 -5.265 17.155 ;
        RECT -5.205 16.895 -4.945 17.155 ;
        RECT -4.885 16.895 -4.625 17.155 ;
        RECT 0.345 16.895 0.605 17.155 ;
        RECT 15.345 16.895 15.605 17.155 ;
        RECT 30.345 16.895 30.605 17.155 ;
        RECT 0.345 2.845 0.605 3.105 ;
        RECT 15.345 2.845 15.605 3.105 ;
        RECT 30.345 2.845 30.605 3.105 ;
        RECT 0.345 -12.155 0.605 -11.895 ;
        RECT 15.345 -12.155 15.605 -11.895 ;
        RECT 30.345 -12.155 30.605 -11.895 ;
        RECT 0.345 -27.155 0.605 -26.895 ;
        RECT 15.345 -27.155 15.605 -26.895 ;
        RECT 30.345 -27.155 30.605 -26.895 ;
      LAYER met2 ;
        RECT 0.300 17.300 0.650 18.000 ;
        RECT 15.300 17.300 15.650 18.000 ;
        RECT 30.300 17.300 30.650 18.000 ;
        RECT -15.000 16.750 -4.450 17.300 ;
        RECT 0.200 16.750 0.750 17.300 ;
        RECT 15.200 16.750 15.750 17.300 ;
        RECT 30.200 16.750 30.750 17.300 ;
        RECT 0.300 -30.000 0.650 16.750 ;
        RECT 15.300 -30.000 15.650 16.750 ;
        RECT 30.300 -30.000 30.650 16.750 ;
    END
  END VREF
  PIN NB2
    ANTENNAGATEAREA 10.349999 ;
    PORT
      LAYER li1 ;
        RECT 5.050 8.450 5.650 9.300 ;
        RECT 20.050 8.450 20.650 9.300 ;
        RECT 35.050 8.450 35.650 9.300 ;
        RECT 5.100 8.050 5.650 8.450 ;
        RECT 20.100 8.050 20.650 8.450 ;
        RECT 35.100 8.050 35.650 8.450 ;
        RECT 5.050 -6.550 5.650 -5.700 ;
        RECT 20.050 -6.550 20.650 -5.700 ;
        RECT 35.050 -6.550 35.650 -5.700 ;
        RECT 5.100 -6.950 5.650 -6.550 ;
        RECT 20.100 -6.950 20.650 -6.550 ;
        RECT 35.100 -6.950 35.650 -6.550 ;
        RECT 5.050 -21.550 5.650 -20.700 ;
        RECT 20.050 -21.550 20.650 -20.700 ;
        RECT 35.050 -21.550 35.650 -20.700 ;
        RECT 5.100 -21.950 5.650 -21.550 ;
        RECT 20.100 -21.950 20.650 -21.550 ;
        RECT 35.100 -21.950 35.650 -21.550 ;
      LAYER mcon ;
        RECT 5.290 8.140 5.460 8.310 ;
        RECT 20.290 8.140 20.460 8.310 ;
        RECT 35.290 8.140 35.460 8.310 ;
        RECT 5.290 -6.860 5.460 -6.690 ;
        RECT 20.290 -6.860 20.460 -6.690 ;
        RECT 35.290 -6.860 35.460 -6.690 ;
        RECT 5.290 -21.860 5.460 -21.690 ;
        RECT 20.290 -21.860 20.460 -21.690 ;
        RECT 35.290 -21.860 35.460 -21.690 ;
      LAYER met1 ;
        RECT 4.950 7.750 5.650 8.450 ;
        RECT 19.950 7.750 20.650 8.450 ;
        RECT 34.950 7.750 35.650 8.450 ;
        RECT 4.950 -7.250 5.650 -6.550 ;
        RECT 19.950 -7.250 20.650 -6.550 ;
        RECT 34.950 -7.250 35.650 -6.550 ;
        RECT 4.950 -22.250 5.650 -21.550 ;
        RECT 19.950 -22.250 20.650 -21.550 ;
        RECT 34.950 -22.250 35.650 -21.550 ;
      LAYER via ;
        RECT 5.170 7.820 5.430 8.080 ;
        RECT 20.170 7.820 20.430 8.080 ;
        RECT 35.170 7.820 35.430 8.080 ;
        RECT 5.170 -7.180 5.430 -6.920 ;
        RECT 20.170 -7.180 20.430 -6.920 ;
        RECT 35.170 -7.180 35.430 -6.920 ;
        RECT 5.170 -22.180 5.430 -21.920 ;
        RECT 20.170 -22.180 20.430 -21.920 ;
        RECT 35.170 -22.180 35.430 -21.920 ;
      LAYER met2 ;
        RECT 0.000 20.200 45.000 20.750 ;
        RECT 5.100 15.000 5.450 20.200 ;
        RECT 20.100 15.000 20.450 20.200 ;
        RECT 35.100 15.000 35.450 20.200 ;
        RECT 5.100 -30.000 5.500 15.000 ;
        RECT 20.100 -30.000 20.500 15.000 ;
        RECT 35.100 -30.000 35.500 15.000 ;
    END
  END NB2
  PIN VDD
    ANTENNADIFFAREA 19.799999 ;
    PORT
      LAYER nwell ;
        RECT 0.000 11.600 45.000 15.000 ;
        RECT 0.000 -3.400 45.000 0.000 ;
        RECT 0.000 -18.400 45.000 -15.000 ;
      LAYER li1 ;
        RECT 5.450 14.550 5.950 14.850 ;
        RECT 14.250 14.800 14.450 14.850 ;
        RECT 14.150 14.600 14.550 14.800 ;
        RECT 5.100 13.550 6.300 14.550 ;
        RECT 14.250 13.400 14.450 14.600 ;
        RECT 20.450 14.550 20.950 14.850 ;
        RECT 29.250 14.800 29.450 14.850 ;
        RECT 29.150 14.600 29.550 14.800 ;
        RECT 20.100 13.550 21.300 14.550 ;
        RECT 29.250 13.400 29.450 14.600 ;
        RECT 35.450 14.550 35.950 14.850 ;
        RECT 44.250 14.800 44.450 14.850 ;
        RECT 44.150 14.600 44.550 14.800 ;
        RECT 35.100 13.550 36.300 14.550 ;
        RECT 44.250 13.400 44.450 14.600 ;
        RECT 4.250 12.050 4.600 12.250 ;
        RECT 19.250 12.050 19.600 12.250 ;
        RECT 34.250 12.050 34.600 12.250 ;
        RECT 4.250 11.250 4.450 12.050 ;
        RECT 19.250 11.250 19.450 12.050 ;
        RECT 34.250 11.250 34.450 12.050 ;
        RECT 4.100 11.000 5.000 11.250 ;
        RECT 19.100 11.000 20.000 11.250 ;
        RECT 34.100 11.000 35.000 11.250 ;
        RECT 9.800 10.400 10.150 10.950 ;
        RECT 24.800 10.400 25.150 10.950 ;
        RECT 39.800 10.400 40.150 10.950 ;
        RECT 9.800 10.100 10.700 10.400 ;
        RECT 24.800 10.100 25.700 10.400 ;
        RECT 39.800 10.100 40.700 10.400 ;
        RECT 5.450 -0.450 5.950 -0.150 ;
        RECT 14.250 -0.200 14.450 -0.150 ;
        RECT 14.150 -0.400 14.550 -0.200 ;
        RECT 5.100 -1.450 6.300 -0.450 ;
        RECT 14.250 -1.600 14.450 -0.400 ;
        RECT 20.450 -0.450 20.950 -0.150 ;
        RECT 29.250 -0.200 29.450 -0.150 ;
        RECT 29.150 -0.400 29.550 -0.200 ;
        RECT 20.100 -1.450 21.300 -0.450 ;
        RECT 29.250 -1.600 29.450 -0.400 ;
        RECT 35.450 -0.450 35.950 -0.150 ;
        RECT 44.250 -0.200 44.450 -0.150 ;
        RECT 44.150 -0.400 44.550 -0.200 ;
        RECT 35.100 -1.450 36.300 -0.450 ;
        RECT 44.250 -1.600 44.450 -0.400 ;
        RECT 4.250 -2.950 4.600 -2.750 ;
        RECT 19.250 -2.950 19.600 -2.750 ;
        RECT 34.250 -2.950 34.600 -2.750 ;
        RECT 4.250 -3.750 4.450 -2.950 ;
        RECT 19.250 -3.750 19.450 -2.950 ;
        RECT 34.250 -3.750 34.450 -2.950 ;
        RECT 4.100 -4.000 5.000 -3.750 ;
        RECT 19.100 -4.000 20.000 -3.750 ;
        RECT 34.100 -4.000 35.000 -3.750 ;
        RECT 9.800 -4.600 10.150 -4.050 ;
        RECT 24.800 -4.600 25.150 -4.050 ;
        RECT 39.800 -4.600 40.150 -4.050 ;
        RECT 9.800 -4.900 10.700 -4.600 ;
        RECT 24.800 -4.900 25.700 -4.600 ;
        RECT 39.800 -4.900 40.700 -4.600 ;
        RECT 5.450 -15.450 5.950 -15.150 ;
        RECT 14.250 -15.200 14.450 -15.150 ;
        RECT 14.150 -15.400 14.550 -15.200 ;
        RECT 5.100 -16.450 6.300 -15.450 ;
        RECT 14.250 -16.600 14.450 -15.400 ;
        RECT 20.450 -15.450 20.950 -15.150 ;
        RECT 29.250 -15.200 29.450 -15.150 ;
        RECT 29.150 -15.400 29.550 -15.200 ;
        RECT 20.100 -16.450 21.300 -15.450 ;
        RECT 29.250 -16.600 29.450 -15.400 ;
        RECT 35.450 -15.450 35.950 -15.150 ;
        RECT 44.250 -15.200 44.450 -15.150 ;
        RECT 44.150 -15.400 44.550 -15.200 ;
        RECT 35.100 -16.450 36.300 -15.450 ;
        RECT 44.250 -16.600 44.450 -15.400 ;
        RECT 4.250 -17.950 4.600 -17.750 ;
        RECT 19.250 -17.950 19.600 -17.750 ;
        RECT 34.250 -17.950 34.600 -17.750 ;
        RECT 4.250 -18.750 4.450 -17.950 ;
        RECT 19.250 -18.750 19.450 -17.950 ;
        RECT 34.250 -18.750 34.450 -17.950 ;
        RECT 4.100 -19.000 5.000 -18.750 ;
        RECT 19.100 -19.000 20.000 -18.750 ;
        RECT 34.100 -19.000 35.000 -18.750 ;
        RECT 9.800 -19.600 10.150 -19.050 ;
        RECT 24.800 -19.600 25.150 -19.050 ;
        RECT 39.800 -19.600 40.150 -19.050 ;
        RECT 9.800 -19.900 10.700 -19.600 ;
        RECT 24.800 -19.900 25.700 -19.600 ;
        RECT 39.800 -19.900 40.700 -19.600 ;
      LAYER mcon ;
        RECT 5.615 14.590 5.785 14.760 ;
        RECT 14.265 14.615 14.435 14.785 ;
        RECT 20.615 14.590 20.785 14.760 ;
        RECT 29.265 14.615 29.435 14.785 ;
        RECT 35.615 14.590 35.785 14.760 ;
        RECT 44.265 14.615 44.435 14.785 ;
        RECT 4.340 12.065 4.510 12.235 ;
        RECT 19.340 12.065 19.510 12.235 ;
        RECT 34.340 12.065 34.510 12.235 ;
        RECT 9.890 10.670 10.060 10.840 ;
        RECT 9.890 10.310 10.060 10.480 ;
        RECT 24.890 10.670 25.060 10.840 ;
        RECT 24.890 10.310 25.060 10.480 ;
        RECT 39.890 10.670 40.060 10.840 ;
        RECT 39.890 10.310 40.060 10.480 ;
        RECT 5.615 -0.410 5.785 -0.240 ;
        RECT 14.265 -0.385 14.435 -0.215 ;
        RECT 20.615 -0.410 20.785 -0.240 ;
        RECT 29.265 -0.385 29.435 -0.215 ;
        RECT 35.615 -0.410 35.785 -0.240 ;
        RECT 44.265 -0.385 44.435 -0.215 ;
        RECT 4.340 -2.935 4.510 -2.765 ;
        RECT 19.340 -2.935 19.510 -2.765 ;
        RECT 34.340 -2.935 34.510 -2.765 ;
        RECT 9.890 -4.330 10.060 -4.160 ;
        RECT 9.890 -4.690 10.060 -4.520 ;
        RECT 24.890 -4.330 25.060 -4.160 ;
        RECT 24.890 -4.690 25.060 -4.520 ;
        RECT 39.890 -4.330 40.060 -4.160 ;
        RECT 39.890 -4.690 40.060 -4.520 ;
        RECT 5.615 -15.410 5.785 -15.240 ;
        RECT 14.265 -15.385 14.435 -15.215 ;
        RECT 20.615 -15.410 20.785 -15.240 ;
        RECT 29.265 -15.385 29.435 -15.215 ;
        RECT 35.615 -15.410 35.785 -15.240 ;
        RECT 44.265 -15.385 44.435 -15.215 ;
        RECT 4.340 -17.935 4.510 -17.765 ;
        RECT 19.340 -17.935 19.510 -17.765 ;
        RECT 34.340 -17.935 34.510 -17.765 ;
        RECT 9.890 -19.330 10.060 -19.160 ;
        RECT 9.890 -19.690 10.060 -19.520 ;
        RECT 24.890 -19.330 25.060 -19.160 ;
        RECT 24.890 -19.690 25.060 -19.520 ;
        RECT 39.890 -19.330 40.060 -19.160 ;
        RECT 39.890 -19.690 40.060 -19.520 ;
      LAYER met1 ;
        RECT -10.000 14.850 -9.000 14.950 ;
        RECT -10.000 14.100 45.000 14.850 ;
        RECT -10.000 -0.150 -9.000 14.100 ;
        RECT 4.550 12.350 5.050 14.100 ;
        RECT 4.150 12.000 5.050 12.350 ;
        RECT 9.800 10.150 10.150 14.100 ;
        RECT 19.550 12.350 20.050 14.100 ;
        RECT 19.150 12.000 20.050 12.350 ;
        RECT 24.800 10.150 25.150 14.100 ;
        RECT 34.550 12.350 35.050 14.100 ;
        RECT 34.150 12.000 35.050 12.350 ;
        RECT 39.800 10.150 40.150 14.100 ;
        RECT -10.000 -0.900 45.000 -0.150 ;
        RECT -10.000 -15.150 -9.000 -0.900 ;
        RECT 4.550 -2.650 5.050 -0.900 ;
        RECT 4.150 -3.000 5.050 -2.650 ;
        RECT 9.800 -4.850 10.150 -0.900 ;
        RECT 19.550 -2.650 20.050 -0.900 ;
        RECT 19.150 -3.000 20.050 -2.650 ;
        RECT 24.800 -4.850 25.150 -0.900 ;
        RECT 34.550 -2.650 35.050 -0.900 ;
        RECT 34.150 -3.000 35.050 -2.650 ;
        RECT 39.800 -4.850 40.150 -0.900 ;
        RECT -10.000 -15.900 45.000 -15.150 ;
        RECT -10.000 -30.000 -9.000 -15.900 ;
        RECT 4.550 -17.650 5.050 -15.900 ;
        RECT 4.150 -18.000 5.050 -17.650 ;
        RECT 9.800 -19.850 10.150 -15.900 ;
        RECT 19.550 -17.650 20.050 -15.900 ;
        RECT 19.150 -18.000 20.050 -17.650 ;
        RECT 24.800 -19.850 25.150 -15.900 ;
        RECT 34.550 -17.650 35.050 -15.900 ;
        RECT 34.150 -18.000 35.050 -17.650 ;
        RECT 39.800 -19.850 40.150 -15.900 ;
    END
  END VDD
  PIN SF_IB
    ANTENNAGATEAREA 9.000000 ;
    PORT
      LAYER li1 ;
        RECT 13.700 12.800 14.600 13.050 ;
        RECT 28.700 12.800 29.600 13.050 ;
        RECT 43.700 12.800 44.600 13.050 ;
        RECT 13.700 -2.200 14.600 -1.950 ;
        RECT 28.700 -2.200 29.600 -1.950 ;
        RECT 43.700 -2.200 44.600 -1.950 ;
        RECT 13.700 -17.200 14.600 -16.950 ;
        RECT 28.700 -17.200 29.600 -16.950 ;
        RECT 43.700 -17.200 44.600 -16.950 ;
      LAYER mcon ;
        RECT 14.415 12.840 14.585 13.010 ;
        RECT 29.415 12.840 29.585 13.010 ;
        RECT 44.415 12.840 44.585 13.010 ;
        RECT 14.415 -2.160 14.585 -1.990 ;
        RECT 29.415 -2.160 29.585 -1.990 ;
        RECT 44.415 -2.160 44.585 -1.990 ;
        RECT 14.415 -17.160 14.585 -16.990 ;
        RECT 29.415 -17.160 29.585 -16.990 ;
        RECT 44.415 -17.160 44.585 -16.990 ;
      LAYER met1 ;
        RECT 14.300 12.750 14.950 13.100 ;
        RECT 29.300 12.750 29.950 13.100 ;
        RECT 44.300 12.750 44.950 13.100 ;
        RECT 14.300 -2.250 14.950 -1.900 ;
        RECT 29.300 -2.250 29.950 -1.900 ;
        RECT 44.300 -2.250 44.950 -1.900 ;
        RECT 14.300 -17.250 14.950 -16.900 ;
        RECT 29.300 -17.250 29.950 -16.900 ;
        RECT 44.300 -17.250 44.950 -16.900 ;
      LAYER via ;
        RECT 14.620 12.795 14.880 13.055 ;
        RECT 29.620 12.795 29.880 13.055 ;
        RECT 44.620 12.795 44.880 13.055 ;
        RECT 14.620 -2.205 14.880 -1.945 ;
        RECT 29.620 -2.205 29.880 -1.945 ;
        RECT 44.620 -2.205 44.880 -1.945 ;
        RECT 14.620 -17.205 14.880 -16.945 ;
        RECT 29.620 -17.205 29.880 -16.945 ;
        RECT 44.620 -17.205 44.880 -16.945 ;
      LAYER met2 ;
        RECT 14.600 12.650 14.900 14.150 ;
        RECT 29.600 12.650 29.900 14.150 ;
        RECT 44.600 12.650 44.900 14.150 ;
        RECT 14.600 -2.350 14.900 -0.850 ;
        RECT 29.600 -2.350 29.900 -0.850 ;
        RECT 44.600 -2.350 44.900 -0.850 ;
        RECT 14.600 -17.350 14.900 -15.850 ;
        RECT 29.600 -17.350 29.900 -15.850 ;
        RECT 44.600 -17.350 44.900 -15.850 ;
      LAYER via2 ;
        RECT 14.610 13.810 14.890 14.090 ;
        RECT 29.610 13.810 29.890 14.090 ;
        RECT 44.610 13.810 44.890 14.090 ;
        RECT 14.610 -1.190 14.890 -0.910 ;
        RECT 29.610 -1.190 29.890 -0.910 ;
        RECT 44.610 -1.190 44.890 -0.910 ;
        RECT 14.610 -16.190 14.890 -15.910 ;
        RECT 29.610 -16.190 29.890 -15.910 ;
        RECT 44.610 -16.190 44.890 -15.910 ;
      LAYER met3 ;
        RECT -6.000 14.200 -5.550 25.000 ;
        RECT -6.000 14.100 1.000 14.200 ;
        RECT 14.550 14.100 14.950 14.150 ;
        RECT 29.550 14.100 29.950 14.150 ;
        RECT 44.550 14.100 44.950 14.150 ;
        RECT -6.000 13.750 45.000 14.100 ;
        RECT -6.000 -0.800 -5.550 13.750 ;
        RECT 14.550 13.700 14.950 13.750 ;
        RECT 29.550 13.700 29.950 13.750 ;
        RECT 44.550 13.700 44.950 13.750 ;
        RECT -6.000 -0.900 1.000 -0.800 ;
        RECT 14.550 -0.900 14.950 -0.850 ;
        RECT 29.550 -0.900 29.950 -0.850 ;
        RECT 44.550 -0.900 44.950 -0.850 ;
        RECT -6.000 -1.250 45.000 -0.900 ;
        RECT -6.000 -15.800 -5.550 -1.250 ;
        RECT 14.550 -1.300 14.950 -1.250 ;
        RECT 29.550 -1.300 29.950 -1.250 ;
        RECT 44.550 -1.300 44.950 -1.250 ;
        RECT -6.000 -15.900 1.000 -15.800 ;
        RECT 14.550 -15.900 14.950 -15.850 ;
        RECT 29.550 -15.900 29.950 -15.850 ;
        RECT 44.550 -15.900 44.950 -15.850 ;
        RECT -6.000 -16.250 45.000 -15.900 ;
        RECT -6.000 -20.000 -5.550 -16.250 ;
        RECT 14.550 -16.300 14.950 -16.250 ;
        RECT 29.550 -16.300 29.950 -16.250 ;
        RECT 44.550 -16.300 44.950 -16.250 ;
    END
  END SF_IB
  PIN CSA_VREF
    ANTENNAGATEAREA 30.240000 ;
    PORT
      LAYER li1 ;
        RECT 13.600 11.350 14.050 11.650 ;
        RECT 28.600 11.350 29.050 11.650 ;
        RECT 43.600 11.350 44.050 11.650 ;
        RECT 13.150 11.100 14.100 11.350 ;
        RECT 28.150 11.100 29.100 11.350 ;
        RECT 43.150 11.100 44.100 11.350 ;
        RECT 13.600 -3.650 14.050 -3.350 ;
        RECT 28.600 -3.650 29.050 -3.350 ;
        RECT 43.600 -3.650 44.050 -3.350 ;
        RECT 13.150 -3.900 14.100 -3.650 ;
        RECT 28.150 -3.900 29.100 -3.650 ;
        RECT 43.150 -3.900 44.100 -3.650 ;
        RECT 13.600 -18.650 14.050 -18.350 ;
        RECT 28.600 -18.650 29.050 -18.350 ;
        RECT 43.600 -18.650 44.050 -18.350 ;
        RECT 13.150 -18.900 14.100 -18.650 ;
        RECT 28.150 -18.900 29.100 -18.650 ;
        RECT 43.150 -18.900 44.100 -18.650 ;
      LAYER mcon ;
        RECT 13.190 11.140 13.360 11.310 ;
        RECT 28.190 11.140 28.360 11.310 ;
        RECT 43.190 11.140 43.360 11.310 ;
        RECT 13.190 -3.860 13.360 -3.690 ;
        RECT 28.190 -3.860 28.360 -3.690 ;
        RECT 43.190 -3.860 43.360 -3.690 ;
        RECT 13.190 -18.860 13.360 -18.690 ;
        RECT 28.190 -18.860 28.360 -18.690 ;
        RECT 43.190 -18.860 43.360 -18.690 ;
      LAYER met1 ;
        RECT 13.050 11.000 13.500 11.500 ;
        RECT 28.050 11.000 28.500 11.500 ;
        RECT 43.050 11.000 43.500 11.500 ;
        RECT 13.050 -4.000 13.500 -3.500 ;
        RECT 28.050 -4.000 28.500 -3.500 ;
        RECT 43.050 -4.000 43.500 -3.500 ;
        RECT 13.050 -19.000 13.500 -18.500 ;
        RECT 28.050 -19.000 28.500 -18.500 ;
        RECT 43.050 -19.000 43.500 -18.500 ;
      LAYER via ;
        RECT 13.145 11.120 13.405 11.380 ;
        RECT 28.145 11.120 28.405 11.380 ;
        RECT 43.145 11.120 43.405 11.380 ;
        RECT 13.145 -3.880 13.405 -3.620 ;
        RECT 28.145 -3.880 28.405 -3.620 ;
        RECT 43.145 -3.880 43.405 -3.620 ;
        RECT 13.145 -18.880 13.405 -18.620 ;
        RECT 28.145 -18.880 28.405 -18.620 ;
        RECT 43.145 -18.880 43.405 -18.620 ;
      LAYER met2 ;
        RECT 13.100 10.950 13.450 12.750 ;
        RECT 28.100 10.950 28.450 12.750 ;
        RECT 43.100 10.950 43.450 12.750 ;
        RECT 13.100 -4.050 13.450 -2.250 ;
        RECT 28.100 -4.050 28.450 -2.250 ;
        RECT 43.100 -4.050 43.450 -2.250 ;
        RECT 13.100 -19.050 13.450 -17.250 ;
        RECT 28.100 -19.050 28.450 -17.250 ;
        RECT 43.100 -19.050 43.450 -17.250 ;
      LAYER via2 ;
        RECT 13.135 12.335 13.415 12.615 ;
        RECT 28.135 12.335 28.415 12.615 ;
        RECT 43.135 12.335 43.415 12.615 ;
        RECT 13.135 -2.665 13.415 -2.385 ;
        RECT 28.135 -2.665 28.415 -2.385 ;
        RECT 43.135 -2.665 43.415 -2.385 ;
        RECT 13.135 -17.665 13.415 -17.385 ;
        RECT 28.135 -17.665 28.415 -17.385 ;
        RECT 43.135 -17.665 43.415 -17.385 ;
      LAYER met3 ;
        RECT -2.400 12.750 -1.850 12.800 ;
        RECT -2.800 12.650 2.600 12.750 ;
        RECT 13.050 12.650 13.500 12.700 ;
        RECT 28.050 12.650 28.500 12.700 ;
        RECT 43.050 12.650 43.500 12.700 ;
        RECT -2.800 12.300 45.800 12.650 ;
        RECT -2.400 12.250 -1.850 12.300 ;
        RECT 13.050 12.250 13.500 12.300 ;
        RECT 28.050 12.250 28.500 12.300 ;
        RECT 43.050 12.250 43.500 12.300 ;
        RECT -2.400 -2.250 -1.850 -2.200 ;
        RECT -2.800 -2.350 2.600 -2.250 ;
        RECT 13.050 -2.350 13.500 -2.300 ;
        RECT 28.050 -2.350 28.500 -2.300 ;
        RECT 43.050 -2.350 43.500 -2.300 ;
        RECT -2.800 -2.700 45.800 -2.350 ;
        RECT -2.400 -2.750 -1.850 -2.700 ;
        RECT 13.050 -2.750 13.500 -2.700 ;
        RECT 28.050 -2.750 28.500 -2.700 ;
        RECT 43.050 -2.750 43.500 -2.700 ;
        RECT -2.400 -17.250 -1.850 -17.200 ;
        RECT -2.800 -17.350 2.600 -17.250 ;
        RECT 13.050 -17.350 13.500 -17.300 ;
        RECT 28.050 -17.350 28.500 -17.300 ;
        RECT 43.050 -17.350 43.500 -17.300 ;
        RECT -2.800 -17.700 45.800 -17.350 ;
        RECT -2.400 -17.750 -1.850 -17.700 ;
        RECT 13.050 -17.750 13.500 -17.700 ;
        RECT 28.050 -17.750 28.500 -17.700 ;
        RECT 43.050 -17.750 43.500 -17.700 ;
      LAYER via3 ;
        RECT -2.285 12.365 -1.965 12.685 ;
        RECT -2.285 -2.635 -1.965 -2.315 ;
        RECT -2.285 -17.635 -1.965 -17.315 ;
      LAYER met4 ;
        RECT -2.400 -38.000 -1.850 13.000 ;
    END
  END CSA_VREF
  PIN NB1
    ANTENNAGATEAREA 10.800000 ;
    PORT
      LAYER li1 ;
        RECT 3.550 1.150 4.000 1.450 ;
        RECT 18.550 1.150 19.000 1.450 ;
        RECT 33.550 1.150 34.000 1.450 ;
        RECT 3.550 0.750 3.900 1.150 ;
        RECT 18.550 0.750 18.900 1.150 ;
        RECT 33.550 0.750 33.900 1.150 ;
        RECT 3.550 -13.850 4.000 -13.550 ;
        RECT 18.550 -13.850 19.000 -13.550 ;
        RECT 33.550 -13.850 34.000 -13.550 ;
        RECT 3.550 -14.250 3.900 -13.850 ;
        RECT 18.550 -14.250 18.900 -13.850 ;
        RECT 33.550 -14.250 33.900 -13.850 ;
        RECT 3.550 -28.850 4.000 -28.550 ;
        RECT 18.550 -28.850 19.000 -28.550 ;
        RECT 33.550 -28.850 34.000 -28.550 ;
        RECT 3.550 -29.250 3.900 -28.850 ;
        RECT 18.550 -29.250 18.900 -28.850 ;
        RECT 33.550 -29.250 33.900 -28.850 ;
      LAYER mcon ;
        RECT 3.690 1.215 3.860 1.385 ;
        RECT 18.690 1.215 18.860 1.385 ;
        RECT 33.690 1.215 33.860 1.385 ;
        RECT 3.690 -13.785 3.860 -13.615 ;
        RECT 18.690 -13.785 18.860 -13.615 ;
        RECT 33.690 -13.785 33.860 -13.615 ;
        RECT 3.690 -28.785 3.860 -28.615 ;
        RECT 18.690 -28.785 18.860 -28.615 ;
        RECT 33.690 -28.785 33.860 -28.615 ;
      LAYER met1 ;
        RECT 3.500 1.150 4.500 1.450 ;
        RECT 18.500 1.150 19.500 1.450 ;
        RECT 33.500 1.150 34.500 1.450 ;
        RECT 3.500 -13.850 4.500 -13.550 ;
        RECT 18.500 -13.850 19.500 -13.550 ;
        RECT 33.500 -13.850 34.500 -13.550 ;
        RECT 3.500 -28.850 4.500 -28.550 ;
        RECT 18.500 -28.850 19.500 -28.550 ;
        RECT 33.500 -28.850 34.500 -28.550 ;
      LAYER via ;
        RECT 4.145 1.170 4.405 1.430 ;
        RECT 19.145 1.170 19.405 1.430 ;
        RECT 34.145 1.170 34.405 1.430 ;
        RECT 4.145 -13.830 4.405 -13.570 ;
        RECT 19.145 -13.830 19.405 -13.570 ;
        RECT 34.145 -13.830 34.405 -13.570 ;
        RECT 4.145 -28.830 4.405 -28.570 ;
        RECT 19.145 -28.830 19.405 -28.570 ;
        RECT 34.145 -28.830 34.405 -28.570 ;
      LAYER met2 ;
        RECT -3.750 -30.000 -3.200 20.000 ;
        RECT 4.100 0.650 4.500 1.500 ;
        RECT 19.100 0.650 19.500 1.500 ;
        RECT 34.100 0.650 34.500 1.500 ;
        RECT 4.100 -14.350 4.500 -13.500 ;
        RECT 19.100 -14.350 19.500 -13.500 ;
        RECT 34.100 -14.350 34.500 -13.500 ;
        RECT 4.100 -29.350 4.500 -28.500 ;
        RECT 19.100 -29.350 19.500 -28.500 ;
        RECT 34.100 -29.350 34.500 -28.500 ;
      LAYER via2 ;
        RECT -3.615 0.835 -3.335 1.115 ;
        RECT 4.160 0.785 4.440 1.065 ;
        RECT 19.160 0.785 19.440 1.065 ;
        RECT 34.160 0.785 34.440 1.065 ;
        RECT -3.615 -14.165 -3.335 -13.885 ;
        RECT 4.160 -14.215 4.440 -13.935 ;
        RECT 19.160 -14.215 19.440 -13.935 ;
        RECT 34.160 -14.215 34.440 -13.935 ;
        RECT -3.615 -29.165 -3.335 -28.885 ;
        RECT 4.160 -29.215 4.440 -28.935 ;
        RECT 19.160 -29.215 19.440 -28.935 ;
        RECT 34.160 -29.215 34.440 -28.935 ;
      LAYER met3 ;
        RECT -3.800 1.150 0.200 1.250 ;
        RECT -3.800 0.800 45.000 1.150 ;
        RECT -3.750 0.700 -3.200 0.800 ;
        RECT 4.100 0.700 4.500 0.800 ;
        RECT 19.100 0.700 19.500 0.800 ;
        RECT 34.100 0.700 34.500 0.800 ;
        RECT -3.800 -13.850 0.200 -13.750 ;
        RECT -3.800 -14.200 45.000 -13.850 ;
        RECT -3.750 -14.300 -3.200 -14.200 ;
        RECT 4.100 -14.300 4.500 -14.200 ;
        RECT 19.100 -14.300 19.500 -14.200 ;
        RECT 34.100 -14.300 34.500 -14.200 ;
        RECT -3.800 -28.850 0.200 -28.750 ;
        RECT -3.800 -29.200 45.000 -28.850 ;
        RECT -3.750 -29.300 -3.200 -29.200 ;
        RECT 4.100 -29.300 4.500 -29.200 ;
        RECT 19.100 -29.300 19.500 -29.200 ;
        RECT 34.100 -29.300 34.500 -29.200 ;
    END
  END NB1
  PIN GND
    ANTENNADIFFAREA 15.750000 ;
    PORT
      LAYER pwell ;
        RECT 0.170 9.620 2.730 11.380 ;
        RECT 15.170 9.620 17.730 11.380 ;
        RECT 30.170 9.620 32.730 11.380 ;
        RECT 0.720 2.270 2.180 9.620 ;
        RECT 15.720 2.270 17.180 9.620 ;
        RECT 30.720 2.270 32.180 9.620 ;
        RECT 1.120 1.880 2.180 2.270 ;
        RECT 16.120 1.880 17.180 2.270 ;
        RECT 31.120 1.880 32.180 2.270 ;
        RECT 1.120 0.420 3.480 1.880 ;
        RECT 16.120 0.420 18.480 1.880 ;
        RECT 31.120 0.420 33.480 1.880 ;
        RECT 0.170 -5.380 2.730 -3.620 ;
        RECT 15.170 -5.380 17.730 -3.620 ;
        RECT 30.170 -5.380 32.730 -3.620 ;
        RECT 0.720 -12.730 2.180 -5.380 ;
        RECT 15.720 -12.730 17.180 -5.380 ;
        RECT 30.720 -12.730 32.180 -5.380 ;
        RECT 1.120 -13.120 2.180 -12.730 ;
        RECT 16.120 -13.120 17.180 -12.730 ;
        RECT 31.120 -13.120 32.180 -12.730 ;
        RECT 1.120 -14.580 3.480 -13.120 ;
        RECT 16.120 -14.580 18.480 -13.120 ;
        RECT 31.120 -14.580 33.480 -13.120 ;
        RECT 0.170 -20.380 2.730 -18.620 ;
        RECT 15.170 -20.380 17.730 -18.620 ;
        RECT 30.170 -20.380 32.730 -18.620 ;
        RECT 0.720 -27.730 2.180 -20.380 ;
        RECT 15.720 -27.730 17.180 -20.380 ;
        RECT 30.720 -27.730 32.180 -20.380 ;
        RECT 1.120 -28.120 2.180 -27.730 ;
        RECT 16.120 -28.120 17.180 -27.730 ;
        RECT 31.120 -28.120 32.180 -27.730 ;
        RECT 1.120 -29.580 3.480 -28.120 ;
        RECT 16.120 -29.580 18.480 -28.120 ;
        RECT 31.120 -29.580 33.480 -28.120 ;
      LAYER li1 ;
        RECT 11.150 13.400 11.550 14.400 ;
        RECT 26.150 13.400 26.550 14.400 ;
        RECT 41.150 13.400 41.550 14.400 ;
        RECT 11.150 12.250 11.400 13.400 ;
        RECT 26.150 12.250 26.400 13.400 ;
        RECT 41.150 12.250 41.400 13.400 ;
        RECT 10.350 11.900 11.400 12.250 ;
        RECT 25.350 11.900 26.400 12.250 ;
        RECT 40.350 11.900 41.400 12.250 ;
        RECT 4.000 7.800 4.900 8.250 ;
        RECT 19.000 7.800 19.900 8.250 ;
        RECT 34.000 7.800 34.900 8.250 ;
        RECT 4.000 5.600 4.500 7.800 ;
        RECT 19.000 5.600 19.500 7.800 ;
        RECT 34.000 5.600 34.500 7.800 ;
        RECT 2.650 0.550 3.350 1.750 ;
        RECT 17.650 0.550 18.350 1.750 ;
        RECT 32.650 0.550 33.350 1.750 ;
        RECT 2.900 0.150 3.150 0.550 ;
        RECT 17.900 0.150 18.150 0.550 ;
        RECT 32.900 0.150 33.150 0.550 ;
        RECT 11.150 -1.600 11.550 -0.600 ;
        RECT 26.150 -1.600 26.550 -0.600 ;
        RECT 41.150 -1.600 41.550 -0.600 ;
        RECT 11.150 -2.750 11.400 -1.600 ;
        RECT 26.150 -2.750 26.400 -1.600 ;
        RECT 41.150 -2.750 41.400 -1.600 ;
        RECT 10.350 -3.100 11.400 -2.750 ;
        RECT 25.350 -3.100 26.400 -2.750 ;
        RECT 40.350 -3.100 41.400 -2.750 ;
        RECT 4.000 -7.200 4.900 -6.750 ;
        RECT 19.000 -7.200 19.900 -6.750 ;
        RECT 34.000 -7.200 34.900 -6.750 ;
        RECT 4.000 -9.400 4.500 -7.200 ;
        RECT 19.000 -9.400 19.500 -7.200 ;
        RECT 34.000 -9.400 34.500 -7.200 ;
        RECT 2.650 -14.450 3.350 -13.250 ;
        RECT 17.650 -14.450 18.350 -13.250 ;
        RECT 32.650 -14.450 33.350 -13.250 ;
        RECT 2.900 -14.850 3.150 -14.450 ;
        RECT 17.900 -14.850 18.150 -14.450 ;
        RECT 32.900 -14.850 33.150 -14.450 ;
        RECT 11.150 -16.600 11.550 -15.600 ;
        RECT 26.150 -16.600 26.550 -15.600 ;
        RECT 41.150 -16.600 41.550 -15.600 ;
        RECT 11.150 -17.750 11.400 -16.600 ;
        RECT 26.150 -17.750 26.400 -16.600 ;
        RECT 41.150 -17.750 41.400 -16.600 ;
        RECT 10.350 -18.100 11.400 -17.750 ;
        RECT 25.350 -18.100 26.400 -17.750 ;
        RECT 40.350 -18.100 41.400 -17.750 ;
        RECT 4.000 -22.200 4.900 -21.750 ;
        RECT 19.000 -22.200 19.900 -21.750 ;
        RECT 34.000 -22.200 34.900 -21.750 ;
        RECT 4.000 -24.400 4.500 -22.200 ;
        RECT 19.000 -24.400 19.500 -22.200 ;
        RECT 34.000 -24.400 34.500 -22.200 ;
        RECT 2.650 -29.450 3.350 -28.250 ;
        RECT 17.650 -29.450 18.350 -28.250 ;
        RECT 32.650 -29.450 33.350 -28.250 ;
        RECT 2.900 -29.850 3.150 -29.450 ;
        RECT 17.900 -29.850 18.150 -29.450 ;
        RECT 32.900 -29.850 33.150 -29.450 ;
      LAYER mcon ;
        RECT 10.540 12.015 10.710 12.185 ;
        RECT 25.540 12.015 25.710 12.185 ;
        RECT 40.540 12.015 40.710 12.185 ;
        RECT 4.165 5.765 4.335 5.935 ;
        RECT 19.165 5.765 19.335 5.935 ;
        RECT 34.165 5.765 34.335 5.935 ;
        RECT 2.915 0.215 3.085 0.385 ;
        RECT 17.915 0.215 18.085 0.385 ;
        RECT 32.915 0.215 33.085 0.385 ;
        RECT 10.540 -2.985 10.710 -2.815 ;
        RECT 25.540 -2.985 25.710 -2.815 ;
        RECT 40.540 -2.985 40.710 -2.815 ;
        RECT 4.165 -9.235 4.335 -9.065 ;
        RECT 19.165 -9.235 19.335 -9.065 ;
        RECT 34.165 -9.235 34.335 -9.065 ;
        RECT 2.915 -14.785 3.085 -14.615 ;
        RECT 17.915 -14.785 18.085 -14.615 ;
        RECT 32.915 -14.785 33.085 -14.615 ;
        RECT 10.540 -17.985 10.710 -17.815 ;
        RECT 25.540 -17.985 25.710 -17.815 ;
        RECT 40.540 -17.985 40.710 -17.815 ;
        RECT 4.165 -24.235 4.335 -24.065 ;
        RECT 19.165 -24.235 19.335 -24.065 ;
        RECT 34.165 -24.235 34.335 -24.065 ;
        RECT 2.915 -29.785 3.085 -29.615 ;
        RECT 17.915 -29.785 18.085 -29.615 ;
        RECT 32.915 -29.785 33.085 -29.615 ;
      LAYER met1 ;
        RECT 10.350 11.900 10.950 12.350 ;
        RECT 25.350 11.900 25.950 12.350 ;
        RECT 40.350 11.900 40.950 12.350 ;
        RECT 3.950 5.600 6.500 6.100 ;
        RECT 5.950 0.900 6.500 5.600 ;
        RECT 10.350 0.900 10.850 11.900 ;
        RECT 18.950 5.600 21.500 6.100 ;
        RECT 20.950 0.900 21.500 5.600 ;
        RECT 25.350 0.900 25.850 11.900 ;
        RECT 33.950 5.600 36.500 6.100 ;
        RECT 35.950 0.900 36.500 5.600 ;
        RECT 40.350 0.900 40.850 11.900 ;
        RECT 47.000 0.900 48.000 15.150 ;
        RECT 0.000 0.150 48.000 0.900 ;
        RECT 10.350 -3.100 10.950 -2.650 ;
        RECT 25.350 -3.100 25.950 -2.650 ;
        RECT 40.350 -3.100 40.950 -2.650 ;
        RECT 3.950 -9.400 6.500 -8.900 ;
        RECT 5.950 -14.100 6.500 -9.400 ;
        RECT 10.350 -14.100 10.850 -3.100 ;
        RECT 18.950 -9.400 21.500 -8.900 ;
        RECT 20.950 -14.100 21.500 -9.400 ;
        RECT 25.350 -14.100 25.850 -3.100 ;
        RECT 33.950 -9.400 36.500 -8.900 ;
        RECT 35.950 -14.100 36.500 -9.400 ;
        RECT 40.350 -14.100 40.850 -3.100 ;
        RECT 47.000 -14.100 48.000 0.150 ;
        RECT 0.000 -14.850 48.000 -14.100 ;
        RECT 10.350 -18.100 10.950 -17.650 ;
        RECT 25.350 -18.100 25.950 -17.650 ;
        RECT 40.350 -18.100 40.950 -17.650 ;
        RECT 3.950 -24.400 6.500 -23.900 ;
        RECT 5.950 -29.100 6.500 -24.400 ;
        RECT 10.350 -29.100 10.850 -18.100 ;
        RECT 18.950 -24.400 21.500 -23.900 ;
        RECT 20.950 -29.100 21.500 -24.400 ;
        RECT 25.350 -29.100 25.850 -18.100 ;
        RECT 33.950 -24.400 36.500 -23.900 ;
        RECT 35.950 -29.100 36.500 -24.400 ;
        RECT 40.350 -29.100 40.850 -18.100 ;
        RECT 47.000 -29.100 48.000 -14.850 ;
        RECT 0.000 -29.850 48.000 -29.100 ;
      LAYER via ;
        RECT 7.420 0.245 7.680 0.505 ;
        RECT 22.420 0.245 22.680 0.505 ;
        RECT 37.420 0.245 37.680 0.505 ;
        RECT 7.420 -14.755 7.680 -14.495 ;
        RECT 22.420 -14.755 22.680 -14.495 ;
        RECT 37.420 -14.755 37.680 -14.495 ;
        RECT 7.420 -29.755 7.680 -29.495 ;
        RECT 22.420 -29.755 22.680 -29.495 ;
        RECT 37.420 -29.755 37.680 -29.495 ;
      LAYER met2 ;
        RECT 7.350 0.150 7.750 2.100 ;
        RECT 22.350 0.150 22.750 2.100 ;
        RECT 37.350 0.150 37.750 2.100 ;
        RECT 7.350 -14.850 7.750 -12.900 ;
        RECT 22.350 -14.850 22.750 -12.900 ;
        RECT 37.350 -14.850 37.750 -12.900 ;
        RECT 7.350 -29.850 7.750 -27.900 ;
        RECT 22.350 -29.850 22.750 -27.900 ;
        RECT 37.350 -29.850 37.750 -27.900 ;
      LAYER via2 ;
        RECT 7.410 1.685 7.690 1.965 ;
        RECT 22.410 1.685 22.690 1.965 ;
        RECT 37.410 1.685 37.690 1.965 ;
        RECT 7.410 -13.315 7.690 -13.035 ;
        RECT 22.410 -13.315 22.690 -13.035 ;
        RECT 37.410 -13.315 37.690 -13.035 ;
        RECT 7.410 -28.315 7.690 -28.035 ;
        RECT 22.410 -28.315 22.690 -28.035 ;
        RECT 37.410 -28.315 37.690 -28.035 ;
      LAYER met3 ;
        RECT 7.250 1.500 8.750 2.100 ;
        RECT 22.250 1.500 23.750 2.100 ;
        RECT 37.250 1.500 38.750 2.100 ;
        RECT 7.250 -13.500 8.750 -12.900 ;
        RECT 22.250 -13.500 23.750 -12.900 ;
        RECT 37.250 -13.500 38.750 -12.900 ;
        RECT 7.250 -28.500 8.750 -27.900 ;
        RECT 22.250 -28.500 23.750 -27.900 ;
        RECT 37.250 -28.500 38.750 -27.900 ;
      LAYER via3 ;
        RECT 8.265 1.640 8.585 1.960 ;
        RECT 23.265 1.640 23.585 1.960 ;
        RECT 38.265 1.640 38.585 1.960 ;
        RECT 8.265 -13.360 8.585 -13.040 ;
        RECT 23.265 -13.360 23.585 -13.040 ;
        RECT 38.265 -13.360 38.585 -13.040 ;
        RECT 8.265 -28.360 8.585 -28.040 ;
        RECT 23.265 -28.360 23.585 -28.040 ;
        RECT 38.265 -28.360 38.585 -28.040 ;
      LAYER met4 ;
        RECT 2.400 7.250 12.600 7.900 ;
        RECT 17.400 7.250 27.600 7.900 ;
        RECT 32.400 7.250 42.600 7.900 ;
        RECT 6.500 2.550 11.650 7.250 ;
        RECT 21.500 2.550 26.650 7.250 ;
        RECT 36.500 2.550 41.650 7.250 ;
        RECT 8.100 0.150 8.950 2.550 ;
        RECT 23.100 0.150 23.950 2.550 ;
        RECT 38.100 0.150 38.950 2.550 ;
        RECT 2.400 -7.750 12.600 -7.100 ;
        RECT 17.400 -7.750 27.600 -7.100 ;
        RECT 32.400 -7.750 42.600 -7.100 ;
        RECT 6.500 -12.450 11.650 -7.750 ;
        RECT 21.500 -12.450 26.650 -7.750 ;
        RECT 36.500 -12.450 41.650 -7.750 ;
        RECT 8.100 -14.850 8.950 -12.450 ;
        RECT 23.100 -14.850 23.950 -12.450 ;
        RECT 38.100 -14.850 38.950 -12.450 ;
        RECT 2.400 -22.750 12.600 -22.100 ;
        RECT 17.400 -22.750 27.600 -22.100 ;
        RECT 32.400 -22.750 42.600 -22.100 ;
        RECT 6.500 -27.450 11.650 -22.750 ;
        RECT 21.500 -27.450 26.650 -22.750 ;
        RECT 36.500 -27.450 41.650 -22.750 ;
        RECT 8.100 -29.850 8.950 -27.450 ;
        RECT 23.100 -29.850 23.950 -27.450 ;
        RECT 38.100 -29.850 38.950 -27.450 ;
    END
  END GND
  PIN ROW_SEL0
    ANTENNAGATEAREA 6.000000 ;
    PORT
      LAYER li1 ;
        RECT 12.000 7.950 12.250 9.000 ;
        RECT 27.000 7.950 27.250 9.000 ;
        RECT 42.000 7.950 42.250 9.000 ;
      LAYER mcon ;
        RECT 12.040 8.140 12.210 8.310 ;
        RECT 27.040 8.140 27.210 8.310 ;
        RECT 42.040 8.140 42.210 8.310 ;
      LAYER met1 ;
        RECT -8.000 7.400 0.000 7.850 ;
        RECT 11.950 7.500 12.300 8.500 ;
        RECT 26.950 7.500 27.300 8.500 ;
        RECT 41.950 7.500 42.300 8.500 ;
      LAYER via ;
        RECT -7.830 7.495 -7.570 7.755 ;
        RECT -7.510 7.495 -7.250 7.755 ;
        RECT -7.190 7.495 -6.930 7.755 ;
        RECT -6.870 7.495 -6.610 7.755 ;
        RECT -6.550 7.495 -6.290 7.755 ;
        RECT -6.230 7.495 -5.970 7.755 ;
        RECT -2.610 7.495 -2.350 7.755 ;
        RECT -2.290 7.495 -2.030 7.755 ;
        RECT -1.970 7.495 -1.710 7.755 ;
        RECT -1.650 7.495 -1.390 7.755 ;
        RECT 11.995 7.645 12.255 7.905 ;
        RECT 26.995 7.645 27.255 7.905 ;
        RECT 41.995 7.645 42.255 7.905 ;
      LAYER met2 ;
        RECT -15.000 7.400 -5.000 7.850 ;
        RECT -2.800 7.400 -1.300 7.850 ;
        RECT 11.950 7.750 12.300 8.050 ;
        RECT 26.950 7.750 27.300 8.050 ;
        RECT 41.950 7.750 42.300 8.050 ;
        RECT 11.950 7.400 12.850 7.750 ;
        RECT 26.950 7.400 27.850 7.750 ;
        RECT 41.950 7.400 42.850 7.750 ;
      LAYER via2 ;
        RECT -2.540 7.485 -2.260 7.765 ;
        RECT -2.140 7.485 -1.860 7.765 ;
        RECT -1.740 7.485 -1.460 7.765 ;
        RECT 12.435 7.435 12.715 7.715 ;
        RECT 27.435 7.435 27.715 7.715 ;
        RECT 42.435 7.435 42.715 7.715 ;
      LAYER met3 ;
        RECT -2.800 7.750 2.200 7.850 ;
        RECT 12.300 7.750 12.850 7.800 ;
        RECT 27.300 7.750 27.850 7.800 ;
        RECT 42.300 7.750 42.850 7.800 ;
        RECT -2.800 7.400 45.000 7.750 ;
        RECT 12.300 7.350 12.850 7.400 ;
        RECT 27.300 7.350 27.850 7.400 ;
        RECT 42.300 7.350 42.850 7.400 ;
    END
  END ROW_SEL0
  PIN ROW_SEL1
    ANTENNAGATEAREA 6.000000 ;
    PORT
      LAYER li1 ;
        RECT 12.000 -7.050 12.250 -6.000 ;
        RECT 27.000 -7.050 27.250 -6.000 ;
        RECT 42.000 -7.050 42.250 -6.000 ;
      LAYER mcon ;
        RECT 12.040 -6.860 12.210 -6.690 ;
        RECT 27.040 -6.860 27.210 -6.690 ;
        RECT 42.040 -6.860 42.210 -6.690 ;
      LAYER met1 ;
        RECT -8.000 -7.600 0.000 -7.150 ;
        RECT 11.950 -7.500 12.300 -6.500 ;
        RECT 26.950 -7.500 27.300 -6.500 ;
        RECT 41.950 -7.500 42.300 -6.500 ;
      LAYER via ;
        RECT -7.830 -7.505 -7.570 -7.245 ;
        RECT -7.510 -7.505 -7.250 -7.245 ;
        RECT -7.190 -7.505 -6.930 -7.245 ;
        RECT -6.870 -7.505 -6.610 -7.245 ;
        RECT -6.550 -7.505 -6.290 -7.245 ;
        RECT -6.230 -7.505 -5.970 -7.245 ;
        RECT -2.610 -7.505 -2.350 -7.245 ;
        RECT -2.290 -7.505 -2.030 -7.245 ;
        RECT -1.970 -7.505 -1.710 -7.245 ;
        RECT -1.650 -7.505 -1.390 -7.245 ;
        RECT 11.995 -7.355 12.255 -7.095 ;
        RECT 26.995 -7.355 27.255 -7.095 ;
        RECT 41.995 -7.355 42.255 -7.095 ;
      LAYER met2 ;
        RECT -15.000 -7.600 -5.000 -7.150 ;
        RECT -2.800 -7.600 -1.300 -7.150 ;
        RECT 11.950 -7.250 12.300 -6.950 ;
        RECT 26.950 -7.250 27.300 -6.950 ;
        RECT 41.950 -7.250 42.300 -6.950 ;
        RECT 11.950 -7.600 12.850 -7.250 ;
        RECT 26.950 -7.600 27.850 -7.250 ;
        RECT 41.950 -7.600 42.850 -7.250 ;
      LAYER via2 ;
        RECT -2.540 -7.515 -2.260 -7.235 ;
        RECT -2.140 -7.515 -1.860 -7.235 ;
        RECT -1.740 -7.515 -1.460 -7.235 ;
        RECT 12.435 -7.565 12.715 -7.285 ;
        RECT 27.435 -7.565 27.715 -7.285 ;
        RECT 42.435 -7.565 42.715 -7.285 ;
      LAYER met3 ;
        RECT -2.800 -7.250 2.200 -7.150 ;
        RECT 12.300 -7.250 12.850 -7.200 ;
        RECT 27.300 -7.250 27.850 -7.200 ;
        RECT 42.300 -7.250 42.850 -7.200 ;
        RECT -2.800 -7.600 45.000 -7.250 ;
        RECT 12.300 -7.650 12.850 -7.600 ;
        RECT 27.300 -7.650 27.850 -7.600 ;
        RECT 42.300 -7.650 42.850 -7.600 ;
    END
  END ROW_SEL1
  PIN ROW_SEL2
    ANTENNAGATEAREA 6.000000 ;
    PORT
      LAYER li1 ;
        RECT 12.000 -22.050 12.250 -21.000 ;
        RECT 27.000 -22.050 27.250 -21.000 ;
        RECT 42.000 -22.050 42.250 -21.000 ;
      LAYER mcon ;
        RECT 12.040 -21.860 12.210 -21.690 ;
        RECT 27.040 -21.860 27.210 -21.690 ;
        RECT 42.040 -21.860 42.210 -21.690 ;
      LAYER met1 ;
        RECT -8.000 -22.600 0.000 -22.150 ;
        RECT 11.950 -22.500 12.300 -21.500 ;
        RECT 26.950 -22.500 27.300 -21.500 ;
        RECT 41.950 -22.500 42.300 -21.500 ;
      LAYER via ;
        RECT -7.830 -22.505 -7.570 -22.245 ;
        RECT -7.510 -22.505 -7.250 -22.245 ;
        RECT -7.190 -22.505 -6.930 -22.245 ;
        RECT -6.870 -22.505 -6.610 -22.245 ;
        RECT -6.550 -22.505 -6.290 -22.245 ;
        RECT -6.230 -22.505 -5.970 -22.245 ;
        RECT -2.610 -22.505 -2.350 -22.245 ;
        RECT -2.290 -22.505 -2.030 -22.245 ;
        RECT -1.970 -22.505 -1.710 -22.245 ;
        RECT -1.650 -22.505 -1.390 -22.245 ;
        RECT 11.995 -22.355 12.255 -22.095 ;
        RECT 26.995 -22.355 27.255 -22.095 ;
        RECT 41.995 -22.355 42.255 -22.095 ;
      LAYER met2 ;
        RECT -15.000 -22.600 -5.000 -22.150 ;
        RECT -2.800 -22.600 -1.300 -22.150 ;
        RECT 11.950 -22.250 12.300 -21.950 ;
        RECT 26.950 -22.250 27.300 -21.950 ;
        RECT 41.950 -22.250 42.300 -21.950 ;
        RECT 11.950 -22.600 12.850 -22.250 ;
        RECT 26.950 -22.600 27.850 -22.250 ;
        RECT 41.950 -22.600 42.850 -22.250 ;
      LAYER via2 ;
        RECT -2.540 -22.515 -2.260 -22.235 ;
        RECT -2.140 -22.515 -1.860 -22.235 ;
        RECT -1.740 -22.515 -1.460 -22.235 ;
        RECT 12.435 -22.565 12.715 -22.285 ;
        RECT 27.435 -22.565 27.715 -22.285 ;
        RECT 42.435 -22.565 42.715 -22.285 ;
      LAYER met3 ;
        RECT -2.800 -22.250 2.200 -22.150 ;
        RECT 12.300 -22.250 12.850 -22.200 ;
        RECT 27.300 -22.250 27.850 -22.200 ;
        RECT 42.300 -22.250 42.850 -22.200 ;
        RECT -2.800 -22.600 45.000 -22.250 ;
        RECT 12.300 -22.650 12.850 -22.600 ;
        RECT 27.300 -22.650 27.850 -22.600 ;
        RECT 42.300 -22.650 42.850 -22.600 ;
    END
  END ROW_SEL2
  PIN PIX0_IN
    ANTENNAGATEAREA 1.050000 ;
    ANTENNADIFFAREA 0.294000 ;
    PORT
      LAYER li1 ;
        RECT 14.200 11.950 14.650 12.320 ;
        RECT 14.350 10.600 14.650 11.950 ;
        RECT 13.000 10.350 14.650 10.600 ;
        RECT 13.000 10.050 13.650 10.350 ;
        RECT 3.200 2.450 3.900 3.100 ;
        RECT 2.450 2.150 3.900 2.450 ;
      LAYER mcon ;
        RECT 13.060 10.240 13.230 10.410 ;
        RECT 13.420 10.240 13.590 10.410 ;
        RECT 3.465 2.870 3.635 3.040 ;
        RECT 3.465 2.510 3.635 2.680 ;
      LAYER met1 ;
        RECT 11.300 10.050 13.700 10.600 ;
        RECT 3.200 2.400 3.900 3.750 ;
      LAYER via ;
        RECT 11.400 10.195 11.660 10.455 ;
        RECT 11.720 10.195 11.980 10.455 ;
        RECT 12.040 10.195 12.300 10.455 ;
        RECT 3.260 3.270 3.520 3.530 ;
        RECT 3.580 3.270 3.840 3.530 ;
      LAYER met2 ;
        RECT 10.350 9.950 12.450 11.300 ;
        RECT 3.200 3.100 4.650 3.750 ;
      LAYER via2 ;
        RECT 10.435 10.060 11.115 11.140 ;
        RECT 3.385 3.335 3.665 3.615 ;
        RECT 3.785 3.335 4.065 3.615 ;
        RECT 4.185 3.335 4.465 3.615 ;
      LAYER met3 ;
        RECT 10.250 9.850 12.500 11.400 ;
        RECT 3.200 3.250 4.650 5.100 ;
      LAYER via3 ;
        RECT 10.390 10.065 11.110 11.185 ;
        RECT 3.590 3.365 4.310 4.885 ;
      LAYER met4 ;
        RECT 8.300 9.650 12.100 11.950 ;
        RECT 3.200 3.250 4.650 5.100 ;
      LAYER via4 ;
        RECT 10.060 10.035 11.240 11.215 ;
        RECT 3.360 3.785 4.540 4.965 ;
      LAYER met5 ;
        RECT 2.400 2.400 12.600 12.600 ;
    END
  END PIX0_IN
  PIN PIX1_IN
    ANTENNAGATEAREA 1.050000 ;
    ANTENNADIFFAREA 0.294000 ;
    PORT
      LAYER li1 ;
        RECT 29.200 11.950 29.650 12.320 ;
        RECT 29.350 10.600 29.650 11.950 ;
        RECT 28.000 10.350 29.650 10.600 ;
        RECT 28.000 10.050 28.650 10.350 ;
        RECT 18.200 2.450 18.900 3.100 ;
        RECT 17.450 2.150 18.900 2.450 ;
      LAYER mcon ;
        RECT 28.060 10.240 28.230 10.410 ;
        RECT 28.420 10.240 28.590 10.410 ;
        RECT 18.465 2.870 18.635 3.040 ;
        RECT 18.465 2.510 18.635 2.680 ;
      LAYER met1 ;
        RECT 26.300 10.050 28.700 10.600 ;
        RECT 18.200 2.400 18.900 3.750 ;
      LAYER via ;
        RECT 26.400 10.195 26.660 10.455 ;
        RECT 26.720 10.195 26.980 10.455 ;
        RECT 27.040 10.195 27.300 10.455 ;
        RECT 18.260 3.270 18.520 3.530 ;
        RECT 18.580 3.270 18.840 3.530 ;
      LAYER met2 ;
        RECT 25.350 9.950 27.450 11.300 ;
        RECT 18.200 3.100 19.650 3.750 ;
      LAYER via2 ;
        RECT 25.435 10.060 26.115 11.140 ;
        RECT 18.385 3.335 18.665 3.615 ;
        RECT 18.785 3.335 19.065 3.615 ;
        RECT 19.185 3.335 19.465 3.615 ;
      LAYER met3 ;
        RECT 25.250 9.850 27.500 11.400 ;
        RECT 18.200 3.250 19.650 5.100 ;
      LAYER via3 ;
        RECT 25.390 10.065 26.110 11.185 ;
        RECT 18.590 3.365 19.310 4.885 ;
      LAYER met4 ;
        RECT 23.300 9.650 27.100 11.950 ;
        RECT 18.200 3.250 19.650 5.100 ;
      LAYER via4 ;
        RECT 25.060 10.035 26.240 11.215 ;
        RECT 18.360 3.785 19.540 4.965 ;
      LAYER met5 ;
        RECT 17.400 2.400 27.600 12.600 ;
    END
  END PIX1_IN
  PIN PIX2_IN
    ANTENNAGATEAREA 1.050000 ;
    ANTENNADIFFAREA 0.294000 ;
    PORT
      LAYER li1 ;
        RECT 44.200 11.950 44.650 12.320 ;
        RECT 44.350 10.600 44.650 11.950 ;
        RECT 43.000 10.350 44.650 10.600 ;
        RECT 43.000 10.050 43.650 10.350 ;
        RECT 33.200 2.450 33.900 3.100 ;
        RECT 32.450 2.150 33.900 2.450 ;
      LAYER mcon ;
        RECT 43.060 10.240 43.230 10.410 ;
        RECT 43.420 10.240 43.590 10.410 ;
        RECT 33.465 2.870 33.635 3.040 ;
        RECT 33.465 2.510 33.635 2.680 ;
      LAYER met1 ;
        RECT 41.300 10.050 43.700 10.600 ;
        RECT 33.200 2.400 33.900 3.750 ;
      LAYER via ;
        RECT 41.400 10.195 41.660 10.455 ;
        RECT 41.720 10.195 41.980 10.455 ;
        RECT 42.040 10.195 42.300 10.455 ;
        RECT 33.260 3.270 33.520 3.530 ;
        RECT 33.580 3.270 33.840 3.530 ;
      LAYER met2 ;
        RECT 40.350 9.950 42.450 11.300 ;
        RECT 33.200 3.100 34.650 3.750 ;
      LAYER via2 ;
        RECT 40.435 10.060 41.115 11.140 ;
        RECT 33.385 3.335 33.665 3.615 ;
        RECT 33.785 3.335 34.065 3.615 ;
        RECT 34.185 3.335 34.465 3.615 ;
      LAYER met3 ;
        RECT 40.250 9.850 42.500 11.400 ;
        RECT 33.200 3.250 34.650 5.100 ;
      LAYER via3 ;
        RECT 40.390 10.065 41.110 11.185 ;
        RECT 33.590 3.365 34.310 4.885 ;
      LAYER met4 ;
        RECT 38.300 9.650 42.100 11.950 ;
        RECT 33.200 3.250 34.650 5.100 ;
      LAYER via4 ;
        RECT 40.060 10.035 41.240 11.215 ;
        RECT 33.360 3.785 34.540 4.965 ;
      LAYER met5 ;
        RECT 32.400 2.400 42.600 12.600 ;
    END
  END PIX2_IN
  PIN PIX3_IN
    ANTENNAGATEAREA 1.050000 ;
    ANTENNADIFFAREA 0.294000 ;
    PORT
      LAYER li1 ;
        RECT 14.200 -3.050 14.650 -2.680 ;
        RECT 14.350 -4.400 14.650 -3.050 ;
        RECT 13.000 -4.650 14.650 -4.400 ;
        RECT 13.000 -4.950 13.650 -4.650 ;
        RECT 3.200 -12.550 3.900 -11.900 ;
        RECT 2.450 -12.850 3.900 -12.550 ;
      LAYER mcon ;
        RECT 13.060 -4.760 13.230 -4.590 ;
        RECT 13.420 -4.760 13.590 -4.590 ;
        RECT 3.465 -12.130 3.635 -11.960 ;
        RECT 3.465 -12.490 3.635 -12.320 ;
      LAYER met1 ;
        RECT 11.300 -4.950 13.700 -4.400 ;
        RECT 3.200 -12.600 3.900 -11.250 ;
      LAYER via ;
        RECT 11.400 -4.805 11.660 -4.545 ;
        RECT 11.720 -4.805 11.980 -4.545 ;
        RECT 12.040 -4.805 12.300 -4.545 ;
        RECT 3.260 -11.730 3.520 -11.470 ;
        RECT 3.580 -11.730 3.840 -11.470 ;
      LAYER met2 ;
        RECT 10.350 -5.050 12.450 -3.700 ;
        RECT 3.200 -11.900 4.650 -11.250 ;
      LAYER via2 ;
        RECT 10.435 -4.940 11.115 -3.860 ;
        RECT 3.385 -11.665 3.665 -11.385 ;
        RECT 3.785 -11.665 4.065 -11.385 ;
        RECT 4.185 -11.665 4.465 -11.385 ;
      LAYER met3 ;
        RECT 10.250 -5.150 12.500 -3.600 ;
        RECT 3.200 -11.750 4.650 -9.900 ;
      LAYER via3 ;
        RECT 10.390 -4.935 11.110 -3.815 ;
        RECT 3.590 -11.635 4.310 -10.115 ;
      LAYER met4 ;
        RECT 8.300 -5.350 12.100 -3.050 ;
        RECT 3.200 -11.750 4.650 -9.900 ;
      LAYER via4 ;
        RECT 10.060 -4.965 11.240 -3.785 ;
        RECT 3.360 -11.215 4.540 -10.035 ;
      LAYER met5 ;
        RECT 2.400 -12.600 12.600 -2.400 ;
    END
  END PIX3_IN
  PIN PIX4_IN
    ANTENNAGATEAREA 1.050000 ;
    ANTENNADIFFAREA 0.294000 ;
    PORT
      LAYER li1 ;
        RECT 29.200 -3.050 29.650 -2.680 ;
        RECT 29.350 -4.400 29.650 -3.050 ;
        RECT 28.000 -4.650 29.650 -4.400 ;
        RECT 28.000 -4.950 28.650 -4.650 ;
        RECT 18.200 -12.550 18.900 -11.900 ;
        RECT 17.450 -12.850 18.900 -12.550 ;
      LAYER mcon ;
        RECT 28.060 -4.760 28.230 -4.590 ;
        RECT 28.420 -4.760 28.590 -4.590 ;
        RECT 18.465 -12.130 18.635 -11.960 ;
        RECT 18.465 -12.490 18.635 -12.320 ;
      LAYER met1 ;
        RECT 26.300 -4.950 28.700 -4.400 ;
        RECT 18.200 -12.600 18.900 -11.250 ;
      LAYER via ;
        RECT 26.400 -4.805 26.660 -4.545 ;
        RECT 26.720 -4.805 26.980 -4.545 ;
        RECT 27.040 -4.805 27.300 -4.545 ;
        RECT 18.260 -11.730 18.520 -11.470 ;
        RECT 18.580 -11.730 18.840 -11.470 ;
      LAYER met2 ;
        RECT 25.350 -5.050 27.450 -3.700 ;
        RECT 18.200 -11.900 19.650 -11.250 ;
      LAYER via2 ;
        RECT 25.435 -4.940 26.115 -3.860 ;
        RECT 18.385 -11.665 18.665 -11.385 ;
        RECT 18.785 -11.665 19.065 -11.385 ;
        RECT 19.185 -11.665 19.465 -11.385 ;
      LAYER met3 ;
        RECT 25.250 -5.150 27.500 -3.600 ;
        RECT 18.200 -11.750 19.650 -9.900 ;
      LAYER via3 ;
        RECT 25.390 -4.935 26.110 -3.815 ;
        RECT 18.590 -11.635 19.310 -10.115 ;
      LAYER met4 ;
        RECT 23.300 -5.350 27.100 -3.050 ;
        RECT 18.200 -11.750 19.650 -9.900 ;
      LAYER via4 ;
        RECT 25.060 -4.965 26.240 -3.785 ;
        RECT 18.360 -11.215 19.540 -10.035 ;
      LAYER met5 ;
        RECT 17.400 -12.600 27.600 -2.400 ;
    END
  END PIX4_IN
  PIN PIX5_IN
    ANTENNAGATEAREA 1.050000 ;
    ANTENNADIFFAREA 0.294000 ;
    PORT
      LAYER li1 ;
        RECT 44.200 -3.050 44.650 -2.680 ;
        RECT 44.350 -4.400 44.650 -3.050 ;
        RECT 43.000 -4.650 44.650 -4.400 ;
        RECT 43.000 -4.950 43.650 -4.650 ;
        RECT 33.200 -12.550 33.900 -11.900 ;
        RECT 32.450 -12.850 33.900 -12.550 ;
      LAYER mcon ;
        RECT 43.060 -4.760 43.230 -4.590 ;
        RECT 43.420 -4.760 43.590 -4.590 ;
        RECT 33.465 -12.130 33.635 -11.960 ;
        RECT 33.465 -12.490 33.635 -12.320 ;
      LAYER met1 ;
        RECT 41.300 -4.950 43.700 -4.400 ;
        RECT 33.200 -12.600 33.900 -11.250 ;
      LAYER via ;
        RECT 41.400 -4.805 41.660 -4.545 ;
        RECT 41.720 -4.805 41.980 -4.545 ;
        RECT 42.040 -4.805 42.300 -4.545 ;
        RECT 33.260 -11.730 33.520 -11.470 ;
        RECT 33.580 -11.730 33.840 -11.470 ;
      LAYER met2 ;
        RECT 40.350 -5.050 42.450 -3.700 ;
        RECT 33.200 -11.900 34.650 -11.250 ;
      LAYER via2 ;
        RECT 40.435 -4.940 41.115 -3.860 ;
        RECT 33.385 -11.665 33.665 -11.385 ;
        RECT 33.785 -11.665 34.065 -11.385 ;
        RECT 34.185 -11.665 34.465 -11.385 ;
      LAYER met3 ;
        RECT 40.250 -5.150 42.500 -3.600 ;
        RECT 33.200 -11.750 34.650 -9.900 ;
      LAYER via3 ;
        RECT 40.390 -4.935 41.110 -3.815 ;
        RECT 33.590 -11.635 34.310 -10.115 ;
      LAYER met4 ;
        RECT 38.300 -5.350 42.100 -3.050 ;
        RECT 33.200 -11.750 34.650 -9.900 ;
      LAYER via4 ;
        RECT 40.060 -4.965 41.240 -3.785 ;
        RECT 33.360 -11.215 34.540 -10.035 ;
      LAYER met5 ;
        RECT 32.400 -12.600 42.600 -2.400 ;
    END
  END PIX5_IN
  PIN PIX6_IN
    ANTENNAGATEAREA 1.050000 ;
    ANTENNADIFFAREA 0.294000 ;
    PORT
      LAYER li1 ;
        RECT 14.200 -18.050 14.650 -17.680 ;
        RECT 14.350 -19.400 14.650 -18.050 ;
        RECT 13.000 -19.650 14.650 -19.400 ;
        RECT 13.000 -19.950 13.650 -19.650 ;
        RECT 3.200 -27.550 3.900 -26.900 ;
        RECT 2.450 -27.850 3.900 -27.550 ;
      LAYER mcon ;
        RECT 13.060 -19.760 13.230 -19.590 ;
        RECT 13.420 -19.760 13.590 -19.590 ;
        RECT 3.465 -27.130 3.635 -26.960 ;
        RECT 3.465 -27.490 3.635 -27.320 ;
      LAYER met1 ;
        RECT 11.300 -19.950 13.700 -19.400 ;
        RECT 3.200 -27.600 3.900 -26.250 ;
      LAYER via ;
        RECT 11.400 -19.805 11.660 -19.545 ;
        RECT 11.720 -19.805 11.980 -19.545 ;
        RECT 12.040 -19.805 12.300 -19.545 ;
        RECT 3.260 -26.730 3.520 -26.470 ;
        RECT 3.580 -26.730 3.840 -26.470 ;
      LAYER met2 ;
        RECT 10.350 -20.050 12.450 -18.700 ;
        RECT 3.200 -26.900 4.650 -26.250 ;
      LAYER via2 ;
        RECT 10.435 -19.940 11.115 -18.860 ;
        RECT 3.385 -26.665 3.665 -26.385 ;
        RECT 3.785 -26.665 4.065 -26.385 ;
        RECT 4.185 -26.665 4.465 -26.385 ;
      LAYER met3 ;
        RECT 10.250 -20.150 12.500 -18.600 ;
        RECT 3.200 -26.750 4.650 -24.900 ;
      LAYER via3 ;
        RECT 10.390 -19.935 11.110 -18.815 ;
        RECT 3.590 -26.635 4.310 -25.115 ;
      LAYER met4 ;
        RECT 8.300 -20.350 12.100 -18.050 ;
        RECT 3.200 -26.750 4.650 -24.900 ;
      LAYER via4 ;
        RECT 10.060 -19.965 11.240 -18.785 ;
        RECT 3.360 -26.215 4.540 -25.035 ;
      LAYER met5 ;
        RECT 2.400 -27.600 12.600 -17.400 ;
    END
  END PIX6_IN
  PIN PIX_OUT0
    ANTENNADIFFAREA 6.400000 ;
    PORT
      LAYER li1 ;
        RECT 9.750 7.450 11.700 7.800 ;
        RECT 10.950 6.050 11.700 7.450 ;
        RECT 10.950 5.300 13.950 6.050 ;
        RECT 9.750 -7.550 11.700 -7.200 ;
        RECT 10.950 -8.950 11.700 -7.550 ;
        RECT 10.950 -9.700 13.950 -8.950 ;
        RECT 9.750 -22.550 11.700 -22.200 ;
        RECT 10.950 -23.950 11.700 -22.550 ;
        RECT 10.950 -24.700 13.950 -23.950 ;
        RECT 2.700 -31.900 10.700 -31.150 ;
      LAYER mcon ;
        RECT 13.260 5.410 13.790 5.940 ;
        RECT 13.260 -9.590 13.790 -9.060 ;
        RECT 13.260 -24.590 13.790 -24.060 ;
        RECT 2.835 -31.385 3.005 -31.215 ;
        RECT 3.195 -31.385 3.365 -31.215 ;
        RECT 3.555 -31.385 3.725 -31.215 ;
        RECT 3.915 -31.385 4.085 -31.215 ;
        RECT 4.275 -31.385 4.445 -31.215 ;
        RECT 4.635 -31.385 4.805 -31.215 ;
        RECT 4.995 -31.385 5.165 -31.215 ;
        RECT 5.355 -31.385 5.525 -31.215 ;
        RECT 5.715 -31.385 5.885 -31.215 ;
        RECT 6.075 -31.385 6.245 -31.215 ;
        RECT 6.435 -31.385 6.605 -31.215 ;
        RECT 6.795 -31.385 6.965 -31.215 ;
        RECT 7.155 -31.385 7.325 -31.215 ;
        RECT 7.515 -31.385 7.685 -31.215 ;
        RECT 7.875 -31.385 8.045 -31.215 ;
        RECT 8.235 -31.385 8.405 -31.215 ;
        RECT 8.595 -31.385 8.765 -31.215 ;
        RECT 8.955 -31.385 9.125 -31.215 ;
        RECT 9.315 -31.385 9.485 -31.215 ;
        RECT 9.675 -31.385 9.845 -31.215 ;
        RECT 10.035 -31.385 10.205 -31.215 ;
        RECT 10.395 -31.385 10.565 -31.215 ;
      LAYER met1 ;
        RECT 13.100 5.300 13.950 6.050 ;
        RECT 13.100 -9.700 13.950 -8.950 ;
        RECT 13.100 -24.700 13.950 -23.950 ;
        RECT 2.700 -31.500 10.700 -30.650 ;
      LAYER via ;
        RECT 13.235 5.385 13.815 5.965 ;
        RECT 13.235 -9.615 13.815 -9.035 ;
        RECT 13.235 -24.615 13.815 -24.035 ;
        RECT 2.890 -30.955 3.150 -30.695 ;
        RECT 3.210 -30.955 3.470 -30.695 ;
        RECT 3.530 -30.955 3.790 -30.695 ;
        RECT 3.850 -30.955 4.110 -30.695 ;
        RECT 4.170 -30.955 4.430 -30.695 ;
        RECT 4.490 -30.955 4.750 -30.695 ;
        RECT 4.810 -30.955 5.070 -30.695 ;
        RECT 5.130 -30.955 5.390 -30.695 ;
        RECT 5.450 -30.955 5.710 -30.695 ;
        RECT 5.770 -30.955 6.030 -30.695 ;
        RECT 6.090 -30.955 6.350 -30.695 ;
        RECT 6.410 -30.955 6.670 -30.695 ;
        RECT 6.730 -30.955 6.990 -30.695 ;
        RECT 7.050 -30.955 7.310 -30.695 ;
        RECT 7.370 -30.955 7.630 -30.695 ;
        RECT 7.690 -30.955 7.950 -30.695 ;
        RECT 8.010 -30.955 8.270 -30.695 ;
        RECT 8.330 -30.955 8.590 -30.695 ;
        RECT 8.650 -30.955 8.910 -30.695 ;
        RECT 8.970 -30.955 9.230 -30.695 ;
        RECT 9.290 -30.955 9.550 -30.695 ;
        RECT 9.610 -30.955 9.870 -30.695 ;
        RECT 9.930 -30.955 10.190 -30.695 ;
        RECT 10.250 -30.955 10.510 -30.695 ;
      LAYER met2 ;
        RECT 13.100 5.250 13.950 6.100 ;
        RECT 13.100 -9.750 13.950 -8.900 ;
        RECT 13.100 -24.750 13.950 -23.900 ;
        RECT 2.700 -31.000 13.900 -30.300 ;
      LAYER via2 ;
        RECT 13.185 5.335 13.865 6.015 ;
        RECT 13.185 -9.665 13.865 -8.985 ;
        RECT 13.185 -24.665 13.865 -23.985 ;
        RECT 2.960 -30.790 3.240 -30.510 ;
        RECT 3.360 -30.790 3.640 -30.510 ;
        RECT 3.760 -30.790 4.040 -30.510 ;
        RECT 4.160 -30.790 4.440 -30.510 ;
        RECT 4.560 -30.790 4.840 -30.510 ;
        RECT 4.960 -30.790 5.240 -30.510 ;
        RECT 5.360 -30.790 5.640 -30.510 ;
        RECT 5.760 -30.790 6.040 -30.510 ;
        RECT 6.160 -30.790 6.440 -30.510 ;
        RECT 6.560 -30.790 6.840 -30.510 ;
        RECT 6.960 -30.790 7.240 -30.510 ;
        RECT 7.360 -30.790 7.640 -30.510 ;
        RECT 7.760 -30.790 8.040 -30.510 ;
        RECT 8.160 -30.790 8.440 -30.510 ;
        RECT 8.560 -30.790 8.840 -30.510 ;
        RECT 8.960 -30.790 9.240 -30.510 ;
        RECT 9.360 -30.790 9.640 -30.510 ;
        RECT 9.760 -30.790 10.040 -30.510 ;
        RECT 10.160 -30.790 10.440 -30.510 ;
        RECT 10.560 -30.790 10.840 -30.510 ;
        RECT 10.960 -30.790 11.240 -30.510 ;
        RECT 11.360 -30.790 11.640 -30.510 ;
        RECT 11.760 -30.790 12.040 -30.510 ;
        RECT 12.160 -30.790 12.440 -30.510 ;
        RECT 12.560 -30.790 12.840 -30.510 ;
        RECT 12.960 -30.790 13.240 -30.510 ;
        RECT 13.360 -30.790 13.640 -30.510 ;
      LAYER met3 ;
        RECT 13.100 5.200 13.950 6.150 ;
        RECT 13.100 -9.800 13.950 -8.850 ;
        RECT 13.100 -24.800 13.950 -23.850 ;
        RECT 2.700 -31.000 13.900 -30.300 ;
      LAYER via3 ;
        RECT 13.165 5.315 13.885 6.035 ;
        RECT 13.165 -9.685 13.885 -8.965 ;
        RECT 13.165 -24.685 13.885 -23.965 ;
        RECT 2.940 -30.810 3.260 -30.490 ;
        RECT 3.340 -30.810 3.660 -30.490 ;
        RECT 3.740 -30.810 4.060 -30.490 ;
        RECT 4.140 -30.810 4.460 -30.490 ;
        RECT 4.540 -30.810 4.860 -30.490 ;
        RECT 4.940 -30.810 5.260 -30.490 ;
        RECT 5.340 -30.810 5.660 -30.490 ;
        RECT 5.740 -30.810 6.060 -30.490 ;
        RECT 6.140 -30.810 6.460 -30.490 ;
        RECT 6.540 -30.810 6.860 -30.490 ;
        RECT 6.940 -30.810 7.260 -30.490 ;
        RECT 7.340 -30.810 7.660 -30.490 ;
        RECT 7.740 -30.810 8.060 -30.490 ;
        RECT 8.140 -30.810 8.460 -30.490 ;
        RECT 8.540 -30.810 8.860 -30.490 ;
        RECT 8.940 -30.810 9.260 -30.490 ;
        RECT 9.340 -30.810 9.660 -30.490 ;
        RECT 9.740 -30.810 10.060 -30.490 ;
        RECT 10.140 -30.810 10.460 -30.490 ;
        RECT 10.540 -30.810 10.860 -30.490 ;
        RECT 10.940 -30.810 11.260 -30.490 ;
        RECT 11.340 -30.810 11.660 -30.490 ;
        RECT 11.740 -30.810 12.060 -30.490 ;
        RECT 12.140 -30.810 12.460 -30.490 ;
        RECT 12.540 -30.810 12.860 -30.490 ;
        RECT 12.940 -30.810 13.260 -30.490 ;
        RECT 13.340 -30.810 13.660 -30.490 ;
      LAYER met4 ;
        RECT 13.150 6.100 13.900 15.800 ;
        RECT 13.100 5.250 13.950 6.100 ;
        RECT 13.150 -8.900 13.900 5.250 ;
        RECT 13.100 -9.750 13.950 -8.900 ;
        RECT 13.150 -23.900 13.900 -9.750 ;
        RECT 13.100 -24.750 13.950 -23.900 ;
        RECT 13.150 -30.300 13.900 -24.750 ;
        RECT 2.700 -31.000 13.900 -30.300 ;
    END
  END PIX_OUT0
  PIN COL_SEL0
    ANTENNAGATEAREA 16.000000 ;
    PORT
      LAYER li1 ;
        RECT 1.100 -33.550 2.200 -32.450 ;
      LAYER mcon ;
        RECT 1.205 -33.445 2.095 -32.555 ;
      LAYER met1 ;
        RECT 1.100 -33.550 2.200 -32.450 ;
      LAYER via ;
        RECT 1.200 -33.450 2.100 -32.550 ;
      LAYER met2 ;
        RECT 1.100 -33.550 2.200 -32.450 ;
      LAYER via2 ;
        RECT 1.310 -33.340 1.990 -32.660 ;
      LAYER met3 ;
        RECT 1.100 -33.550 2.200 -32.450 ;
      LAYER via3 ;
        RECT 1.290 -33.360 2.010 -32.640 ;
      LAYER met4 ;
        RECT 1.100 -35.500 2.200 -32.450 ;
    END
  END COL_SEL0
  PIN PIX7_IN
    ANTENNAGATEAREA 1.050000 ;
    ANTENNADIFFAREA 0.294000 ;
    PORT
      LAYER li1 ;
        RECT 29.200 -18.050 29.650 -17.680 ;
        RECT 29.350 -19.400 29.650 -18.050 ;
        RECT 28.000 -19.650 29.650 -19.400 ;
        RECT 28.000 -19.950 28.650 -19.650 ;
        RECT 18.200 -27.550 18.900 -26.900 ;
        RECT 17.450 -27.850 18.900 -27.550 ;
      LAYER mcon ;
        RECT 28.060 -19.760 28.230 -19.590 ;
        RECT 28.420 -19.760 28.590 -19.590 ;
        RECT 18.465 -27.130 18.635 -26.960 ;
        RECT 18.465 -27.490 18.635 -27.320 ;
      LAYER met1 ;
        RECT 26.300 -19.950 28.700 -19.400 ;
        RECT 18.200 -27.600 18.900 -26.250 ;
      LAYER via ;
        RECT 26.400 -19.805 26.660 -19.545 ;
        RECT 26.720 -19.805 26.980 -19.545 ;
        RECT 27.040 -19.805 27.300 -19.545 ;
        RECT 18.260 -26.730 18.520 -26.470 ;
        RECT 18.580 -26.730 18.840 -26.470 ;
      LAYER met2 ;
        RECT 25.350 -20.050 27.450 -18.700 ;
        RECT 18.200 -26.900 19.650 -26.250 ;
      LAYER via2 ;
        RECT 25.435 -19.940 26.115 -18.860 ;
        RECT 18.385 -26.665 18.665 -26.385 ;
        RECT 18.785 -26.665 19.065 -26.385 ;
        RECT 19.185 -26.665 19.465 -26.385 ;
      LAYER met3 ;
        RECT 25.250 -20.150 27.500 -18.600 ;
        RECT 18.200 -26.750 19.650 -24.900 ;
      LAYER via3 ;
        RECT 25.390 -19.935 26.110 -18.815 ;
        RECT 18.590 -26.635 19.310 -25.115 ;
      LAYER met4 ;
        RECT 23.300 -20.350 27.100 -18.050 ;
        RECT 18.200 -26.750 19.650 -24.900 ;
      LAYER via4 ;
        RECT 25.060 -19.965 26.240 -18.785 ;
        RECT 18.360 -26.215 19.540 -25.035 ;
      LAYER met5 ;
        RECT 17.400 -27.600 27.600 -17.400 ;
    END
  END PIX7_IN
  PIN PIX_OUT1
    ANTENNADIFFAREA 6.400000 ;
    PORT
      LAYER li1 ;
        RECT 24.750 7.450 26.700 7.800 ;
        RECT 25.950 6.050 26.700 7.450 ;
        RECT 25.950 5.300 28.950 6.050 ;
        RECT 24.750 -7.550 26.700 -7.200 ;
        RECT 25.950 -8.950 26.700 -7.550 ;
        RECT 25.950 -9.700 28.950 -8.950 ;
        RECT 24.750 -22.550 26.700 -22.200 ;
        RECT 25.950 -23.950 26.700 -22.550 ;
        RECT 25.950 -24.700 28.950 -23.950 ;
        RECT 17.700 -31.900 25.700 -31.150 ;
      LAYER mcon ;
        RECT 28.260 5.410 28.790 5.940 ;
        RECT 28.260 -9.590 28.790 -9.060 ;
        RECT 28.260 -24.590 28.790 -24.060 ;
        RECT 17.835 -31.385 18.005 -31.215 ;
        RECT 18.195 -31.385 18.365 -31.215 ;
        RECT 18.555 -31.385 18.725 -31.215 ;
        RECT 18.915 -31.385 19.085 -31.215 ;
        RECT 19.275 -31.385 19.445 -31.215 ;
        RECT 19.635 -31.385 19.805 -31.215 ;
        RECT 19.995 -31.385 20.165 -31.215 ;
        RECT 20.355 -31.385 20.525 -31.215 ;
        RECT 20.715 -31.385 20.885 -31.215 ;
        RECT 21.075 -31.385 21.245 -31.215 ;
        RECT 21.435 -31.385 21.605 -31.215 ;
        RECT 21.795 -31.385 21.965 -31.215 ;
        RECT 22.155 -31.385 22.325 -31.215 ;
        RECT 22.515 -31.385 22.685 -31.215 ;
        RECT 22.875 -31.385 23.045 -31.215 ;
        RECT 23.235 -31.385 23.405 -31.215 ;
        RECT 23.595 -31.385 23.765 -31.215 ;
        RECT 23.955 -31.385 24.125 -31.215 ;
        RECT 24.315 -31.385 24.485 -31.215 ;
        RECT 24.675 -31.385 24.845 -31.215 ;
        RECT 25.035 -31.385 25.205 -31.215 ;
        RECT 25.395 -31.385 25.565 -31.215 ;
      LAYER met1 ;
        RECT 28.100 5.300 28.950 6.050 ;
        RECT 28.100 -9.700 28.950 -8.950 ;
        RECT 28.100 -24.700 28.950 -23.950 ;
        RECT 17.700 -31.500 25.700 -30.650 ;
      LAYER via ;
        RECT 28.235 5.385 28.815 5.965 ;
        RECT 28.235 -9.615 28.815 -9.035 ;
        RECT 28.235 -24.615 28.815 -24.035 ;
        RECT 17.890 -30.955 18.150 -30.695 ;
        RECT 18.210 -30.955 18.470 -30.695 ;
        RECT 18.530 -30.955 18.790 -30.695 ;
        RECT 18.850 -30.955 19.110 -30.695 ;
        RECT 19.170 -30.955 19.430 -30.695 ;
        RECT 19.490 -30.955 19.750 -30.695 ;
        RECT 19.810 -30.955 20.070 -30.695 ;
        RECT 20.130 -30.955 20.390 -30.695 ;
        RECT 20.450 -30.955 20.710 -30.695 ;
        RECT 20.770 -30.955 21.030 -30.695 ;
        RECT 21.090 -30.955 21.350 -30.695 ;
        RECT 21.410 -30.955 21.670 -30.695 ;
        RECT 21.730 -30.955 21.990 -30.695 ;
        RECT 22.050 -30.955 22.310 -30.695 ;
        RECT 22.370 -30.955 22.630 -30.695 ;
        RECT 22.690 -30.955 22.950 -30.695 ;
        RECT 23.010 -30.955 23.270 -30.695 ;
        RECT 23.330 -30.955 23.590 -30.695 ;
        RECT 23.650 -30.955 23.910 -30.695 ;
        RECT 23.970 -30.955 24.230 -30.695 ;
        RECT 24.290 -30.955 24.550 -30.695 ;
        RECT 24.610 -30.955 24.870 -30.695 ;
        RECT 24.930 -30.955 25.190 -30.695 ;
        RECT 25.250 -30.955 25.510 -30.695 ;
      LAYER met2 ;
        RECT 28.100 5.250 28.950 6.100 ;
        RECT 28.100 -9.750 28.950 -8.900 ;
        RECT 28.100 -24.750 28.950 -23.900 ;
        RECT 17.700 -31.000 28.900 -30.300 ;
      LAYER via2 ;
        RECT 28.185 5.335 28.865 6.015 ;
        RECT 28.185 -9.665 28.865 -8.985 ;
        RECT 28.185 -24.665 28.865 -23.985 ;
        RECT 17.960 -30.790 18.240 -30.510 ;
        RECT 18.360 -30.790 18.640 -30.510 ;
        RECT 18.760 -30.790 19.040 -30.510 ;
        RECT 19.160 -30.790 19.440 -30.510 ;
        RECT 19.560 -30.790 19.840 -30.510 ;
        RECT 19.960 -30.790 20.240 -30.510 ;
        RECT 20.360 -30.790 20.640 -30.510 ;
        RECT 20.760 -30.790 21.040 -30.510 ;
        RECT 21.160 -30.790 21.440 -30.510 ;
        RECT 21.560 -30.790 21.840 -30.510 ;
        RECT 21.960 -30.790 22.240 -30.510 ;
        RECT 22.360 -30.790 22.640 -30.510 ;
        RECT 22.760 -30.790 23.040 -30.510 ;
        RECT 23.160 -30.790 23.440 -30.510 ;
        RECT 23.560 -30.790 23.840 -30.510 ;
        RECT 23.960 -30.790 24.240 -30.510 ;
        RECT 24.360 -30.790 24.640 -30.510 ;
        RECT 24.760 -30.790 25.040 -30.510 ;
        RECT 25.160 -30.790 25.440 -30.510 ;
        RECT 25.560 -30.790 25.840 -30.510 ;
        RECT 25.960 -30.790 26.240 -30.510 ;
        RECT 26.360 -30.790 26.640 -30.510 ;
        RECT 26.760 -30.790 27.040 -30.510 ;
        RECT 27.160 -30.790 27.440 -30.510 ;
        RECT 27.560 -30.790 27.840 -30.510 ;
        RECT 27.960 -30.790 28.240 -30.510 ;
        RECT 28.360 -30.790 28.640 -30.510 ;
      LAYER met3 ;
        RECT 28.100 5.200 28.950 6.150 ;
        RECT 28.100 -9.800 28.950 -8.850 ;
        RECT 28.100 -24.800 28.950 -23.850 ;
        RECT 17.700 -31.000 28.900 -30.300 ;
      LAYER via3 ;
        RECT 28.165 5.315 28.885 6.035 ;
        RECT 28.165 -9.685 28.885 -8.965 ;
        RECT 28.165 -24.685 28.885 -23.965 ;
        RECT 17.940 -30.810 18.260 -30.490 ;
        RECT 18.340 -30.810 18.660 -30.490 ;
        RECT 18.740 -30.810 19.060 -30.490 ;
        RECT 19.140 -30.810 19.460 -30.490 ;
        RECT 19.540 -30.810 19.860 -30.490 ;
        RECT 19.940 -30.810 20.260 -30.490 ;
        RECT 20.340 -30.810 20.660 -30.490 ;
        RECT 20.740 -30.810 21.060 -30.490 ;
        RECT 21.140 -30.810 21.460 -30.490 ;
        RECT 21.540 -30.810 21.860 -30.490 ;
        RECT 21.940 -30.810 22.260 -30.490 ;
        RECT 22.340 -30.810 22.660 -30.490 ;
        RECT 22.740 -30.810 23.060 -30.490 ;
        RECT 23.140 -30.810 23.460 -30.490 ;
        RECT 23.540 -30.810 23.860 -30.490 ;
        RECT 23.940 -30.810 24.260 -30.490 ;
        RECT 24.340 -30.810 24.660 -30.490 ;
        RECT 24.740 -30.810 25.060 -30.490 ;
        RECT 25.140 -30.810 25.460 -30.490 ;
        RECT 25.540 -30.810 25.860 -30.490 ;
        RECT 25.940 -30.810 26.260 -30.490 ;
        RECT 26.340 -30.810 26.660 -30.490 ;
        RECT 26.740 -30.810 27.060 -30.490 ;
        RECT 27.140 -30.810 27.460 -30.490 ;
        RECT 27.540 -30.810 27.860 -30.490 ;
        RECT 27.940 -30.810 28.260 -30.490 ;
        RECT 28.340 -30.810 28.660 -30.490 ;
      LAYER met4 ;
        RECT 28.150 6.100 28.900 15.800 ;
        RECT 28.100 5.250 28.950 6.100 ;
        RECT 28.150 -8.900 28.900 5.250 ;
        RECT 28.100 -9.750 28.950 -8.900 ;
        RECT 28.150 -23.900 28.900 -9.750 ;
        RECT 28.100 -24.750 28.950 -23.900 ;
        RECT 28.150 -30.300 28.900 -24.750 ;
        RECT 17.700 -31.000 28.900 -30.300 ;
    END
  END PIX_OUT1
  PIN COL_SEL1
    ANTENNAGATEAREA 16.000000 ;
    PORT
      LAYER li1 ;
        RECT 16.100 -33.550 17.200 -32.450 ;
      LAYER mcon ;
        RECT 16.205 -33.445 17.095 -32.555 ;
      LAYER met1 ;
        RECT 16.100 -33.550 17.200 -32.450 ;
      LAYER via ;
        RECT 16.200 -33.450 17.100 -32.550 ;
      LAYER met2 ;
        RECT 16.100 -33.550 17.200 -32.450 ;
      LAYER via2 ;
        RECT 16.310 -33.340 16.990 -32.660 ;
      LAYER met3 ;
        RECT 16.100 -33.550 17.200 -32.450 ;
      LAYER via3 ;
        RECT 16.290 -33.360 17.010 -32.640 ;
      LAYER met4 ;
        RECT 16.100 -35.500 17.200 -32.450 ;
    END
  END COL_SEL1
  PIN PIX8_IN
    ANTENNAGATEAREA 1.050000 ;
    ANTENNADIFFAREA 0.294000 ;
    PORT
      LAYER li1 ;
        RECT 44.200 -18.050 44.650 -17.680 ;
        RECT 44.350 -19.400 44.650 -18.050 ;
        RECT 43.000 -19.650 44.650 -19.400 ;
        RECT 43.000 -19.950 43.650 -19.650 ;
        RECT 33.200 -27.550 33.900 -26.900 ;
        RECT 32.450 -27.850 33.900 -27.550 ;
      LAYER mcon ;
        RECT 43.060 -19.760 43.230 -19.590 ;
        RECT 43.420 -19.760 43.590 -19.590 ;
        RECT 33.465 -27.130 33.635 -26.960 ;
        RECT 33.465 -27.490 33.635 -27.320 ;
      LAYER met1 ;
        RECT 41.300 -19.950 43.700 -19.400 ;
        RECT 33.200 -27.600 33.900 -26.250 ;
      LAYER via ;
        RECT 41.400 -19.805 41.660 -19.545 ;
        RECT 41.720 -19.805 41.980 -19.545 ;
        RECT 42.040 -19.805 42.300 -19.545 ;
        RECT 33.260 -26.730 33.520 -26.470 ;
        RECT 33.580 -26.730 33.840 -26.470 ;
      LAYER met2 ;
        RECT 40.350 -20.050 42.450 -18.700 ;
        RECT 33.200 -26.900 34.650 -26.250 ;
      LAYER via2 ;
        RECT 40.435 -19.940 41.115 -18.860 ;
        RECT 33.385 -26.665 33.665 -26.385 ;
        RECT 33.785 -26.665 34.065 -26.385 ;
        RECT 34.185 -26.665 34.465 -26.385 ;
      LAYER met3 ;
        RECT 40.250 -20.150 42.500 -18.600 ;
        RECT 33.200 -26.750 34.650 -24.900 ;
      LAYER via3 ;
        RECT 40.390 -19.935 41.110 -18.815 ;
        RECT 33.590 -26.635 34.310 -25.115 ;
      LAYER met4 ;
        RECT 38.300 -20.350 42.100 -18.050 ;
        RECT 33.200 -26.750 34.650 -24.900 ;
      LAYER via4 ;
        RECT 40.060 -19.965 41.240 -18.785 ;
        RECT 33.360 -26.215 34.540 -25.035 ;
      LAYER met5 ;
        RECT 32.400 -27.600 42.600 -17.400 ;
    END
  END PIX8_IN
  PIN PIX_OUT2
    ANTENNADIFFAREA 6.400000 ;
    PORT
      LAYER li1 ;
        RECT 39.750 7.450 41.700 7.800 ;
        RECT 40.950 6.050 41.700 7.450 ;
        RECT 40.950 5.300 43.950 6.050 ;
        RECT 39.750 -7.550 41.700 -7.200 ;
        RECT 40.950 -8.950 41.700 -7.550 ;
        RECT 40.950 -9.700 43.950 -8.950 ;
        RECT 39.750 -22.550 41.700 -22.200 ;
        RECT 40.950 -23.950 41.700 -22.550 ;
        RECT 40.950 -24.700 43.950 -23.950 ;
        RECT 32.700 -31.900 40.700 -31.150 ;
      LAYER mcon ;
        RECT 43.260 5.410 43.790 5.940 ;
        RECT 43.260 -9.590 43.790 -9.060 ;
        RECT 43.260 -24.590 43.790 -24.060 ;
        RECT 32.835 -31.385 33.005 -31.215 ;
        RECT 33.195 -31.385 33.365 -31.215 ;
        RECT 33.555 -31.385 33.725 -31.215 ;
        RECT 33.915 -31.385 34.085 -31.215 ;
        RECT 34.275 -31.385 34.445 -31.215 ;
        RECT 34.635 -31.385 34.805 -31.215 ;
        RECT 34.995 -31.385 35.165 -31.215 ;
        RECT 35.355 -31.385 35.525 -31.215 ;
        RECT 35.715 -31.385 35.885 -31.215 ;
        RECT 36.075 -31.385 36.245 -31.215 ;
        RECT 36.435 -31.385 36.605 -31.215 ;
        RECT 36.795 -31.385 36.965 -31.215 ;
        RECT 37.155 -31.385 37.325 -31.215 ;
        RECT 37.515 -31.385 37.685 -31.215 ;
        RECT 37.875 -31.385 38.045 -31.215 ;
        RECT 38.235 -31.385 38.405 -31.215 ;
        RECT 38.595 -31.385 38.765 -31.215 ;
        RECT 38.955 -31.385 39.125 -31.215 ;
        RECT 39.315 -31.385 39.485 -31.215 ;
        RECT 39.675 -31.385 39.845 -31.215 ;
        RECT 40.035 -31.385 40.205 -31.215 ;
        RECT 40.395 -31.385 40.565 -31.215 ;
      LAYER met1 ;
        RECT 43.100 5.300 43.950 6.050 ;
        RECT 43.100 -9.700 43.950 -8.950 ;
        RECT 43.100 -24.700 43.950 -23.950 ;
        RECT 32.700 -31.500 40.700 -30.650 ;
      LAYER via ;
        RECT 43.235 5.385 43.815 5.965 ;
        RECT 43.235 -9.615 43.815 -9.035 ;
        RECT 43.235 -24.615 43.815 -24.035 ;
        RECT 32.890 -30.955 33.150 -30.695 ;
        RECT 33.210 -30.955 33.470 -30.695 ;
        RECT 33.530 -30.955 33.790 -30.695 ;
        RECT 33.850 -30.955 34.110 -30.695 ;
        RECT 34.170 -30.955 34.430 -30.695 ;
        RECT 34.490 -30.955 34.750 -30.695 ;
        RECT 34.810 -30.955 35.070 -30.695 ;
        RECT 35.130 -30.955 35.390 -30.695 ;
        RECT 35.450 -30.955 35.710 -30.695 ;
        RECT 35.770 -30.955 36.030 -30.695 ;
        RECT 36.090 -30.955 36.350 -30.695 ;
        RECT 36.410 -30.955 36.670 -30.695 ;
        RECT 36.730 -30.955 36.990 -30.695 ;
        RECT 37.050 -30.955 37.310 -30.695 ;
        RECT 37.370 -30.955 37.630 -30.695 ;
        RECT 37.690 -30.955 37.950 -30.695 ;
        RECT 38.010 -30.955 38.270 -30.695 ;
        RECT 38.330 -30.955 38.590 -30.695 ;
        RECT 38.650 -30.955 38.910 -30.695 ;
        RECT 38.970 -30.955 39.230 -30.695 ;
        RECT 39.290 -30.955 39.550 -30.695 ;
        RECT 39.610 -30.955 39.870 -30.695 ;
        RECT 39.930 -30.955 40.190 -30.695 ;
        RECT 40.250 -30.955 40.510 -30.695 ;
      LAYER met2 ;
        RECT 43.100 5.250 43.950 6.100 ;
        RECT 43.100 -9.750 43.950 -8.900 ;
        RECT 43.100 -24.750 43.950 -23.900 ;
        RECT 32.700 -31.000 43.900 -30.300 ;
      LAYER via2 ;
        RECT 43.185 5.335 43.865 6.015 ;
        RECT 43.185 -9.665 43.865 -8.985 ;
        RECT 43.185 -24.665 43.865 -23.985 ;
        RECT 32.960 -30.790 33.240 -30.510 ;
        RECT 33.360 -30.790 33.640 -30.510 ;
        RECT 33.760 -30.790 34.040 -30.510 ;
        RECT 34.160 -30.790 34.440 -30.510 ;
        RECT 34.560 -30.790 34.840 -30.510 ;
        RECT 34.960 -30.790 35.240 -30.510 ;
        RECT 35.360 -30.790 35.640 -30.510 ;
        RECT 35.760 -30.790 36.040 -30.510 ;
        RECT 36.160 -30.790 36.440 -30.510 ;
        RECT 36.560 -30.790 36.840 -30.510 ;
        RECT 36.960 -30.790 37.240 -30.510 ;
        RECT 37.360 -30.790 37.640 -30.510 ;
        RECT 37.760 -30.790 38.040 -30.510 ;
        RECT 38.160 -30.790 38.440 -30.510 ;
        RECT 38.560 -30.790 38.840 -30.510 ;
        RECT 38.960 -30.790 39.240 -30.510 ;
        RECT 39.360 -30.790 39.640 -30.510 ;
        RECT 39.760 -30.790 40.040 -30.510 ;
        RECT 40.160 -30.790 40.440 -30.510 ;
        RECT 40.560 -30.790 40.840 -30.510 ;
        RECT 40.960 -30.790 41.240 -30.510 ;
        RECT 41.360 -30.790 41.640 -30.510 ;
        RECT 41.760 -30.790 42.040 -30.510 ;
        RECT 42.160 -30.790 42.440 -30.510 ;
        RECT 42.560 -30.790 42.840 -30.510 ;
        RECT 42.960 -30.790 43.240 -30.510 ;
        RECT 43.360 -30.790 43.640 -30.510 ;
      LAYER met3 ;
        RECT 43.100 5.200 43.950 6.150 ;
        RECT 43.100 -9.800 43.950 -8.850 ;
        RECT 43.100 -24.800 43.950 -23.850 ;
        RECT 32.700 -31.000 43.900 -30.300 ;
      LAYER via3 ;
        RECT 43.165 5.315 43.885 6.035 ;
        RECT 43.165 -9.685 43.885 -8.965 ;
        RECT 43.165 -24.685 43.885 -23.965 ;
        RECT 32.940 -30.810 33.260 -30.490 ;
        RECT 33.340 -30.810 33.660 -30.490 ;
        RECT 33.740 -30.810 34.060 -30.490 ;
        RECT 34.140 -30.810 34.460 -30.490 ;
        RECT 34.540 -30.810 34.860 -30.490 ;
        RECT 34.940 -30.810 35.260 -30.490 ;
        RECT 35.340 -30.810 35.660 -30.490 ;
        RECT 35.740 -30.810 36.060 -30.490 ;
        RECT 36.140 -30.810 36.460 -30.490 ;
        RECT 36.540 -30.810 36.860 -30.490 ;
        RECT 36.940 -30.810 37.260 -30.490 ;
        RECT 37.340 -30.810 37.660 -30.490 ;
        RECT 37.740 -30.810 38.060 -30.490 ;
        RECT 38.140 -30.810 38.460 -30.490 ;
        RECT 38.540 -30.810 38.860 -30.490 ;
        RECT 38.940 -30.810 39.260 -30.490 ;
        RECT 39.340 -30.810 39.660 -30.490 ;
        RECT 39.740 -30.810 40.060 -30.490 ;
        RECT 40.140 -30.810 40.460 -30.490 ;
        RECT 40.540 -30.810 40.860 -30.490 ;
        RECT 40.940 -30.810 41.260 -30.490 ;
        RECT 41.340 -30.810 41.660 -30.490 ;
        RECT 41.740 -30.810 42.060 -30.490 ;
        RECT 42.140 -30.810 42.460 -30.490 ;
        RECT 42.540 -30.810 42.860 -30.490 ;
        RECT 42.940 -30.810 43.260 -30.490 ;
        RECT 43.340 -30.810 43.660 -30.490 ;
      LAYER met4 ;
        RECT 43.150 6.100 43.900 15.800 ;
        RECT 43.100 5.250 43.950 6.100 ;
        RECT 43.150 -8.900 43.900 5.250 ;
        RECT 43.100 -9.750 43.950 -8.900 ;
        RECT 43.150 -23.900 43.900 -9.750 ;
        RECT 43.100 -24.750 43.950 -23.900 ;
        RECT 43.150 -30.300 43.900 -24.750 ;
        RECT 32.700 -31.000 43.900 -30.300 ;
    END
  END PIX_OUT2
  PIN ARRAY_OUT
    ANTENNADIFFAREA 9.599999 ;
    PORT
      LAYER li1 ;
        RECT 2.700 -35.000 10.700 -34.000 ;
        RECT 17.700 -35.000 25.700 -34.000 ;
        RECT 32.700 -35.000 40.700 -34.000 ;
      LAYER mcon ;
        RECT 2.835 -34.835 3.005 -34.665 ;
        RECT 3.195 -34.835 3.365 -34.665 ;
        RECT 3.555 -34.835 3.725 -34.665 ;
        RECT 3.915 -34.835 4.085 -34.665 ;
        RECT 4.275 -34.835 4.445 -34.665 ;
        RECT 4.635 -34.835 4.805 -34.665 ;
        RECT 4.995 -34.835 5.165 -34.665 ;
        RECT 5.355 -34.835 5.525 -34.665 ;
        RECT 5.715 -34.835 5.885 -34.665 ;
        RECT 6.075 -34.835 6.245 -34.665 ;
        RECT 6.435 -34.835 6.605 -34.665 ;
        RECT 6.795 -34.835 6.965 -34.665 ;
        RECT 7.155 -34.835 7.325 -34.665 ;
        RECT 7.515 -34.835 7.685 -34.665 ;
        RECT 7.875 -34.835 8.045 -34.665 ;
        RECT 8.235 -34.835 8.405 -34.665 ;
        RECT 8.595 -34.835 8.765 -34.665 ;
        RECT 8.955 -34.835 9.125 -34.665 ;
        RECT 9.315 -34.835 9.485 -34.665 ;
        RECT 9.675 -34.835 9.845 -34.665 ;
        RECT 10.035 -34.835 10.205 -34.665 ;
        RECT 10.395 -34.835 10.565 -34.665 ;
        RECT 17.835 -34.835 18.005 -34.665 ;
        RECT 18.195 -34.835 18.365 -34.665 ;
        RECT 18.555 -34.835 18.725 -34.665 ;
        RECT 18.915 -34.835 19.085 -34.665 ;
        RECT 19.275 -34.835 19.445 -34.665 ;
        RECT 19.635 -34.835 19.805 -34.665 ;
        RECT 19.995 -34.835 20.165 -34.665 ;
        RECT 20.355 -34.835 20.525 -34.665 ;
        RECT 20.715 -34.835 20.885 -34.665 ;
        RECT 21.075 -34.835 21.245 -34.665 ;
        RECT 21.435 -34.835 21.605 -34.665 ;
        RECT 21.795 -34.835 21.965 -34.665 ;
        RECT 22.155 -34.835 22.325 -34.665 ;
        RECT 22.515 -34.835 22.685 -34.665 ;
        RECT 22.875 -34.835 23.045 -34.665 ;
        RECT 23.235 -34.835 23.405 -34.665 ;
        RECT 23.595 -34.835 23.765 -34.665 ;
        RECT 23.955 -34.835 24.125 -34.665 ;
        RECT 24.315 -34.835 24.485 -34.665 ;
        RECT 24.675 -34.835 24.845 -34.665 ;
        RECT 25.035 -34.835 25.205 -34.665 ;
        RECT 25.395 -34.835 25.565 -34.665 ;
        RECT 32.835 -34.835 33.005 -34.665 ;
        RECT 33.195 -34.835 33.365 -34.665 ;
        RECT 33.555 -34.835 33.725 -34.665 ;
        RECT 33.915 -34.835 34.085 -34.665 ;
        RECT 34.275 -34.835 34.445 -34.665 ;
        RECT 34.635 -34.835 34.805 -34.665 ;
        RECT 34.995 -34.835 35.165 -34.665 ;
        RECT 35.355 -34.835 35.525 -34.665 ;
        RECT 35.715 -34.835 35.885 -34.665 ;
        RECT 36.075 -34.835 36.245 -34.665 ;
        RECT 36.435 -34.835 36.605 -34.665 ;
        RECT 36.795 -34.835 36.965 -34.665 ;
        RECT 37.155 -34.835 37.325 -34.665 ;
        RECT 37.515 -34.835 37.685 -34.665 ;
        RECT 37.875 -34.835 38.045 -34.665 ;
        RECT 38.235 -34.835 38.405 -34.665 ;
        RECT 38.595 -34.835 38.765 -34.665 ;
        RECT 38.955 -34.835 39.125 -34.665 ;
        RECT 39.315 -34.835 39.485 -34.665 ;
        RECT 39.675 -34.835 39.845 -34.665 ;
        RECT 40.035 -34.835 40.205 -34.665 ;
        RECT 40.395 -34.835 40.565 -34.665 ;
      LAYER met1 ;
        RECT 2.700 -35.500 48.700 -34.500 ;
      LAYER via ;
        RECT 2.900 -35.290 48.600 -34.710 ;
      LAYER met2 ;
        RECT 2.700 -35.500 48.700 -34.500 ;
    END
  END ARRAY_OUT
  PIN COL_SEL2
    ANTENNAGATEAREA 16.000000 ;
    PORT
      LAYER li1 ;
        RECT 31.100 -33.550 32.200 -32.450 ;
      LAYER mcon ;
        RECT 31.205 -33.445 32.095 -32.555 ;
      LAYER met1 ;
        RECT 31.100 -33.550 32.200 -32.450 ;
      LAYER via ;
        RECT 31.200 -33.450 32.100 -32.550 ;
      LAYER met2 ;
        RECT 31.100 -33.550 32.200 -32.450 ;
      LAYER via2 ;
        RECT 31.310 -33.340 31.990 -32.660 ;
      LAYER met3 ;
        RECT 31.100 -33.550 32.200 -32.450 ;
      LAYER via3 ;
        RECT 31.290 -33.360 32.010 -32.640 ;
      LAYER met4 ;
        RECT 31.100 -35.500 32.200 -32.450 ;
    END
  END COL_SEL2
  OBS
      LAYER pwell ;
        RECT 3.870 7.670 5.130 11.380 ;
        RECT 9.620 9.280 10.880 10.480 ;
        RECT 9.620 7.370 11.880 9.280 ;
        RECT 18.870 7.670 20.130 11.380 ;
        RECT 24.620 9.280 25.880 10.480 ;
        RECT 24.620 7.370 26.880 9.280 ;
        RECT 33.870 7.670 35.130 11.380 ;
        RECT 39.620 9.280 40.880 10.480 ;
        RECT 39.620 7.370 41.880 9.280 ;
        RECT 3.870 -7.330 5.130 -3.620 ;
        RECT 9.620 -5.720 10.880 -4.520 ;
        RECT 9.620 -7.630 11.880 -5.720 ;
        RECT 18.870 -7.330 20.130 -3.620 ;
        RECT 24.620 -5.720 25.880 -4.520 ;
        RECT 24.620 -7.630 26.880 -5.720 ;
        RECT 33.870 -7.330 35.130 -3.620 ;
        RECT 39.620 -5.720 40.880 -4.520 ;
        RECT 39.620 -7.630 41.880 -5.720 ;
        RECT 3.870 -22.330 5.130 -18.620 ;
        RECT 9.620 -20.720 10.880 -19.520 ;
        RECT 9.620 -22.630 11.880 -20.720 ;
        RECT 18.870 -22.330 20.130 -18.620 ;
        RECT 24.620 -20.720 25.880 -19.520 ;
        RECT 24.620 -22.630 26.880 -20.720 ;
        RECT 33.870 -22.330 35.130 -18.620 ;
        RECT 39.620 -20.720 40.880 -19.520 ;
        RECT 39.620 -22.630 41.880 -20.720 ;
        RECT 2.570 -34.530 10.830 -31.370 ;
        RECT 17.570 -34.530 25.830 -31.370 ;
        RECT 32.570 -34.530 40.830 -31.370 ;
      LAYER li1 ;
        RECT 0.400 13.350 0.650 14.350 ;
        RECT 1.050 13.350 1.400 13.450 ;
        RECT 0.300 13.150 1.400 13.350 ;
        RECT 2.850 13.350 3.050 14.550 ;
        RECT 3.400 13.350 3.750 13.450 ;
        RECT 2.850 13.150 3.750 13.350 ;
        RECT 0.300 11.250 0.500 13.150 ;
        RECT 1.050 13.000 1.400 13.150 ;
        RECT 3.400 13.000 3.750 13.150 ;
        RECT 10.750 12.650 10.950 14.550 ;
        RECT 11.600 12.700 12.100 13.100 ;
        RECT 12.750 12.900 13.050 14.350 ;
        RECT 15.400 13.350 15.650 14.350 ;
        RECT 16.050 13.350 16.400 13.450 ;
        RECT 2.400 12.450 10.950 12.650 ;
        RECT 11.650 12.550 12.050 12.700 ;
        RECT 12.600 12.600 13.050 12.900 ;
        RECT 15.300 13.150 16.400 13.350 ;
        RECT 17.850 13.350 18.050 14.550 ;
        RECT 18.400 13.350 18.750 13.450 ;
        RECT 17.850 13.150 18.750 13.350 ;
        RECT 2.400 12.100 2.600 12.450 ;
        RECT 2.400 11.850 3.850 12.100 ;
        RECT 2.400 11.250 2.600 11.850 ;
        RECT 0.300 10.950 1.300 11.250 ;
        RECT 1.600 10.950 2.600 11.250 ;
        RECT 3.600 10.950 3.850 11.850 ;
        RECT 3.500 10.050 3.850 10.950 ;
        RECT 5.450 11.900 6.050 12.250 ;
        RECT 5.450 11.500 5.800 11.900 ;
        RECT 11.700 11.500 11.900 12.550 ;
        RECT 5.450 11.300 11.900 11.500 ;
        RECT 5.450 9.900 5.800 11.300 ;
        RECT 12.600 10.850 12.800 12.600 ;
        RECT 15.300 11.250 15.500 13.150 ;
        RECT 16.050 13.000 16.400 13.150 ;
        RECT 18.400 13.000 18.750 13.150 ;
        RECT 25.750 12.650 25.950 14.550 ;
        RECT 26.600 12.700 27.100 13.100 ;
        RECT 27.750 12.900 28.050 14.350 ;
        RECT 30.400 13.350 30.650 14.350 ;
        RECT 31.050 13.350 31.400 13.450 ;
        RECT 17.400 12.450 25.950 12.650 ;
        RECT 26.650 12.550 27.050 12.700 ;
        RECT 27.600 12.600 28.050 12.900 ;
        RECT 30.300 13.150 31.400 13.350 ;
        RECT 32.850 13.350 33.050 14.550 ;
        RECT 33.400 13.350 33.750 13.450 ;
        RECT 32.850 13.150 33.750 13.350 ;
        RECT 17.400 12.100 17.600 12.450 ;
        RECT 17.400 11.850 18.850 12.100 ;
        RECT 17.400 11.250 17.600 11.850 ;
        RECT 15.300 10.950 16.300 11.250 ;
        RECT 16.600 10.950 17.600 11.250 ;
        RECT 18.600 10.950 18.850 11.850 ;
        RECT 10.950 10.650 12.800 10.850 ;
        RECT 10.950 10.100 11.200 10.650 ;
        RECT 4.100 9.850 5.800 9.900 ;
        RECT 4.000 9.550 5.800 9.850 ;
        RECT 10.900 9.750 11.250 10.100 ;
        RECT 18.500 10.050 18.850 10.950 ;
        RECT 20.450 11.900 21.050 12.250 ;
        RECT 20.450 11.500 20.800 11.900 ;
        RECT 26.700 11.500 26.900 12.550 ;
        RECT 20.450 11.300 26.900 11.500 ;
        RECT 20.450 9.900 20.800 11.300 ;
        RECT 27.600 10.850 27.800 12.600 ;
        RECT 30.300 11.250 30.500 13.150 ;
        RECT 31.050 13.000 31.400 13.150 ;
        RECT 33.400 13.000 33.750 13.150 ;
        RECT 40.750 12.650 40.950 14.550 ;
        RECT 41.600 12.700 42.100 13.100 ;
        RECT 42.750 12.900 43.050 14.350 ;
        RECT 32.400 12.450 40.950 12.650 ;
        RECT 41.650 12.550 42.050 12.700 ;
        RECT 42.600 12.600 43.050 12.900 ;
        RECT 32.400 12.100 32.600 12.450 ;
        RECT 32.400 11.850 33.850 12.100 ;
        RECT 32.400 11.250 32.600 11.850 ;
        RECT 30.300 10.950 31.300 11.250 ;
        RECT 31.600 10.950 32.600 11.250 ;
        RECT 33.600 10.950 33.850 11.850 ;
        RECT 25.950 10.650 27.800 10.850 ;
        RECT 25.950 10.100 26.200 10.650 ;
        RECT 19.100 9.850 20.800 9.900 ;
        RECT 10.950 9.650 11.200 9.750 ;
        RECT 19.000 9.550 20.800 9.850 ;
        RECT 25.900 9.750 26.250 10.100 ;
        RECT 33.500 10.050 33.850 10.950 ;
        RECT 35.450 11.900 36.050 12.250 ;
        RECT 35.450 11.500 35.800 11.900 ;
        RECT 41.700 11.500 41.900 12.550 ;
        RECT 35.450 11.300 41.900 11.500 ;
        RECT 35.450 9.900 35.800 11.300 ;
        RECT 42.600 10.850 42.800 12.600 ;
        RECT 40.950 10.650 42.800 10.850 ;
        RECT 40.950 10.100 41.200 10.650 ;
        RECT 34.100 9.850 35.800 9.900 ;
        RECT 25.950 9.650 26.200 9.750 ;
        RECT 34.000 9.550 35.800 9.850 ;
        RECT 40.900 9.750 41.250 10.100 ;
        RECT 40.950 9.650 41.200 9.750 ;
        RECT 4.100 9.500 5.800 9.550 ;
        RECT 19.100 9.500 20.800 9.550 ;
        RECT 34.100 9.500 35.800 9.550 ;
        RECT 1.300 2.400 1.600 9.400 ;
        RECT 16.300 2.400 16.600 9.400 ;
        RECT 31.300 2.400 31.600 9.400 ;
        RECT 1.300 1.750 1.550 2.400 ;
        RECT 16.300 1.750 16.550 2.400 ;
        RECT 31.300 1.750 31.550 2.400 ;
        RECT 1.250 0.550 1.550 1.750 ;
        RECT 16.250 0.550 16.550 1.750 ;
        RECT 31.250 0.550 31.550 1.750 ;
        RECT 0.400 -1.650 0.650 -0.650 ;
        RECT 1.050 -1.650 1.400 -1.550 ;
        RECT 0.300 -1.850 1.400 -1.650 ;
        RECT 2.850 -1.650 3.050 -0.450 ;
        RECT 3.400 -1.650 3.750 -1.550 ;
        RECT 2.850 -1.850 3.750 -1.650 ;
        RECT 0.300 -3.750 0.500 -1.850 ;
        RECT 1.050 -2.000 1.400 -1.850 ;
        RECT 3.400 -2.000 3.750 -1.850 ;
        RECT 10.750 -2.350 10.950 -0.450 ;
        RECT 11.600 -2.300 12.100 -1.900 ;
        RECT 12.750 -2.100 13.050 -0.650 ;
        RECT 15.400 -1.650 15.650 -0.650 ;
        RECT 16.050 -1.650 16.400 -1.550 ;
        RECT 2.400 -2.550 10.950 -2.350 ;
        RECT 11.650 -2.450 12.050 -2.300 ;
        RECT 12.600 -2.400 13.050 -2.100 ;
        RECT 15.300 -1.850 16.400 -1.650 ;
        RECT 17.850 -1.650 18.050 -0.450 ;
        RECT 18.400 -1.650 18.750 -1.550 ;
        RECT 17.850 -1.850 18.750 -1.650 ;
        RECT 2.400 -2.900 2.600 -2.550 ;
        RECT 2.400 -3.150 3.850 -2.900 ;
        RECT 2.400 -3.750 2.600 -3.150 ;
        RECT 0.300 -4.050 1.300 -3.750 ;
        RECT 1.600 -4.050 2.600 -3.750 ;
        RECT 3.600 -4.050 3.850 -3.150 ;
        RECT 3.500 -4.950 3.850 -4.050 ;
        RECT 5.450 -3.100 6.050 -2.750 ;
        RECT 5.450 -3.500 5.800 -3.100 ;
        RECT 11.700 -3.500 11.900 -2.450 ;
        RECT 5.450 -3.700 11.900 -3.500 ;
        RECT 5.450 -5.100 5.800 -3.700 ;
        RECT 12.600 -4.150 12.800 -2.400 ;
        RECT 15.300 -3.750 15.500 -1.850 ;
        RECT 16.050 -2.000 16.400 -1.850 ;
        RECT 18.400 -2.000 18.750 -1.850 ;
        RECT 25.750 -2.350 25.950 -0.450 ;
        RECT 26.600 -2.300 27.100 -1.900 ;
        RECT 27.750 -2.100 28.050 -0.650 ;
        RECT 30.400 -1.650 30.650 -0.650 ;
        RECT 31.050 -1.650 31.400 -1.550 ;
        RECT 17.400 -2.550 25.950 -2.350 ;
        RECT 26.650 -2.450 27.050 -2.300 ;
        RECT 27.600 -2.400 28.050 -2.100 ;
        RECT 30.300 -1.850 31.400 -1.650 ;
        RECT 32.850 -1.650 33.050 -0.450 ;
        RECT 33.400 -1.650 33.750 -1.550 ;
        RECT 32.850 -1.850 33.750 -1.650 ;
        RECT 17.400 -2.900 17.600 -2.550 ;
        RECT 17.400 -3.150 18.850 -2.900 ;
        RECT 17.400 -3.750 17.600 -3.150 ;
        RECT 15.300 -4.050 16.300 -3.750 ;
        RECT 16.600 -4.050 17.600 -3.750 ;
        RECT 18.600 -4.050 18.850 -3.150 ;
        RECT 10.950 -4.350 12.800 -4.150 ;
        RECT 10.950 -4.900 11.200 -4.350 ;
        RECT 4.100 -5.150 5.800 -5.100 ;
        RECT 4.000 -5.450 5.800 -5.150 ;
        RECT 10.900 -5.250 11.250 -4.900 ;
        RECT 18.500 -4.950 18.850 -4.050 ;
        RECT 20.450 -3.100 21.050 -2.750 ;
        RECT 20.450 -3.500 20.800 -3.100 ;
        RECT 26.700 -3.500 26.900 -2.450 ;
        RECT 20.450 -3.700 26.900 -3.500 ;
        RECT 20.450 -5.100 20.800 -3.700 ;
        RECT 27.600 -4.150 27.800 -2.400 ;
        RECT 30.300 -3.750 30.500 -1.850 ;
        RECT 31.050 -2.000 31.400 -1.850 ;
        RECT 33.400 -2.000 33.750 -1.850 ;
        RECT 40.750 -2.350 40.950 -0.450 ;
        RECT 41.600 -2.300 42.100 -1.900 ;
        RECT 42.750 -2.100 43.050 -0.650 ;
        RECT 32.400 -2.550 40.950 -2.350 ;
        RECT 41.650 -2.450 42.050 -2.300 ;
        RECT 42.600 -2.400 43.050 -2.100 ;
        RECT 32.400 -2.900 32.600 -2.550 ;
        RECT 32.400 -3.150 33.850 -2.900 ;
        RECT 32.400 -3.750 32.600 -3.150 ;
        RECT 30.300 -4.050 31.300 -3.750 ;
        RECT 31.600 -4.050 32.600 -3.750 ;
        RECT 33.600 -4.050 33.850 -3.150 ;
        RECT 25.950 -4.350 27.800 -4.150 ;
        RECT 25.950 -4.900 26.200 -4.350 ;
        RECT 19.100 -5.150 20.800 -5.100 ;
        RECT 10.950 -5.350 11.200 -5.250 ;
        RECT 19.000 -5.450 20.800 -5.150 ;
        RECT 25.900 -5.250 26.250 -4.900 ;
        RECT 33.500 -4.950 33.850 -4.050 ;
        RECT 35.450 -3.100 36.050 -2.750 ;
        RECT 35.450 -3.500 35.800 -3.100 ;
        RECT 41.700 -3.500 41.900 -2.450 ;
        RECT 35.450 -3.700 41.900 -3.500 ;
        RECT 35.450 -5.100 35.800 -3.700 ;
        RECT 42.600 -4.150 42.800 -2.400 ;
        RECT 40.950 -4.350 42.800 -4.150 ;
        RECT 40.950 -4.900 41.200 -4.350 ;
        RECT 34.100 -5.150 35.800 -5.100 ;
        RECT 25.950 -5.350 26.200 -5.250 ;
        RECT 34.000 -5.450 35.800 -5.150 ;
        RECT 40.900 -5.250 41.250 -4.900 ;
        RECT 40.950 -5.350 41.200 -5.250 ;
        RECT 4.100 -5.500 5.800 -5.450 ;
        RECT 19.100 -5.500 20.800 -5.450 ;
        RECT 34.100 -5.500 35.800 -5.450 ;
        RECT 1.300 -12.600 1.600 -5.600 ;
        RECT 16.300 -12.600 16.600 -5.600 ;
        RECT 31.300 -12.600 31.600 -5.600 ;
        RECT 1.300 -13.250 1.550 -12.600 ;
        RECT 16.300 -13.250 16.550 -12.600 ;
        RECT 31.300 -13.250 31.550 -12.600 ;
        RECT 1.250 -14.450 1.550 -13.250 ;
        RECT 16.250 -14.450 16.550 -13.250 ;
        RECT 31.250 -14.450 31.550 -13.250 ;
        RECT 0.400 -16.650 0.650 -15.650 ;
        RECT 1.050 -16.650 1.400 -16.550 ;
        RECT 0.300 -16.850 1.400 -16.650 ;
        RECT 2.850 -16.650 3.050 -15.450 ;
        RECT 3.400 -16.650 3.750 -16.550 ;
        RECT 2.850 -16.850 3.750 -16.650 ;
        RECT 0.300 -18.750 0.500 -16.850 ;
        RECT 1.050 -17.000 1.400 -16.850 ;
        RECT 3.400 -17.000 3.750 -16.850 ;
        RECT 10.750 -17.350 10.950 -15.450 ;
        RECT 11.600 -17.300 12.100 -16.900 ;
        RECT 12.750 -17.100 13.050 -15.650 ;
        RECT 15.400 -16.650 15.650 -15.650 ;
        RECT 16.050 -16.650 16.400 -16.550 ;
        RECT 2.400 -17.550 10.950 -17.350 ;
        RECT 11.650 -17.450 12.050 -17.300 ;
        RECT 12.600 -17.400 13.050 -17.100 ;
        RECT 15.300 -16.850 16.400 -16.650 ;
        RECT 17.850 -16.650 18.050 -15.450 ;
        RECT 18.400 -16.650 18.750 -16.550 ;
        RECT 17.850 -16.850 18.750 -16.650 ;
        RECT 2.400 -17.900 2.600 -17.550 ;
        RECT 2.400 -18.150 3.850 -17.900 ;
        RECT 2.400 -18.750 2.600 -18.150 ;
        RECT 0.300 -19.050 1.300 -18.750 ;
        RECT 1.600 -19.050 2.600 -18.750 ;
        RECT 3.600 -19.050 3.850 -18.150 ;
        RECT 3.500 -19.950 3.850 -19.050 ;
        RECT 5.450 -18.100 6.050 -17.750 ;
        RECT 5.450 -18.500 5.800 -18.100 ;
        RECT 11.700 -18.500 11.900 -17.450 ;
        RECT 5.450 -18.700 11.900 -18.500 ;
        RECT 5.450 -20.100 5.800 -18.700 ;
        RECT 12.600 -19.150 12.800 -17.400 ;
        RECT 15.300 -18.750 15.500 -16.850 ;
        RECT 16.050 -17.000 16.400 -16.850 ;
        RECT 18.400 -17.000 18.750 -16.850 ;
        RECT 25.750 -17.350 25.950 -15.450 ;
        RECT 26.600 -17.300 27.100 -16.900 ;
        RECT 27.750 -17.100 28.050 -15.650 ;
        RECT 30.400 -16.650 30.650 -15.650 ;
        RECT 31.050 -16.650 31.400 -16.550 ;
        RECT 17.400 -17.550 25.950 -17.350 ;
        RECT 26.650 -17.450 27.050 -17.300 ;
        RECT 27.600 -17.400 28.050 -17.100 ;
        RECT 30.300 -16.850 31.400 -16.650 ;
        RECT 32.850 -16.650 33.050 -15.450 ;
        RECT 33.400 -16.650 33.750 -16.550 ;
        RECT 32.850 -16.850 33.750 -16.650 ;
        RECT 17.400 -17.900 17.600 -17.550 ;
        RECT 17.400 -18.150 18.850 -17.900 ;
        RECT 17.400 -18.750 17.600 -18.150 ;
        RECT 15.300 -19.050 16.300 -18.750 ;
        RECT 16.600 -19.050 17.600 -18.750 ;
        RECT 18.600 -19.050 18.850 -18.150 ;
        RECT 10.950 -19.350 12.800 -19.150 ;
        RECT 10.950 -19.900 11.200 -19.350 ;
        RECT 4.100 -20.150 5.800 -20.100 ;
        RECT 4.000 -20.450 5.800 -20.150 ;
        RECT 10.900 -20.250 11.250 -19.900 ;
        RECT 18.500 -19.950 18.850 -19.050 ;
        RECT 20.450 -18.100 21.050 -17.750 ;
        RECT 20.450 -18.500 20.800 -18.100 ;
        RECT 26.700 -18.500 26.900 -17.450 ;
        RECT 20.450 -18.700 26.900 -18.500 ;
        RECT 20.450 -20.100 20.800 -18.700 ;
        RECT 27.600 -19.150 27.800 -17.400 ;
        RECT 30.300 -18.750 30.500 -16.850 ;
        RECT 31.050 -17.000 31.400 -16.850 ;
        RECT 33.400 -17.000 33.750 -16.850 ;
        RECT 40.750 -17.350 40.950 -15.450 ;
        RECT 41.600 -17.300 42.100 -16.900 ;
        RECT 42.750 -17.100 43.050 -15.650 ;
        RECT 32.400 -17.550 40.950 -17.350 ;
        RECT 41.650 -17.450 42.050 -17.300 ;
        RECT 42.600 -17.400 43.050 -17.100 ;
        RECT 32.400 -17.900 32.600 -17.550 ;
        RECT 32.400 -18.150 33.850 -17.900 ;
        RECT 32.400 -18.750 32.600 -18.150 ;
        RECT 30.300 -19.050 31.300 -18.750 ;
        RECT 31.600 -19.050 32.600 -18.750 ;
        RECT 33.600 -19.050 33.850 -18.150 ;
        RECT 25.950 -19.350 27.800 -19.150 ;
        RECT 25.950 -19.900 26.200 -19.350 ;
        RECT 19.100 -20.150 20.800 -20.100 ;
        RECT 10.950 -20.350 11.200 -20.250 ;
        RECT 19.000 -20.450 20.800 -20.150 ;
        RECT 25.900 -20.250 26.250 -19.900 ;
        RECT 33.500 -19.950 33.850 -19.050 ;
        RECT 35.450 -18.100 36.050 -17.750 ;
        RECT 35.450 -18.500 35.800 -18.100 ;
        RECT 41.700 -18.500 41.900 -17.450 ;
        RECT 35.450 -18.700 41.900 -18.500 ;
        RECT 35.450 -20.100 35.800 -18.700 ;
        RECT 42.600 -19.150 42.800 -17.400 ;
        RECT 40.950 -19.350 42.800 -19.150 ;
        RECT 40.950 -19.900 41.200 -19.350 ;
        RECT 34.100 -20.150 35.800 -20.100 ;
        RECT 25.950 -20.350 26.200 -20.250 ;
        RECT 34.000 -20.450 35.800 -20.150 ;
        RECT 40.900 -20.250 41.250 -19.900 ;
        RECT 40.950 -20.350 41.200 -20.250 ;
        RECT 4.100 -20.500 5.800 -20.450 ;
        RECT 19.100 -20.500 20.800 -20.450 ;
        RECT 34.100 -20.500 35.800 -20.450 ;
        RECT 1.300 -27.600 1.600 -20.600 ;
        RECT 16.300 -27.600 16.600 -20.600 ;
        RECT 31.300 -27.600 31.600 -20.600 ;
        RECT 1.300 -28.250 1.550 -27.600 ;
        RECT 16.300 -28.250 16.550 -27.600 ;
        RECT 31.300 -28.250 31.550 -27.600 ;
        RECT 1.250 -29.450 1.550 -28.250 ;
        RECT 16.250 -29.450 16.550 -28.250 ;
        RECT 31.250 -29.450 31.550 -28.250 ;
      LAYER mcon ;
        RECT 5.540 10.590 5.710 10.760 ;
        RECT 20.540 10.590 20.710 10.760 ;
        RECT 35.540 10.590 35.710 10.760 ;
        RECT 5.540 -4.410 5.710 -4.240 ;
        RECT 20.540 -4.410 20.710 -4.240 ;
        RECT 35.540 -4.410 35.710 -4.240 ;
        RECT 5.540 -19.410 5.710 -19.240 ;
        RECT 20.540 -19.410 20.710 -19.240 ;
        RECT 35.540 -19.410 35.710 -19.240 ;
      LAYER met1 ;
        RECT 5.450 10.800 5.800 10.900 ;
        RECT 6.400 10.800 6.800 10.900 ;
        RECT 5.450 10.550 6.800 10.800 ;
        RECT 20.450 10.800 20.800 10.900 ;
        RECT 21.400 10.800 21.800 10.900 ;
        RECT 20.450 10.550 21.800 10.800 ;
        RECT 35.450 10.800 35.800 10.900 ;
        RECT 36.400 10.800 36.800 10.900 ;
        RECT 35.450 10.550 36.800 10.800 ;
        RECT 5.450 10.450 5.800 10.550 ;
        RECT 20.450 10.450 20.800 10.550 ;
        RECT 35.450 10.450 35.800 10.550 ;
        RECT 5.450 -4.200 5.800 -4.100 ;
        RECT 6.400 -4.200 6.800 -4.100 ;
        RECT 5.450 -4.450 6.800 -4.200 ;
        RECT 20.450 -4.200 20.800 -4.100 ;
        RECT 21.400 -4.200 21.800 -4.100 ;
        RECT 20.450 -4.450 21.800 -4.200 ;
        RECT 35.450 -4.200 35.800 -4.100 ;
        RECT 36.400 -4.200 36.800 -4.100 ;
        RECT 35.450 -4.450 36.800 -4.200 ;
        RECT 5.450 -4.550 5.800 -4.450 ;
        RECT 20.450 -4.550 20.800 -4.450 ;
        RECT 35.450 -4.550 35.800 -4.450 ;
        RECT 5.450 -19.200 5.800 -19.100 ;
        RECT 6.400 -19.200 6.800 -19.100 ;
        RECT 5.450 -19.450 6.800 -19.200 ;
        RECT 20.450 -19.200 20.800 -19.100 ;
        RECT 21.400 -19.200 21.800 -19.100 ;
        RECT 20.450 -19.450 21.800 -19.200 ;
        RECT 35.450 -19.200 35.800 -19.100 ;
        RECT 36.400 -19.200 36.800 -19.100 ;
        RECT 35.450 -19.450 36.800 -19.200 ;
        RECT 5.450 -19.550 5.800 -19.450 ;
        RECT 20.450 -19.550 20.800 -19.450 ;
        RECT 35.450 -19.550 35.800 -19.450 ;
      LAYER via ;
        RECT 6.470 10.620 6.730 10.880 ;
        RECT 21.470 10.620 21.730 10.880 ;
        RECT 36.470 10.620 36.730 10.880 ;
        RECT 6.470 -4.380 6.730 -4.120 ;
        RECT 21.470 -4.380 21.730 -4.120 ;
        RECT 36.470 -4.380 36.730 -4.120 ;
        RECT 6.470 -19.380 6.730 -19.120 ;
        RECT 21.470 -19.380 21.730 -19.120 ;
        RECT 36.470 -19.380 36.730 -19.120 ;
      LAYER met2 ;
        RECT 6.400 10.500 6.800 11.500 ;
        RECT 21.400 10.500 21.800 11.500 ;
        RECT 36.400 10.500 36.800 11.500 ;
        RECT 6.400 -4.500 6.800 -3.500 ;
        RECT 21.400 -4.500 21.800 -3.500 ;
        RECT 36.400 -4.500 36.800 -3.500 ;
        RECT 6.400 -19.500 6.800 -18.500 ;
        RECT 21.400 -19.500 21.800 -18.500 ;
        RECT 36.400 -19.500 36.800 -18.500 ;
      LAYER via2 ;
        RECT 6.485 11.110 6.765 11.390 ;
        RECT 21.485 11.110 21.765 11.390 ;
        RECT 36.485 11.110 36.765 11.390 ;
        RECT 6.485 -3.890 6.765 -3.610 ;
        RECT 21.485 -3.890 21.765 -3.610 ;
        RECT 36.485 -3.890 36.765 -3.610 ;
        RECT 6.485 -18.890 6.765 -18.610 ;
        RECT 21.485 -18.890 21.765 -18.610 ;
        RECT 36.485 -18.890 36.765 -18.610 ;
      LAYER met3 ;
        RECT 7.550 11.450 9.850 11.600 ;
        RECT 22.550 11.450 24.850 11.600 ;
        RECT 37.550 11.450 39.850 11.600 ;
        RECT 6.400 11.400 9.850 11.450 ;
        RECT 21.400 11.400 24.850 11.450 ;
        RECT 36.400 11.400 39.850 11.450 ;
        RECT 6.350 11.050 9.850 11.400 ;
        RECT 21.350 11.050 24.850 11.400 ;
        RECT 36.350 11.050 39.850 11.400 ;
        RECT 6.400 11.000 9.850 11.050 ;
        RECT 21.400 11.000 24.850 11.050 ;
        RECT 36.400 11.000 39.850 11.050 ;
        RECT 7.550 9.300 9.850 11.000 ;
        RECT 22.550 9.300 24.850 11.000 ;
        RECT 37.550 9.300 39.850 11.000 ;
        RECT 7.550 -3.550 9.850 -3.400 ;
        RECT 22.550 -3.550 24.850 -3.400 ;
        RECT 37.550 -3.550 39.850 -3.400 ;
        RECT 6.400 -3.600 9.850 -3.550 ;
        RECT 21.400 -3.600 24.850 -3.550 ;
        RECT 36.400 -3.600 39.850 -3.550 ;
        RECT 6.350 -3.950 9.850 -3.600 ;
        RECT 21.350 -3.950 24.850 -3.600 ;
        RECT 36.350 -3.950 39.850 -3.600 ;
        RECT 6.400 -4.000 9.850 -3.950 ;
        RECT 21.400 -4.000 24.850 -3.950 ;
        RECT 36.400 -4.000 39.850 -3.950 ;
        RECT 7.550 -5.700 9.850 -4.000 ;
        RECT 22.550 -5.700 24.850 -4.000 ;
        RECT 37.550 -5.700 39.850 -4.000 ;
        RECT 7.550 -18.550 9.850 -18.400 ;
        RECT 22.550 -18.550 24.850 -18.400 ;
        RECT 37.550 -18.550 39.850 -18.400 ;
        RECT 6.400 -18.600 9.850 -18.550 ;
        RECT 21.400 -18.600 24.850 -18.550 ;
        RECT 36.400 -18.600 39.850 -18.550 ;
        RECT 6.350 -18.950 9.850 -18.600 ;
        RECT 21.350 -18.950 24.850 -18.600 ;
        RECT 36.350 -18.950 39.850 -18.600 ;
        RECT 6.400 -19.000 9.850 -18.950 ;
        RECT 21.400 -19.000 24.850 -18.950 ;
        RECT 36.400 -19.000 39.850 -18.950 ;
        RECT 7.550 -20.700 9.850 -19.000 ;
        RECT 22.550 -20.700 24.850 -19.000 ;
        RECT 37.550 -20.700 39.850 -19.000 ;
      LAYER met5 ;
        RECT -10.000 14.200 45.800 15.800 ;
        RECT -0.800 0.800 0.800 14.200 ;
        RECT 14.200 0.800 15.800 14.200 ;
        RECT 29.200 0.800 30.800 14.200 ;
        RECT 44.200 0.800 45.800 14.200 ;
        RECT -0.800 -0.800 45.800 0.800 ;
        RECT -0.800 -14.200 0.800 -0.800 ;
        RECT 14.200 -14.200 15.800 -0.800 ;
        RECT 29.200 -14.200 30.800 -0.800 ;
        RECT 44.200 -14.200 45.800 -0.800 ;
        RECT -0.800 -15.800 45.800 -14.200 ;
        RECT -0.800 -29.200 0.800 -15.800 ;
        RECT 14.200 -29.200 15.800 -15.800 ;
        RECT 29.200 -29.200 30.800 -15.800 ;
        RECT 44.200 -29.200 45.800 -15.800 ;
        RECT -0.800 -30.800 45.800 -29.200 ;
  END
END pixel_array#0
END LIBRARY

