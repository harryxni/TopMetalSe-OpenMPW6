magic
tech sky130A
magscale 1 2
timestamp 1654648307
<< error_p >>
rect 21517 15656 21551 16232
rect 21635 15656 21669 16232
rect 21753 15656 21787 16232
rect 21871 15656 21905 16232
rect 21989 15656 22023 16232
rect 22107 15656 22141 16232
rect 22225 15656 22259 16232
rect 22343 15656 22377 16232
rect 22461 15656 22495 16232
rect 22579 15656 22613 16232
rect 22697 15656 22731 16232
rect 22815 15656 22849 16232
rect 22933 15656 22967 16232
rect 23051 15656 23085 16232
rect 23169 15656 23203 16232
rect 23287 15656 23321 16232
rect 23405 15656 23439 16232
rect 23523 15656 23557 16232
rect 23641 15656 23675 16232
rect 23759 15656 23793 16232
rect 23877 15656 23911 16232
rect 23995 15656 24029 16232
rect 24113 15656 24147 16232
rect 24231 15656 24265 16232
rect 25640 15656 25674 16232
rect 25758 15656 25792 16232
rect 25876 15656 25910 16232
rect 25994 15656 26028 16232
rect 26112 15656 26146 16232
rect 26230 15656 26264 16232
rect 26348 15656 26382 16232
rect 26466 15656 26500 16232
rect 26584 15656 26618 16232
rect 26702 15656 26736 16232
rect 26820 15656 26854 16232
rect 26938 15656 26972 16232
rect 27056 15656 27090 16232
rect 27174 15656 27208 16232
rect 27292 15656 27326 16232
rect 27410 15656 27444 16232
rect 27528 15656 27562 16232
rect 27646 15656 27680 16232
rect 27764 15656 27798 16232
rect 27882 15656 27916 16232
rect 28000 15656 28034 16232
rect 28118 15656 28152 16232
rect 28236 15656 28270 16232
rect 28354 15656 28388 16232
rect 29763 15656 29797 16232
rect 29881 15656 29915 16232
rect 29999 15656 30033 16232
rect 30117 15656 30151 16232
rect 30235 15656 30269 16232
rect 30353 15656 30387 16232
rect 30471 15656 30505 16232
rect 30589 15656 30623 16232
rect 30707 15656 30741 16232
rect 30825 15656 30859 16232
rect 30943 15656 30977 16232
rect 31061 15656 31095 16232
rect 31179 15656 31213 16232
rect 31297 15656 31331 16232
rect 31415 15656 31449 16232
rect 31533 15656 31567 16232
rect 31651 15656 31685 16232
rect 31769 15656 31803 16232
rect 31887 15656 31921 16232
rect 32005 15656 32039 16232
rect 32123 15656 32157 16232
rect 32241 15656 32275 16232
rect 32359 15656 32393 16232
rect 32477 15656 32511 16232
rect 16704 14897 19543 14931
rect 16777 14160 16811 14736
rect 16895 14160 16929 14736
rect 17013 14160 17047 14736
rect 17131 14160 17165 14736
rect 17249 14160 17283 14736
rect 17367 14160 17401 14736
rect 17485 14160 17519 14736
rect 17603 14160 17637 14736
rect 17721 14160 17755 14736
rect 17839 14160 17873 14736
rect 17957 14160 17991 14736
rect 18075 14160 18109 14736
rect 18193 14160 18227 14736
rect 18311 14160 18345 14736
rect 18429 14160 18463 14736
rect 18547 14160 18581 14736
rect 18665 14160 18699 14736
rect 18783 14160 18817 14736
rect 18901 14160 18935 14736
rect 19019 14160 19053 14736
rect 19137 14160 19171 14736
rect 19255 14160 19289 14736
rect 19373 14160 19407 14736
rect 19491 14160 19525 14736
rect 16777 13324 16811 13900
rect 16895 13324 16929 13900
rect 17013 13324 17047 13900
rect 17131 13324 17165 13900
rect 17249 13324 17283 13900
rect 17367 13324 17401 13900
rect 17485 13324 17519 13900
rect 17603 13324 17637 13900
rect 17721 13324 17755 13900
rect 17839 13324 17873 13900
rect 17957 13324 17991 13900
rect 18075 13324 18109 13900
rect 18193 13324 18227 13900
rect 18311 13324 18345 13900
rect 18429 13324 18463 13900
rect 18547 13324 18581 13900
rect 18665 13324 18699 13900
rect 18783 13324 18817 13900
rect 18901 13324 18935 13900
rect 19019 13324 19053 13900
rect 19137 13324 19171 13900
rect 19255 13324 19289 13900
rect 19373 13324 19407 13900
rect 19491 13324 19525 13900
rect 19605 13225 19639 14835
rect 21281 14820 21315 15396
rect 21399 14820 21433 15396
rect 21517 14820 21551 15396
rect 21635 14820 21669 15396
rect 21753 14820 21787 15396
rect 21871 14820 21905 15396
rect 21989 14820 22023 15396
rect 22107 14820 22141 15396
rect 22225 14820 22259 15396
rect 22343 14820 22377 15396
rect 22461 14820 22495 15396
rect 22579 14820 22613 15396
rect 22697 14820 22731 15396
rect 22815 14820 22849 15396
rect 22933 14820 22967 15396
rect 23051 14820 23085 15396
rect 23169 14820 23203 15396
rect 23287 14820 23321 15396
rect 23405 14820 23439 15396
rect 23523 14820 23557 15396
rect 23641 14820 23675 15396
rect 23759 14820 23793 15396
rect 23877 14820 23911 15396
rect 23995 14820 24029 15396
rect 24113 14820 24147 15396
rect 24231 14820 24265 15396
rect 25404 14820 25438 15396
rect 25522 14820 25556 15396
rect 25640 14820 25674 15396
rect 25758 14820 25792 15396
rect 25876 14820 25910 15396
rect 25994 14820 26028 15396
rect 26112 14820 26146 15396
rect 26230 14820 26264 15396
rect 26348 14820 26382 15396
rect 26466 14820 26500 15396
rect 26584 14820 26618 15396
rect 26702 14820 26736 15396
rect 26820 14820 26854 15396
rect 26938 14820 26972 15396
rect 27056 14820 27090 15396
rect 27174 14820 27208 15396
rect 27292 14820 27326 15396
rect 27410 14820 27444 15396
rect 27528 14820 27562 15396
rect 27646 14820 27680 15396
rect 27764 14820 27798 15396
rect 27882 14820 27916 15396
rect 28000 14820 28034 15396
rect 28118 14820 28152 15396
rect 28236 14820 28270 15396
rect 28354 14820 28388 15396
rect 29527 14820 29561 15396
rect 29645 14820 29679 15396
rect 29763 14820 29797 15396
rect 29881 14820 29915 15396
rect 29999 14820 30033 15396
rect 30117 14820 30151 15396
rect 30235 14820 30269 15396
rect 30353 14820 30387 15396
rect 30471 14820 30505 15396
rect 30589 14820 30623 15396
rect 30707 14820 30741 15396
rect 30825 14820 30859 15396
rect 30943 14820 30977 15396
rect 31061 14820 31095 15396
rect 31179 14820 31213 15396
rect 31297 14820 31331 15396
rect 31415 14820 31449 15396
rect 31533 14820 31567 15396
rect 31651 14820 31685 15396
rect 31769 14820 31803 15396
rect 31887 14820 31921 15396
rect 32005 14820 32039 15396
rect 32123 14820 32157 15396
rect 32241 14820 32275 15396
rect 32359 14820 32393 15396
rect 32477 14820 32511 15396
rect 16704 13129 19543 13163
rect 16704 12847 19543 12881
rect 17367 12110 17401 12686
rect 17485 12110 17519 12686
rect 17603 12110 17637 12686
rect 17721 12110 17755 12686
rect 17839 12110 17873 12686
rect 17957 12110 17991 12686
rect 18075 12110 18109 12686
rect 18193 12110 18227 12686
rect 18311 12110 18345 12686
rect 18429 12110 18463 12686
rect 18547 12110 18581 12686
rect 18665 12110 18699 12686
rect 18783 12110 18817 12686
rect 18901 12110 18935 12686
rect 19019 12110 19053 12686
rect 19137 12110 19171 12686
rect 19255 12110 19289 12686
rect 19373 12110 19407 12686
rect 19491 12110 19525 12686
rect 17367 11274 17401 11850
rect 17485 11274 17519 11850
rect 17603 11274 17637 11850
rect 17721 11274 17755 11850
rect 17839 11274 17873 11850
rect 17957 11274 17991 11850
rect 18075 11274 18109 11850
rect 18193 11274 18227 11850
rect 18311 11274 18345 11850
rect 18429 11274 18463 11850
rect 18547 11274 18581 11850
rect 18665 11274 18699 11850
rect 18783 11274 18817 11850
rect 18901 11274 18935 11850
rect 19019 11274 19053 11850
rect 19137 11274 19171 11850
rect 19255 11274 19289 11850
rect 19373 11274 19407 11850
rect 19491 11274 19525 11850
rect 19605 11175 19639 12785
rect 17344 11079 19543 11113
rect 17344 10797 19543 10831
rect 17367 10060 17401 10636
rect 17485 10060 17519 10636
rect 17603 10060 17637 10636
rect 17721 10060 17755 10636
rect 17839 10060 17873 10636
rect 17957 10060 17991 10636
rect 18075 10060 18109 10636
rect 18193 10060 18227 10636
rect 18311 10060 18345 10636
rect 18429 10060 18463 10636
rect 18547 10060 18581 10636
rect 18665 10060 18699 10636
rect 18783 10060 18817 10636
rect 18901 10060 18935 10636
rect 19019 10060 19053 10636
rect 19137 10060 19171 10636
rect 19255 10060 19289 10636
rect 19373 10060 19407 10636
rect 19491 10060 19525 10636
rect 17367 9224 17401 9800
rect 17485 9224 17519 9800
rect 17603 9224 17637 9800
rect 17721 9224 17755 9800
rect 17839 9224 17873 9800
rect 17957 9224 17991 9800
rect 18075 9224 18109 9800
rect 18193 9224 18227 9800
rect 18311 9224 18345 9800
rect 18429 9224 18463 9800
rect 18547 9224 18581 9800
rect 18665 9224 18699 9800
rect 18783 9224 18817 9800
rect 18901 9224 18935 9800
rect 19019 9224 19053 9800
rect 19137 9224 19171 9800
rect 19255 9224 19289 9800
rect 19373 9224 19407 9800
rect 19491 9224 19525 9800
rect 19605 9125 19639 10735
rect 17344 9029 19543 9063
rect 17367 8010 17401 8586
rect 17485 8010 17519 8586
rect 17603 8010 17637 8586
rect 17721 8010 17755 8586
rect 17839 8010 17873 8586
rect 17957 8010 17991 8586
rect 18075 8010 18109 8586
rect 18193 8010 18227 8586
rect 18311 8010 18345 8586
rect 18429 8010 18463 8586
rect 18547 8010 18581 8586
rect 18665 8010 18699 8586
rect 18783 8010 18817 8586
rect 18901 8010 18935 8586
rect 19019 8010 19053 8586
rect 19137 8010 19171 8586
rect 19255 8010 19289 8586
rect 19373 8010 19407 8586
rect 19491 8010 19525 8586
rect 17367 7174 17401 7750
rect 17485 7174 17519 7750
rect 17603 7174 17637 7750
rect 17721 7174 17755 7750
rect 17839 7174 17873 7750
rect 17957 7174 17991 7750
rect 18075 7174 18109 7750
rect 18193 7174 18227 7750
rect 18311 7174 18345 7750
rect 18429 7174 18463 7750
rect 18547 7174 18581 7750
rect 18665 7174 18699 7750
rect 18783 7174 18817 7750
rect 18901 7174 18935 7750
rect 19019 7174 19053 7750
rect 19137 7174 19171 7750
rect 19255 7174 19289 7750
rect 19373 7174 19407 7750
rect 19491 7174 19525 7750
rect 17363 5767 17397 6343
rect 17481 5767 17515 6343
rect 17599 5767 17633 6343
rect 17717 5767 17751 6343
rect 17835 5767 17869 6343
rect 17953 5767 17987 6343
rect 18071 5767 18105 6343
rect 18189 5767 18223 6343
rect 18307 5767 18341 6343
rect 18425 5767 18459 6343
rect 19518 5965 19552 6271
rect 19632 6055 19666 6181
rect 19720 6055 19754 6181
rect 19834 5965 19868 6271
rect 19948 6055 19982 6181
rect 20036 6055 20070 6181
rect 20150 5965 20184 6271
rect 20264 6055 20298 6181
rect 20352 6055 20386 6181
rect 20466 5965 20500 6271
rect 20580 6055 20614 6181
rect 20668 6055 20702 6181
rect 20782 5965 20816 6271
rect 20896 6055 20930 6181
rect 20984 6055 21018 6181
rect 21098 5965 21132 6271
rect 17363 4949 17397 5525
rect 17481 4949 17515 5525
rect 17599 4949 17633 5525
rect 17717 4949 17751 5525
rect 17835 4949 17869 5525
rect 17953 4949 17987 5525
rect 18071 4949 18105 5525
rect 18189 4949 18223 5525
rect 18307 4949 18341 5525
rect 18425 4949 18459 5525
rect 21315 5467 21349 6343
rect 21463 5467 21497 6343
rect 21611 5467 21645 6343
rect 21759 5467 21793 6343
rect 21907 5467 21941 6343
rect 22055 5467 22089 6343
rect 22203 5467 22237 6343
rect 22351 5467 22385 6343
rect 22499 5467 22533 6343
rect 22647 5467 22681 6343
rect 22795 5467 22829 6343
rect 22943 5467 22977 6343
rect 23091 5467 23125 6343
rect 23239 5467 23273 6343
rect 23387 5467 23421 6343
rect 23535 5467 23569 6343
rect 23683 5467 23717 6343
rect 23831 5467 23865 6343
rect 23979 5467 24013 6343
rect 24127 5467 24161 6343
rect 24275 5467 24309 6343
rect 24423 5467 24457 6343
rect 24571 5467 24605 6343
rect 24719 5467 24753 6343
rect 24867 5467 24901 6343
rect 25015 5467 25049 6343
rect 25163 5467 25197 6343
rect 25311 5467 25345 6343
rect 25459 5467 25493 6343
rect 25607 5467 25641 6343
rect 25755 5467 25789 6343
rect 25903 5467 25937 6343
rect 26051 5467 26085 6343
rect 26199 5467 26233 6343
rect 26347 5467 26381 6343
rect 26495 5467 26529 6343
rect 26643 5467 26677 6343
rect 26791 5467 26825 6343
rect 26939 5467 26973 6343
rect 27087 5467 27121 6343
rect 27235 5467 27269 6343
rect 27383 5467 27417 6343
rect 27531 5467 27565 6343
rect 27679 5467 27713 6343
rect 27827 5467 27861 6343
rect 27975 5467 28009 6343
rect 28123 5467 28157 6343
rect 28271 5467 28305 6343
rect 28419 5467 28453 6343
rect 28567 5467 28601 6343
rect 28715 5467 28749 6343
rect 28863 5467 28897 6343
rect 29011 5467 29045 6343
rect 29159 5467 29193 6343
rect 29307 5467 29341 6343
rect 29455 5467 29489 6343
rect 29603 5467 29637 6343
rect 29751 5467 29785 6343
rect 29899 5467 29933 6343
rect 30047 5467 30081 6343
rect 30195 5467 30229 6343
rect 30343 5467 30377 6343
rect 30491 5467 30525 6343
rect 30639 5467 30673 6343
rect 30787 5467 30821 6343
rect 30935 5467 30969 6343
rect 31083 5467 31117 6343
rect 31231 5467 31265 6343
rect 31379 5467 31413 6343
rect 31527 5467 31561 6343
rect 31675 5467 31709 6343
rect 31823 5467 31857 6343
rect 31971 5467 32005 6343
rect 32119 5467 32153 6343
rect 32415 5467 32449 6343
rect 21525 5383 21583 5417
rect 21673 5383 21731 5417
rect 21821 5383 21879 5417
rect 21969 5383 22027 5417
rect 22117 5383 22175 5417
rect 22265 5383 22323 5417
rect 22413 5383 22471 5417
rect 22561 5383 22619 5417
rect 22709 5383 22767 5417
rect 22857 5383 22915 5417
rect 23005 5383 23063 5417
rect 23153 5383 23211 5417
rect 23301 5383 23359 5417
rect 23449 5383 23507 5417
rect 23597 5383 23655 5417
rect 23745 5383 23803 5417
rect 23893 5383 23951 5417
rect 24041 5383 24099 5417
rect 24189 5383 24247 5417
rect 24337 5383 24395 5417
rect 24485 5383 24543 5417
rect 24633 5383 24691 5417
rect 24781 5383 24839 5417
rect 24929 5383 24987 5417
rect 25077 5383 25135 5417
rect 25225 5383 25283 5417
rect 25373 5383 25431 5417
rect 25521 5383 25579 5417
rect 25669 5383 25727 5417
rect 25817 5383 25875 5417
rect 25965 5383 26023 5417
rect 26113 5383 26171 5417
rect 26261 5383 26319 5417
rect 26409 5383 26467 5417
rect 26557 5383 26615 5417
rect 26705 5383 26763 5417
rect 26853 5383 26911 5417
rect 27001 5383 27059 5417
rect 27149 5383 27207 5417
rect 27297 5383 27355 5417
rect 27445 5383 27503 5417
rect 27593 5383 27651 5417
rect 27741 5383 27799 5417
rect 27889 5383 27947 5417
rect 28037 5383 28095 5417
rect 28185 5383 28243 5417
rect 28333 5383 28391 5417
rect 28481 5383 28539 5417
rect 28629 5383 28687 5417
rect 28777 5383 28835 5417
rect 28925 5383 28983 5417
rect 29073 5383 29131 5417
rect 29221 5383 29279 5417
rect 29369 5383 29427 5417
rect 29517 5383 29575 5417
rect 29665 5383 29723 5417
rect 29813 5383 29871 5417
rect 29961 5383 30019 5417
rect 30109 5383 30167 5417
rect 30257 5383 30315 5417
rect 30405 5383 30463 5417
rect 30553 5383 30611 5417
rect 30701 5383 30759 5417
rect 30849 5383 30907 5417
rect 30997 5383 31055 5417
rect 31145 5383 31203 5417
rect 31293 5383 31351 5417
rect 31441 5383 31499 5417
rect 31589 5383 31647 5417
rect 31737 5383 31795 5417
rect 31885 5383 31943 5417
rect 32033 5383 32091 5417
rect 32181 5383 32239 5417
rect 32329 5383 32387 5417
rect 21525 5275 21583 5309
rect 21673 5275 21731 5309
rect 21821 5275 21879 5309
rect 21969 5275 22027 5309
rect 22117 5275 22175 5309
rect 22265 5275 22323 5309
rect 22413 5275 22471 5309
rect 22561 5275 22619 5309
rect 22709 5275 22767 5309
rect 22857 5275 22915 5309
rect 23005 5275 23063 5309
rect 23153 5275 23211 5309
rect 23301 5275 23359 5309
rect 23449 5275 23507 5309
rect 23597 5275 23655 5309
rect 23745 5275 23803 5309
rect 23893 5275 23951 5309
rect 24041 5275 24099 5309
rect 24189 5275 24247 5309
rect 24337 5275 24395 5309
rect 24485 5275 24543 5309
rect 24633 5275 24691 5309
rect 24781 5275 24839 5309
rect 24929 5275 24987 5309
rect 25077 5275 25135 5309
rect 25225 5275 25283 5309
rect 25373 5275 25431 5309
rect 25521 5275 25579 5309
rect 25669 5275 25727 5309
rect 25817 5275 25875 5309
rect 25965 5275 26023 5309
rect 26113 5275 26171 5309
rect 26261 5275 26319 5309
rect 26409 5275 26467 5309
rect 26557 5275 26615 5309
rect 26705 5275 26763 5309
rect 26853 5275 26911 5309
rect 27001 5275 27059 5309
rect 27149 5275 27207 5309
rect 27297 5275 27355 5309
rect 27445 5275 27503 5309
rect 27593 5275 27651 5309
rect 27741 5275 27799 5309
rect 27889 5275 27947 5309
rect 28037 5275 28095 5309
rect 28185 5275 28243 5309
rect 28333 5275 28391 5309
rect 28481 5275 28539 5309
rect 28629 5275 28687 5309
rect 28777 5275 28835 5309
rect 28925 5275 28983 5309
rect 29073 5275 29131 5309
rect 29221 5275 29279 5309
rect 29369 5275 29427 5309
rect 29517 5275 29575 5309
rect 29665 5275 29723 5309
rect 29813 5275 29871 5309
rect 29961 5275 30019 5309
rect 30109 5275 30167 5309
rect 30257 5275 30315 5309
rect 30405 5275 30463 5309
rect 30553 5275 30611 5309
rect 30701 5275 30759 5309
rect 30849 5275 30907 5309
rect 30997 5275 31055 5309
rect 31145 5275 31203 5309
rect 31293 5275 31351 5309
rect 31441 5275 31499 5309
rect 31589 5275 31647 5309
rect 31737 5275 31795 5309
rect 31885 5275 31943 5309
rect 32033 5275 32091 5309
rect 32181 5275 32239 5309
rect 32329 5275 32387 5309
rect 21315 4349 21349 5225
rect 21463 4349 21497 5225
rect 21611 4349 21645 5225
rect 21759 4349 21793 5225
rect 21907 4349 21941 5225
rect 22055 4349 22089 5225
rect 22203 4349 22237 5225
rect 22351 4349 22385 5225
rect 22499 4349 22533 5225
rect 22647 4349 22681 5225
rect 22795 4349 22829 5225
rect 22943 4349 22977 5225
rect 23091 4349 23125 5225
rect 23239 4349 23273 5225
rect 23387 4349 23421 5225
rect 23535 4349 23569 5225
rect 23683 4349 23717 5225
rect 23831 4349 23865 5225
rect 23979 4349 24013 5225
rect 24127 4349 24161 5225
rect 24275 4349 24309 5225
rect 24423 4349 24457 5225
rect 24571 4349 24605 5225
rect 24719 4349 24753 5225
rect 24867 4349 24901 5225
rect 25015 4349 25049 5225
rect 25163 4349 25197 5225
rect 25311 4349 25345 5225
rect 25459 4349 25493 5225
rect 25607 4349 25641 5225
rect 25755 4349 25789 5225
rect 25903 4349 25937 5225
rect 26051 4349 26085 5225
rect 26199 4349 26233 5225
rect 26347 4349 26381 5225
rect 26495 4349 26529 5225
rect 26643 4349 26677 5225
rect 26791 4349 26825 5225
rect 26939 4349 26973 5225
rect 27087 4349 27121 5225
rect 27235 4349 27269 5225
rect 27383 4349 27417 5225
rect 27531 4349 27565 5225
rect 27679 4349 27713 5225
rect 27827 4349 27861 5225
rect 27975 4349 28009 5225
rect 28123 4349 28157 5225
rect 28271 4349 28305 5225
rect 28419 4349 28453 5225
rect 28567 4349 28601 5225
rect 28715 4349 28749 5225
rect 28863 4349 28897 5225
rect 29011 4349 29045 5225
rect 29159 4349 29193 5225
rect 29307 4349 29341 5225
rect 29455 4349 29489 5225
rect 29603 4349 29637 5225
rect 29751 4349 29785 5225
rect 29899 4349 29933 5225
rect 30047 4349 30081 5225
rect 30195 4349 30229 5225
rect 30343 4349 30377 5225
rect 30491 4349 30525 5225
rect 30639 4349 30673 5225
rect 30787 4349 30821 5225
rect 30935 4349 30969 5225
rect 31083 4349 31117 5225
rect 31231 4349 31265 5225
rect 31379 4349 31413 5225
rect 31527 4349 31561 5225
rect 31675 4349 31709 5225
rect 31823 4349 31857 5225
rect 31971 4349 32005 5225
rect 32119 4349 32153 5225
<< error_ps >>
rect 16179 15657 16213 16233
rect 13573 14897 16704 14931
rect 13477 13225 13511 14835
rect 13591 14160 13625 14736
rect 13709 14160 13743 14736
rect 13827 14160 13861 14736
rect 13945 14160 13979 14736
rect 14063 14160 14097 14736
rect 14181 14160 14215 14736
rect 14299 14160 14333 14736
rect 14417 14160 14451 14736
rect 14535 14160 14569 14736
rect 14653 14160 14687 14736
rect 14771 14160 14805 14736
rect 14889 14160 14923 14736
rect 15007 14160 15041 14736
rect 15125 14160 15159 14736
rect 15243 14160 15277 14736
rect 15361 14160 15395 14736
rect 15479 14160 15513 14736
rect 15597 14160 15631 14736
rect 15715 14160 15749 14736
rect 15833 14160 15867 14736
rect 15951 14160 15985 14736
rect 16069 14160 16103 14736
rect 16187 14160 16221 14736
rect 16305 14160 16339 14736
rect 16423 14160 16457 14736
rect 16541 14160 16575 14736
rect 16659 14160 16693 14736
rect 13591 13324 13625 13900
rect 13709 13324 13743 13900
rect 13827 13324 13861 13900
rect 13945 13324 13979 13900
rect 14063 13324 14097 13900
rect 14181 13324 14215 13900
rect 14299 13324 14333 13900
rect 14417 13324 14451 13900
rect 14535 13324 14569 13900
rect 14653 13324 14687 13900
rect 14771 13324 14805 13900
rect 14889 13324 14923 13900
rect 15007 13324 15041 13900
rect 15125 13324 15159 13900
rect 15243 13324 15277 13900
rect 15361 13324 15395 13900
rect 15479 13324 15513 13900
rect 15597 13324 15631 13900
rect 15715 13324 15749 13900
rect 15833 13324 15867 13900
rect 15951 13324 15985 13900
rect 16069 13324 16103 13900
rect 16187 13324 16221 13900
rect 16305 13324 16339 13900
rect 16423 13324 16457 13900
rect 16541 13324 16575 13900
rect 16659 13324 16693 13900
rect 13573 13129 16704 13163
rect 13573 12847 16704 12881
rect 13477 11175 13511 12785
rect 13591 12110 13625 12686
rect 13709 12110 13743 12686
rect 13827 12110 13861 12686
rect 13945 12110 13979 12686
rect 14063 12110 14097 12686
rect 14181 12110 14215 12686
rect 14299 12110 14333 12686
rect 14417 12110 14451 12686
rect 14535 12110 14569 12686
rect 14653 12110 14687 12686
rect 14771 12110 14805 12686
rect 14889 12110 14923 12686
rect 15007 12110 15041 12686
rect 15125 12110 15159 12686
rect 15243 12110 15277 12686
rect 15361 12110 15395 12686
rect 15479 12110 15513 12686
rect 15597 12110 15631 12686
rect 15715 12110 15749 12686
rect 15833 12110 15867 12686
rect 15951 12110 15985 12686
rect 16069 12110 16103 12686
rect 16187 12110 16221 12686
rect 16305 12110 16339 12686
rect 16423 12110 16457 12686
rect 16541 12110 16575 12686
rect 16659 12110 16693 12686
rect 16777 12110 16811 12686
rect 16895 12110 16929 12686
rect 17013 12110 17047 12686
rect 17131 12110 17165 12686
rect 17249 12110 17283 12686
rect 13591 11274 13625 11850
rect 13709 11274 13743 11850
rect 13827 11274 13861 11850
rect 13945 11274 13979 11850
rect 14063 11274 14097 11850
rect 14181 11274 14215 11850
rect 14299 11274 14333 11850
rect 14417 11274 14451 11850
rect 14535 11274 14569 11850
rect 14653 11274 14687 11850
rect 14771 11274 14805 11850
rect 14889 11274 14923 11850
rect 15007 11274 15041 11850
rect 15125 11274 15159 11850
rect 15243 11274 15277 11850
rect 15361 11274 15395 11850
rect 15479 11274 15513 11850
rect 15597 11274 15631 11850
rect 15715 11274 15749 11850
rect 15833 11274 15867 11850
rect 15951 11274 15985 11850
rect 16069 11274 16103 11850
rect 16187 11274 16221 11850
rect 16305 11274 16339 11850
rect 16423 11274 16457 11850
rect 16541 11274 16575 11850
rect 16659 11274 16693 11850
rect 16777 11274 16811 11850
rect 16895 11274 16929 11850
rect 17013 11274 17047 11850
rect 17131 11274 17165 11850
rect 17249 11274 17283 11850
rect 13573 11079 17344 11113
rect 13573 10797 17344 10831
rect 13477 9125 13511 10735
rect 13591 10060 13625 10636
rect 13709 10060 13743 10636
rect 13827 10060 13861 10636
rect 13945 10060 13979 10636
rect 14063 10060 14097 10636
rect 14181 10060 14215 10636
rect 14299 10060 14333 10636
rect 14417 10060 14451 10636
rect 14535 10060 14569 10636
rect 14653 10060 14687 10636
rect 14771 10060 14805 10636
rect 14889 10060 14923 10636
rect 15007 10060 15041 10636
rect 15125 10060 15159 10636
rect 15243 10060 15277 10636
rect 15361 10060 15395 10636
rect 15479 10060 15513 10636
rect 15597 10060 15631 10636
rect 15715 10060 15749 10636
rect 15833 10060 15867 10636
rect 15951 10060 15985 10636
rect 16069 10060 16103 10636
rect 16187 10060 16221 10636
rect 16305 10060 16339 10636
rect 16423 10060 16457 10636
rect 16541 10060 16575 10636
rect 16659 10060 16693 10636
rect 16777 10060 16811 10636
rect 16895 10060 16929 10636
rect 17013 10060 17047 10636
rect 17131 10060 17165 10636
rect 17249 10060 17283 10636
rect 13591 9224 13625 9800
rect 13709 9224 13743 9800
rect 13827 9224 13861 9800
rect 13945 9224 13979 9800
rect 14063 9224 14097 9800
rect 14181 9224 14215 9800
rect 14299 9224 14333 9800
rect 14417 9224 14451 9800
rect 14535 9224 14569 9800
rect 14653 9224 14687 9800
rect 14771 9224 14805 9800
rect 14889 9224 14923 9800
rect 15007 9224 15041 9800
rect 15125 9224 15159 9800
rect 15243 9224 15277 9800
rect 15361 9224 15395 9800
rect 15479 9224 15513 9800
rect 15597 9224 15631 9800
rect 15715 9224 15749 9800
rect 15833 9224 15867 9800
rect 15951 9224 15985 9800
rect 16069 9224 16103 9800
rect 16187 9224 16221 9800
rect 16305 9224 16339 9800
rect 16423 9224 16457 9800
rect 16541 9224 16575 9800
rect 16659 9224 16693 9800
rect 16777 9224 16811 9800
rect 16895 9224 16929 9800
rect 17013 9224 17047 9800
rect 17131 9224 17165 9800
rect 17249 9224 17283 9800
rect 13573 9029 17344 9063
rect 13827 8010 13861 8586
rect 13945 8010 13979 8586
rect 14063 8010 14097 8586
rect 14181 8010 14215 8586
rect 14299 8010 14333 8586
rect 14417 8010 14451 8586
rect 14535 8010 14569 8586
rect 14653 8010 14687 8586
rect 14771 8010 14805 8586
rect 14889 8010 14923 8586
rect 15007 8010 15041 8586
rect 15125 8010 15159 8586
rect 15243 8010 15277 8586
rect 15361 8010 15395 8586
rect 15479 8010 15513 8586
rect 15597 8010 15631 8586
rect 15715 8010 15749 8586
rect 15833 8010 15867 8586
rect 15951 8010 15985 8586
rect 16069 8010 16103 8586
rect 16187 8010 16221 8586
rect 16305 8010 16339 8586
rect 16423 8010 16457 8586
rect 16541 8010 16575 8586
rect 16659 8010 16693 8586
rect 16777 8010 16811 8586
rect 16895 8010 16929 8586
rect 17013 8010 17047 8586
rect 17131 8010 17165 8586
rect 17249 8010 17283 8586
rect 13591 7174 13625 7750
rect 13709 7174 13743 7750
rect 13827 7174 13861 7750
rect 13945 7174 13979 7750
rect 14063 7174 14097 7750
rect 14181 7174 14215 7750
rect 14299 7174 14333 7750
rect 14417 7174 14451 7750
rect 14535 7174 14569 7750
rect 14653 7174 14687 7750
rect 14771 7174 14805 7750
rect 14889 7174 14923 7750
rect 15007 7174 15041 7750
rect 15125 7174 15159 7750
rect 15243 7174 15277 7750
rect 15361 7174 15395 7750
rect 15479 7174 15513 7750
rect 15597 7174 15631 7750
rect 15715 7174 15749 7750
rect 15833 7174 15867 7750
rect 15951 7174 15985 7750
rect 16069 7174 16103 7750
rect 16187 7174 16221 7750
rect 16305 7174 16339 7750
rect 16423 7174 16457 7750
rect 16541 7174 16575 7750
rect 16659 7174 16693 7750
rect 16777 7174 16811 7750
rect 16895 7174 16929 7750
rect 17013 7174 17047 7750
rect 17131 7174 17165 7750
rect 17249 7174 17283 7750
rect 14893 5767 14927 6343
rect 15011 5767 15045 6343
rect 15129 5767 15163 6343
rect 15247 5767 15281 6343
rect 15365 5767 15399 6343
rect 15483 5767 15517 6343
rect 15601 5767 15635 6343
rect 15719 5767 15753 6343
rect 15837 5767 15871 6343
rect 15955 5767 15989 6343
rect 16073 5767 16107 6343
rect 16191 5767 16225 6343
rect 16309 5767 16343 6343
rect 16427 5767 16461 6343
rect 16655 5767 16689 6343
rect 16773 5767 16807 6343
rect 16891 5767 16925 6343
rect 17009 5767 17043 6343
rect 17127 5767 17161 6343
rect 17245 5767 17279 6343
rect 14657 4949 14691 5525
rect 14775 4949 14809 5525
rect 14893 4949 14927 5525
rect 15011 4949 15045 5525
rect 15129 4949 15163 5525
rect 15247 4949 15281 5525
rect 15365 4949 15399 5525
rect 15483 4949 15517 5525
rect 15601 4949 15635 5525
rect 15719 4949 15753 5525
rect 15837 4949 15871 5525
rect 15955 4949 15989 5525
rect 16073 4949 16107 5525
rect 16191 4949 16225 5525
rect 16309 4949 16343 5525
rect 16427 4949 16461 5525
rect 16655 4949 16689 5525
rect 16773 4949 16807 5525
rect 16891 4949 16925 5525
rect 17009 4949 17043 5525
rect 17127 4949 17161 5525
rect 17245 4949 17279 5525
<< metal1 >>
rect 3270 17968 7575 18001
rect 3270 17852 3294 17968
rect 7570 17852 7575 17968
rect 3270 17819 7575 17852
rect 2275 17185 6745 17205
rect 2269 17170 6751 17185
rect 2269 16990 2276 17170
rect 6744 16990 6751 17170
rect 2269 16975 6751 16990
rect 6515 14295 6745 16975
rect 7405 15230 7575 17819
rect 7405 15060 8390 15230
rect 6515 14065 7695 14295
rect 7465 6285 7695 14065
rect 7465 6055 9310 6285
rect 9080 4975 9310 6055
rect 9080 4970 9558 4975
rect 9080 4967 9560 4970
rect 9080 4723 9312 4967
rect 9556 4723 9560 4967
rect 9080 4720 9560 4723
rect 9310 4715 9558 4720
rect 37180 3600 38650 3900
<< via1 >>
rect 3294 17852 7570 17968
rect 2276 16990 6744 17170
rect 9312 4723 9556 4967
<< metal2 >>
rect -3150 19580 -2820 19680
rect -1650 16075 -1560 18571
rect -4300 15965 -1560 16075
rect -4300 15315 -4190 15965
rect -1140 15470 -1050 18581
rect 1300 17115 1410 18621
rect 3300 18000 3410 18621
rect 3270 17995 3650 18000
rect 3270 17968 7581 17995
rect 3270 17852 3294 17968
rect 7570 17852 7581 17968
rect 3270 17825 7581 17852
rect 3270 17820 3650 17825
rect 2275 17170 6745 17191
rect 2275 17115 2276 17170
rect 1300 17005 2276 17115
rect 2275 16990 2276 17005
rect 6744 16990 6745 17170
rect 2275 16969 6745 16990
rect -6725 14780 -6405 14890
rect -6815 12910 -6445 13000
rect -6885 9910 -6415 10000
rect 7150 8781 9060 9029
rect -6785 6910 -6460 7000
rect 7150 4598 7398 8781
rect 9304 4967 9564 4969
rect 9304 4723 9312 4967
rect 9556 4723 9564 4967
rect 9304 4721 9564 4723
rect 5990 4480 7398 4598
rect 5984 4232 7398 4480
<< metal3 >>
rect -1380 20090 -1180 20620
rect -870 20146 -670 20610
rect 150 19916 270 20280
rect 2220 19916 2340 20380
rect -1900 16385 -1810 18570
rect -4745 16295 -1810 16385
<< metal4 >>
rect -6705 14980 -6435 15090
rect 36260 12000 39290 12860
rect -4030 3675 -3920 3940
rect -3330 3840 -3110 4560
rect -330 3940 -110 4700
rect 2670 3690 2890 4690
<< metal5 >>
rect -6700 14270 -4950 14590
use bias#0  bias_0
timestamp 1654643737
transform 1 0 -3740 0 1 20716
box 790 -2236 7180 -220
use opamp_wrapper  opamp_wrapper_0
timestamp 1654646295
transform 1 0 10500 0 1 5170
box -2280 -1609 26995 13665
use pixel_array#0  pixel_array_0
timestamp 1654643737
transform 1 0 -3550 0 1 11430
box -3000 -7600 9740 5000
<< labels >>
rlabel metal1 s 38350 3600 38650 3900 4 GND
port 1 nsew
rlabel metal3 s 230 20230 230 20230 4 OUT_IB
port 2 nsew
rlabel metal3 s 2220 20260 2340 20380 4 AMP_Ib
port 3 nsew
rlabel metal3 s -870 20410 -670 20610 4 NB2
port 4 nsew
rlabel metal3 s -1380 20420 -1180 20620 4 NB1
port 5 nsew
rlabel metal2 s -3150 19580 -2820 19680 4 SF_IB
port 6 nsew
rlabel metal4 s 38430 12000 39290 12860 4 AOUT
port 7 nsew
rlabel metal4 s -6705 14980 -6595 15090 4 VBIAS
port 8 nsew
rlabel metal2 s -6725 14780 -6615 14890 4 VREF
port 9 nsew
rlabel metal4 s -4030 3675 -3920 3785 4 CSA_VREF
port 10 nsew
rlabel metal4 s -3330 3840 -3110 4060 4 COL_SEL0
port 11 nsew
rlabel metal4 s -330 3940 -110 4160 4 COL_SEL1
port 12 nsew
rlabel metal4 s 2670 3690 2890 3910 4 COL_SEL2
port 13 nsew
rlabel metal2 s -6785 6910 -6695 7000 4 ROW_SEL2
port 14 nsew
rlabel metal2 s -6885 9910 -6795 10000 4 ROW_SEL1
port 15 nsew
rlabel metal2 s -6815 12910 -6725 13000 4 ROW_SEL0
port 16 nsew
rlabel metal5 s -6700 14270 -6380 14590 4 GRING
port 17 nsew
<< end >>
