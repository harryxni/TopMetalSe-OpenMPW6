magic
tech sky130A
magscale 1 2
timestamp 1654648307
<< nwell >>
rect 3800 -380 6800 300
<< pwell >>
rect 3834 -776 4346 -424
rect 3944 -2246 4236 -776
rect 4574 -1166 4826 -424
rect 5724 -844 5976 -604
rect 5724 -1226 6176 -844
rect 4024 -2324 4236 -2246
rect 4024 -2616 4496 -2324
<< pmoslvt >>
rect 3950 10 4350 210
rect 4420 10 4820 210
rect 5060 10 5460 210
rect 5530 10 5930 210
rect 6130 -20 6330 180
rect 6430 -20 6630 180
rect 5020 -320 6620 -236
<< nmoslvt >>
rect 3860 -680 4060 -520
rect 4120 -680 4320 -520
rect 4600 -710 4800 -510
rect 5750 -730 5950 -700
rect 4020 -2220 4050 -820
rect 4130 -2220 4160 -820
rect 4600 -1040 4800 -810
rect 5750 -1120 6150 -920
rect 4120 -2590 4320 -2350
<< ndiff >>
rect 3860 -463 4060 -450
rect 3860 -497 3909 -463
rect 3943 -497 3977 -463
rect 4011 -497 4060 -463
rect 3860 -520 4060 -497
rect 4120 -463 4320 -450
rect 4120 -497 4169 -463
rect 4203 -497 4237 -463
rect 4271 -497 4320 -463
rect 4120 -520 4320 -497
rect 4600 -461 4800 -450
rect 4600 -495 4643 -461
rect 4677 -495 4723 -461
rect 4757 -495 4800 -461
rect 4600 -510 4800 -495
rect 3860 -750 4060 -680
rect 4120 -750 4320 -680
rect 5750 -643 5950 -630
rect 5750 -677 5783 -643
rect 5817 -677 5863 -643
rect 5897 -677 5950 -643
rect 5750 -700 5950 -677
rect 4600 -743 4800 -710
rect 3970 -820 4000 -750
rect 4180 -820 4210 -750
rect 4600 -777 4659 -743
rect 4693 -777 4727 -743
rect 4761 -777 4800 -743
rect 4600 -810 4800 -777
rect 5750 -760 5950 -730
rect 3970 -2220 4020 -820
rect 4050 -881 4130 -820
rect 4050 -915 4073 -881
rect 4107 -915 4130 -881
rect 4050 -949 4130 -915
rect 4050 -983 4073 -949
rect 4107 -983 4130 -949
rect 4050 -1017 4130 -983
rect 4050 -1051 4073 -1017
rect 4107 -1051 4130 -1017
rect 4050 -1085 4130 -1051
rect 4050 -1119 4073 -1085
rect 4107 -1119 4130 -1085
rect 4050 -1153 4130 -1119
rect 4050 -1187 4073 -1153
rect 4107 -1187 4130 -1153
rect 4050 -1221 4130 -1187
rect 4050 -1255 4073 -1221
rect 4107 -1255 4130 -1221
rect 4050 -1289 4130 -1255
rect 4050 -1323 4073 -1289
rect 4107 -1323 4130 -1289
rect 4050 -1357 4130 -1323
rect 4050 -1391 4073 -1357
rect 4107 -1391 4130 -1357
rect 4050 -1425 4130 -1391
rect 4050 -1459 4073 -1425
rect 4107 -1459 4130 -1425
rect 4050 -1493 4130 -1459
rect 4050 -1527 4073 -1493
rect 4107 -1527 4130 -1493
rect 4050 -1561 4130 -1527
rect 4050 -1595 4073 -1561
rect 4107 -1595 4130 -1561
rect 4050 -1629 4130 -1595
rect 4050 -1663 4073 -1629
rect 4107 -1663 4130 -1629
rect 4050 -1697 4130 -1663
rect 4050 -1731 4073 -1697
rect 4107 -1731 4130 -1697
rect 4050 -1765 4130 -1731
rect 4050 -1799 4073 -1765
rect 4107 -1799 4130 -1765
rect 4050 -1833 4130 -1799
rect 4050 -1867 4073 -1833
rect 4107 -1867 4130 -1833
rect 4050 -1901 4130 -1867
rect 4050 -1935 4073 -1901
rect 4107 -1935 4130 -1901
rect 4050 -1969 4130 -1935
rect 4050 -2003 4073 -1969
rect 4107 -2003 4130 -1969
rect 4050 -2037 4130 -2003
rect 4050 -2071 4073 -2037
rect 4107 -2071 4130 -2037
rect 4050 -2105 4130 -2071
rect 4050 -2139 4073 -2105
rect 4107 -2139 4130 -2105
rect 4050 -2220 4130 -2139
rect 4160 -2220 4210 -820
rect 5750 -870 5840 -760
rect 5750 -920 6150 -870
rect 4600 -1078 4800 -1040
rect 4600 -1112 4644 -1078
rect 4678 -1112 4712 -1078
rect 4746 -1112 4800 -1078
rect 4600 -1140 4800 -1112
rect 5750 -1148 6150 -1120
rect 5750 -1182 5782 -1148
rect 5816 -1182 5850 -1148
rect 5884 -1182 5918 -1148
rect 5952 -1182 5986 -1148
rect 6020 -1182 6054 -1148
rect 6088 -1182 6150 -1148
rect 5750 -1200 6150 -1182
rect 4050 -2380 4120 -2350
rect 4050 -2414 4063 -2380
rect 4097 -2414 4120 -2380
rect 4050 -2448 4120 -2414
rect 4050 -2482 4063 -2448
rect 4097 -2482 4120 -2448
rect 4050 -2516 4120 -2482
rect 4050 -2550 4063 -2516
rect 4097 -2550 4120 -2516
rect 4050 -2590 4120 -2550
rect 4320 -2380 4390 -2350
rect 4320 -2414 4343 -2380
rect 4377 -2414 4390 -2380
rect 4320 -2448 4390 -2414
rect 4320 -2482 4343 -2448
rect 4377 -2482 4390 -2448
rect 4320 -2516 4390 -2482
rect 4320 -2550 4343 -2516
rect 4377 -2550 4390 -2516
rect 4320 -2590 4390 -2550
<< pdiff >>
rect 3880 141 3950 210
rect 3880 107 3893 141
rect 3927 107 3950 141
rect 3880 73 3950 107
rect 3880 39 3893 73
rect 3927 39 3950 73
rect 3880 10 3950 39
rect 4350 134 4420 210
rect 4350 100 4370 134
rect 4404 100 4420 134
rect 4350 54 4420 100
rect 4350 20 4370 54
rect 4404 20 4420 54
rect 4350 10 4420 20
rect 4820 161 4890 210
rect 4990 161 5060 210
rect 4820 127 4843 161
rect 4877 127 4890 161
rect 4990 127 5003 161
rect 5037 127 5060 161
rect 4820 93 4890 127
rect 4990 93 5060 127
rect 4820 59 4843 93
rect 4877 59 4890 93
rect 4990 59 5003 93
rect 5037 59 5060 93
rect 4820 10 4890 59
rect 4990 10 5060 59
rect 5460 10 5530 210
rect 5930 134 6000 210
rect 5930 100 5950 134
rect 5984 100 6000 134
rect 5930 54 6000 100
rect 5930 20 5950 54
rect 5984 20 6000 54
rect 5930 10 6000 20
rect 6060 129 6130 180
rect 6060 95 6076 129
rect 6110 95 6130 129
rect 6060 61 6130 95
rect 6060 27 6076 61
rect 6110 27 6130 61
rect 6060 -20 6130 27
rect 6330 121 6430 180
rect 6330 87 6363 121
rect 6397 87 6430 121
rect 6330 53 6430 87
rect 6330 19 6363 53
rect 6397 19 6430 53
rect 6330 -20 6430 19
rect 6630 131 6700 180
rect 6630 97 6653 131
rect 6687 97 6700 131
rect 6630 63 6700 97
rect 6630 29 6653 63
rect 6687 29 6700 63
rect 6630 -20 6700 29
rect 4890 -268 5020 -236
rect 4890 -302 4933 -268
rect 4967 -302 5020 -268
rect 4890 -320 5020 -302
rect 6620 -255 6760 -236
rect 6620 -289 6668 -255
rect 6702 -289 6760 -255
rect 6620 -320 6760 -289
<< ndiffc >>
rect 3909 -497 3943 -463
rect 3977 -497 4011 -463
rect 4169 -497 4203 -463
rect 4237 -497 4271 -463
rect 4643 -495 4677 -461
rect 4723 -495 4757 -461
rect 5783 -677 5817 -643
rect 5863 -677 5897 -643
rect 4659 -777 4693 -743
rect 4727 -777 4761 -743
rect 4073 -915 4107 -881
rect 4073 -983 4107 -949
rect 4073 -1051 4107 -1017
rect 4073 -1119 4107 -1085
rect 4073 -1187 4107 -1153
rect 4073 -1255 4107 -1221
rect 4073 -1323 4107 -1289
rect 4073 -1391 4107 -1357
rect 4073 -1459 4107 -1425
rect 4073 -1527 4107 -1493
rect 4073 -1595 4107 -1561
rect 4073 -1663 4107 -1629
rect 4073 -1731 4107 -1697
rect 4073 -1799 4107 -1765
rect 4073 -1867 4107 -1833
rect 4073 -1935 4107 -1901
rect 4073 -2003 4107 -1969
rect 4073 -2071 4107 -2037
rect 4073 -2139 4107 -2105
rect 4644 -1112 4678 -1078
rect 4712 -1112 4746 -1078
rect 5782 -1182 5816 -1148
rect 5850 -1182 5884 -1148
rect 5918 -1182 5952 -1148
rect 5986 -1182 6020 -1148
rect 6054 -1182 6088 -1148
rect 4063 -2414 4097 -2380
rect 4063 -2482 4097 -2448
rect 4063 -2550 4097 -2516
rect 4343 -2414 4377 -2380
rect 4343 -2482 4377 -2448
rect 4343 -2550 4377 -2516
<< pdiffc >>
rect 3893 107 3927 141
rect 3893 39 3927 73
rect 4370 100 4404 134
rect 4370 20 4404 54
rect 4843 127 4877 161
rect 5003 127 5037 161
rect 4843 59 4877 93
rect 5003 59 5037 93
rect 5950 100 5984 134
rect 5950 20 5984 54
rect 6076 95 6110 129
rect 6076 27 6110 61
rect 6363 87 6397 121
rect 6363 19 6397 53
rect 6653 97 6687 131
rect 6653 29 6687 63
rect 4933 -302 4967 -268
rect 6668 -289 6702 -255
<< psubdiff >>
rect 4390 -2385 4470 -2350
rect 4390 -2419 4423 -2385
rect 4457 -2419 4470 -2385
rect 4390 -2453 4470 -2419
rect 4390 -2487 4423 -2453
rect 4457 -2487 4470 -2453
rect 4390 -2521 4470 -2487
rect 4390 -2555 4423 -2521
rect 4457 -2555 4470 -2521
rect 4390 -2590 4470 -2555
<< nsubdiff >>
rect 4890 161 4990 210
rect 4890 127 4923 161
rect 4957 127 4990 161
rect 4890 93 4990 127
rect 4890 59 4923 93
rect 4957 59 4990 93
rect 4890 10 4990 59
<< psubdiffcont >>
rect 4423 -2419 4457 -2385
rect 4423 -2487 4457 -2453
rect 4423 -2555 4457 -2521
<< nsubdiffcont >>
rect 4923 127 4957 161
rect 4923 59 4957 93
<< poly >>
rect 3950 210 4350 240
rect 4420 210 4820 240
rect 5060 210 5460 240
rect 5530 210 5930 240
rect 6130 180 6330 210
rect 6430 180 6630 210
rect 3950 -20 4350 10
rect 4420 -20 4820 10
rect 5060 -20 5460 10
rect 5530 -20 5930 10
rect 4010 -43 4080 -20
rect 4010 -77 4033 -43
rect 4067 -77 4080 -43
rect 4010 -100 4080 -77
rect 4300 -150 4350 -20
rect 4480 -43 4550 -20
rect 4480 -77 4503 -43
rect 4537 -77 4550 -43
rect 4770 -50 5110 -20
rect 4480 -100 4550 -77
rect 5530 -100 5580 -20
rect 4600 -140 5580 -100
rect 6130 -50 6330 -20
rect 6430 -50 6630 -20
rect 6130 -98 6210 -50
rect 6130 -132 6153 -98
rect 6187 -132 6210 -98
rect 4600 -150 4630 -140
rect 4300 -180 4630 -150
rect 6130 -160 6210 -132
rect 6550 -98 6630 -50
rect 6550 -132 6573 -98
rect 6607 -132 6630 -98
rect 6550 -160 6630 -132
rect 5020 -236 6620 -208
rect 5020 -350 6620 -320
rect 6510 -413 6620 -350
rect 6510 -447 6548 -413
rect 6582 -447 6620 -413
rect 6510 -480 6620 -447
rect 3830 -680 3860 -520
rect 4060 -680 4120 -520
rect 4320 -550 4350 -520
rect 4500 -544 4600 -510
rect 4320 -583 4420 -550
rect 4320 -617 4363 -583
rect 4397 -617 4420 -583
rect 4320 -650 4420 -617
rect 4500 -578 4518 -544
rect 4552 -578 4600 -544
rect 4500 -612 4600 -578
rect 4500 -646 4518 -612
rect 4552 -646 4600 -612
rect 4320 -680 4350 -650
rect 4500 -710 4600 -646
rect 4800 -710 4830 -510
rect 5970 -698 6060 -680
rect 5970 -700 5998 -698
rect 5720 -730 5750 -700
rect 5950 -730 5998 -700
rect 4020 -820 4050 -790
rect 4130 -820 4160 -790
rect 5970 -732 5998 -730
rect 6032 -732 6060 -698
rect 5970 -750 6060 -732
rect 3850 -2238 3940 -2210
rect 4560 -1040 4600 -810
rect 4800 -840 4840 -810
rect 4800 -874 4930 -840
rect 4800 -908 4873 -874
rect 4907 -908 4930 -874
rect 4800 -942 4930 -908
rect 6190 -920 6270 -910
rect 4800 -976 4873 -942
rect 4907 -976 4930 -942
rect 4800 -1010 4930 -976
rect 4800 -1040 4840 -1010
rect 5720 -1120 5750 -920
rect 6150 -933 6270 -920
rect 6150 -967 6208 -933
rect 6242 -967 6270 -933
rect 6150 -990 6270 -967
rect 6150 -1120 6180 -990
rect 3850 -2272 3878 -2238
rect 3912 -2240 3940 -2238
rect 4020 -2240 4050 -2220
rect 3912 -2270 4050 -2240
rect 4130 -2240 4160 -2220
rect 4280 -2223 4570 -2210
rect 4280 -2240 4311 -2223
rect 4130 -2257 4311 -2240
rect 4345 -2257 4379 -2223
rect 4413 -2257 4447 -2223
rect 4481 -2257 4515 -2223
rect 4549 -2257 4570 -2223
rect 4130 -2270 4570 -2257
rect 3912 -2272 3940 -2270
rect 3850 -2300 3940 -2272
rect 4120 -2350 4320 -2320
rect 4500 -2488 4590 -2470
rect 4500 -2522 4528 -2488
rect 4562 -2522 4590 -2488
rect 4500 -2540 4590 -2522
rect 4510 -2550 4580 -2540
rect 4120 -2620 4320 -2590
rect 4530 -2620 4560 -2550
rect 4290 -2650 4560 -2620
<< polycont >>
rect 4033 -77 4067 -43
rect 4503 -77 4537 -43
rect 6153 -132 6187 -98
rect 6573 -132 6607 -98
rect 6548 -447 6582 -413
rect 4363 -617 4397 -583
rect 4518 -578 4552 -544
rect 4518 -646 4552 -612
rect 5998 -732 6032 -698
rect 4873 -908 4907 -874
rect 4873 -976 4907 -942
rect 6208 -967 6242 -933
rect 3878 -2272 3912 -2238
rect 4311 -2257 4345 -2223
rect 4379 -2257 4413 -2223
rect 4447 -2257 4481 -2223
rect 4515 -2257 4549 -2223
rect 4528 -2522 4562 -2488
<< locali >>
rect 4890 252 4990 270
rect 6650 260 6690 270
rect 4890 218 4923 252
rect 4957 218 4990 252
rect 6630 257 6710 260
rect 6630 223 6653 257
rect 6687 223 6710 257
rect 6630 220 6710 223
rect 4890 210 4990 218
rect 3880 141 3930 170
rect 3880 107 3893 141
rect 3927 107 3930 141
rect 3880 73 3930 107
rect 3880 39 3893 73
rect 3927 39 3930 73
rect 3880 -30 3930 39
rect 4370 134 4410 210
rect 4404 100 4410 134
rect 4370 54 4410 100
rect 4404 20 4410 54
rect 4010 -30 4080 -10
rect 3860 -43 4080 -30
rect 3860 -70 4033 -43
rect 3860 -450 3900 -70
rect 4010 -77 4033 -70
rect 4067 -77 4080 -43
rect 4370 -30 4410 20
rect 4820 161 5060 210
rect 4820 127 4843 161
rect 4877 127 4923 161
rect 4957 127 5003 161
rect 5037 127 5060 161
rect 4820 93 5060 127
rect 4820 59 4843 93
rect 4877 59 4923 93
rect 4957 59 5003 93
rect 5037 59 5060 93
rect 4820 10 5060 59
rect 5950 134 5990 210
rect 5984 100 5990 134
rect 5950 54 5990 100
rect 5984 20 5990 54
rect 4480 -30 4550 -10
rect 4370 -43 4550 -30
rect 4370 -70 4503 -43
rect 4010 -100 4080 -77
rect 4480 -77 4503 -70
rect 4537 -77 4550 -43
rect 4480 -100 4550 -77
rect 5950 -170 5990 20
rect 4280 -210 5990 -170
rect 6030 129 6110 180
rect 6030 95 6076 129
rect 6030 61 6110 95
rect 6030 27 6076 61
rect 6030 -20 6110 27
rect 6350 121 6410 170
rect 6350 87 6363 121
rect 6397 87 6410 121
rect 6350 53 6410 87
rect 6350 19 6363 53
rect 6397 19 6410 53
rect 4280 -280 4320 -210
rect 6030 -250 6080 -20
rect 6120 -98 6220 -80
rect 6120 -132 6153 -98
rect 6187 -132 6220 -98
rect 6350 -120 6410 19
rect 6650 131 6690 220
rect 6650 97 6653 131
rect 6687 97 6690 131
rect 6650 63 6690 97
rect 6650 29 6653 63
rect 6687 29 6690 63
rect 6650 -20 6690 29
rect 6120 -160 6220 -132
rect 6130 -190 6210 -160
rect 6320 -180 6410 -120
rect 6540 -98 6720 -90
rect 6540 -132 6573 -98
rect 6607 -132 6683 -98
rect 6717 -132 6720 -98
rect 6540 -140 6720 -132
rect 4650 -253 4720 -250
rect 4280 -330 4570 -280
rect 4280 -450 4320 -330
rect 3860 -463 4060 -450
rect 3860 -497 3909 -463
rect 3943 -497 3977 -463
rect 4011 -497 4060 -463
rect 3860 -510 4060 -497
rect 4120 -463 4320 -450
rect 4120 -497 4169 -463
rect 4203 -497 4237 -463
rect 4271 -497 4320 -463
rect 4120 -510 4320 -497
rect 4370 -483 4420 -460
rect 4370 -517 4378 -483
rect 4412 -517 4420 -483
rect 4520 -510 4570 -330
rect 4650 -287 4668 -253
rect 4702 -287 4720 -253
rect 4650 -290 4720 -287
rect 4890 -268 5010 -250
rect 4650 -450 4690 -290
rect 4890 -302 4933 -268
rect 4967 -302 5010 -268
rect 4890 -320 5010 -302
rect 5870 -263 6080 -250
rect 5870 -297 5908 -263
rect 5942 -297 6080 -263
rect 5870 -320 6080 -297
rect 4890 -400 4960 -320
rect 6140 -400 6180 -190
rect 4890 -440 6180 -400
rect 4620 -461 4800 -450
rect 4620 -495 4643 -461
rect 4677 -495 4723 -461
rect 4757 -495 4800 -461
rect 4620 -500 4800 -495
rect 4370 -550 4420 -517
rect 4340 -583 4420 -550
rect 4340 -617 4363 -583
rect 4397 -617 4420 -583
rect 4340 -650 4420 -617
rect 4500 -544 4570 -510
rect 4500 -578 4518 -544
rect 4552 -578 4570 -544
rect 4500 -612 4570 -578
rect 4500 -646 4518 -612
rect 4552 -646 4570 -612
rect 4500 -690 4570 -646
rect 4890 -548 4960 -440
rect 4890 -582 4908 -548
rect 4942 -582 4960 -548
rect 4890 -720 4960 -582
rect 5760 -532 5830 -510
rect 6320 -530 6360 -180
rect 6640 -255 6730 -236
rect 6640 -289 6668 -255
rect 6702 -289 6730 -255
rect 6640 -310 6730 -289
rect 6520 -413 6610 -370
rect 6520 -430 6548 -413
rect 6430 -438 6548 -430
rect 6430 -472 6438 -438
rect 6472 -447 6548 -438
rect 6582 -430 6610 -413
rect 6582 -447 6620 -430
rect 6472 -472 6620 -447
rect 6430 -480 6620 -472
rect 5760 -566 5778 -532
rect 5812 -566 5830 -532
rect 5760 -604 5830 -566
rect 5760 -638 5778 -604
rect 5812 -620 5830 -604
rect 5990 -570 6360 -530
rect 5812 -638 5940 -620
rect 5760 -643 5940 -638
rect 5760 -677 5783 -643
rect 5817 -677 5863 -643
rect 5897 -677 5940 -643
rect 5760 -680 5940 -677
rect 5990 -680 6040 -570
rect 6670 -580 6730 -310
rect 6400 -618 6730 -580
rect 6400 -652 6412 -618
rect 6446 -652 6484 -618
rect 6518 -630 6730 -618
rect 6518 -652 6530 -630
rect 4620 -730 4960 -720
rect 4600 -743 4960 -730
rect 4600 -777 4659 -743
rect 4693 -777 4727 -743
rect 4761 -777 4960 -743
rect 5980 -698 6050 -680
rect 6400 -690 6530 -652
rect 5980 -732 5998 -698
rect 6032 -732 6050 -698
rect 5980 -750 6050 -732
rect 5990 -770 6040 -750
rect 4600 -790 4960 -777
rect 4620 -800 4960 -790
rect 4060 -881 4120 -820
rect 4060 -915 4073 -881
rect 4107 -915 4120 -881
rect 4060 -949 4120 -915
rect 4060 -983 4073 -949
rect 4107 -983 4120 -949
rect 4060 -1017 4120 -983
rect 4810 -874 4930 -840
rect 4810 -908 4873 -874
rect 4907 -908 4930 -874
rect 4810 -942 4930 -908
rect 4810 -976 4873 -942
rect 4907 -976 4930 -942
rect 4810 -1010 4930 -976
rect 4060 -1051 4073 -1017
rect 4107 -1051 4120 -1017
rect 4820 -1038 4930 -1010
rect 4060 -1085 4120 -1051
rect 4060 -1119 4073 -1085
rect 4107 -1119 4120 -1085
rect 4060 -1153 4120 -1119
rect 4060 -1187 4073 -1153
rect 4107 -1187 4120 -1153
rect 4060 -1221 4120 -1187
rect 4060 -1255 4073 -1221
rect 4107 -1255 4120 -1221
rect 4060 -1289 4120 -1255
rect 4060 -1323 4073 -1289
rect 4107 -1323 4120 -1289
rect 4060 -1357 4120 -1323
rect 4060 -1391 4073 -1357
rect 4107 -1391 4120 -1357
rect 4060 -1425 4120 -1391
rect 4060 -1459 4073 -1425
rect 4107 -1459 4120 -1425
rect 4060 -1493 4120 -1459
rect 4060 -1527 4073 -1493
rect 4107 -1527 4120 -1493
rect 4060 -1561 4120 -1527
rect 4060 -1595 4073 -1561
rect 4107 -1595 4120 -1561
rect 4600 -1078 4780 -1050
rect 4600 -1112 4644 -1078
rect 4678 -1112 4712 -1078
rect 4746 -1112 4780 -1078
rect 4820 -1072 4858 -1038
rect 4892 -1072 4930 -1038
rect 4820 -1090 4930 -1072
rect 6200 -933 6250 -900
rect 6200 -967 6208 -933
rect 6242 -967 6250 -933
rect 6200 -1038 6250 -967
rect 6200 -1072 6208 -1038
rect 6242 -1072 6250 -1038
rect 6200 -1110 6250 -1072
rect 4600 -1140 4780 -1112
rect 4600 -1513 4700 -1140
rect 5750 -1148 6140 -1140
rect 5750 -1182 5782 -1148
rect 5816 -1182 5850 -1148
rect 5884 -1182 5918 -1148
rect 5952 -1182 5986 -1148
rect 6020 -1182 6054 -1148
rect 6088 -1182 6140 -1148
rect 5750 -1210 6140 -1182
rect 4600 -1547 4633 -1513
rect 4667 -1547 4700 -1513
rect 4600 -1580 4700 -1547
rect 5990 -1490 6140 -1210
rect 5990 -1512 6590 -1490
rect 4060 -1629 4120 -1595
rect 4060 -1663 4073 -1629
rect 4107 -1663 4120 -1629
rect 5990 -1618 6452 -1512
rect 6558 -1618 6590 -1512
rect 5990 -1640 6590 -1618
rect 4060 -1697 4120 -1663
rect 4060 -1731 4073 -1697
rect 4107 -1731 4120 -1697
rect 4060 -1765 4120 -1731
rect 4060 -1799 4073 -1765
rect 4107 -1799 4120 -1765
rect 4060 -1833 4120 -1799
rect 4060 -1867 4073 -1833
rect 4107 -1867 4120 -1833
rect 4060 -1901 4120 -1867
rect 4060 -1935 4073 -1901
rect 4107 -1935 4120 -1901
rect 4060 -1969 4120 -1935
rect 4060 -2003 4073 -1969
rect 4107 -2003 4120 -1969
rect 4060 -2037 4120 -2003
rect 4060 -2071 4073 -2037
rect 4107 -2071 4120 -2037
rect 4060 -2105 4120 -2071
rect 4060 -2139 4073 -2105
rect 4107 -2139 4120 -2105
rect 3850 -2158 3940 -2150
rect 3850 -2192 3878 -2158
rect 3912 -2192 3940 -2158
rect 3850 -2238 3940 -2192
rect 3850 -2272 3878 -2238
rect 3912 -2272 3940 -2238
rect 3850 -2300 3940 -2272
rect 4060 -2220 4120 -2139
rect 4440 -2092 4580 -2080
rect 4440 -2126 4493 -2092
rect 4527 -2126 4580 -2092
rect 4440 -2164 4580 -2126
rect 4440 -2198 4493 -2164
rect 4527 -2198 4580 -2164
rect 4440 -2210 4580 -2198
rect 4060 -2350 4110 -2220
rect 4290 -2223 4580 -2210
rect 4290 -2257 4311 -2223
rect 4345 -2257 4379 -2223
rect 4413 -2257 4447 -2223
rect 4481 -2257 4515 -2223
rect 4549 -2257 4580 -2223
rect 4290 -2270 4580 -2257
rect 4050 -2380 4110 -2350
rect 4050 -2414 4063 -2380
rect 4097 -2414 4110 -2380
rect 4050 -2448 4110 -2414
rect 4050 -2482 4063 -2448
rect 4097 -2482 4110 -2448
rect 4050 -2516 4110 -2482
rect 4050 -2550 4063 -2516
rect 4097 -2550 4110 -2516
rect 4050 -2590 4110 -2550
rect 4330 -2380 4470 -2350
rect 4330 -2414 4343 -2380
rect 4377 -2385 4470 -2380
rect 4377 -2414 4423 -2385
rect 4330 -2419 4423 -2414
rect 4457 -2419 4470 -2385
rect 4330 -2448 4470 -2419
rect 4330 -2482 4343 -2448
rect 4377 -2453 4470 -2448
rect 4377 -2482 4423 -2453
rect 4330 -2487 4423 -2482
rect 4457 -2487 4470 -2453
rect 4330 -2516 4470 -2487
rect 4330 -2550 4343 -2516
rect 4377 -2521 4470 -2516
rect 4377 -2550 4423 -2521
rect 4330 -2555 4423 -2550
rect 4457 -2555 4470 -2521
rect 4510 -2423 4600 -2410
rect 4510 -2457 4538 -2423
rect 4572 -2457 4600 -2423
rect 4510 -2470 4600 -2457
rect 4510 -2488 4580 -2470
rect 4510 -2522 4528 -2488
rect 4562 -2522 4580 -2488
rect 4510 -2550 4580 -2522
rect 4330 -2590 4470 -2555
rect 4380 -2623 4430 -2590
rect 4380 -2657 4383 -2623
rect 4417 -2657 4430 -2623
rect 4380 -2670 4430 -2657
<< viali >>
rect 4923 218 4957 252
rect 6653 223 6687 257
rect 6683 -132 6717 -98
rect 4378 -517 4412 -483
rect 4668 -287 4702 -253
rect 5908 -297 5942 -263
rect 4908 -582 4942 -548
rect 6438 -472 6472 -438
rect 5778 -566 5812 -532
rect 5778 -638 5812 -604
rect 6412 -652 6446 -618
rect 6484 -652 6518 -618
rect 4858 -1072 4892 -1038
rect 6208 -1072 6242 -1038
rect 4633 -1547 4667 -1513
rect 6452 -1618 6558 -1512
rect 3878 -2192 3912 -2158
rect 4493 -2126 4527 -2092
rect 4493 -2198 4527 -2164
rect 4538 -2457 4572 -2423
rect 4383 -2657 4417 -2623
<< metal1 >>
rect 3800 257 6800 270
rect 3800 252 6653 257
rect 3800 218 4923 252
rect 4957 223 6653 252
rect 6687 223 6800 257
rect 4957 218 6800 223
rect 3800 120 6800 218
rect 4710 -230 4810 120
rect 4630 -253 4810 -230
rect 4630 -287 4668 -253
rect 4702 -287 4810 -253
rect 4630 -300 4810 -287
rect 4280 -394 4430 -390
rect 4280 -446 4299 -394
rect 4351 -446 4430 -394
rect 4280 -460 4430 -446
rect 4360 -483 4430 -460
rect 4360 -517 4378 -483
rect 4412 -517 4430 -483
rect 4360 -550 4430 -517
rect 4890 -540 4960 -520
rect 5080 -524 5160 -520
rect 5080 -540 5094 -524
rect 4890 -548 5094 -540
rect 4370 -610 4420 -550
rect 4890 -582 4908 -548
rect 4942 -576 5094 -548
rect 5146 -576 5160 -524
rect 4942 -582 5160 -576
rect 4890 -590 5160 -582
rect 5760 -532 5830 120
rect 6660 -89 6790 -80
rect 6660 -98 6724 -89
rect 6660 -132 6683 -98
rect 6717 -132 6724 -98
rect 6660 -141 6724 -132
rect 6776 -141 6790 -89
rect 6660 -150 6790 -141
rect 5760 -566 5778 -532
rect 5812 -566 5830 -532
rect 4890 -610 4960 -590
rect 5760 -604 5830 -566
rect 5760 -638 5778 -604
rect 5812 -638 5830 -604
rect 5760 -670 5830 -638
rect 5870 -263 5990 -230
rect 5870 -297 5908 -263
rect 5942 -297 5990 -263
rect 5870 -320 5990 -297
rect 4790 -1038 4930 -1010
rect 4790 -1072 4858 -1038
rect 4892 -1072 4930 -1038
rect 4790 -1084 4930 -1072
rect 4790 -1136 4834 -1084
rect 4886 -1136 4930 -1084
rect 4790 -1150 4930 -1136
rect 4590 -1513 5100 -1480
rect 4590 -1547 4633 -1513
rect 4667 -1547 5100 -1513
rect 4590 -1580 5100 -1547
rect 4440 -1994 4580 -1950
rect 4440 -2046 4452 -1994
rect 4504 -2046 4516 -1994
rect 4568 -2046 4580 -1994
rect 3850 -2079 3940 -2060
rect 3850 -2131 3869 -2079
rect 3921 -2131 3940 -2079
rect 3850 -2158 3940 -2131
rect 3850 -2192 3878 -2158
rect 3912 -2192 3940 -2158
rect 3850 -2210 3940 -2192
rect 4440 -2092 4580 -2046
rect 4440 -2126 4493 -2092
rect 4527 -2126 4580 -2092
rect 4440 -2164 4580 -2126
rect 4440 -2198 4493 -2164
rect 4527 -2198 4580 -2164
rect 4440 -2220 4580 -2198
rect 4500 -2414 4700 -2410
rect 4500 -2423 4629 -2414
rect 4500 -2457 4538 -2423
rect 4572 -2457 4629 -2423
rect 4500 -2466 4629 -2457
rect 4681 -2466 4700 -2414
rect 4500 -2470 4700 -2466
rect 4990 -2520 5100 -1580
rect 5870 -2520 5970 -320
rect 6410 -424 6500 -400
rect 6410 -476 6429 -424
rect 6481 -476 6500 -424
rect 6410 -500 6500 -476
rect 6060 -609 6540 -580
rect 6060 -661 6080 -609
rect 6132 -661 6144 -609
rect 6196 -661 6208 -609
rect 6260 -618 6540 -609
rect 6260 -652 6412 -618
rect 6446 -652 6484 -618
rect 6518 -652 6540 -618
rect 6260 -661 6540 -652
rect 6060 -690 6540 -661
rect 6190 -1038 6260 -1000
rect 6190 -1072 6208 -1038
rect 6242 -1072 6260 -1038
rect 6190 -1119 6260 -1072
rect 6190 -1171 6199 -1119
rect 6251 -1171 6260 -1119
rect 6190 -1200 6260 -1171
rect 6420 -1507 6590 -1490
rect 6420 -1623 6447 -1507
rect 6563 -1623 6590 -1507
rect 6420 -1640 6590 -1623
rect 3800 -2599 6800 -2520
rect 3800 -2623 5284 -2599
rect 3800 -2657 4383 -2623
rect 4417 -2651 5284 -2623
rect 5336 -2651 6800 -2599
rect 4417 -2657 6800 -2651
rect 3800 -2670 6800 -2657
<< via1 >>
rect 4299 -446 4351 -394
rect 5094 -576 5146 -524
rect 6724 -141 6776 -89
rect 4834 -1136 4886 -1084
rect 4452 -2046 4504 -1994
rect 4516 -2046 4568 -1994
rect 3869 -2131 3921 -2079
rect 4629 -2466 4681 -2414
rect 6429 -438 6481 -424
rect 6429 -472 6438 -438
rect 6438 -472 6472 -438
rect 6472 -472 6481 -438
rect 6429 -476 6481 -472
rect 6080 -661 6132 -609
rect 6144 -661 6196 -609
rect 6208 -661 6260 -609
rect 6199 -1171 6251 -1119
rect 6447 -1512 6563 -1507
rect 6447 -1618 6452 -1512
rect 6452 -1618 6558 -1512
rect 6558 -1618 6563 -1512
rect 6447 -1623 6563 -1618
rect 5284 -2651 5336 -2599
<< metal2 >>
rect 3860 -2079 3930 300
rect 4300 -390 4370 300
rect 4280 -394 4380 -390
rect 4280 -446 4299 -394
rect 4351 -446 4380 -394
rect 4280 -460 4380 -446
rect 3860 -2131 3869 -2079
rect 3921 -2131 3930 -2079
rect 3860 -2700 3930 -2131
rect 4300 -2700 4370 -460
rect 4820 -1084 4900 300
rect 6720 118 6780 130
rect 6720 62 6722 118
rect 6778 62 6780 118
rect 6720 -89 6780 62
rect 6720 -141 6724 -89
rect 6776 -141 6780 -89
rect 6420 -177 6490 -150
rect 6720 -170 6780 -141
rect 6420 -233 6427 -177
rect 6483 -233 6490 -177
rect 5080 -422 5160 -400
rect 5080 -478 5097 -422
rect 5153 -478 5160 -422
rect 6420 -424 6490 -233
rect 5080 -524 5160 -478
rect 5080 -576 5094 -524
rect 5146 -576 5160 -524
rect 5080 -600 5160 -576
rect 5870 -472 6290 -440
rect 5870 -688 5887 -472
rect 6023 -609 6290 -472
rect 6420 -476 6429 -424
rect 6481 -476 6490 -424
rect 6420 -510 6490 -476
rect 6023 -661 6080 -609
rect 6132 -661 6144 -609
rect 6196 -661 6208 -609
rect 6260 -661 6290 -609
rect 6023 -688 6290 -661
rect 5870 -710 6290 -688
rect 4820 -1136 4834 -1084
rect 4886 -1136 4900 -1084
rect 4440 -1977 4730 -1950
rect 4440 -1994 4477 -1977
rect 4533 -1994 4557 -1977
rect 4440 -2046 4452 -1994
rect 4613 -2033 4637 -1977
rect 4693 -2033 4730 -1977
rect 4504 -2046 4516 -2033
rect 4568 -2046 4730 -2033
rect 4440 -2080 4730 -2046
rect 4620 -2414 4700 -2400
rect 4620 -2466 4629 -2414
rect 4681 -2466 4700 -2414
rect 4620 -2487 4700 -2466
rect 4620 -2543 4632 -2487
rect 4688 -2543 4700 -2487
rect 4620 -2570 4700 -2543
rect 4820 -2700 4900 -1136
rect 6190 -1119 6260 -1090
rect 6190 -1171 6199 -1119
rect 6251 -1150 6260 -1119
rect 6251 -1157 6370 -1150
rect 6251 -1171 6287 -1157
rect 6190 -1213 6287 -1171
rect 6343 -1213 6370 -1157
rect 6190 -1220 6370 -1213
rect 6420 -1497 6590 -1480
rect 6420 -1633 6437 -1497
rect 6573 -1633 6590 -1497
rect 6420 -1650 6590 -1633
rect 5270 -2307 5350 -2280
rect 5270 -2363 5282 -2307
rect 5338 -2363 5350 -2307
rect 5270 -2599 5350 -2363
rect 5270 -2651 5284 -2599
rect 5336 -2651 5350 -2599
rect 5270 -2670 5350 -2651
<< via2 >>
rect 6722 62 6778 118
rect 6427 -233 6483 -177
rect 5097 -478 5153 -422
rect 5887 -688 6023 -472
rect 4477 -1994 4533 -1977
rect 4557 -1994 4613 -1977
rect 4477 -2033 4504 -1994
rect 4504 -2033 4516 -1994
rect 4516 -2033 4533 -1994
rect 4557 -2033 4568 -1994
rect 4568 -2033 4613 -1994
rect 4637 -2033 4693 -1977
rect 4632 -2543 4688 -2487
rect 6287 -1213 6343 -1157
rect 6437 -1507 6573 -1497
rect 6437 -1623 6447 -1507
rect 6447 -1623 6563 -1507
rect 6563 -1623 6573 -1507
rect 6437 -1633 6573 -1623
rect 5282 -2363 5338 -2307
<< metal3 >>
rect 6710 120 6790 130
rect 3800 118 6800 120
rect 3800 62 6722 118
rect 6778 62 6800 118
rect 3800 50 6800 62
rect 6710 40 6790 50
rect 6410 -170 6500 -160
rect 3740 -177 6960 -170
rect 3740 -233 6427 -177
rect 6483 -233 6960 -177
rect 3740 -240 6960 -233
rect 6410 -250 6500 -240
rect 5310 -410 5770 -380
rect 5080 -420 5770 -410
rect 5070 -422 5770 -420
rect 5070 -478 5097 -422
rect 5153 -478 5770 -422
rect 5070 -490 5770 -478
rect 5080 -500 5770 -490
rect 5310 -840 5770 -500
rect 5850 -463 6300 -420
rect 5850 -687 5878 -463
rect 6022 -472 6300 -463
rect 5850 -688 5887 -687
rect 6023 -688 6300 -472
rect 5850 -730 6300 -688
rect 6260 -1150 6370 -1140
rect 3800 -1157 6800 -1150
rect 3800 -1213 6287 -1157
rect 6343 -1213 6800 -1157
rect 3800 -1220 6800 -1213
rect 6260 -1230 6370 -1220
rect 6420 -1493 6590 -1470
rect 6420 -1637 6433 -1493
rect 6577 -1637 6590 -1493
rect 6420 -1660 6590 -1637
rect 4440 -1723 4730 -1680
rect 4440 -1977 4518 -1723
rect 4662 -1977 4730 -1723
rect 4440 -2033 4477 -1977
rect 4533 -2033 4557 -2027
rect 4613 -2033 4637 -2027
rect 4693 -2033 4730 -1977
rect 4440 -2050 4730 -2033
rect 5250 -2307 5550 -2280
rect 5250 -2363 5282 -2307
rect 5338 -2308 5550 -2307
rect 5338 -2363 5453 -2308
rect 5250 -2372 5453 -2363
rect 5517 -2372 5550 -2308
rect 5250 -2400 5550 -2372
rect 3800 -2487 6800 -2470
rect 3800 -2540 4632 -2487
rect 4620 -2543 4632 -2540
rect 4688 -2540 6800 -2487
rect 4688 -2543 4700 -2540
rect 4620 -2560 4700 -2543
<< via3 >>
rect 5878 -472 6022 -463
rect 5878 -687 5887 -472
rect 5887 -687 6022 -472
rect 6433 -1497 6577 -1493
rect 6433 -1633 6437 -1497
rect 6437 -1633 6573 -1497
rect 6573 -1633 6577 -1497
rect 6433 -1637 6577 -1633
rect 4518 -1977 4662 -1723
rect 4518 -2027 4533 -1977
rect 4533 -2027 4557 -1977
rect 4557 -2027 4613 -1977
rect 4613 -2027 4637 -1977
rect 4637 -2027 4662 -1977
rect 5453 -2372 5517 -2308
<< mimcap >>
rect 5340 -508 5740 -410
rect 5340 -732 5513 -508
rect 5657 -732 5740 -508
rect 5340 -810 5740 -732
<< mimcapcontact >>
rect 5513 -732 5657 -508
<< metal4 >>
rect 5460 -457 6220 -310
rect 5460 -508 5812 -457
rect 5460 -732 5513 -508
rect 5657 -693 5812 -508
rect 6048 -693 6220 -457
rect 5657 -732 6220 -693
rect 5460 -770 6220 -732
rect 4280 -1250 6320 -1120
rect 4440 -1707 4730 -1680
rect 4440 -1943 4472 -1707
rect 4708 -1943 4730 -1707
rect 4440 -2027 4518 -1943
rect 4662 -2027 4730 -1943
rect 4440 -2050 4730 -2027
rect 5100 -2190 6130 -1250
rect 6430 -1480 6580 460
rect 6420 -1493 6590 -1480
rect 6420 -1637 6433 -1493
rect 6577 -1637 6590 -1493
rect 6420 -1650 6590 -1637
rect 5420 -2308 5590 -2190
rect 5420 -2372 5453 -2308
rect 5517 -2372 5590 -2308
rect 5420 -2670 5590 -2372
rect 6430 -2860 6580 -1650
<< via4 >>
rect 5812 -463 6048 -457
rect 5812 -687 5878 -463
rect 5878 -687 6022 -463
rect 6022 -687 6048 -463
rect 5812 -693 6048 -687
rect 4472 -1723 4708 -1707
rect 4472 -1943 4518 -1723
rect 4518 -1943 4662 -1723
rect 4662 -1943 4708 -1723
<< metal5 >>
rect 3640 140 6960 460
rect 3640 -2540 3960 140
rect 4280 -457 6320 -180
rect 4280 -693 5812 -457
rect 6048 -693 6320 -457
rect 4280 -1707 6320 -693
rect 4280 -1943 4472 -1707
rect 4708 -1943 6320 -1707
rect 4280 -2220 6320 -1943
rect 6640 -2540 6960 140
rect 3640 -2860 6960 -2540
<< glass >>
rect 4480 -2020 6120 -380
<< labels >>
rlabel metal5 s 6700 -1680 6700 -1680 4 gring
port 2 nsew
rlabel metal4 s 5570 -2360 5570 -2360 4 shield
port 4 nsew
rlabel locali s 6340 -500 6340 -500 4 test_net
port 5 nsew
rlabel metal1 s 3830 240 3830 240 4 VDD
port 7 nsew
rlabel metal1 s 3910 -2620 3910 -2620 4 GND
port 8 nsew
rlabel metal2 s 3870 290 3870 290 4 VREF
port 9 nsew
rlabel metal3 s 6780 -1180 6780 -1180 4 ROW_SEL
port 10 nsew
rlabel metal3 s 6770 -2510 6770 -2510 4 NB1
port 11 nsew
rlabel metal2 s 4330 290 4330 290 4 VBIAS
port 12 nsew
rlabel metal2 s 4860 280 4860 280 4 NB2
port 13 nsew
rlabel metal5 s 5690 -1950 5690 -1950 4 AMP_IN
port 14 nsew
rlabel metal3 s 6790 100 6790 100 4 SF_IB
port 15 nsew
rlabel metal4 s 6510 -2850 6510 -2850 4 PIX_OUT
port 16 nsew
rlabel metal3 s 3800 -200 3800 -200 4 CSA_VREF
port 17 nsew
<< end >>
