VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO /home/damic/CMOS/TopmetalSe/magic/pixel_array
  CLASS BLOCK ;
  FOREIGN /home/damic/CMOS/TopmetalSe/magic/pixel_array ;
  ORIGIN 2.800 35.500 ;
  SIZE 50.800 BY 53.500 ;
  PIN PIX0_IN
    ANTENNAGATEAREA 1.050000 ;
    ANTENNADIFFAREA 0.294000 ;
    PORT
      LAYER li1 ;
        RECT 14.200 11.950 14.650 12.320 ;
        RECT 14.350 10.600 14.650 11.950 ;
        RECT 13.000 10.350 14.650 10.600 ;
        RECT 13.000 10.050 13.650 10.350 ;
        RECT 3.200 2.450 3.900 3.100 ;
        RECT 2.450 2.150 3.900 2.450 ;
      LAYER mcon ;
        RECT 13.050 10.100 13.600 10.550 ;
        RECT 3.300 2.500 3.800 3.050 ;
      LAYER met1 ;
        RECT 11.300 10.050 13.700 10.600 ;
        RECT 3.200 2.400 3.900 3.750 ;
      LAYER via ;
        RECT 11.350 10.050 12.350 10.600 ;
        RECT 3.250 3.150 3.850 3.650 ;
      LAYER met2 ;
        RECT 10.350 9.950 12.450 11.300 ;
        RECT 3.200 3.100 4.650 3.750 ;
      LAYER via2 ;
        RECT 10.400 10.000 11.150 11.200 ;
        RECT 3.250 3.300 4.600 3.650 ;
      LAYER met3 ;
        RECT 10.250 9.850 12.500 11.400 ;
        RECT 3.200 3.250 4.650 5.100 ;
      LAYER via3 ;
        RECT 10.350 9.950 11.150 11.300 ;
        RECT 3.400 4.350 4.500 4.900 ;
        RECT 3.350 3.750 4.500 4.350 ;
        RECT 3.400 3.350 4.500 3.750 ;
      LAYER met4 ;
        RECT 8.300 9.650 12.100 11.950 ;
        RECT 3.200 3.250 4.650 5.100 ;
      LAYER via4 ;
        RECT 10.050 9.850 11.250 11.400 ;
        RECT 3.350 3.750 4.550 5.000 ;
      LAYER met5 ;
        RECT 2.400 2.400 12.600 12.600 ;
    END
  END PIX0_IN
  PIN VBIAS
    ANTENNAGATEAREA 4.800000 ;
    PORT
      LAYER li1 ;
        RECT 2.850 10.750 3.100 11.200 ;
        RECT 2.700 10.250 3.100 10.750 ;
        RECT 2.850 -4.250 3.100 -3.800 ;
        RECT 2.700 -4.750 3.100 -4.250 ;
        RECT 2.850 -19.250 3.100 -18.800 ;
        RECT 2.700 -19.750 3.100 -19.250 ;
      LAYER mcon ;
        RECT 2.850 10.800 3.100 11.200 ;
        RECT 2.850 -4.200 3.100 -3.800 ;
        RECT 2.850 -19.200 3.100 -18.800 ;
      LAYER met1 ;
        RECT 2.400 11.200 3.150 11.550 ;
        RECT 2.800 10.750 3.150 11.200 ;
        RECT 2.850 10.450 3.100 10.750 ;
        RECT 2.400 -3.800 3.150 -3.450 ;
        RECT 2.800 -4.250 3.150 -3.800 ;
        RECT 2.850 -4.550 3.100 -4.250 ;
        RECT 2.400 -18.800 3.150 -18.450 ;
        RECT 2.800 -19.250 3.150 -18.800 ;
        RECT 2.850 -19.550 3.100 -19.250 ;
      LAYER via ;
        RECT 2.450 11.250 2.800 11.550 ;
        RECT 2.450 -3.750 2.800 -3.450 ;
        RECT 2.450 -18.750 2.800 -18.450 ;
      LAYER met2 ;
        RECT 2.500 11.550 2.850 18.000 ;
        RECT 2.400 11.200 2.900 11.550 ;
        RECT 2.500 -3.450 2.850 11.200 ;
        RECT 2.400 -3.800 2.900 -3.450 ;
        RECT 2.500 -18.450 2.850 -3.800 ;
        RECT 2.400 -18.800 2.900 -18.450 ;
        RECT 2.500 -30.000 2.850 -18.800 ;
    END
  END VBIAS
  PIN VREF
    ANTENNAGATEAREA 3.150000 ;
    PORT
      LAYER li1 ;
        RECT 0.250 2.000 0.700 2.750 ;
        RECT 0.250 -13.000 0.700 -12.250 ;
        RECT 0.250 -28.000 0.700 -27.250 ;
      LAYER mcon ;
        RECT 0.350 2.500 0.600 2.750 ;
        RECT 0.350 -12.500 0.600 -12.250 ;
        RECT 0.350 -27.500 0.600 -27.250 ;
      LAYER met1 ;
        RECT 0.250 2.450 0.700 3.200 ;
        RECT 0.250 -12.550 0.700 -11.800 ;
        RECT 0.250 -27.550 0.700 -26.800 ;
      LAYER via ;
        RECT 0.300 2.800 0.650 3.150 ;
        RECT 0.300 -12.200 0.650 -11.850 ;
        RECT 0.300 -27.200 0.650 -26.850 ;
      LAYER met2 ;
        RECT 0.300 -30.000 0.650 18.000 ;
    END
  END VREF
  PIN NB2
    ANTENNAGATEAREA 3.450000 ;
    PORT
      LAYER li1 ;
        RECT 5.050 8.450 5.650 9.300 ;
        RECT 5.100 8.050 5.650 8.450 ;
        RECT 5.050 -6.550 5.650 -5.700 ;
        RECT 5.100 -6.950 5.650 -6.550 ;
        RECT 5.050 -21.550 5.650 -20.700 ;
        RECT 5.100 -21.950 5.650 -21.550 ;
      LAYER mcon ;
        RECT 5.150 8.100 5.600 8.350 ;
        RECT 5.150 -6.900 5.600 -6.650 ;
        RECT 5.150 -21.900 5.600 -21.650 ;
      LAYER met1 ;
        RECT 4.950 7.750 5.650 8.450 ;
        RECT 4.950 -7.250 5.650 -6.550 ;
        RECT 4.950 -22.250 5.650 -21.550 ;
      LAYER via ;
        RECT 5.100 7.800 5.500 8.100 ;
        RECT 5.100 -7.200 5.500 -6.900 ;
        RECT 5.100 -22.200 5.500 -21.900 ;
      LAYER met2 ;
        RECT 5.100 15.000 5.450 18.000 ;
        RECT 5.100 -30.000 5.500 15.000 ;
    END
  END NB2
  PIN VDD
    ANTENNADIFFAREA 6.600000 ;
    PORT
      LAYER nwell ;
        RECT 0.000 11.600 45.000 15.000 ;
      LAYER li1 ;
        RECT 5.450 14.550 5.950 14.850 ;
        RECT 14.250 14.800 14.450 14.850 ;
        RECT 14.150 14.600 14.550 14.800 ;
        RECT 5.100 13.550 6.300 14.550 ;
        RECT 14.250 13.400 14.450 14.600 ;
        RECT 20.450 14.550 20.950 14.850 ;
        RECT 29.250 14.800 29.450 14.850 ;
        RECT 29.150 14.600 29.550 14.800 ;
        RECT 20.100 13.550 21.300 14.550 ;
        RECT 29.250 13.400 29.450 14.600 ;
        RECT 35.450 14.550 35.950 14.850 ;
        RECT 44.250 14.800 44.450 14.850 ;
        RECT 44.150 14.600 44.550 14.800 ;
        RECT 35.100 13.550 36.300 14.550 ;
        RECT 44.250 13.400 44.450 14.600 ;
        RECT 4.250 12.050 4.600 12.250 ;
        RECT 19.250 12.050 19.600 12.250 ;
        RECT 34.250 12.050 34.600 12.250 ;
        RECT 4.250 11.250 4.450 12.050 ;
        RECT 19.250 11.250 19.450 12.050 ;
        RECT 34.250 11.250 34.450 12.050 ;
        RECT 4.100 11.000 5.000 11.250 ;
        RECT 19.100 11.000 20.000 11.250 ;
        RECT 34.100 11.000 35.000 11.250 ;
        RECT 9.800 10.400 10.150 10.950 ;
        RECT 24.800 10.400 25.150 10.950 ;
        RECT 39.800 10.400 40.150 10.950 ;
        RECT 9.800 10.100 10.700 10.400 ;
        RECT 24.800 10.100 25.700 10.400 ;
        RECT 39.800 10.100 40.700 10.400 ;
      LAYER mcon ;
        RECT 5.500 14.550 5.900 14.800 ;
        RECT 20.500 14.550 20.900 14.800 ;
        RECT 35.500 14.550 35.900 14.800 ;
        RECT 9.850 10.250 10.100 10.900 ;
        RECT 24.850 10.250 25.100 10.900 ;
        RECT 39.850 10.250 40.100 10.900 ;
      LAYER met1 ;
        RECT -2.800 14.400 45.000 14.850 ;
        RECT 0.000 14.100 45.000 14.400 ;
        RECT 4.550 12.350 5.050 14.100 ;
        RECT 4.150 12.000 5.050 12.350 ;
        RECT 9.800 10.150 10.150 14.100 ;
        RECT 19.550 12.350 20.050 14.100 ;
        RECT 19.150 12.000 20.050 12.350 ;
        RECT 24.800 10.150 25.150 14.100 ;
        RECT 34.550 12.350 35.050 14.100 ;
        RECT 34.150 12.000 35.050 12.350 ;
        RECT 39.800 10.150 40.150 14.100 ;
    END
  END VDD
  PIN SF_IB
    ANTENNAGATEAREA 3.000000 ;
    PORT
      LAYER li1 ;
        RECT 13.700 12.800 14.600 13.050 ;
        RECT 28.700 12.800 29.600 13.050 ;
        RECT 43.700 12.800 44.600 13.050 ;
      LAYER mcon ;
        RECT 14.400 12.800 14.600 13.050 ;
        RECT 29.400 12.800 29.600 13.050 ;
        RECT 44.400 12.800 44.600 13.050 ;
      LAYER met1 ;
        RECT 14.300 12.750 14.950 13.100 ;
        RECT 29.300 12.750 29.950 13.100 ;
        RECT 44.300 12.750 44.950 13.100 ;
      LAYER via ;
        RECT 14.600 12.750 14.900 13.100 ;
        RECT 29.600 12.750 29.900 13.100 ;
        RECT 44.600 12.750 44.900 13.100 ;
      LAYER met2 ;
        RECT 14.600 12.650 14.900 14.150 ;
        RECT 29.600 12.650 29.900 14.150 ;
        RECT 44.600 12.650 44.900 14.150 ;
      LAYER via2 ;
        RECT 14.600 13.800 14.900 14.100 ;
        RECT 29.600 13.800 29.900 14.100 ;
        RECT 44.600 13.800 44.900 14.100 ;
      LAYER met3 ;
        RECT -2.800 14.100 0.200 14.200 ;
        RECT 14.550 14.100 14.950 14.150 ;
        RECT 29.550 14.100 29.950 14.150 ;
        RECT 44.550 14.100 44.950 14.150 ;
        RECT -2.800 13.750 45.000 14.100 ;
        RECT 14.550 13.700 14.950 13.750 ;
        RECT 29.550 13.700 29.950 13.750 ;
        RECT 44.550 13.700 44.950 13.750 ;
    END
  END SF_IB
  PIN CSA_VREF
    ANTENNAGATEAREA 10.080000 ;
    PORT
      LAYER li1 ;
        RECT 13.600 11.350 14.050 11.650 ;
        RECT 28.600 11.350 29.050 11.650 ;
        RECT 43.600 11.350 44.050 11.650 ;
        RECT 13.150 11.100 14.100 11.350 ;
        RECT 28.150 11.100 29.100 11.350 ;
        RECT 43.150 11.100 44.100 11.350 ;
      LAYER met1 ;
        RECT 13.050 11.000 13.500 11.500 ;
        RECT 28.050 11.000 28.500 11.500 ;
        RECT 43.050 11.000 43.500 11.500 ;
      LAYER via ;
        RECT 13.100 11.000 13.450 11.500 ;
        RECT 28.100 11.000 28.450 11.500 ;
        RECT 43.100 11.000 43.450 11.500 ;
      LAYER met2 ;
        RECT 13.100 10.950 13.450 12.750 ;
        RECT 28.100 10.950 28.450 12.750 ;
        RECT 43.100 10.950 43.450 12.750 ;
      LAYER via2 ;
        RECT 13.100 12.300 13.450 12.650 ;
        RECT 28.100 12.300 28.450 12.650 ;
        RECT 43.100 12.300 43.450 12.650 ;
      LAYER met3 ;
        RECT -2.800 12.650 0.200 12.750 ;
        RECT 13.050 12.650 13.500 12.700 ;
        RECT 28.050 12.650 28.500 12.700 ;
        RECT 43.050 12.650 43.500 12.700 ;
        RECT -2.800 12.300 45.800 12.650 ;
        RECT 13.050 12.250 13.500 12.300 ;
        RECT 28.050 12.250 28.500 12.300 ;
        RECT 43.050 12.250 43.500 12.300 ;
    END
  END CSA_VREF
  PIN NB1
    ANTENNAGATEAREA 3.600000 ;
    PORT
      LAYER li1 ;
        RECT 3.550 1.150 4.000 1.450 ;
        RECT 18.550 1.150 19.000 1.450 ;
        RECT 33.550 1.150 34.000 1.450 ;
        RECT 3.550 0.750 3.900 1.150 ;
        RECT 18.550 0.750 18.900 1.150 ;
        RECT 33.550 0.750 33.900 1.150 ;
      LAYER mcon ;
        RECT 3.600 1.200 3.950 1.400 ;
        RECT 18.600 1.200 18.950 1.400 ;
        RECT 33.600 1.200 33.950 1.400 ;
      LAYER met1 ;
        RECT 3.500 1.150 4.500 1.450 ;
        RECT 18.500 1.150 19.500 1.450 ;
        RECT 33.500 1.150 34.500 1.450 ;
      LAYER via ;
        RECT 4.100 1.150 4.450 1.450 ;
        RECT 19.100 1.150 19.450 1.450 ;
        RECT 34.100 1.150 34.450 1.450 ;
      LAYER met2 ;
        RECT 4.100 0.650 4.500 1.500 ;
        RECT 19.100 0.650 19.500 1.500 ;
        RECT 34.100 0.650 34.500 1.500 ;
      LAYER via2 ;
        RECT 4.150 0.750 4.450 1.100 ;
        RECT 19.150 0.750 19.450 1.100 ;
        RECT 34.150 0.750 34.450 1.100 ;
      LAYER met3 ;
        RECT -2.800 1.150 0.200 1.250 ;
        RECT -2.800 0.800 45.000 1.150 ;
        RECT 4.100 0.700 4.500 0.800 ;
        RECT 19.100 0.700 19.500 0.800 ;
        RECT 34.100 0.700 34.500 0.800 ;
    END
  END NB1
  PIN ROW_SEL0
    ANTENNAGATEAREA 6.000000 ;
    PORT
      LAYER li1 ;
        RECT 12.000 7.950 12.250 9.000 ;
        RECT 27.000 7.950 27.250 9.000 ;
        RECT 42.000 7.950 42.250 9.000 ;
      LAYER mcon ;
        RECT 12.000 8.050 12.250 8.400 ;
        RECT 27.000 8.050 27.250 8.400 ;
        RECT 42.000 8.050 42.250 8.400 ;
      LAYER met1 ;
        RECT 11.950 7.500 12.300 8.500 ;
        RECT 26.950 7.500 27.300 8.500 ;
        RECT 41.950 7.500 42.300 8.500 ;
      LAYER via ;
        RECT 11.950 7.550 12.300 8.000 ;
        RECT 26.950 7.550 27.300 8.000 ;
        RECT 41.950 7.550 42.300 8.000 ;
      LAYER met2 ;
        RECT 11.950 7.750 12.300 8.050 ;
        RECT 26.950 7.750 27.300 8.050 ;
        RECT 41.950 7.750 42.300 8.050 ;
        RECT 11.950 7.400 12.850 7.750 ;
        RECT 26.950 7.400 27.850 7.750 ;
        RECT 41.950 7.400 42.850 7.750 ;
      LAYER via2 ;
        RECT 12.350 7.400 12.800 7.750 ;
        RECT 27.350 7.400 27.800 7.750 ;
        RECT 42.350 7.400 42.800 7.750 ;
      LAYER met3 ;
        RECT -2.800 7.750 0.200 7.850 ;
        RECT 12.300 7.750 12.850 7.800 ;
        RECT 27.300 7.750 27.850 7.800 ;
        RECT 42.300 7.750 42.850 7.800 ;
        RECT -2.800 7.400 45.000 7.750 ;
        RECT 12.300 7.350 12.850 7.400 ;
        RECT 27.300 7.350 27.850 7.400 ;
        RECT 42.300 7.350 42.850 7.400 ;
    END
  END ROW_SEL0
  PIN PIX1_IN
    ANTENNAGATEAREA 1.050000 ;
    ANTENNADIFFAREA 0.294000 ;
    PORT
      LAYER li1 ;
        RECT 29.200 11.950 29.650 12.320 ;
        RECT 29.350 10.600 29.650 11.950 ;
        RECT 28.000 10.350 29.650 10.600 ;
        RECT 28.000 10.050 28.650 10.350 ;
        RECT 18.200 2.450 18.900 3.100 ;
        RECT 17.450 2.150 18.900 2.450 ;
      LAYER mcon ;
        RECT 28.050 10.100 28.600 10.550 ;
        RECT 18.300 2.500 18.800 3.050 ;
      LAYER met1 ;
        RECT 26.300 10.050 28.700 10.600 ;
        RECT 18.200 2.400 18.900 3.750 ;
      LAYER via ;
        RECT 26.350 10.050 27.350 10.600 ;
        RECT 18.250 3.150 18.850 3.650 ;
      LAYER met2 ;
        RECT 25.350 9.950 27.450 11.300 ;
        RECT 18.200 3.100 19.650 3.750 ;
      LAYER via2 ;
        RECT 25.400 10.000 26.150 11.200 ;
        RECT 18.250 3.300 19.600 3.650 ;
      LAYER met3 ;
        RECT 25.250 9.850 27.500 11.400 ;
        RECT 18.200 3.250 19.650 5.100 ;
      LAYER via3 ;
        RECT 25.350 9.950 26.150 11.300 ;
        RECT 18.400 4.350 19.500 4.900 ;
        RECT 18.350 3.750 19.500 4.350 ;
        RECT 18.400 3.350 19.500 3.750 ;
      LAYER met4 ;
        RECT 23.300 9.650 27.100 11.950 ;
        RECT 18.200 3.250 19.650 5.100 ;
      LAYER via4 ;
        RECT 25.050 9.850 26.250 11.400 ;
        RECT 18.350 3.750 19.550 5.000 ;
      LAYER met5 ;
        RECT 17.400 2.400 27.600 12.600 ;
    END
  END PIX1_IN
  PIN PIX2_IN
    ANTENNAGATEAREA 1.050000 ;
    ANTENNADIFFAREA 0.294000 ;
    PORT
      LAYER li1 ;
        RECT 44.200 11.950 44.650 12.320 ;
        RECT 44.350 10.600 44.650 11.950 ;
        RECT 43.000 10.350 44.650 10.600 ;
        RECT 43.000 10.050 43.650 10.350 ;
        RECT 33.200 2.450 33.900 3.100 ;
        RECT 32.450 2.150 33.900 2.450 ;
      LAYER mcon ;
        RECT 43.050 10.100 43.600 10.550 ;
        RECT 33.300 2.500 33.800 3.050 ;
      LAYER met1 ;
        RECT 41.300 10.050 43.700 10.600 ;
        RECT 33.200 2.400 33.900 3.750 ;
      LAYER via ;
        RECT 41.350 10.050 42.350 10.600 ;
        RECT 33.250 3.150 33.850 3.650 ;
      LAYER met2 ;
        RECT 40.350 9.950 42.450 11.300 ;
        RECT 33.200 3.100 34.650 3.750 ;
      LAYER via2 ;
        RECT 40.400 10.000 41.150 11.200 ;
        RECT 33.250 3.300 34.600 3.650 ;
      LAYER met3 ;
        RECT 40.250 9.850 42.500 11.400 ;
        RECT 33.200 3.250 34.650 5.100 ;
      LAYER via3 ;
        RECT 40.350 9.950 41.150 11.300 ;
        RECT 33.400 4.350 34.500 4.900 ;
        RECT 33.350 3.750 34.500 4.350 ;
        RECT 33.400 3.350 34.500 3.750 ;
      LAYER met4 ;
        RECT 38.300 9.650 42.100 11.950 ;
        RECT 33.200 3.250 34.650 5.100 ;
      LAYER via4 ;
        RECT 40.050 9.850 41.250 11.400 ;
        RECT 33.350 3.750 34.550 5.000 ;
      LAYER met5 ;
        RECT 32.400 2.400 42.600 12.600 ;
    END
  END PIX2_IN
  PIN GND
    ANTENNADIFFAREA 5.250000 ;
    PORT
      LAYER li1 ;
        RECT 11.150 13.400 11.550 14.400 ;
        RECT 26.150 13.400 26.550 14.400 ;
        RECT 41.150 13.400 41.550 14.400 ;
        RECT 11.150 12.250 11.400 13.400 ;
        RECT 26.150 12.250 26.400 13.400 ;
        RECT 41.150 12.250 41.400 13.400 ;
        RECT 10.350 11.900 11.400 12.250 ;
        RECT 25.350 11.900 26.400 12.250 ;
        RECT 40.350 11.900 41.400 12.250 ;
        RECT 4.000 7.800 4.900 8.250 ;
        RECT 19.000 7.800 19.900 8.250 ;
        RECT 34.000 7.800 34.900 8.250 ;
        RECT 4.000 5.600 4.500 7.800 ;
        RECT 19.000 5.600 19.500 7.800 ;
        RECT 34.000 5.600 34.500 7.800 ;
        RECT 2.650 0.550 3.350 1.750 ;
        RECT 17.650 0.550 18.350 1.750 ;
        RECT 32.650 0.550 33.350 1.750 ;
        RECT 2.900 0.150 3.150 0.550 ;
        RECT 17.900 0.150 18.150 0.550 ;
        RECT 32.900 0.150 33.150 0.550 ;
      LAYER mcon ;
        RECT 10.400 11.950 10.850 12.250 ;
        RECT 25.400 11.950 25.850 12.250 ;
        RECT 40.400 11.950 40.850 12.250 ;
        RECT 4.050 5.650 4.450 6.050 ;
        RECT 19.050 5.650 19.450 6.050 ;
        RECT 34.050 5.650 34.450 6.050 ;
        RECT 2.900 0.200 3.100 0.400 ;
        RECT 17.900 0.200 18.100 0.400 ;
        RECT 32.900 0.200 33.100 0.400 ;
      LAYER met1 ;
        RECT 10.350 11.900 10.950 12.350 ;
        RECT 25.350 11.900 25.950 12.350 ;
        RECT 40.350 11.900 40.950 12.350 ;
        RECT 3.950 5.600 6.500 6.100 ;
        RECT 5.950 0.900 6.500 5.600 ;
        RECT 10.350 0.900 10.850 11.900 ;
        RECT 18.950 5.600 21.500 6.100 ;
        RECT 20.950 0.900 21.500 5.600 ;
        RECT 25.350 0.900 25.850 11.900 ;
        RECT 33.950 5.600 36.500 6.100 ;
        RECT 35.950 0.900 36.500 5.600 ;
        RECT 40.350 0.900 40.850 11.900 ;
        RECT 0.000 0.600 45.000 0.900 ;
        RECT 0.000 0.150 48.000 0.600 ;
      LAYER via ;
        RECT 7.350 0.200 7.750 0.550 ;
        RECT 22.350 0.200 22.750 0.550 ;
        RECT 37.350 0.200 37.750 0.550 ;
      LAYER met2 ;
        RECT 7.350 0.150 7.750 2.100 ;
        RECT 22.350 0.150 22.750 2.100 ;
        RECT 37.350 0.150 37.750 2.100 ;
      LAYER via2 ;
        RECT 7.400 1.600 7.700 2.050 ;
        RECT 22.400 1.600 22.700 2.050 ;
        RECT 37.400 1.600 37.700 2.050 ;
      LAYER met3 ;
        RECT 7.250 1.500 8.750 2.100 ;
        RECT 22.250 1.500 23.750 2.100 ;
        RECT 37.250 1.500 38.750 2.100 ;
      LAYER via3 ;
        RECT 8.150 1.550 8.700 2.050 ;
        RECT 23.150 1.550 23.700 2.050 ;
        RECT 38.150 1.550 38.700 2.050 ;
      LAYER met4 ;
        RECT 2.400 7.250 12.600 7.900 ;
        RECT 17.400 7.250 27.600 7.900 ;
        RECT 32.400 7.250 42.600 7.900 ;
        RECT 6.500 2.550 11.650 7.250 ;
        RECT 21.500 2.550 26.650 7.250 ;
        RECT 36.500 2.550 41.650 7.250 ;
        RECT 8.100 0.150 8.950 2.550 ;
        RECT 23.100 0.150 23.950 2.550 ;
        RECT 38.100 0.150 38.950 2.550 ;
    END
  END GND
  PIN PIX3_IN
    ANTENNAGATEAREA 1.050000 ;
    ANTENNADIFFAREA 0.294000 ;
    PORT
      LAYER li1 ;
        RECT 14.200 -3.050 14.650 -2.680 ;
        RECT 14.350 -4.400 14.650 -3.050 ;
        RECT 13.000 -4.650 14.650 -4.400 ;
        RECT 13.000 -4.950 13.650 -4.650 ;
        RECT 3.200 -12.550 3.900 -11.900 ;
        RECT 2.450 -12.850 3.900 -12.550 ;
      LAYER mcon ;
        RECT 13.050 -4.900 13.600 -4.450 ;
        RECT 3.300 -12.500 3.800 -11.950 ;
      LAYER met1 ;
        RECT 11.300 -4.950 13.700 -4.400 ;
        RECT 3.200 -12.600 3.900 -11.250 ;
      LAYER via ;
        RECT 11.350 -4.950 12.350 -4.400 ;
        RECT 3.250 -11.850 3.850 -11.350 ;
      LAYER met2 ;
        RECT 10.350 -5.050 12.450 -3.700 ;
        RECT 3.200 -11.900 4.650 -11.250 ;
      LAYER via2 ;
        RECT 10.400 -5.000 11.150 -3.800 ;
        RECT 3.250 -11.700 4.600 -11.350 ;
      LAYER met3 ;
        RECT 10.250 -5.150 12.500 -3.600 ;
        RECT 3.200 -11.750 4.650 -9.900 ;
      LAYER via3 ;
        RECT 10.350 -5.050 11.150 -3.700 ;
        RECT 3.400 -10.650 4.500 -10.100 ;
        RECT 3.350 -11.250 4.500 -10.650 ;
        RECT 3.400 -11.650 4.500 -11.250 ;
      LAYER met4 ;
        RECT 8.300 -5.350 12.100 -3.050 ;
        RECT 3.200 -11.750 4.650 -9.900 ;
      LAYER via4 ;
        RECT 10.050 -5.150 11.250 -3.600 ;
        RECT 3.350 -11.250 4.550 -10.000 ;
      LAYER met5 ;
        RECT 2.400 -12.600 12.600 -2.400 ;
    END
  END PIX3_IN
  PIN ROW_SEL1
    ANTENNAGATEAREA 6.000000 ;
    PORT
      LAYER li1 ;
        RECT 12.000 -7.050 12.250 -6.000 ;
        RECT 27.000 -7.050 27.250 -6.000 ;
        RECT 42.000 -7.050 42.250 -6.000 ;
      LAYER mcon ;
        RECT 12.000 -6.950 12.250 -6.600 ;
        RECT 27.000 -6.950 27.250 -6.600 ;
        RECT 42.000 -6.950 42.250 -6.600 ;
      LAYER met1 ;
        RECT 11.950 -7.500 12.300 -6.500 ;
        RECT 26.950 -7.500 27.300 -6.500 ;
        RECT 41.950 -7.500 42.300 -6.500 ;
      LAYER via ;
        RECT 11.950 -7.450 12.300 -7.000 ;
        RECT 26.950 -7.450 27.300 -7.000 ;
        RECT 41.950 -7.450 42.300 -7.000 ;
      LAYER met2 ;
        RECT 11.950 -7.250 12.300 -6.950 ;
        RECT 26.950 -7.250 27.300 -6.950 ;
        RECT 41.950 -7.250 42.300 -6.950 ;
        RECT 11.950 -7.600 12.850 -7.250 ;
        RECT 26.950 -7.600 27.850 -7.250 ;
        RECT 41.950 -7.600 42.850 -7.250 ;
      LAYER via2 ;
        RECT 12.350 -7.600 12.800 -7.250 ;
        RECT 27.350 -7.600 27.800 -7.250 ;
        RECT 42.350 -7.600 42.800 -7.250 ;
      LAYER met3 ;
        RECT -2.800 -7.250 0.200 -7.150 ;
        RECT 12.300 -7.250 12.850 -7.200 ;
        RECT 27.300 -7.250 27.850 -7.200 ;
        RECT 42.300 -7.250 42.850 -7.200 ;
        RECT -2.800 -7.600 45.000 -7.250 ;
        RECT 12.300 -7.650 12.850 -7.600 ;
        RECT 27.300 -7.650 27.850 -7.600 ;
        RECT 42.300 -7.650 42.850 -7.600 ;
    END
  END ROW_SEL1
  PIN PIX4_IN
    ANTENNAGATEAREA 1.050000 ;
    ANTENNADIFFAREA 0.294000 ;
    PORT
      LAYER li1 ;
        RECT 29.200 -3.050 29.650 -2.680 ;
        RECT 29.350 -4.400 29.650 -3.050 ;
        RECT 28.000 -4.650 29.650 -4.400 ;
        RECT 28.000 -4.950 28.650 -4.650 ;
        RECT 18.200 -12.550 18.900 -11.900 ;
        RECT 17.450 -12.850 18.900 -12.550 ;
      LAYER mcon ;
        RECT 28.050 -4.900 28.600 -4.450 ;
        RECT 18.300 -12.500 18.800 -11.950 ;
      LAYER met1 ;
        RECT 26.300 -4.950 28.700 -4.400 ;
        RECT 18.200 -12.600 18.900 -11.250 ;
      LAYER via ;
        RECT 26.350 -4.950 27.350 -4.400 ;
        RECT 18.250 -11.850 18.850 -11.350 ;
      LAYER met2 ;
        RECT 25.350 -5.050 27.450 -3.700 ;
        RECT 18.200 -11.900 19.650 -11.250 ;
      LAYER via2 ;
        RECT 25.400 -5.000 26.150 -3.800 ;
        RECT 18.250 -11.700 19.600 -11.350 ;
      LAYER met3 ;
        RECT 25.250 -5.150 27.500 -3.600 ;
        RECT 18.200 -11.750 19.650 -9.900 ;
      LAYER via3 ;
        RECT 25.350 -5.050 26.150 -3.700 ;
        RECT 18.400 -10.650 19.500 -10.100 ;
        RECT 18.350 -11.250 19.500 -10.650 ;
        RECT 18.400 -11.650 19.500 -11.250 ;
      LAYER met4 ;
        RECT 23.300 -5.350 27.100 -3.050 ;
        RECT 18.200 -11.750 19.650 -9.900 ;
      LAYER via4 ;
        RECT 25.050 -5.150 26.250 -3.600 ;
        RECT 18.350 -11.250 19.550 -10.000 ;
      LAYER met5 ;
        RECT 17.400 -12.600 27.600 -2.400 ;
    END
  END PIX4_IN
  PIN PIX5_IN
    ANTENNAGATEAREA 1.050000 ;
    ANTENNADIFFAREA 0.294000 ;
    PORT
      LAYER li1 ;
        RECT 44.200 -3.050 44.650 -2.680 ;
        RECT 44.350 -4.400 44.650 -3.050 ;
        RECT 43.000 -4.650 44.650 -4.400 ;
        RECT 43.000 -4.950 43.650 -4.650 ;
        RECT 33.200 -12.550 33.900 -11.900 ;
        RECT 32.450 -12.850 33.900 -12.550 ;
      LAYER mcon ;
        RECT 43.050 -4.900 43.600 -4.450 ;
        RECT 33.300 -12.500 33.800 -11.950 ;
      LAYER met1 ;
        RECT 41.300 -4.950 43.700 -4.400 ;
        RECT 33.200 -12.600 33.900 -11.250 ;
      LAYER via ;
        RECT 41.350 -4.950 42.350 -4.400 ;
        RECT 33.250 -11.850 33.850 -11.350 ;
      LAYER met2 ;
        RECT 40.350 -5.050 42.450 -3.700 ;
        RECT 33.200 -11.900 34.650 -11.250 ;
      LAYER via2 ;
        RECT 40.400 -5.000 41.150 -3.800 ;
        RECT 33.250 -11.700 34.600 -11.350 ;
      LAYER met3 ;
        RECT 40.250 -5.150 42.500 -3.600 ;
        RECT 33.200 -11.750 34.650 -9.900 ;
      LAYER via3 ;
        RECT 40.350 -5.050 41.150 -3.700 ;
        RECT 33.400 -10.650 34.500 -10.100 ;
        RECT 33.350 -11.250 34.500 -10.650 ;
        RECT 33.400 -11.650 34.500 -11.250 ;
      LAYER met4 ;
        RECT 38.300 -5.350 42.100 -3.050 ;
        RECT 33.200 -11.750 34.650 -9.900 ;
      LAYER via4 ;
        RECT 40.050 -5.150 41.250 -3.600 ;
        RECT 33.350 -11.250 34.550 -10.000 ;
      LAYER met5 ;
        RECT 32.400 -12.600 42.600 -2.400 ;
    END
  END PIX5_IN
  PIN PIX6_IN
    ANTENNAGATEAREA 1.050000 ;
    ANTENNADIFFAREA 0.294000 ;
    PORT
      LAYER li1 ;
        RECT 14.200 -18.050 14.650 -17.680 ;
        RECT 14.350 -19.400 14.650 -18.050 ;
        RECT 13.000 -19.650 14.650 -19.400 ;
        RECT 13.000 -19.950 13.650 -19.650 ;
        RECT 3.200 -27.550 3.900 -26.900 ;
        RECT 2.450 -27.850 3.900 -27.550 ;
      LAYER mcon ;
        RECT 13.050 -19.900 13.600 -19.450 ;
        RECT 3.300 -27.500 3.800 -26.950 ;
      LAYER met1 ;
        RECT 11.300 -19.950 13.700 -19.400 ;
        RECT 3.200 -27.600 3.900 -26.250 ;
      LAYER via ;
        RECT 11.350 -19.950 12.350 -19.400 ;
        RECT 3.250 -26.850 3.850 -26.350 ;
      LAYER met2 ;
        RECT 10.350 -20.050 12.450 -18.700 ;
        RECT 3.200 -26.900 4.650 -26.250 ;
      LAYER via2 ;
        RECT 10.400 -20.000 11.150 -18.800 ;
        RECT 3.250 -26.700 4.600 -26.350 ;
      LAYER met3 ;
        RECT 10.250 -20.150 12.500 -18.600 ;
        RECT 3.200 -26.750 4.650 -24.900 ;
      LAYER via3 ;
        RECT 10.350 -20.050 11.150 -18.700 ;
        RECT 3.400 -25.650 4.500 -25.100 ;
        RECT 3.350 -26.250 4.500 -25.650 ;
        RECT 3.400 -26.650 4.500 -26.250 ;
      LAYER met4 ;
        RECT 8.300 -20.350 12.100 -18.050 ;
        RECT 3.200 -26.750 4.650 -24.900 ;
      LAYER via4 ;
        RECT 10.050 -20.150 11.250 -18.600 ;
        RECT 3.350 -26.250 4.550 -25.000 ;
      LAYER met5 ;
        RECT 2.400 -27.600 12.600 -17.400 ;
    END
  END PIX6_IN
  PIN PIX_OUT0
    ANTENNADIFFAREA 6.400000 ;
    PORT
      LAYER li1 ;
        RECT 9.750 7.450 11.700 7.800 ;
        RECT 10.950 6.050 11.700 7.450 ;
        RECT 10.950 5.300 13.950 6.050 ;
        RECT 9.750 -7.550 11.700 -7.200 ;
        RECT 10.950 -8.950 11.700 -7.550 ;
        RECT 10.950 -9.700 13.950 -8.950 ;
        RECT 9.750 -22.550 11.700 -22.200 ;
        RECT 10.950 -23.950 11.700 -22.550 ;
        RECT 10.950 -24.700 13.950 -23.950 ;
        RECT 2.700 -31.900 10.700 -31.150 ;
      LAYER mcon ;
        RECT 13.200 5.350 13.850 6.000 ;
        RECT 13.200 -9.650 13.850 -9.000 ;
        RECT 13.200 -24.650 13.850 -24.000 ;
        RECT 2.800 -31.450 10.600 -31.150 ;
      LAYER met1 ;
        RECT 13.100 5.300 13.950 6.050 ;
        RECT 13.100 -9.700 13.950 -8.950 ;
        RECT 13.100 -24.700 13.950 -23.950 ;
        RECT 2.700 -31.500 10.700 -30.650 ;
      LAYER via ;
        RECT 13.150 5.300 13.900 6.050 ;
        RECT 13.150 -9.700 13.900 -8.950 ;
        RECT 13.150 -24.700 13.900 -23.950 ;
        RECT 2.800 -31.000 10.600 -30.650 ;
      LAYER met2 ;
        RECT 13.100 5.250 13.950 6.100 ;
        RECT 13.100 -9.750 13.950 -8.900 ;
        RECT 13.100 -24.750 13.950 -23.900 ;
        RECT 2.700 -31.000 13.900 -30.300 ;
      LAYER via2 ;
        RECT 13.150 5.300 13.900 6.050 ;
        RECT 13.150 -9.700 13.900 -8.950 ;
        RECT 13.150 -24.700 13.900 -23.950 ;
        RECT 2.800 -30.900 13.800 -30.400 ;
      LAYER met3 ;
        RECT 13.100 5.200 13.950 6.150 ;
        RECT 13.100 -9.800 13.950 -8.850 ;
        RECT 13.100 -24.800 13.950 -23.850 ;
        RECT 2.700 -31.000 13.900 -30.300 ;
      LAYER via3 ;
        RECT 13.150 5.300 13.900 6.050 ;
        RECT 13.150 -9.700 13.900 -8.950 ;
        RECT 13.150 -24.700 13.900 -23.950 ;
        RECT 2.800 -30.900 13.800 -30.400 ;
      LAYER met4 ;
        RECT 13.150 6.100 13.900 15.800 ;
        RECT 13.100 5.250 13.950 6.100 ;
        RECT 13.150 -8.900 13.900 5.250 ;
        RECT 13.100 -9.750 13.950 -8.900 ;
        RECT 13.150 -23.900 13.900 -9.750 ;
        RECT 13.100 -24.750 13.950 -23.900 ;
        RECT 13.150 -30.300 13.900 -24.750 ;
        RECT 2.700 -31.000 13.900 -30.300 ;
    END
  END PIX_OUT0
  PIN COL_SEL0
    ANTENNAGATEAREA 16.000000 ;
    PORT
      LAYER li1 ;
        RECT 1.100 -33.550 2.200 -32.450 ;
      LAYER mcon ;
        RECT 1.200 -33.500 2.100 -32.500 ;
      LAYER met1 ;
        RECT 1.100 -33.550 2.200 -32.450 ;
      LAYER via ;
        RECT 1.200 -33.500 2.100 -32.500 ;
      LAYER met2 ;
        RECT 1.100 -33.550 2.200 -32.450 ;
      LAYER via2 ;
        RECT 1.200 -33.500 2.100 -32.500 ;
      LAYER met3 ;
        RECT 1.100 -33.550 2.200 -32.450 ;
      LAYER via3 ;
        RECT 1.200 -33.500 2.100 -32.500 ;
      LAYER met4 ;
        RECT 1.100 -35.500 2.200 -32.450 ;
    END
  END COL_SEL0
  PIN ROW_SEL2
    ANTENNAGATEAREA 6.000000 ;
    PORT
      LAYER li1 ;
        RECT 12.000 -22.050 12.250 -21.000 ;
        RECT 27.000 -22.050 27.250 -21.000 ;
        RECT 42.000 -22.050 42.250 -21.000 ;
      LAYER mcon ;
        RECT 12.000 -21.950 12.250 -21.600 ;
        RECT 27.000 -21.950 27.250 -21.600 ;
        RECT 42.000 -21.950 42.250 -21.600 ;
      LAYER met1 ;
        RECT 11.950 -22.500 12.300 -21.500 ;
        RECT 26.950 -22.500 27.300 -21.500 ;
        RECT 41.950 -22.500 42.300 -21.500 ;
      LAYER via ;
        RECT 11.950 -22.450 12.300 -22.000 ;
        RECT 26.950 -22.450 27.300 -22.000 ;
        RECT 41.950 -22.450 42.300 -22.000 ;
      LAYER met2 ;
        RECT 11.950 -22.250 12.300 -21.950 ;
        RECT 26.950 -22.250 27.300 -21.950 ;
        RECT 41.950 -22.250 42.300 -21.950 ;
        RECT 11.950 -22.600 12.850 -22.250 ;
        RECT 26.950 -22.600 27.850 -22.250 ;
        RECT 41.950 -22.600 42.850 -22.250 ;
      LAYER via2 ;
        RECT 12.350 -22.600 12.800 -22.250 ;
        RECT 27.350 -22.600 27.800 -22.250 ;
        RECT 42.350 -22.600 42.800 -22.250 ;
      LAYER met3 ;
        RECT -2.800 -22.250 0.200 -22.150 ;
        RECT 12.300 -22.250 12.850 -22.200 ;
        RECT 27.300 -22.250 27.850 -22.200 ;
        RECT 42.300 -22.250 42.850 -22.200 ;
        RECT -2.800 -22.600 45.000 -22.250 ;
        RECT 12.300 -22.650 12.850 -22.600 ;
        RECT 27.300 -22.650 27.850 -22.600 ;
        RECT 42.300 -22.650 42.850 -22.600 ;
    END
  END ROW_SEL2
  PIN PIX7_IN
    ANTENNAGATEAREA 1.050000 ;
    ANTENNADIFFAREA 0.294000 ;
    PORT
      LAYER li1 ;
        RECT 29.200 -18.050 29.650 -17.680 ;
        RECT 29.350 -19.400 29.650 -18.050 ;
        RECT 28.000 -19.650 29.650 -19.400 ;
        RECT 28.000 -19.950 28.650 -19.650 ;
        RECT 18.200 -27.550 18.900 -26.900 ;
        RECT 17.450 -27.850 18.900 -27.550 ;
      LAYER mcon ;
        RECT 28.050 -19.900 28.600 -19.450 ;
        RECT 18.300 -27.500 18.800 -26.950 ;
      LAYER met1 ;
        RECT 26.300 -19.950 28.700 -19.400 ;
        RECT 18.200 -27.600 18.900 -26.250 ;
      LAYER via ;
        RECT 26.350 -19.950 27.350 -19.400 ;
        RECT 18.250 -26.850 18.850 -26.350 ;
      LAYER met2 ;
        RECT 25.350 -20.050 27.450 -18.700 ;
        RECT 18.200 -26.900 19.650 -26.250 ;
      LAYER via2 ;
        RECT 25.400 -20.000 26.150 -18.800 ;
        RECT 18.250 -26.700 19.600 -26.350 ;
      LAYER met3 ;
        RECT 25.250 -20.150 27.500 -18.600 ;
        RECT 18.200 -26.750 19.650 -24.900 ;
      LAYER via3 ;
        RECT 25.350 -20.050 26.150 -18.700 ;
        RECT 18.400 -25.650 19.500 -25.100 ;
        RECT 18.350 -26.250 19.500 -25.650 ;
        RECT 18.400 -26.650 19.500 -26.250 ;
      LAYER met4 ;
        RECT 23.300 -20.350 27.100 -18.050 ;
        RECT 18.200 -26.750 19.650 -24.900 ;
      LAYER via4 ;
        RECT 25.050 -20.150 26.250 -18.600 ;
        RECT 18.350 -26.250 19.550 -25.000 ;
      LAYER met5 ;
        RECT 17.400 -27.600 27.600 -17.400 ;
    END
  END PIX7_IN
  PIN PIX_OUT1
    ANTENNADIFFAREA 6.400000 ;
    PORT
      LAYER li1 ;
        RECT 24.750 7.450 26.700 7.800 ;
        RECT 25.950 6.050 26.700 7.450 ;
        RECT 25.950 5.300 28.950 6.050 ;
        RECT 24.750 -7.550 26.700 -7.200 ;
        RECT 25.950 -8.950 26.700 -7.550 ;
        RECT 25.950 -9.700 28.950 -8.950 ;
        RECT 24.750 -22.550 26.700 -22.200 ;
        RECT 25.950 -23.950 26.700 -22.550 ;
        RECT 25.950 -24.700 28.950 -23.950 ;
        RECT 17.700 -31.900 25.700 -31.150 ;
      LAYER mcon ;
        RECT 28.200 5.350 28.850 6.000 ;
        RECT 28.200 -9.650 28.850 -9.000 ;
        RECT 28.200 -24.650 28.850 -24.000 ;
        RECT 17.800 -31.450 25.600 -31.150 ;
      LAYER met1 ;
        RECT 28.100 5.300 28.950 6.050 ;
        RECT 28.100 -9.700 28.950 -8.950 ;
        RECT 28.100 -24.700 28.950 -23.950 ;
        RECT 17.700 -31.500 25.700 -30.650 ;
      LAYER via ;
        RECT 28.150 5.300 28.900 6.050 ;
        RECT 28.150 -9.700 28.900 -8.950 ;
        RECT 28.150 -24.700 28.900 -23.950 ;
        RECT 17.800 -31.000 25.600 -30.650 ;
      LAYER met2 ;
        RECT 28.100 5.250 28.950 6.100 ;
        RECT 28.100 -9.750 28.950 -8.900 ;
        RECT 28.100 -24.750 28.950 -23.900 ;
        RECT 17.700 -31.000 28.900 -30.300 ;
      LAYER via2 ;
        RECT 28.150 5.300 28.900 6.050 ;
        RECT 28.150 -9.700 28.900 -8.950 ;
        RECT 28.150 -24.700 28.900 -23.950 ;
        RECT 17.800 -30.900 28.800 -30.400 ;
      LAYER met3 ;
        RECT 28.100 5.200 28.950 6.150 ;
        RECT 28.100 -9.800 28.950 -8.850 ;
        RECT 28.100 -24.800 28.950 -23.850 ;
        RECT 17.700 -31.000 28.900 -30.300 ;
      LAYER via3 ;
        RECT 28.150 5.300 28.900 6.050 ;
        RECT 28.150 -9.700 28.900 -8.950 ;
        RECT 28.150 -24.700 28.900 -23.950 ;
        RECT 17.800 -30.900 28.800 -30.400 ;
      LAYER met4 ;
        RECT 28.150 6.100 28.900 15.800 ;
        RECT 28.100 5.250 28.950 6.100 ;
        RECT 28.150 -8.900 28.900 5.250 ;
        RECT 28.100 -9.750 28.950 -8.900 ;
        RECT 28.150 -23.900 28.900 -9.750 ;
        RECT 28.100 -24.750 28.950 -23.900 ;
        RECT 28.150 -30.300 28.900 -24.750 ;
        RECT 17.700 -31.000 28.900 -30.300 ;
    END
  END PIX_OUT1
  PIN COL_SEL1
    ANTENNAGATEAREA 16.000000 ;
    PORT
      LAYER li1 ;
        RECT 16.100 -33.550 17.200 -32.450 ;
      LAYER mcon ;
        RECT 16.200 -33.500 17.100 -32.500 ;
      LAYER met1 ;
        RECT 16.100 -33.550 17.200 -32.450 ;
      LAYER via ;
        RECT 16.200 -33.500 17.100 -32.500 ;
      LAYER met2 ;
        RECT 16.100 -33.550 17.200 -32.450 ;
      LAYER via2 ;
        RECT 16.200 -33.500 17.100 -32.500 ;
      LAYER met3 ;
        RECT 16.100 -33.550 17.200 -32.450 ;
      LAYER via3 ;
        RECT 16.200 -33.500 17.100 -32.500 ;
      LAYER met4 ;
        RECT 16.100 -35.500 17.200 -32.450 ;
    END
  END COL_SEL1
  PIN PIX8_IN
    ANTENNAGATEAREA 1.050000 ;
    ANTENNADIFFAREA 0.294000 ;
    PORT
      LAYER li1 ;
        RECT 44.200 -18.050 44.650 -17.680 ;
        RECT 44.350 -19.400 44.650 -18.050 ;
        RECT 43.000 -19.650 44.650 -19.400 ;
        RECT 43.000 -19.950 43.650 -19.650 ;
        RECT 33.200 -27.550 33.900 -26.900 ;
        RECT 32.450 -27.850 33.900 -27.550 ;
      LAYER mcon ;
        RECT 43.050 -19.900 43.600 -19.450 ;
        RECT 33.300 -27.500 33.800 -26.950 ;
      LAYER met1 ;
        RECT 41.300 -19.950 43.700 -19.400 ;
        RECT 33.200 -27.600 33.900 -26.250 ;
      LAYER via ;
        RECT 41.350 -19.950 42.350 -19.400 ;
        RECT 33.250 -26.850 33.850 -26.350 ;
      LAYER met2 ;
        RECT 40.350 -20.050 42.450 -18.700 ;
        RECT 33.200 -26.900 34.650 -26.250 ;
      LAYER via2 ;
        RECT 40.400 -20.000 41.150 -18.800 ;
        RECT 33.250 -26.700 34.600 -26.350 ;
      LAYER met3 ;
        RECT 40.250 -20.150 42.500 -18.600 ;
        RECT 33.200 -26.750 34.650 -24.900 ;
      LAYER via3 ;
        RECT 40.350 -20.050 41.150 -18.700 ;
        RECT 33.400 -25.650 34.500 -25.100 ;
        RECT 33.350 -26.250 34.500 -25.650 ;
        RECT 33.400 -26.650 34.500 -26.250 ;
      LAYER met4 ;
        RECT 38.300 -20.350 42.100 -18.050 ;
        RECT 33.200 -26.750 34.650 -24.900 ;
      LAYER via4 ;
        RECT 40.050 -20.150 41.250 -18.600 ;
        RECT 33.350 -26.250 34.550 -25.000 ;
      LAYER met5 ;
        RECT 32.400 -27.600 42.600 -17.400 ;
    END
  END PIX8_IN
  PIN PIX_OUT2
    ANTENNADIFFAREA 6.400000 ;
    PORT
      LAYER li1 ;
        RECT 39.750 7.450 41.700 7.800 ;
        RECT 40.950 6.050 41.700 7.450 ;
        RECT 40.950 5.300 43.950 6.050 ;
        RECT 39.750 -7.550 41.700 -7.200 ;
        RECT 40.950 -8.950 41.700 -7.550 ;
        RECT 40.950 -9.700 43.950 -8.950 ;
        RECT 39.750 -22.550 41.700 -22.200 ;
        RECT 40.950 -23.950 41.700 -22.550 ;
        RECT 40.950 -24.700 43.950 -23.950 ;
        RECT 32.700 -31.900 40.700 -31.150 ;
      LAYER mcon ;
        RECT 43.200 5.350 43.850 6.000 ;
        RECT 43.200 -9.650 43.850 -9.000 ;
        RECT 43.200 -24.650 43.850 -24.000 ;
        RECT 32.800 -31.450 40.600 -31.150 ;
      LAYER met1 ;
        RECT 43.100 5.300 43.950 6.050 ;
        RECT 43.100 -9.700 43.950 -8.950 ;
        RECT 43.100 -24.700 43.950 -23.950 ;
        RECT 32.700 -31.500 40.700 -30.650 ;
      LAYER via ;
        RECT 43.150 5.300 43.900 6.050 ;
        RECT 43.150 -9.700 43.900 -8.950 ;
        RECT 43.150 -24.700 43.900 -23.950 ;
        RECT 32.800 -31.000 40.600 -30.650 ;
      LAYER met2 ;
        RECT 43.100 5.250 43.950 6.100 ;
        RECT 43.100 -9.750 43.950 -8.900 ;
        RECT 43.100 -24.750 43.950 -23.900 ;
        RECT 32.700 -31.000 43.900 -30.300 ;
      LAYER via2 ;
        RECT 43.150 5.300 43.900 6.050 ;
        RECT 43.150 -9.700 43.900 -8.950 ;
        RECT 43.150 -24.700 43.900 -23.950 ;
        RECT 32.800 -30.900 43.800 -30.400 ;
      LAYER met3 ;
        RECT 43.100 5.200 43.950 6.150 ;
        RECT 43.100 -9.800 43.950 -8.850 ;
        RECT 43.100 -24.800 43.950 -23.850 ;
        RECT 32.700 -31.000 43.900 -30.300 ;
      LAYER via3 ;
        RECT 43.150 5.300 43.900 6.050 ;
        RECT 43.150 -9.700 43.900 -8.950 ;
        RECT 43.150 -24.700 43.900 -23.950 ;
        RECT 32.800 -30.900 43.800 -30.400 ;
      LAYER met4 ;
        RECT 43.150 6.100 43.900 15.800 ;
        RECT 43.100 5.250 43.950 6.100 ;
        RECT 43.150 -8.900 43.900 5.250 ;
        RECT 43.100 -9.750 43.950 -8.900 ;
        RECT 43.150 -23.900 43.900 -9.750 ;
        RECT 43.100 -24.750 43.950 -23.900 ;
        RECT 43.150 -30.300 43.900 -24.750 ;
        RECT 32.700 -31.000 43.900 -30.300 ;
    END
  END PIX_OUT2
  PIN COL_SEL2
    ANTENNAGATEAREA 16.000000 ;
    PORT
      LAYER li1 ;
        RECT 31.100 -33.550 32.200 -32.450 ;
      LAYER mcon ;
        RECT 31.200 -33.500 32.100 -32.500 ;
      LAYER met1 ;
        RECT 31.100 -33.550 32.200 -32.450 ;
      LAYER via ;
        RECT 31.200 -33.500 32.100 -32.500 ;
      LAYER met2 ;
        RECT 31.100 -33.550 32.200 -32.450 ;
      LAYER via2 ;
        RECT 31.200 -33.500 32.100 -32.500 ;
      LAYER met3 ;
        RECT 31.100 -33.550 32.200 -32.450 ;
      LAYER via3 ;
        RECT 31.200 -33.500 32.100 -32.500 ;
      LAYER met4 ;
        RECT 31.100 -35.500 32.200 -32.450 ;
    END
  END COL_SEL2
  OBS
      LAYER nwell ;
        RECT 0.000 -3.400 45.000 0.000 ;
        RECT 0.000 -18.400 45.000 -15.000 ;
      LAYER li1 ;
        RECT 0.400 13.350 0.650 14.350 ;
        RECT 1.050 13.350 1.400 13.450 ;
        RECT 0.300 13.150 1.400 13.350 ;
        RECT 2.850 13.350 3.050 14.550 ;
        RECT 3.400 13.350 3.750 13.450 ;
        RECT 2.850 13.150 3.750 13.350 ;
        RECT 0.300 11.250 0.500 13.150 ;
        RECT 1.050 13.000 1.400 13.150 ;
        RECT 3.400 13.000 3.750 13.150 ;
        RECT 10.750 12.650 10.950 14.550 ;
        RECT 11.600 12.700 12.100 13.100 ;
        RECT 12.750 12.900 13.050 14.350 ;
        RECT 15.400 13.350 15.650 14.350 ;
        RECT 16.050 13.350 16.400 13.450 ;
        RECT 2.400 12.450 10.950 12.650 ;
        RECT 11.650 12.550 12.050 12.700 ;
        RECT 12.600 12.600 13.050 12.900 ;
        RECT 15.300 13.150 16.400 13.350 ;
        RECT 17.850 13.350 18.050 14.550 ;
        RECT 18.400 13.350 18.750 13.450 ;
        RECT 17.850 13.150 18.750 13.350 ;
        RECT 2.400 12.100 2.600 12.450 ;
        RECT 2.400 11.850 3.850 12.100 ;
        RECT 2.400 11.250 2.600 11.850 ;
        RECT 0.300 10.950 1.300 11.250 ;
        RECT 1.600 10.950 2.600 11.250 ;
        RECT 3.600 10.950 3.850 11.850 ;
        RECT 3.500 10.050 3.850 10.950 ;
        RECT 5.450 11.900 6.050 12.250 ;
        RECT 5.450 11.500 5.800 11.900 ;
        RECT 11.700 11.500 11.900 12.550 ;
        RECT 5.450 11.300 11.900 11.500 ;
        RECT 5.450 9.900 5.800 11.300 ;
        RECT 12.600 10.850 12.800 12.600 ;
        RECT 15.300 11.250 15.500 13.150 ;
        RECT 16.050 13.000 16.400 13.150 ;
        RECT 18.400 13.000 18.750 13.150 ;
        RECT 25.750 12.650 25.950 14.550 ;
        RECT 26.600 12.700 27.100 13.100 ;
        RECT 27.750 12.900 28.050 14.350 ;
        RECT 30.400 13.350 30.650 14.350 ;
        RECT 31.050 13.350 31.400 13.450 ;
        RECT 17.400 12.450 25.950 12.650 ;
        RECT 26.650 12.550 27.050 12.700 ;
        RECT 27.600 12.600 28.050 12.900 ;
        RECT 30.300 13.150 31.400 13.350 ;
        RECT 32.850 13.350 33.050 14.550 ;
        RECT 33.400 13.350 33.750 13.450 ;
        RECT 32.850 13.150 33.750 13.350 ;
        RECT 17.400 12.100 17.600 12.450 ;
        RECT 17.400 11.850 18.850 12.100 ;
        RECT 17.400 11.250 17.600 11.850 ;
        RECT 15.300 10.950 16.300 11.250 ;
        RECT 16.600 10.950 17.600 11.250 ;
        RECT 10.950 10.650 12.800 10.850 ;
        RECT 17.850 10.750 18.100 11.200 ;
        RECT 18.600 10.950 18.850 11.850 ;
        RECT 10.950 10.100 11.200 10.650 ;
        RECT 17.700 10.250 18.100 10.750 ;
        RECT 4.100 9.850 5.800 9.900 ;
        RECT 4.000 9.550 5.800 9.850 ;
        RECT 10.900 9.750 11.250 10.100 ;
        RECT 18.500 10.050 18.850 10.950 ;
        RECT 20.450 11.900 21.050 12.250 ;
        RECT 20.450 11.500 20.800 11.900 ;
        RECT 26.700 11.500 26.900 12.550 ;
        RECT 20.450 11.300 26.900 11.500 ;
        RECT 20.450 9.900 20.800 11.300 ;
        RECT 27.600 10.850 27.800 12.600 ;
        RECT 30.300 11.250 30.500 13.150 ;
        RECT 31.050 13.000 31.400 13.150 ;
        RECT 33.400 13.000 33.750 13.150 ;
        RECT 40.750 12.650 40.950 14.550 ;
        RECT 41.600 12.700 42.100 13.100 ;
        RECT 42.750 12.900 43.050 14.350 ;
        RECT 32.400 12.450 40.950 12.650 ;
        RECT 41.650 12.550 42.050 12.700 ;
        RECT 42.600 12.600 43.050 12.900 ;
        RECT 32.400 12.100 32.600 12.450 ;
        RECT 32.400 11.850 33.850 12.100 ;
        RECT 32.400 11.250 32.600 11.850 ;
        RECT 30.300 10.950 31.300 11.250 ;
        RECT 31.600 10.950 32.600 11.250 ;
        RECT 25.950 10.650 27.800 10.850 ;
        RECT 32.850 10.750 33.100 11.200 ;
        RECT 33.600 10.950 33.850 11.850 ;
        RECT 25.950 10.100 26.200 10.650 ;
        RECT 32.700 10.250 33.100 10.750 ;
        RECT 19.100 9.850 20.800 9.900 ;
        RECT 10.950 9.650 11.200 9.750 ;
        RECT 19.000 9.550 20.800 9.850 ;
        RECT 25.900 9.750 26.250 10.100 ;
        RECT 33.500 10.050 33.850 10.950 ;
        RECT 35.450 11.900 36.050 12.250 ;
        RECT 35.450 11.500 35.800 11.900 ;
        RECT 41.700 11.500 41.900 12.550 ;
        RECT 35.450 11.300 41.900 11.500 ;
        RECT 35.450 9.900 35.800 11.300 ;
        RECT 42.600 10.850 42.800 12.600 ;
        RECT 40.950 10.650 42.800 10.850 ;
        RECT 40.950 10.100 41.200 10.650 ;
        RECT 34.100 9.850 35.800 9.900 ;
        RECT 25.950 9.650 26.200 9.750 ;
        RECT 34.000 9.550 35.800 9.850 ;
        RECT 40.900 9.750 41.250 10.100 ;
        RECT 40.950 9.650 41.200 9.750 ;
        RECT 4.100 9.500 5.800 9.550 ;
        RECT 19.100 9.500 20.800 9.550 ;
        RECT 34.100 9.500 35.800 9.550 ;
        RECT 1.300 2.400 1.600 9.400 ;
        RECT 1.300 1.750 1.550 2.400 ;
        RECT 15.250 2.000 15.700 2.750 ;
        RECT 16.300 2.400 16.600 9.400 ;
        RECT 20.050 8.450 20.650 9.300 ;
        RECT 20.100 8.050 20.650 8.450 ;
        RECT 16.300 1.750 16.550 2.400 ;
        RECT 30.250 2.000 30.700 2.750 ;
        RECT 31.300 2.400 31.600 9.400 ;
        RECT 35.050 8.450 35.650 9.300 ;
        RECT 35.100 8.050 35.650 8.450 ;
        RECT 31.300 1.750 31.550 2.400 ;
        RECT 1.250 0.550 1.550 1.750 ;
        RECT 16.250 0.550 16.550 1.750 ;
        RECT 31.250 0.550 31.550 1.750 ;
        RECT 5.450 -0.450 5.950 -0.150 ;
        RECT 14.250 -0.200 14.450 -0.150 ;
        RECT 14.150 -0.400 14.550 -0.200 ;
        RECT 0.400 -1.650 0.650 -0.650 ;
        RECT 1.050 -1.650 1.400 -1.550 ;
        RECT 0.300 -1.850 1.400 -1.650 ;
        RECT 2.850 -1.650 3.050 -0.450 ;
        RECT 5.100 -1.450 6.300 -0.450 ;
        RECT 3.400 -1.650 3.750 -1.550 ;
        RECT 2.850 -1.850 3.750 -1.650 ;
        RECT 0.300 -3.750 0.500 -1.850 ;
        RECT 1.050 -2.000 1.400 -1.850 ;
        RECT 3.400 -2.000 3.750 -1.850 ;
        RECT 10.750 -2.350 10.950 -0.450 ;
        RECT 2.400 -2.550 10.950 -2.350 ;
        RECT 11.150 -1.600 11.550 -0.600 ;
        RECT 2.400 -2.900 2.600 -2.550 ;
        RECT 11.150 -2.750 11.400 -1.600 ;
        RECT 11.600 -2.300 12.100 -1.900 ;
        RECT 12.750 -2.100 13.050 -0.650 ;
        RECT 14.250 -1.600 14.450 -0.400 ;
        RECT 20.450 -0.450 20.950 -0.150 ;
        RECT 29.250 -0.200 29.450 -0.150 ;
        RECT 29.150 -0.400 29.550 -0.200 ;
        RECT 15.400 -1.650 15.650 -0.650 ;
        RECT 16.050 -1.650 16.400 -1.550 ;
        RECT 15.300 -1.850 16.400 -1.650 ;
        RECT 17.850 -1.650 18.050 -0.450 ;
        RECT 20.100 -1.450 21.300 -0.450 ;
        RECT 18.400 -1.650 18.750 -1.550 ;
        RECT 17.850 -1.850 18.750 -1.650 ;
        RECT 11.650 -2.450 12.050 -2.300 ;
        RECT 12.600 -2.400 13.050 -2.100 ;
        RECT 13.700 -2.200 14.600 -1.950 ;
        RECT 2.400 -3.150 3.850 -2.900 ;
        RECT 2.400 -3.750 2.600 -3.150 ;
        RECT 0.300 -4.050 1.300 -3.750 ;
        RECT 1.600 -4.050 2.600 -3.750 ;
        RECT 3.600 -4.050 3.850 -3.150 ;
        RECT 4.250 -2.950 4.600 -2.750 ;
        RECT 4.250 -3.750 4.450 -2.950 ;
        RECT 5.450 -3.100 6.050 -2.750 ;
        RECT 10.350 -3.100 11.400 -2.750 ;
        RECT 5.450 -3.500 5.800 -3.100 ;
        RECT 11.700 -3.500 11.900 -2.450 ;
        RECT 5.450 -3.700 11.900 -3.500 ;
        RECT 4.100 -4.000 5.000 -3.750 ;
        RECT 3.500 -4.950 3.850 -4.050 ;
        RECT 5.450 -5.100 5.800 -3.700 ;
        RECT 9.800 -4.600 10.150 -4.050 ;
        RECT 12.600 -4.150 12.800 -2.400 ;
        RECT 13.600 -3.650 14.050 -3.350 ;
        RECT 13.150 -3.900 14.100 -3.650 ;
        RECT 15.300 -3.750 15.500 -1.850 ;
        RECT 16.050 -2.000 16.400 -1.850 ;
        RECT 18.400 -2.000 18.750 -1.850 ;
        RECT 25.750 -2.350 25.950 -0.450 ;
        RECT 17.400 -2.550 25.950 -2.350 ;
        RECT 26.150 -1.600 26.550 -0.600 ;
        RECT 17.400 -2.900 17.600 -2.550 ;
        RECT 26.150 -2.750 26.400 -1.600 ;
        RECT 26.600 -2.300 27.100 -1.900 ;
        RECT 27.750 -2.100 28.050 -0.650 ;
        RECT 29.250 -1.600 29.450 -0.400 ;
        RECT 35.450 -0.450 35.950 -0.150 ;
        RECT 44.250 -0.200 44.450 -0.150 ;
        RECT 44.150 -0.400 44.550 -0.200 ;
        RECT 30.400 -1.650 30.650 -0.650 ;
        RECT 31.050 -1.650 31.400 -1.550 ;
        RECT 30.300 -1.850 31.400 -1.650 ;
        RECT 32.850 -1.650 33.050 -0.450 ;
        RECT 35.100 -1.450 36.300 -0.450 ;
        RECT 33.400 -1.650 33.750 -1.550 ;
        RECT 32.850 -1.850 33.750 -1.650 ;
        RECT 26.650 -2.450 27.050 -2.300 ;
        RECT 27.600 -2.400 28.050 -2.100 ;
        RECT 28.700 -2.200 29.600 -1.950 ;
        RECT 17.400 -3.150 18.850 -2.900 ;
        RECT 17.400 -3.750 17.600 -3.150 ;
        RECT 15.300 -4.050 16.300 -3.750 ;
        RECT 16.600 -4.050 17.600 -3.750 ;
        RECT 10.950 -4.350 12.800 -4.150 ;
        RECT 17.850 -4.250 18.100 -3.800 ;
        RECT 18.600 -4.050 18.850 -3.150 ;
        RECT 19.250 -2.950 19.600 -2.750 ;
        RECT 19.250 -3.750 19.450 -2.950 ;
        RECT 20.450 -3.100 21.050 -2.750 ;
        RECT 25.350 -3.100 26.400 -2.750 ;
        RECT 20.450 -3.500 20.800 -3.100 ;
        RECT 26.700 -3.500 26.900 -2.450 ;
        RECT 20.450 -3.700 26.900 -3.500 ;
        RECT 19.100 -4.000 20.000 -3.750 ;
        RECT 9.800 -4.900 10.700 -4.600 ;
        RECT 10.950 -4.900 11.200 -4.350 ;
        RECT 17.700 -4.750 18.100 -4.250 ;
        RECT 4.100 -5.150 5.800 -5.100 ;
        RECT 4.000 -5.450 5.800 -5.150 ;
        RECT 10.900 -5.250 11.250 -4.900 ;
        RECT 18.500 -4.950 18.850 -4.050 ;
        RECT 20.450 -5.100 20.800 -3.700 ;
        RECT 24.800 -4.600 25.150 -4.050 ;
        RECT 27.600 -4.150 27.800 -2.400 ;
        RECT 28.600 -3.650 29.050 -3.350 ;
        RECT 28.150 -3.900 29.100 -3.650 ;
        RECT 30.300 -3.750 30.500 -1.850 ;
        RECT 31.050 -2.000 31.400 -1.850 ;
        RECT 33.400 -2.000 33.750 -1.850 ;
        RECT 40.750 -2.350 40.950 -0.450 ;
        RECT 32.400 -2.550 40.950 -2.350 ;
        RECT 41.150 -1.600 41.550 -0.600 ;
        RECT 32.400 -2.900 32.600 -2.550 ;
        RECT 41.150 -2.750 41.400 -1.600 ;
        RECT 41.600 -2.300 42.100 -1.900 ;
        RECT 42.750 -2.100 43.050 -0.650 ;
        RECT 44.250 -1.600 44.450 -0.400 ;
        RECT 41.650 -2.450 42.050 -2.300 ;
        RECT 42.600 -2.400 43.050 -2.100 ;
        RECT 43.700 -2.200 44.600 -1.950 ;
        RECT 32.400 -3.150 33.850 -2.900 ;
        RECT 32.400 -3.750 32.600 -3.150 ;
        RECT 30.300 -4.050 31.300 -3.750 ;
        RECT 31.600 -4.050 32.600 -3.750 ;
        RECT 25.950 -4.350 27.800 -4.150 ;
        RECT 32.850 -4.250 33.100 -3.800 ;
        RECT 33.600 -4.050 33.850 -3.150 ;
        RECT 34.250 -2.950 34.600 -2.750 ;
        RECT 34.250 -3.750 34.450 -2.950 ;
        RECT 35.450 -3.100 36.050 -2.750 ;
        RECT 40.350 -3.100 41.400 -2.750 ;
        RECT 35.450 -3.500 35.800 -3.100 ;
        RECT 41.700 -3.500 41.900 -2.450 ;
        RECT 35.450 -3.700 41.900 -3.500 ;
        RECT 34.100 -4.000 35.000 -3.750 ;
        RECT 24.800 -4.900 25.700 -4.600 ;
        RECT 25.950 -4.900 26.200 -4.350 ;
        RECT 32.700 -4.750 33.100 -4.250 ;
        RECT 19.100 -5.150 20.800 -5.100 ;
        RECT 10.950 -5.350 11.200 -5.250 ;
        RECT 19.000 -5.450 20.800 -5.150 ;
        RECT 25.900 -5.250 26.250 -4.900 ;
        RECT 33.500 -4.950 33.850 -4.050 ;
        RECT 35.450 -5.100 35.800 -3.700 ;
        RECT 39.800 -4.600 40.150 -4.050 ;
        RECT 42.600 -4.150 42.800 -2.400 ;
        RECT 43.600 -3.650 44.050 -3.350 ;
        RECT 43.150 -3.900 44.100 -3.650 ;
        RECT 40.950 -4.350 42.800 -4.150 ;
        RECT 39.800 -4.900 40.700 -4.600 ;
        RECT 40.950 -4.900 41.200 -4.350 ;
        RECT 34.100 -5.150 35.800 -5.100 ;
        RECT 25.950 -5.350 26.200 -5.250 ;
        RECT 34.000 -5.450 35.800 -5.150 ;
        RECT 40.900 -5.250 41.250 -4.900 ;
        RECT 40.950 -5.350 41.200 -5.250 ;
        RECT 4.100 -5.500 5.800 -5.450 ;
        RECT 19.100 -5.500 20.800 -5.450 ;
        RECT 34.100 -5.500 35.800 -5.450 ;
        RECT 1.300 -12.600 1.600 -5.600 ;
        RECT 4.000 -7.200 4.900 -6.750 ;
        RECT 4.000 -9.400 4.500 -7.200 ;
        RECT 1.300 -13.250 1.550 -12.600 ;
        RECT 15.250 -13.000 15.700 -12.250 ;
        RECT 16.300 -12.600 16.600 -5.600 ;
        RECT 20.050 -6.550 20.650 -5.700 ;
        RECT 19.000 -7.200 19.900 -6.750 ;
        RECT 20.100 -6.950 20.650 -6.550 ;
        RECT 19.000 -9.400 19.500 -7.200 ;
        RECT 16.300 -13.250 16.550 -12.600 ;
        RECT 30.250 -13.000 30.700 -12.250 ;
        RECT 31.300 -12.600 31.600 -5.600 ;
        RECT 35.050 -6.550 35.650 -5.700 ;
        RECT 34.000 -7.200 34.900 -6.750 ;
        RECT 35.100 -6.950 35.650 -6.550 ;
        RECT 34.000 -9.400 34.500 -7.200 ;
        RECT 31.300 -13.250 31.550 -12.600 ;
        RECT 1.250 -14.450 1.550 -13.250 ;
        RECT 2.650 -14.450 3.350 -13.250 ;
        RECT 3.550 -13.850 4.000 -13.550 ;
        RECT 3.550 -14.250 3.900 -13.850 ;
        RECT 16.250 -14.450 16.550 -13.250 ;
        RECT 17.650 -14.450 18.350 -13.250 ;
        RECT 18.550 -13.850 19.000 -13.550 ;
        RECT 18.550 -14.250 18.900 -13.850 ;
        RECT 31.250 -14.450 31.550 -13.250 ;
        RECT 32.650 -14.450 33.350 -13.250 ;
        RECT 33.550 -13.850 34.000 -13.550 ;
        RECT 33.550 -14.250 33.900 -13.850 ;
        RECT 2.900 -14.850 3.150 -14.450 ;
        RECT 17.900 -14.850 18.150 -14.450 ;
        RECT 32.900 -14.850 33.150 -14.450 ;
        RECT 5.450 -15.450 5.950 -15.150 ;
        RECT 14.250 -15.200 14.450 -15.150 ;
        RECT 14.150 -15.400 14.550 -15.200 ;
        RECT 0.400 -16.650 0.650 -15.650 ;
        RECT 1.050 -16.650 1.400 -16.550 ;
        RECT 0.300 -16.850 1.400 -16.650 ;
        RECT 2.850 -16.650 3.050 -15.450 ;
        RECT 5.100 -16.450 6.300 -15.450 ;
        RECT 3.400 -16.650 3.750 -16.550 ;
        RECT 2.850 -16.850 3.750 -16.650 ;
        RECT 0.300 -18.750 0.500 -16.850 ;
        RECT 1.050 -17.000 1.400 -16.850 ;
        RECT 3.400 -17.000 3.750 -16.850 ;
        RECT 10.750 -17.350 10.950 -15.450 ;
        RECT 2.400 -17.550 10.950 -17.350 ;
        RECT 11.150 -16.600 11.550 -15.600 ;
        RECT 2.400 -17.900 2.600 -17.550 ;
        RECT 11.150 -17.750 11.400 -16.600 ;
        RECT 11.600 -17.300 12.100 -16.900 ;
        RECT 12.750 -17.100 13.050 -15.650 ;
        RECT 14.250 -16.600 14.450 -15.400 ;
        RECT 20.450 -15.450 20.950 -15.150 ;
        RECT 29.250 -15.200 29.450 -15.150 ;
        RECT 29.150 -15.400 29.550 -15.200 ;
        RECT 15.400 -16.650 15.650 -15.650 ;
        RECT 16.050 -16.650 16.400 -16.550 ;
        RECT 15.300 -16.850 16.400 -16.650 ;
        RECT 17.850 -16.650 18.050 -15.450 ;
        RECT 20.100 -16.450 21.300 -15.450 ;
        RECT 18.400 -16.650 18.750 -16.550 ;
        RECT 17.850 -16.850 18.750 -16.650 ;
        RECT 11.650 -17.450 12.050 -17.300 ;
        RECT 12.600 -17.400 13.050 -17.100 ;
        RECT 13.700 -17.200 14.600 -16.950 ;
        RECT 2.400 -18.150 3.850 -17.900 ;
        RECT 2.400 -18.750 2.600 -18.150 ;
        RECT 0.300 -19.050 1.300 -18.750 ;
        RECT 1.600 -19.050 2.600 -18.750 ;
        RECT 3.600 -19.050 3.850 -18.150 ;
        RECT 4.250 -17.950 4.600 -17.750 ;
        RECT 4.250 -18.750 4.450 -17.950 ;
        RECT 5.450 -18.100 6.050 -17.750 ;
        RECT 10.350 -18.100 11.400 -17.750 ;
        RECT 5.450 -18.500 5.800 -18.100 ;
        RECT 11.700 -18.500 11.900 -17.450 ;
        RECT 5.450 -18.700 11.900 -18.500 ;
        RECT 4.100 -19.000 5.000 -18.750 ;
        RECT 3.500 -19.950 3.850 -19.050 ;
        RECT 5.450 -20.100 5.800 -18.700 ;
        RECT 9.800 -19.600 10.150 -19.050 ;
        RECT 12.600 -19.150 12.800 -17.400 ;
        RECT 13.600 -18.650 14.050 -18.350 ;
        RECT 13.150 -18.900 14.100 -18.650 ;
        RECT 15.300 -18.750 15.500 -16.850 ;
        RECT 16.050 -17.000 16.400 -16.850 ;
        RECT 18.400 -17.000 18.750 -16.850 ;
        RECT 25.750 -17.350 25.950 -15.450 ;
        RECT 17.400 -17.550 25.950 -17.350 ;
        RECT 26.150 -16.600 26.550 -15.600 ;
        RECT 17.400 -17.900 17.600 -17.550 ;
        RECT 26.150 -17.750 26.400 -16.600 ;
        RECT 26.600 -17.300 27.100 -16.900 ;
        RECT 27.750 -17.100 28.050 -15.650 ;
        RECT 29.250 -16.600 29.450 -15.400 ;
        RECT 35.450 -15.450 35.950 -15.150 ;
        RECT 44.250 -15.200 44.450 -15.150 ;
        RECT 44.150 -15.400 44.550 -15.200 ;
        RECT 30.400 -16.650 30.650 -15.650 ;
        RECT 31.050 -16.650 31.400 -16.550 ;
        RECT 30.300 -16.850 31.400 -16.650 ;
        RECT 32.850 -16.650 33.050 -15.450 ;
        RECT 35.100 -16.450 36.300 -15.450 ;
        RECT 33.400 -16.650 33.750 -16.550 ;
        RECT 32.850 -16.850 33.750 -16.650 ;
        RECT 26.650 -17.450 27.050 -17.300 ;
        RECT 27.600 -17.400 28.050 -17.100 ;
        RECT 28.700 -17.200 29.600 -16.950 ;
        RECT 17.400 -18.150 18.850 -17.900 ;
        RECT 17.400 -18.750 17.600 -18.150 ;
        RECT 15.300 -19.050 16.300 -18.750 ;
        RECT 16.600 -19.050 17.600 -18.750 ;
        RECT 10.950 -19.350 12.800 -19.150 ;
        RECT 17.850 -19.250 18.100 -18.800 ;
        RECT 18.600 -19.050 18.850 -18.150 ;
        RECT 19.250 -17.950 19.600 -17.750 ;
        RECT 19.250 -18.750 19.450 -17.950 ;
        RECT 20.450 -18.100 21.050 -17.750 ;
        RECT 25.350 -18.100 26.400 -17.750 ;
        RECT 20.450 -18.500 20.800 -18.100 ;
        RECT 26.700 -18.500 26.900 -17.450 ;
        RECT 20.450 -18.700 26.900 -18.500 ;
        RECT 19.100 -19.000 20.000 -18.750 ;
        RECT 9.800 -19.900 10.700 -19.600 ;
        RECT 10.950 -19.900 11.200 -19.350 ;
        RECT 17.700 -19.750 18.100 -19.250 ;
        RECT 4.100 -20.150 5.800 -20.100 ;
        RECT 4.000 -20.450 5.800 -20.150 ;
        RECT 10.900 -20.250 11.250 -19.900 ;
        RECT 18.500 -19.950 18.850 -19.050 ;
        RECT 20.450 -20.100 20.800 -18.700 ;
        RECT 24.800 -19.600 25.150 -19.050 ;
        RECT 27.600 -19.150 27.800 -17.400 ;
        RECT 28.600 -18.650 29.050 -18.350 ;
        RECT 28.150 -18.900 29.100 -18.650 ;
        RECT 30.300 -18.750 30.500 -16.850 ;
        RECT 31.050 -17.000 31.400 -16.850 ;
        RECT 33.400 -17.000 33.750 -16.850 ;
        RECT 40.750 -17.350 40.950 -15.450 ;
        RECT 32.400 -17.550 40.950 -17.350 ;
        RECT 41.150 -16.600 41.550 -15.600 ;
        RECT 32.400 -17.900 32.600 -17.550 ;
        RECT 41.150 -17.750 41.400 -16.600 ;
        RECT 41.600 -17.300 42.100 -16.900 ;
        RECT 42.750 -17.100 43.050 -15.650 ;
        RECT 44.250 -16.600 44.450 -15.400 ;
        RECT 41.650 -17.450 42.050 -17.300 ;
        RECT 42.600 -17.400 43.050 -17.100 ;
        RECT 43.700 -17.200 44.600 -16.950 ;
        RECT 32.400 -18.150 33.850 -17.900 ;
        RECT 32.400 -18.750 32.600 -18.150 ;
        RECT 30.300 -19.050 31.300 -18.750 ;
        RECT 31.600 -19.050 32.600 -18.750 ;
        RECT 25.950 -19.350 27.800 -19.150 ;
        RECT 32.850 -19.250 33.100 -18.800 ;
        RECT 33.600 -19.050 33.850 -18.150 ;
        RECT 34.250 -17.950 34.600 -17.750 ;
        RECT 34.250 -18.750 34.450 -17.950 ;
        RECT 35.450 -18.100 36.050 -17.750 ;
        RECT 40.350 -18.100 41.400 -17.750 ;
        RECT 35.450 -18.500 35.800 -18.100 ;
        RECT 41.700 -18.500 41.900 -17.450 ;
        RECT 35.450 -18.700 41.900 -18.500 ;
        RECT 34.100 -19.000 35.000 -18.750 ;
        RECT 24.800 -19.900 25.700 -19.600 ;
        RECT 25.950 -19.900 26.200 -19.350 ;
        RECT 32.700 -19.750 33.100 -19.250 ;
        RECT 19.100 -20.150 20.800 -20.100 ;
        RECT 10.950 -20.350 11.200 -20.250 ;
        RECT 19.000 -20.450 20.800 -20.150 ;
        RECT 25.900 -20.250 26.250 -19.900 ;
        RECT 33.500 -19.950 33.850 -19.050 ;
        RECT 35.450 -20.100 35.800 -18.700 ;
        RECT 39.800 -19.600 40.150 -19.050 ;
        RECT 42.600 -19.150 42.800 -17.400 ;
        RECT 43.600 -18.650 44.050 -18.350 ;
        RECT 43.150 -18.900 44.100 -18.650 ;
        RECT 40.950 -19.350 42.800 -19.150 ;
        RECT 39.800 -19.900 40.700 -19.600 ;
        RECT 40.950 -19.900 41.200 -19.350 ;
        RECT 34.100 -20.150 35.800 -20.100 ;
        RECT 25.950 -20.350 26.200 -20.250 ;
        RECT 34.000 -20.450 35.800 -20.150 ;
        RECT 40.900 -20.250 41.250 -19.900 ;
        RECT 40.950 -20.350 41.200 -20.250 ;
        RECT 4.100 -20.500 5.800 -20.450 ;
        RECT 19.100 -20.500 20.800 -20.450 ;
        RECT 34.100 -20.500 35.800 -20.450 ;
        RECT 1.300 -27.600 1.600 -20.600 ;
        RECT 4.000 -22.200 4.900 -21.750 ;
        RECT 4.000 -24.400 4.500 -22.200 ;
        RECT 1.300 -28.250 1.550 -27.600 ;
        RECT 15.250 -28.000 15.700 -27.250 ;
        RECT 16.300 -27.600 16.600 -20.600 ;
        RECT 20.050 -21.550 20.650 -20.700 ;
        RECT 19.000 -22.200 19.900 -21.750 ;
        RECT 20.100 -21.950 20.650 -21.550 ;
        RECT 19.000 -24.400 19.500 -22.200 ;
        RECT 16.300 -28.250 16.550 -27.600 ;
        RECT 30.250 -28.000 30.700 -27.250 ;
        RECT 31.300 -27.600 31.600 -20.600 ;
        RECT 35.050 -21.550 35.650 -20.700 ;
        RECT 34.000 -22.200 34.900 -21.750 ;
        RECT 35.100 -21.950 35.650 -21.550 ;
        RECT 34.000 -24.400 34.500 -22.200 ;
        RECT 31.300 -28.250 31.550 -27.600 ;
        RECT 1.250 -29.450 1.550 -28.250 ;
        RECT 2.650 -29.450 3.350 -28.250 ;
        RECT 3.550 -28.850 4.000 -28.550 ;
        RECT 3.550 -29.250 3.900 -28.850 ;
        RECT 16.250 -29.450 16.550 -28.250 ;
        RECT 17.650 -29.450 18.350 -28.250 ;
        RECT 18.550 -28.850 19.000 -28.550 ;
        RECT 18.550 -29.250 18.900 -28.850 ;
        RECT 31.250 -29.450 31.550 -28.250 ;
        RECT 32.650 -29.450 33.350 -28.250 ;
        RECT 33.550 -28.850 34.000 -28.550 ;
        RECT 33.550 -29.250 33.900 -28.850 ;
        RECT 2.900 -29.850 3.150 -29.450 ;
        RECT 17.900 -29.850 18.150 -29.450 ;
        RECT 32.900 -29.850 33.150 -29.450 ;
        RECT 2.700 -35.000 10.700 -34.000 ;
        RECT 17.700 -35.000 25.700 -34.000 ;
        RECT 32.700 -35.000 40.700 -34.000 ;
      LAYER mcon ;
        RECT 5.500 10.550 5.750 10.800 ;
        RECT 17.850 10.800 18.100 11.200 ;
        RECT 20.500 10.550 20.750 10.800 ;
        RECT 32.850 10.800 33.100 11.200 ;
        RECT 35.500 10.550 35.750 10.800 ;
        RECT 15.350 2.500 15.600 2.750 ;
        RECT 20.150 8.100 20.600 8.350 ;
        RECT 30.350 2.500 30.600 2.750 ;
        RECT 35.150 8.100 35.600 8.350 ;
        RECT 5.500 -0.450 5.900 -0.200 ;
        RECT 20.500 -0.450 20.900 -0.200 ;
        RECT 14.400 -2.200 14.600 -1.950 ;
        RECT 10.400 -3.050 10.850 -2.750 ;
        RECT 5.500 -4.450 5.750 -4.200 ;
        RECT 9.850 -4.750 10.100 -4.100 ;
        RECT 35.500 -0.450 35.900 -0.200 ;
        RECT 29.400 -2.200 29.600 -1.950 ;
        RECT 17.850 -4.200 18.100 -3.800 ;
        RECT 25.400 -3.050 25.850 -2.750 ;
        RECT 20.500 -4.450 20.750 -4.200 ;
        RECT 24.850 -4.750 25.100 -4.100 ;
        RECT 44.400 -2.200 44.600 -1.950 ;
        RECT 32.850 -4.200 33.100 -3.800 ;
        RECT 40.400 -3.050 40.850 -2.750 ;
        RECT 35.500 -4.450 35.750 -4.200 ;
        RECT 39.850 -4.750 40.100 -4.100 ;
        RECT 4.050 -9.350 4.450 -8.950 ;
        RECT 15.350 -12.500 15.600 -12.250 ;
        RECT 20.150 -6.900 20.600 -6.650 ;
        RECT 19.050 -9.350 19.450 -8.950 ;
        RECT 30.350 -12.500 30.600 -12.250 ;
        RECT 35.150 -6.900 35.600 -6.650 ;
        RECT 34.050 -9.350 34.450 -8.950 ;
        RECT 3.600 -13.800 3.950 -13.600 ;
        RECT 18.600 -13.800 18.950 -13.600 ;
        RECT 33.600 -13.800 33.950 -13.600 ;
        RECT 2.900 -14.800 3.100 -14.600 ;
        RECT 17.900 -14.800 18.100 -14.600 ;
        RECT 32.900 -14.800 33.100 -14.600 ;
        RECT 5.500 -15.450 5.900 -15.200 ;
        RECT 20.500 -15.450 20.900 -15.200 ;
        RECT 14.400 -17.200 14.600 -16.950 ;
        RECT 10.400 -18.050 10.850 -17.750 ;
        RECT 5.500 -19.450 5.750 -19.200 ;
        RECT 9.850 -19.750 10.100 -19.100 ;
        RECT 35.500 -15.450 35.900 -15.200 ;
        RECT 29.400 -17.200 29.600 -16.950 ;
        RECT 17.850 -19.200 18.100 -18.800 ;
        RECT 25.400 -18.050 25.850 -17.750 ;
        RECT 20.500 -19.450 20.750 -19.200 ;
        RECT 24.850 -19.750 25.100 -19.100 ;
        RECT 44.400 -17.200 44.600 -16.950 ;
        RECT 32.850 -19.200 33.100 -18.800 ;
        RECT 40.400 -18.050 40.850 -17.750 ;
        RECT 35.500 -19.450 35.750 -19.200 ;
        RECT 39.850 -19.750 40.100 -19.100 ;
        RECT 4.050 -24.350 4.450 -23.950 ;
        RECT 15.350 -27.500 15.600 -27.250 ;
        RECT 20.150 -21.900 20.600 -21.650 ;
        RECT 19.050 -24.350 19.450 -23.950 ;
        RECT 30.350 -27.500 30.600 -27.250 ;
        RECT 35.150 -21.900 35.600 -21.650 ;
        RECT 34.050 -24.350 34.450 -23.950 ;
        RECT 3.600 -28.800 3.950 -28.600 ;
        RECT 18.600 -28.800 18.950 -28.600 ;
        RECT 33.600 -28.800 33.950 -28.600 ;
        RECT 2.900 -29.800 3.100 -29.600 ;
        RECT 17.900 -29.800 18.100 -29.600 ;
        RECT 32.900 -29.800 33.100 -29.600 ;
        RECT 2.800 -34.900 10.600 -34.600 ;
        RECT 17.800 -34.900 25.600 -34.600 ;
        RECT 32.800 -34.900 40.600 -34.600 ;
      LAYER met1 ;
        RECT 17.400 11.200 18.150 11.550 ;
        RECT 32.400 11.200 33.150 11.550 ;
        RECT 5.450 10.800 5.800 10.900 ;
        RECT 6.400 10.800 6.800 10.900 ;
        RECT 5.450 10.550 6.800 10.800 ;
        RECT 17.800 10.750 18.150 11.200 ;
        RECT 20.450 10.800 20.800 10.900 ;
        RECT 21.400 10.800 21.800 10.900 ;
        RECT 5.450 10.450 5.800 10.550 ;
        RECT 17.850 10.450 18.100 10.750 ;
        RECT 20.450 10.550 21.800 10.800 ;
        RECT 32.800 10.750 33.150 11.200 ;
        RECT 35.450 10.800 35.800 10.900 ;
        RECT 36.400 10.800 36.800 10.900 ;
        RECT 20.450 10.450 20.800 10.550 ;
        RECT 32.850 10.450 33.100 10.750 ;
        RECT 35.450 10.550 36.800 10.800 ;
        RECT 35.450 10.450 35.800 10.550 ;
        RECT 19.950 7.750 20.650 8.450 ;
        RECT 34.950 7.750 35.650 8.450 ;
        RECT 15.250 2.450 15.700 3.200 ;
        RECT 30.250 2.450 30.700 3.200 ;
        RECT -2.800 -0.600 45.000 -0.150 ;
        RECT 0.000 -0.900 45.000 -0.600 ;
        RECT 4.550 -2.650 5.050 -0.900 ;
        RECT 4.150 -3.000 5.050 -2.650 ;
        RECT 5.450 -4.200 5.800 -4.100 ;
        RECT 6.400 -4.200 6.800 -4.100 ;
        RECT 5.450 -4.450 6.800 -4.200 ;
        RECT 5.450 -4.550 5.800 -4.450 ;
        RECT 9.800 -4.850 10.150 -0.900 ;
        RECT 14.300 -2.250 14.950 -1.900 ;
        RECT 19.550 -2.650 20.050 -0.900 ;
        RECT 10.350 -3.100 10.950 -2.650 ;
        RECT 19.150 -3.000 20.050 -2.650 ;
        RECT 3.950 -9.400 6.500 -8.900 ;
        RECT 3.500 -13.850 4.500 -13.550 ;
        RECT 5.950 -14.100 6.500 -9.400 ;
        RECT 10.350 -14.100 10.850 -3.100 ;
        RECT 13.050 -4.000 13.500 -3.500 ;
        RECT 17.400 -3.800 18.150 -3.450 ;
        RECT 17.800 -4.250 18.150 -3.800 ;
        RECT 20.450 -4.200 20.800 -4.100 ;
        RECT 21.400 -4.200 21.800 -4.100 ;
        RECT 17.850 -4.550 18.100 -4.250 ;
        RECT 20.450 -4.450 21.800 -4.200 ;
        RECT 20.450 -4.550 20.800 -4.450 ;
        RECT 24.800 -4.850 25.150 -0.900 ;
        RECT 29.300 -2.250 29.950 -1.900 ;
        RECT 34.550 -2.650 35.050 -0.900 ;
        RECT 25.350 -3.100 25.950 -2.650 ;
        RECT 34.150 -3.000 35.050 -2.650 ;
        RECT 19.950 -7.250 20.650 -6.550 ;
        RECT 18.950 -9.400 21.500 -8.900 ;
        RECT 15.250 -12.550 15.700 -11.800 ;
        RECT 18.500 -13.850 19.500 -13.550 ;
        RECT 20.950 -14.100 21.500 -9.400 ;
        RECT 25.350 -14.100 25.850 -3.100 ;
        RECT 28.050 -4.000 28.500 -3.500 ;
        RECT 32.400 -3.800 33.150 -3.450 ;
        RECT 32.800 -4.250 33.150 -3.800 ;
        RECT 35.450 -4.200 35.800 -4.100 ;
        RECT 36.400 -4.200 36.800 -4.100 ;
        RECT 32.850 -4.550 33.100 -4.250 ;
        RECT 35.450 -4.450 36.800 -4.200 ;
        RECT 35.450 -4.550 35.800 -4.450 ;
        RECT 39.800 -4.850 40.150 -0.900 ;
        RECT 44.300 -2.250 44.950 -1.900 ;
        RECT 40.350 -3.100 40.950 -2.650 ;
        RECT 34.950 -7.250 35.650 -6.550 ;
        RECT 33.950 -9.400 36.500 -8.900 ;
        RECT 30.250 -12.550 30.700 -11.800 ;
        RECT 33.500 -13.850 34.500 -13.550 ;
        RECT 35.950 -14.100 36.500 -9.400 ;
        RECT 40.350 -14.100 40.850 -3.100 ;
        RECT 43.050 -4.000 43.500 -3.500 ;
        RECT 0.000 -14.400 45.000 -14.100 ;
        RECT 0.000 -14.850 47.600 -14.400 ;
        RECT -2.800 -15.600 45.000 -15.150 ;
        RECT 0.000 -15.900 45.000 -15.600 ;
        RECT 4.550 -17.650 5.050 -15.900 ;
        RECT 4.150 -18.000 5.050 -17.650 ;
        RECT 5.450 -19.200 5.800 -19.100 ;
        RECT 6.400 -19.200 6.800 -19.100 ;
        RECT 5.450 -19.450 6.800 -19.200 ;
        RECT 5.450 -19.550 5.800 -19.450 ;
        RECT 9.800 -19.850 10.150 -15.900 ;
        RECT 14.300 -17.250 14.950 -16.900 ;
        RECT 19.550 -17.650 20.050 -15.900 ;
        RECT 10.350 -18.100 10.950 -17.650 ;
        RECT 19.150 -18.000 20.050 -17.650 ;
        RECT 3.950 -24.400 6.500 -23.900 ;
        RECT 3.500 -28.850 4.500 -28.550 ;
        RECT 5.950 -29.100 6.500 -24.400 ;
        RECT 10.350 -29.100 10.850 -18.100 ;
        RECT 13.050 -19.000 13.500 -18.500 ;
        RECT 17.400 -18.800 18.150 -18.450 ;
        RECT 17.800 -19.250 18.150 -18.800 ;
        RECT 20.450 -19.200 20.800 -19.100 ;
        RECT 21.400 -19.200 21.800 -19.100 ;
        RECT 17.850 -19.550 18.100 -19.250 ;
        RECT 20.450 -19.450 21.800 -19.200 ;
        RECT 20.450 -19.550 20.800 -19.450 ;
        RECT 24.800 -19.850 25.150 -15.900 ;
        RECT 29.300 -17.250 29.950 -16.900 ;
        RECT 34.550 -17.650 35.050 -15.900 ;
        RECT 25.350 -18.100 25.950 -17.650 ;
        RECT 34.150 -18.000 35.050 -17.650 ;
        RECT 19.950 -22.250 20.650 -21.550 ;
        RECT 18.950 -24.400 21.500 -23.900 ;
        RECT 15.250 -27.550 15.700 -26.800 ;
        RECT 18.500 -28.850 19.500 -28.550 ;
        RECT 20.950 -29.100 21.500 -24.400 ;
        RECT 25.350 -29.100 25.850 -18.100 ;
        RECT 28.050 -19.000 28.500 -18.500 ;
        RECT 32.400 -18.800 33.150 -18.450 ;
        RECT 32.800 -19.250 33.150 -18.800 ;
        RECT 35.450 -19.200 35.800 -19.100 ;
        RECT 36.400 -19.200 36.800 -19.100 ;
        RECT 32.850 -19.550 33.100 -19.250 ;
        RECT 35.450 -19.450 36.800 -19.200 ;
        RECT 35.450 -19.550 35.800 -19.450 ;
        RECT 39.800 -19.850 40.150 -15.900 ;
        RECT 44.300 -17.250 44.950 -16.900 ;
        RECT 40.350 -18.100 40.950 -17.650 ;
        RECT 34.950 -22.250 35.650 -21.550 ;
        RECT 33.950 -24.400 36.500 -23.900 ;
        RECT 30.250 -27.550 30.700 -26.800 ;
        RECT 33.500 -28.850 34.500 -28.550 ;
        RECT 35.950 -29.100 36.500 -24.400 ;
        RECT 40.350 -29.100 40.850 -18.100 ;
        RECT 43.050 -19.000 43.500 -18.500 ;
        RECT 0.000 -29.400 45.000 -29.100 ;
        RECT 0.000 -29.850 47.600 -29.400 ;
        RECT 2.700 -35.500 47.600 -34.500 ;
      LAYER via ;
        RECT 17.450 11.250 17.800 11.550 ;
        RECT 32.450 11.250 32.800 11.550 ;
        RECT 6.450 10.600 6.750 10.900 ;
        RECT 21.450 10.600 21.750 10.900 ;
        RECT 36.450 10.600 36.750 10.900 ;
        RECT 20.100 7.800 20.500 8.100 ;
        RECT 35.100 7.800 35.500 8.100 ;
        RECT 15.300 2.800 15.650 3.150 ;
        RECT 30.300 2.800 30.650 3.150 ;
        RECT 6.450 -4.400 6.750 -4.100 ;
        RECT 14.600 -2.250 14.900 -1.900 ;
        RECT 4.100 -13.850 4.450 -13.550 ;
        RECT 13.100 -4.000 13.450 -3.500 ;
        RECT 17.450 -3.750 17.800 -3.450 ;
        RECT 21.450 -4.400 21.750 -4.100 ;
        RECT 29.600 -2.250 29.900 -1.900 ;
        RECT 20.100 -7.200 20.500 -6.900 ;
        RECT 15.300 -12.200 15.650 -11.850 ;
        RECT 19.100 -13.850 19.450 -13.550 ;
        RECT 28.100 -4.000 28.450 -3.500 ;
        RECT 32.450 -3.750 32.800 -3.450 ;
        RECT 36.450 -4.400 36.750 -4.100 ;
        RECT 44.600 -2.250 44.900 -1.900 ;
        RECT 35.100 -7.200 35.500 -6.900 ;
        RECT 30.300 -12.200 30.650 -11.850 ;
        RECT 34.100 -13.850 34.450 -13.550 ;
        RECT 43.100 -4.000 43.450 -3.500 ;
        RECT 7.350 -14.800 7.750 -14.450 ;
        RECT 22.350 -14.800 22.750 -14.450 ;
        RECT 37.350 -14.800 37.750 -14.450 ;
        RECT 6.450 -19.400 6.750 -19.100 ;
        RECT 14.600 -17.250 14.900 -16.900 ;
        RECT 4.100 -28.850 4.450 -28.550 ;
        RECT 13.100 -19.000 13.450 -18.500 ;
        RECT 17.450 -18.750 17.800 -18.450 ;
        RECT 21.450 -19.400 21.750 -19.100 ;
        RECT 29.600 -17.250 29.900 -16.900 ;
        RECT 20.100 -22.200 20.500 -21.900 ;
        RECT 15.300 -27.200 15.650 -26.850 ;
        RECT 19.100 -28.850 19.450 -28.550 ;
        RECT 28.100 -19.000 28.450 -18.500 ;
        RECT 32.450 -18.750 32.800 -18.450 ;
        RECT 36.450 -19.400 36.750 -19.100 ;
        RECT 44.600 -17.250 44.900 -16.900 ;
        RECT 35.100 -22.200 35.500 -21.900 ;
        RECT 30.300 -27.200 30.650 -26.850 ;
        RECT 34.100 -28.850 34.450 -28.550 ;
        RECT 43.100 -19.000 43.450 -18.500 ;
        RECT 7.350 -29.800 7.750 -29.450 ;
        RECT 22.350 -29.800 22.750 -29.450 ;
        RECT 37.350 -29.800 37.750 -29.450 ;
        RECT 2.800 -35.400 47.600 -34.600 ;
      LAYER met2 ;
        RECT 6.400 10.500 6.800 11.500 ;
        RECT 6.400 -4.500 6.800 -3.500 ;
        RECT 13.100 -4.050 13.450 -2.250 ;
        RECT 14.600 -2.350 14.900 -0.850 ;
        RECT 4.100 -14.350 4.500 -13.500 ;
        RECT 7.350 -14.850 7.750 -12.900 ;
        RECT 6.400 -19.500 6.800 -18.500 ;
        RECT 13.100 -19.050 13.450 -17.250 ;
        RECT 14.600 -17.350 14.900 -15.850 ;
        RECT 4.100 -29.350 4.500 -28.500 ;
        RECT 7.350 -29.850 7.750 -27.900 ;
        RECT 15.300 -30.000 15.650 18.000 ;
        RECT 17.500 11.550 17.850 18.000 ;
        RECT 20.100 15.000 20.450 18.000 ;
        RECT 17.400 11.200 17.900 11.550 ;
        RECT 17.500 -3.450 17.850 11.200 ;
        RECT 17.400 -3.800 17.900 -3.450 ;
        RECT 17.500 -18.450 17.850 -3.800 ;
        RECT 19.100 -14.350 19.500 -13.500 ;
        RECT 17.400 -18.800 17.900 -18.450 ;
        RECT 17.500 -30.000 17.850 -18.800 ;
        RECT 19.100 -29.350 19.500 -28.500 ;
        RECT 20.100 -30.000 20.500 15.000 ;
        RECT 21.400 10.500 21.800 11.500 ;
        RECT 21.400 -4.500 21.800 -3.500 ;
        RECT 28.100 -4.050 28.450 -2.250 ;
        RECT 29.600 -2.350 29.900 -0.850 ;
        RECT 22.350 -14.850 22.750 -12.900 ;
        RECT 21.400 -19.500 21.800 -18.500 ;
        RECT 28.100 -19.050 28.450 -17.250 ;
        RECT 29.600 -17.350 29.900 -15.850 ;
        RECT 22.350 -29.850 22.750 -27.900 ;
        RECT 30.300 -30.000 30.650 18.000 ;
        RECT 32.500 11.550 32.850 18.000 ;
        RECT 35.100 15.000 35.450 18.000 ;
        RECT 32.400 11.200 32.900 11.550 ;
        RECT 32.500 -3.450 32.850 11.200 ;
        RECT 32.400 -3.800 32.900 -3.450 ;
        RECT 32.500 -18.450 32.850 -3.800 ;
        RECT 34.100 -14.350 34.500 -13.500 ;
        RECT 32.400 -18.800 32.900 -18.450 ;
        RECT 32.500 -30.000 32.850 -18.800 ;
        RECT 34.100 -29.350 34.500 -28.500 ;
        RECT 35.100 -30.000 35.500 15.000 ;
        RECT 36.400 10.500 36.800 11.500 ;
        RECT 36.400 -4.500 36.800 -3.500 ;
        RECT 43.100 -4.050 43.450 -2.250 ;
        RECT 44.600 -2.350 44.900 -0.850 ;
        RECT 37.350 -14.850 37.750 -12.900 ;
        RECT 36.400 -19.500 36.800 -18.500 ;
        RECT 43.100 -19.050 43.450 -17.250 ;
        RECT 44.600 -17.350 44.900 -15.850 ;
        RECT 37.350 -29.850 37.750 -27.900 ;
        RECT 2.700 -35.500 47.600 -34.500 ;
      LAYER via2 ;
        RECT 6.450 11.100 6.800 11.400 ;
        RECT 14.600 -1.200 14.900 -0.900 ;
        RECT 13.100 -2.700 13.450 -2.350 ;
        RECT 6.450 -3.900 6.800 -3.600 ;
        RECT 7.400 -13.400 7.700 -12.950 ;
        RECT 4.150 -14.250 4.450 -13.900 ;
        RECT 14.600 -16.200 14.900 -15.900 ;
        RECT 13.100 -17.700 13.450 -17.350 ;
        RECT 6.450 -18.900 6.800 -18.600 ;
        RECT 7.400 -28.400 7.700 -27.950 ;
        RECT 4.150 -29.250 4.450 -28.900 ;
        RECT 19.150 -14.250 19.450 -13.900 ;
        RECT 19.150 -29.250 19.450 -28.900 ;
        RECT 21.450 11.100 21.800 11.400 ;
        RECT 29.600 -1.200 29.900 -0.900 ;
        RECT 28.100 -2.700 28.450 -2.350 ;
        RECT 21.450 -3.900 21.800 -3.600 ;
        RECT 22.400 -13.400 22.700 -12.950 ;
        RECT 29.600 -16.200 29.900 -15.900 ;
        RECT 28.100 -17.700 28.450 -17.350 ;
        RECT 21.450 -18.900 21.800 -18.600 ;
        RECT 22.400 -28.400 22.700 -27.950 ;
        RECT 34.150 -14.250 34.450 -13.900 ;
        RECT 34.150 -29.250 34.450 -28.900 ;
        RECT 36.450 11.100 36.800 11.400 ;
        RECT 44.600 -1.200 44.900 -0.900 ;
        RECT 43.100 -2.700 43.450 -2.350 ;
        RECT 36.450 -3.900 36.800 -3.600 ;
        RECT 37.400 -13.400 37.700 -12.950 ;
        RECT 44.600 -16.200 44.900 -15.900 ;
        RECT 43.100 -17.700 43.450 -17.350 ;
        RECT 36.450 -18.900 36.800 -18.600 ;
        RECT 37.400 -28.400 37.700 -27.950 ;
      LAYER met3 ;
        RECT 7.550 11.450 9.850 11.600 ;
        RECT 22.550 11.450 24.850 11.600 ;
        RECT 37.550 11.450 39.850 11.600 ;
        RECT 6.400 11.400 9.850 11.450 ;
        RECT 21.400 11.400 24.850 11.450 ;
        RECT 36.400 11.400 39.850 11.450 ;
        RECT 6.350 11.050 9.850 11.400 ;
        RECT 21.350 11.050 24.850 11.400 ;
        RECT 36.350 11.050 39.850 11.400 ;
        RECT 6.400 11.000 9.850 11.050 ;
        RECT 21.400 11.000 24.850 11.050 ;
        RECT 36.400 11.000 39.850 11.050 ;
        RECT 7.550 9.300 9.850 11.000 ;
        RECT 22.550 9.300 24.850 11.000 ;
        RECT 37.550 9.300 39.850 11.000 ;
        RECT -2.800 -0.900 0.200 -0.800 ;
        RECT 14.550 -0.900 14.950 -0.850 ;
        RECT 29.550 -0.900 29.950 -0.850 ;
        RECT 44.550 -0.900 44.950 -0.850 ;
        RECT -2.800 -1.250 45.000 -0.900 ;
        RECT 14.550 -1.300 14.950 -1.250 ;
        RECT 29.550 -1.300 29.950 -1.250 ;
        RECT 44.550 -1.300 44.950 -1.250 ;
        RECT -2.800 -2.350 0.200 -2.250 ;
        RECT 13.050 -2.350 13.500 -2.300 ;
        RECT 28.050 -2.350 28.500 -2.300 ;
        RECT 43.050 -2.350 43.500 -2.300 ;
        RECT -2.800 -2.700 45.800 -2.350 ;
        RECT 13.050 -2.750 13.500 -2.700 ;
        RECT 28.050 -2.750 28.500 -2.700 ;
        RECT 43.050 -2.750 43.500 -2.700 ;
        RECT 7.550 -3.550 9.850 -3.400 ;
        RECT 22.550 -3.550 24.850 -3.400 ;
        RECT 37.550 -3.550 39.850 -3.400 ;
        RECT 6.400 -3.600 9.850 -3.550 ;
        RECT 21.400 -3.600 24.850 -3.550 ;
        RECT 36.400 -3.600 39.850 -3.550 ;
        RECT 6.350 -3.950 9.850 -3.600 ;
        RECT 21.350 -3.950 24.850 -3.600 ;
        RECT 36.350 -3.950 39.850 -3.600 ;
        RECT 6.400 -4.000 9.850 -3.950 ;
        RECT 21.400 -4.000 24.850 -3.950 ;
        RECT 36.400 -4.000 39.850 -3.950 ;
        RECT 7.550 -5.700 9.850 -4.000 ;
        RECT 22.550 -5.700 24.850 -4.000 ;
        RECT 37.550 -5.700 39.850 -4.000 ;
        RECT 7.250 -13.500 8.750 -12.900 ;
        RECT 22.250 -13.500 23.750 -12.900 ;
        RECT 37.250 -13.500 38.750 -12.900 ;
        RECT -2.800 -13.850 0.200 -13.750 ;
        RECT -2.800 -14.200 45.000 -13.850 ;
        RECT 4.100 -14.300 4.500 -14.200 ;
        RECT 19.100 -14.300 19.500 -14.200 ;
        RECT 34.100 -14.300 34.500 -14.200 ;
        RECT -2.800 -15.900 0.200 -15.800 ;
        RECT 14.550 -15.900 14.950 -15.850 ;
        RECT 29.550 -15.900 29.950 -15.850 ;
        RECT 44.550 -15.900 44.950 -15.850 ;
        RECT -2.800 -16.250 45.000 -15.900 ;
        RECT 14.550 -16.300 14.950 -16.250 ;
        RECT 29.550 -16.300 29.950 -16.250 ;
        RECT 44.550 -16.300 44.950 -16.250 ;
        RECT -2.800 -17.350 0.200 -17.250 ;
        RECT 13.050 -17.350 13.500 -17.300 ;
        RECT 28.050 -17.350 28.500 -17.300 ;
        RECT 43.050 -17.350 43.500 -17.300 ;
        RECT -2.800 -17.700 45.800 -17.350 ;
        RECT 13.050 -17.750 13.500 -17.700 ;
        RECT 28.050 -17.750 28.500 -17.700 ;
        RECT 43.050 -17.750 43.500 -17.700 ;
        RECT 7.550 -18.550 9.850 -18.400 ;
        RECT 22.550 -18.550 24.850 -18.400 ;
        RECT 37.550 -18.550 39.850 -18.400 ;
        RECT 6.400 -18.600 9.850 -18.550 ;
        RECT 21.400 -18.600 24.850 -18.550 ;
        RECT 36.400 -18.600 39.850 -18.550 ;
        RECT 6.350 -18.950 9.850 -18.600 ;
        RECT 21.350 -18.950 24.850 -18.600 ;
        RECT 36.350 -18.950 39.850 -18.600 ;
        RECT 6.400 -19.000 9.850 -18.950 ;
        RECT 21.400 -19.000 24.850 -18.950 ;
        RECT 36.400 -19.000 39.850 -18.950 ;
        RECT 7.550 -20.700 9.850 -19.000 ;
        RECT 22.550 -20.700 24.850 -19.000 ;
        RECT 37.550 -20.700 39.850 -19.000 ;
        RECT 7.250 -28.500 8.750 -27.900 ;
        RECT 22.250 -28.500 23.750 -27.900 ;
        RECT 37.250 -28.500 38.750 -27.900 ;
        RECT -2.800 -28.850 0.200 -28.750 ;
        RECT -2.800 -29.200 45.000 -28.850 ;
        RECT 4.100 -29.300 4.500 -29.200 ;
        RECT 19.100 -29.300 19.500 -29.200 ;
        RECT 34.100 -29.300 34.500 -29.200 ;
      LAYER via3 ;
        RECT 8.150 -13.450 8.700 -12.950 ;
        RECT 23.150 -13.450 23.700 -12.950 ;
        RECT 38.150 -13.450 38.700 -12.950 ;
        RECT 8.150 -28.450 8.700 -27.950 ;
        RECT 23.150 -28.450 23.700 -27.950 ;
        RECT 38.150 -28.450 38.700 -27.950 ;
      LAYER met4 ;
        RECT 2.400 -7.750 12.600 -7.100 ;
        RECT 17.400 -7.750 27.600 -7.100 ;
        RECT 32.400 -7.750 42.600 -7.100 ;
        RECT 6.500 -12.450 11.650 -7.750 ;
        RECT 21.500 -12.450 26.650 -7.750 ;
        RECT 36.500 -12.450 41.650 -7.750 ;
        RECT 8.100 -14.850 8.950 -12.450 ;
        RECT 23.100 -14.850 23.950 -12.450 ;
        RECT 38.100 -14.850 38.950 -12.450 ;
        RECT 2.400 -22.750 12.600 -22.100 ;
        RECT 17.400 -22.750 27.600 -22.100 ;
        RECT 32.400 -22.750 42.600 -22.100 ;
        RECT 6.500 -27.450 11.650 -22.750 ;
        RECT 21.500 -27.450 26.650 -22.750 ;
        RECT 36.500 -27.450 41.650 -22.750 ;
        RECT 8.100 -29.850 8.950 -27.450 ;
        RECT 23.100 -29.850 23.950 -27.450 ;
        RECT 38.100 -29.850 38.950 -27.450 ;
      LAYER met5 ;
        RECT -0.800 14.200 45.800 15.800 ;
        RECT -0.800 0.800 0.800 14.200 ;
        RECT 14.200 0.800 15.800 14.200 ;
        RECT 29.200 0.800 30.800 14.200 ;
        RECT 44.200 0.800 45.800 14.200 ;
        RECT -0.800 -0.800 45.800 0.800 ;
        RECT -0.800 -14.200 0.800 -0.800 ;
        RECT 14.200 -14.200 15.800 -0.800 ;
        RECT 29.200 -14.200 30.800 -0.800 ;
        RECT 44.200 -14.200 45.800 -0.800 ;
        RECT -0.800 -15.800 45.800 -14.200 ;
        RECT -0.800 -29.200 0.800 -15.800 ;
        RECT 14.200 -29.200 15.800 -15.800 ;
        RECT 29.200 -29.200 30.800 -15.800 ;
        RECT 44.200 -29.200 45.800 -15.800 ;
        RECT -0.800 -30.800 45.800 -29.200 ;
  END
END /home/damic/CMOS/TopmetalSe/magic/pixel_array
END LIBRARY

