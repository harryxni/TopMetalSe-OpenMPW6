* SPICE3 file created from pixel_array.ext - technology: sky130A

.subckt pixel gring test_net VREF ROW_SEL NB1 VBIAS NB2 AMP_IN SF_IB PIX_OUT CSA_VREF
+ VDD GND
X0 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt ad=2.52844e+13p pd=5.625e+07u as=0p ps=0u w=2e+06u l=2e+06u
X1 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.57e+12p pd=1.23e+07u as=0p ps=0u w=650000u l=650000u
X2 a_4120_n520# VBIAS a_4120_n750# GND sky130_fd_pr__nfet_01v8_lvt ad=3.5e+11p pd=2.7e+06u as=3.99e+12p ps=1.76e+07u w=1e+06u l=800000u
X3 test_net a_4600_n810# GND VDD sky130_fd_pr__pfet_01v8_lvt ad=5e+11p pd=3e+06u as=8.3e+11p ps=5.9e+06u w=1e+06u l=1e+06u
X4 VDD SF_IB test_net VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5 a_5460_10# a_4350_10# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=3.5e+11p pd=2.7e+06u as=0p ps=0u w=1e+06u l=2e+06u
X6 a_3860_n520# VBIAS a_3860_n1150# GND sky130_fd_pr__nfet_01v8_lvt ad=3.5e+11p pd=2.7e+06u as=3.52e+12p ps=1.76e+07u w=1e+06u l=800000u
X7 VDD a_4120_n520# a_4600_n810# GND sky130_fd_pr__nfet_01v8_lvt ad=1.15e+12p pd=8.3e+06u as=5e+11p ps=3e+06u w=1e+06u l=1e+06u
X8 a_4350_10# a_3860_n520# a_3860_n520# VDD sky130_fd_pr__pfet_01v8_lvt ad=3.5e+11p pd=2.7e+06u as=3.5e+11p ps=2.7e+06u w=1e+06u l=2e+06u
X9 a_4120_n750# AMP_IN a_4050_n2590# GND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.22e+12p ps=1.79e+07u w=7e+06u l=150000u
X10 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=3.35e+06u
X11 a_4120_n520# a_3860_n520# a_5460_10# VDD sky130_fd_pr__pfet_01v8_lvt ad=3.5e+11p pd=2.7e+06u as=0p ps=0u w=1e+06u l=2e+06u
X12 GND NB1 a_4050_n2590# GND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.2e+06u l=1e+06u
X13 a_5750_n920# ROW_SEL PIX_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=5.9e+06u as=5.4e+12p ps=9.4e+06u w=2e+06u l=1e+06u
X14 a_4050_n2590# VREF a_3860_n1150# GND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=7e+06u l=150000u
X15 a_4600_n810# NB2 GND GND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1.15e+06u
X16 AMP_IN a_4600_n810# sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X17 VDD a_4350_10# a_4350_10# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X18 VDD test_net a_5750_n920# GND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 AMP_IN CSA_VREF a_4600_n810# VDD sky130_fd_pr__pfet_01v8_lvt ad=2.94e+11p pd=2.24e+06u as=2.73e+11p ps=2.14e+06u w=420000u l=8e+06u
X20 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.6e+06u l=350000u
C0 gring AMP_IN 3.09fF
C1 gring GND 3.59fF
C2 NB1 GND 3.07fF
C3 PIX_OUT GND 2.60fF
C4 AMP_IN GND 5.66fF
C5 VDD GND 8.13fF
.ends

.subckt pixel_array VBIAS VREF NB2 VDD SF_IB CSA_VREF NB1 ROW_SEL0 GND ROW_SEL1 ROW_SEL2
+ PIX0_IN GRING PIX1_IN PIX2_IN PIX3_IN PIX4_IN PIX5_IN PIX6_IN PIX_OUT0 PIX7_IN PIX_OUT1
+ PIX8_IN PIX_OUT2 ARRAY_OUT COL_SEL0 COL_SEl1 COL_SEL2
Xpixel_0 GRING pixel_0/test_net VREF ROW_SEL0 NB1 VBIAS NB2 PIX0_IN SF_IB PIX_OUT0
+ CSA_VREF VDD GND pixel
Xpixel_1 GRING pixel_1/test_net VREF ROW_SEL0 NB1 VBIAS NB2 PIX1_IN SF_IB PIX_OUT1
+ CSA_VREF VDD GND pixel
Xpixel_2 GRING pixel_2/test_net VREF ROW_SEL0 NB1 VBIAS NB2 PIX2_IN SF_IB PIX_OUT2
+ CSA_VREF VDD GND pixel
Xpixel_3 GRING pixel_3/test_net VREF ROW_SEL1 NB1 VBIAS NB2 PIX3_IN SF_IB PIX_OUT0
+ CSA_VREF VDD GND pixel
Xpixel_5 GRING pixel_5/test_net VREF ROW_SEL1 NB1 VBIAS NB2 PIX5_IN SF_IB PIX_OUT2
+ CSA_VREF VDD GND pixel
Xpixel_4 GRING pixel_4/test_net VREF ROW_SEL1 NB1 VBIAS NB2 PIX4_IN SF_IB PIX_OUT1
+ CSA_VREF VDD GND pixel
Xpixel_6 GRING pixel_6/test_net VREF ROW_SEL2 NB1 VBIAS NB2 PIX6_IN SF_IB PIX_OUT0
+ CSA_VREF VDD GND pixel
Xpixel_7 GRING pixel_7/test_net VREF ROW_SEL2 NB1 VBIAS NB2 PIX7_IN SF_IB PIX_OUT1
+ CSA_VREF VDD GND pixel
Xpixel_8 GRING pixel_8/test_net VREF ROW_SEL2 NB1 VBIAS NB2 PIX8_IN SF_IB PIX_OUT2
+ CSA_VREF VDD GND pixel
X0 PIX_OUT2 COL_SEL2 ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=-2.56998e+12p pd=4.52e+07u as=9.6e+12p ps=5.04e+07u w=8e+06u l=2e+06u
X1 PIX_OUT1 COL_SEl1 ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=7.23002e+12p pd=4.52e+07u as=0p ps=0u w=8e+06u l=2e+06u
X2 PIX_OUT0 COL_SEL0 ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=-5.474e+13p pd=4.52e+07u as=0p ps=0u w=8e+06u l=2e+06u
C0 VDD GND 22.79fF
C1 PIX_OUT1 GRING -2.72fF
C2 GND VREF -4.24fF
C3 VDD NB1 2.44fF
C4 SF_IB NB1 4.08fF
C5 PIX_OUT2 GND 3.00fF
C6 VDD SF_IB -6.49fF
C7 GRING GND -8.38fF
C8 PIX_OUT0 GRING -2.16fF
C9 VDD CSA_VREF -7.92fF
C10 VDD GRING -7.03fF
C11 PIX_OUT1 GND 2.63fF
C12 PIX_OUT2 GRING -3.51fF
C13 PIX_OUT0 GND 2.43fF
C14 NB1 GND -10.41fF
C15 ARRAY_OUT 0 8.23fF
C16 GND 0 -73.74fF
C17 PIX8_IN 0 5.01fF
C18 GRING 0 42.58fF
C19 PIX7_IN 0 5.00fF
C20 PIX6_IN 0 5.62fF
C21 CSA_VREF 0 13.14fF
C22 SF_IB 0 -11.22fF
C23 VDD 0 -20.68fF
C24 PIX_OUT1 0 4.15fF
C25 PIX4_IN 0 4.67fF
C26 PIX_OUT2 0 2.37fF
C27 PIX5_IN 0 4.68fF
C28 PIX3_IN 0 5.30fF
C29 PIX2_IN 0 4.91fF
C30 PIX1_IN 0 4.88fF
C31 ROW_SEL0 0 3.23fF
C32 NB2 0 13.98fF
C33 PIX0_IN 0 5.50fF
.ends

