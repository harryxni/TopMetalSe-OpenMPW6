magic
tech sky130A
magscale 1 2
timestamp 1654643737
<< metal3 >>
rect -1941 1552 1941 1600
rect -1941 1488 1857 1552
rect 1921 1488 1941 1552
rect -1941 1472 1941 1488
rect -1941 1408 1857 1472
rect 1921 1408 1941 1472
rect -1941 1392 1941 1408
rect -1941 1328 1857 1392
rect 1921 1328 1941 1392
rect -1941 1312 1941 1328
rect -1941 1248 1857 1312
rect 1921 1248 1941 1312
rect -1941 1232 1941 1248
rect -1941 1168 1857 1232
rect 1921 1168 1941 1232
rect -1941 1152 1941 1168
rect -1941 1088 1857 1152
rect 1921 1088 1941 1152
rect -1941 1072 1941 1088
rect -1941 1008 1857 1072
rect 1921 1008 1941 1072
rect -1941 992 1941 1008
rect -1941 928 1857 992
rect 1921 928 1941 992
rect -1941 912 1941 928
rect -1941 848 1857 912
rect 1921 848 1941 912
rect -1941 832 1941 848
rect -1941 768 1857 832
rect 1921 768 1941 832
rect -1941 752 1941 768
rect -1941 688 1857 752
rect 1921 688 1941 752
rect -1941 672 1941 688
rect -1941 608 1857 672
rect 1921 608 1941 672
rect -1941 592 1941 608
rect -1941 528 1857 592
rect 1921 528 1941 592
rect -1941 512 1941 528
rect -1941 448 1857 512
rect 1921 448 1941 512
rect -1941 432 1941 448
rect -1941 368 1857 432
rect 1921 368 1941 432
rect -1941 352 1941 368
rect -1941 288 1857 352
rect 1921 288 1941 352
rect -1941 272 1941 288
rect -1941 208 1857 272
rect 1921 208 1941 272
rect -1941 192 1941 208
rect -1941 128 1857 192
rect 1921 128 1941 192
rect -1941 112 1941 128
rect -1941 48 1857 112
rect 1921 48 1941 112
rect -1941 32 1941 48
rect -1941 -32 1857 32
rect 1921 -32 1941 32
rect -1941 -48 1941 -32
rect -1941 -112 1857 -48
rect 1921 -112 1941 -48
rect -1941 -128 1941 -112
rect -1941 -192 1857 -128
rect 1921 -192 1941 -128
rect -1941 -208 1941 -192
rect -1941 -272 1857 -208
rect 1921 -272 1941 -208
rect -1941 -288 1941 -272
rect -1941 -352 1857 -288
rect 1921 -352 1941 -288
rect -1941 -368 1941 -352
rect -1941 -432 1857 -368
rect 1921 -432 1941 -368
rect -1941 -448 1941 -432
rect -1941 -512 1857 -448
rect 1921 -512 1941 -448
rect -1941 -528 1941 -512
rect -1941 -592 1857 -528
rect 1921 -592 1941 -528
rect -1941 -608 1941 -592
rect -1941 -672 1857 -608
rect 1921 -672 1941 -608
rect -1941 -688 1941 -672
rect -1941 -752 1857 -688
rect 1921 -752 1941 -688
rect -1941 -768 1941 -752
rect -1941 -832 1857 -768
rect 1921 -832 1941 -768
rect -1941 -848 1941 -832
rect -1941 -912 1857 -848
rect 1921 -912 1941 -848
rect -1941 -928 1941 -912
rect -1941 -992 1857 -928
rect 1921 -992 1941 -928
rect -1941 -1008 1941 -992
rect -1941 -1072 1857 -1008
rect 1921 -1072 1941 -1008
rect -1941 -1088 1941 -1072
rect -1941 -1152 1857 -1088
rect 1921 -1152 1941 -1088
rect -1941 -1168 1941 -1152
rect -1941 -1232 1857 -1168
rect 1921 -1232 1941 -1168
rect -1941 -1248 1941 -1232
rect -1941 -1312 1857 -1248
rect 1921 -1312 1941 -1248
rect -1941 -1328 1941 -1312
rect -1941 -1392 1857 -1328
rect 1921 -1392 1941 -1328
rect -1941 -1408 1941 -1392
rect -1941 -1472 1857 -1408
rect 1921 -1472 1941 -1408
rect -1941 -1488 1941 -1472
rect -1941 -1552 1857 -1488
rect 1921 -1552 1941 -1488
rect -1941 -1600 1941 -1552
<< via3 >>
rect 1857 1488 1921 1552
rect 1857 1408 1921 1472
rect 1857 1328 1921 1392
rect 1857 1248 1921 1312
rect 1857 1168 1921 1232
rect 1857 1088 1921 1152
rect 1857 1008 1921 1072
rect 1857 928 1921 992
rect 1857 848 1921 912
rect 1857 768 1921 832
rect 1857 688 1921 752
rect 1857 608 1921 672
rect 1857 528 1921 592
rect 1857 448 1921 512
rect 1857 368 1921 432
rect 1857 288 1921 352
rect 1857 208 1921 272
rect 1857 128 1921 192
rect 1857 48 1921 112
rect 1857 -32 1921 32
rect 1857 -112 1921 -48
rect 1857 -192 1921 -128
rect 1857 -272 1921 -208
rect 1857 -352 1921 -288
rect 1857 -432 1921 -368
rect 1857 -512 1921 -448
rect 1857 -592 1921 -528
rect 1857 -672 1921 -608
rect 1857 -752 1921 -688
rect 1857 -832 1921 -768
rect 1857 -912 1921 -848
rect 1857 -992 1921 -928
rect 1857 -1072 1921 -1008
rect 1857 -1152 1921 -1088
rect 1857 -1232 1921 -1168
rect 1857 -1312 1921 -1248
rect 1857 -1392 1921 -1328
rect 1857 -1472 1921 -1408
rect 1857 -1552 1921 -1488
<< mimcap >>
rect -1841 1432 1669 1500
rect -1841 -1432 -1798 1432
rect 1626 -1432 1669 1432
rect -1841 -1500 1669 -1432
<< mimcapcontact >>
rect -1798 -1432 1626 1432
<< metal4 >>
rect 1841 1552 1937 1588
rect 1841 1488 1857 1552
rect 1921 1488 1937 1552
rect 1841 1472 1937 1488
rect -1802 1432 1630 1461
rect -1802 -1432 -1798 1432
rect 1626 -1432 1630 1432
rect -1802 -1461 1630 -1432
rect 1841 1408 1857 1472
rect 1921 1408 1937 1472
rect 1841 1392 1937 1408
rect 1841 1328 1857 1392
rect 1921 1328 1937 1392
rect 1841 1312 1937 1328
rect 1841 1248 1857 1312
rect 1921 1248 1937 1312
rect 1841 1232 1937 1248
rect 1841 1168 1857 1232
rect 1921 1168 1937 1232
rect 1841 1152 1937 1168
rect 1841 1088 1857 1152
rect 1921 1088 1937 1152
rect 1841 1072 1937 1088
rect 1841 1008 1857 1072
rect 1921 1008 1937 1072
rect 1841 992 1937 1008
rect 1841 928 1857 992
rect 1921 928 1937 992
rect 1841 912 1937 928
rect 1841 848 1857 912
rect 1921 848 1937 912
rect 1841 832 1937 848
rect 1841 768 1857 832
rect 1921 768 1937 832
rect 1841 752 1937 768
rect 1841 688 1857 752
rect 1921 688 1937 752
rect 1841 672 1937 688
rect 1841 608 1857 672
rect 1921 608 1937 672
rect 1841 592 1937 608
rect 1841 528 1857 592
rect 1921 528 1937 592
rect 1841 512 1937 528
rect 1841 448 1857 512
rect 1921 448 1937 512
rect 1841 432 1937 448
rect 1841 368 1857 432
rect 1921 368 1937 432
rect 1841 352 1937 368
rect 1841 288 1857 352
rect 1921 288 1937 352
rect 1841 272 1937 288
rect 1841 208 1857 272
rect 1921 208 1937 272
rect 1841 192 1937 208
rect 1841 128 1857 192
rect 1921 128 1937 192
rect 1841 112 1937 128
rect 1841 48 1857 112
rect 1921 48 1937 112
rect 1841 32 1937 48
rect 1841 -32 1857 32
rect 1921 -32 1937 32
rect 1841 -48 1937 -32
rect 1841 -112 1857 -48
rect 1921 -112 1937 -48
rect 1841 -128 1937 -112
rect 1841 -192 1857 -128
rect 1921 -192 1937 -128
rect 1841 -208 1937 -192
rect 1841 -272 1857 -208
rect 1921 -272 1937 -208
rect 1841 -288 1937 -272
rect 1841 -352 1857 -288
rect 1921 -352 1937 -288
rect 1841 -368 1937 -352
rect 1841 -432 1857 -368
rect 1921 -432 1937 -368
rect 1841 -448 1937 -432
rect 1841 -512 1857 -448
rect 1921 -512 1937 -448
rect 1841 -528 1937 -512
rect 1841 -592 1857 -528
rect 1921 -592 1937 -528
rect 1841 -608 1937 -592
rect 1841 -672 1857 -608
rect 1921 -672 1937 -608
rect 1841 -688 1937 -672
rect 1841 -752 1857 -688
rect 1921 -752 1937 -688
rect 1841 -768 1937 -752
rect 1841 -832 1857 -768
rect 1921 -832 1937 -768
rect 1841 -848 1937 -832
rect 1841 -912 1857 -848
rect 1921 -912 1937 -848
rect 1841 -928 1937 -912
rect 1841 -992 1857 -928
rect 1921 -992 1937 -928
rect 1841 -1008 1937 -992
rect 1841 -1072 1857 -1008
rect 1921 -1072 1937 -1008
rect 1841 -1088 1937 -1072
rect 1841 -1152 1857 -1088
rect 1921 -1152 1937 -1088
rect 1841 -1168 1937 -1152
rect 1841 -1232 1857 -1168
rect 1921 -1232 1937 -1168
rect 1841 -1248 1937 -1232
rect 1841 -1312 1857 -1248
rect 1921 -1312 1937 -1248
rect 1841 -1328 1937 -1312
rect 1841 -1392 1857 -1328
rect 1921 -1392 1937 -1328
rect 1841 -1408 1937 -1392
rect 1841 -1472 1857 -1408
rect 1921 -1472 1937 -1408
rect 1841 -1488 1937 -1472
rect 1841 -1552 1857 -1488
rect 1921 -1552 1937 -1488
rect 1841 -1588 1937 -1552
<< properties >>
string FIXED_BBOX -1941 -1600 1769 1600
<< end >>
