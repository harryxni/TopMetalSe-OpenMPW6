magic
tech sky130A
magscale 1 2
timestamp 1654742121
<< metal1 >>
rect 302508 324533 302708 324539
rect 302508 320098 302708 324333
rect 108 17947 308 20712
rect 302508 20408 307134 20608
rect -6205 17747 -6199 17947
rect -5999 17747 308 17947
rect 108 15588 308 17747
rect 306934 17175 307134 20408
rect 306934 16969 307134 16975
rect 108 15382 308 15388
<< via1 >>
rect 302508 324333 302708 324533
rect -6199 17747 -5999 17947
rect 306934 16975 307134 17175
rect 108 15388 308 15588
<< metal2 >>
rect 302508 324533 302708 324542
rect 302502 324333 302508 324533
rect 302708 324333 302714 324533
rect 302508 324324 302708 324333
rect -5180 322443 -2033 322533
rect -5132 319402 -2403 319458
rect -5168 316366 -2742 316422
rect -5148 313238 -3102 313294
rect -3535 310258 -3445 310275
rect -5148 310202 -3445 310258
rect -5138 307166 -3932 307222
rect -5158 304038 -4342 304094
rect -4398 302338 -4342 304038
rect -3988 303948 -3932 307166
rect -3535 306948 -3445 310202
rect -3158 309948 -3102 313238
rect -2798 312948 -2742 316366
rect -2459 315930 -2403 319402
rect -2123 318948 -2033 322443
rect -2123 318858 -802 318948
rect -2459 315874 -579 315930
rect -2798 312892 -622 312948
rect -3165 309858 -755 309948
rect -3535 306858 -802 306948
rect -4005 303858 -775 303948
rect -4398 302282 -692 302338
rect -1485 301058 -1005 301065
rect -5128 301002 -1005 301058
rect -1485 300975 -1005 301002
rect -5148 297966 -1542 298022
rect -1635 294948 -1545 297966
rect -1095 297948 -1005 300975
rect -835 300858 -745 302282
rect -1095 297858 -745 297948
rect -5148 294838 -2152 294894
rect -1635 294858 -725 294948
rect -3095 291858 -3005 292055
rect -2208 291918 -2152 294838
rect -2208 291862 -452 291918
rect -5148 291802 -3005 291858
rect -3095 288948 -3005 291802
rect -3095 288858 -785 288948
rect -3915 288730 -3825 288815
rect -5148 288674 -3825 288730
rect -3915 285948 -3825 288674
rect -3915 285858 -765 285948
rect -5138 285638 -4232 285694
rect -4288 284088 -4232 285638
rect -1105 284088 -1015 284105
rect -4288 284032 -962 284088
rect -1105 282948 -1015 284032
rect -1105 282858 -802 282948
rect -2205 282658 -2115 282765
rect -5158 282602 -2115 282658
rect -2205 279948 -2115 282602
rect -2205 279858 -802 279948
rect -5218 279474 -1962 279530
rect -2055 276948 -1965 279474
rect -2055 276858 -785 276948
rect -892 276494 -802 276525
rect -5188 276438 -802 276494
rect -892 273858 -802 276438
rect -3965 273458 -3875 273585
rect -5228 273402 -3875 273458
rect -3965 270948 -3875 273402
rect -3965 270858 -802 270948
rect -5168 270274 -4582 270330
rect -4638 267948 -4582 270274
rect -4638 267882 -802 267948
rect -4615 267858 -802 267882
rect -4285 267294 -4195 267425
rect -5148 267238 -4195 267294
rect -4285 264948 -4195 267238
rect -4285 264858 -802 264948
rect -5148 264110 -1932 264166
rect -1988 261948 -1932 264110
rect -1988 261858 -802 261948
rect -1988 261812 -1932 261858
rect -5178 261074 -1092 261130
rect -1148 258948 -1092 261074
rect -1148 258858 -775 258948
rect -1148 258822 -1092 258858
rect -5218 258038 -1112 258094
rect -1168 255948 -1112 258038
rect -1168 255858 -802 255948
rect -1168 255842 -1112 255858
rect -5168 254910 -1172 254966
rect -1228 252948 -1172 254910
rect -1228 252858 -802 252948
rect -1228 252852 -1172 252858
rect -5208 251874 -1402 251930
rect -1458 249948 -1402 251874
rect -1458 249892 -795 249948
rect -1435 249858 -795 249892
rect -885 248894 -795 249085
rect -5128 248838 -792 248894
rect -885 246858 -795 248838
rect -892 245766 -802 245885
rect -5268 245710 -802 245766
rect -892 243858 -802 245710
rect -5228 242674 -832 242730
rect -888 240852 -832 242674
rect -5158 239638 -812 239694
rect -868 237892 -812 239638
rect -892 236566 -802 236725
rect -5188 236510 -802 236566
rect -892 234858 -802 236510
rect -5168 233474 -892 233530
rect -948 231852 -892 233474
rect -5168 228948 -5112 230402
rect -5168 228892 -785 228948
rect -5155 228858 -785 228892
rect -5138 227310 -612 227366
rect -835 225858 -745 227310
rect -5195 224265 -802 224355
rect -892 222858 -802 224265
rect -5148 221146 -808 221202
rect -864 219882 -808 221146
rect -808 218178 -752 218202
rect -5128 218122 -752 218178
rect -808 216872 -752 218122
rect -5128 215082 -752 215138
rect -808 213858 -752 215082
rect -5135 211915 -802 212005
rect -892 210858 -802 211915
rect -5128 208910 -732 208966
rect -892 207872 -732 208910
rect -892 207858 -765 207872
rect -5168 205782 -802 205838
rect -858 204842 -802 205782
rect -5158 202746 -762 202802
rect -885 201858 -795 202746
rect -5208 199710 -722 199766
rect -778 198852 -722 199710
rect -5145 196582 -1202 196638
rect -1258 195948 -1202 196582
rect -1258 195858 -793 195948
rect -1258 195805 -1202 195858
rect -5145 193552 -4891 193642
rect -4981 192948 -4891 193552
rect -4981 192858 -782 192948
rect -5134 190510 -737 190566
rect -793 189806 -737 190510
rect -5140 186948 -5050 187461
rect -5140 186858 -793 186948
rect -5140 183948 -5050 184425
rect -5140 183858 -578 183948
rect -5185 180948 -5095 181338
rect -5185 180858 -802 180948
rect -5168 177948 -5078 178234
rect -5168 177858 -572 177948
rect -5128 174948 -5072 175202
rect -5128 174858 -691 174948
rect -5128 174790 -5072 174858
rect -5208 171948 -5118 172065
rect -5208 171858 -782 171948
rect -5157 168948 -5067 169080
rect -5157 168858 -802 168948
rect -5145 165948 -5055 166032
rect -5145 165858 -731 165948
rect -5145 162858 -771 162948
rect -3852 159858 -799 159948
rect -5208 159782 -5202 159838
rect -3852 159779 -816 159858
rect -827 156901 -737 156948
rect -5162 156856 -737 156901
rect -5168 156743 -737 156856
rect -883 153678 -793 153948
rect -5134 153588 -793 153678
rect -5242 150585 -5010 150658
rect -892 150585 -802 150948
rect -5242 150568 -802 150585
rect -5100 150495 -802 150568
rect -5123 147429 -5033 147554
rect -883 147429 -793 147948
rect -5123 147339 -793 147429
rect -883 144569 -793 144948
rect -5179 144479 -793 144569
rect -5179 144417 -839 144479
rect -866 141505 -776 141948
rect -5140 141415 -776 141505
rect -5140 141352 -816 141415
rect -861 138338 -771 138948
rect -5179 138248 -771 138338
rect -892 135341 -802 135948
rect -5191 135251 -802 135341
rect -5134 135183 -805 135251
rect -849 132368 -759 132948
rect -5174 132278 -759 132368
rect -5174 132187 -5084 132278
rect -881 129085 -791 129948
rect -5186 128937 -791 129085
rect -853 126085 -763 126948
rect -5198 125938 -763 126085
rect -892 122977 -802 123948
rect -5141 122790 -802 122977
rect -5128 120948 -5072 121158
rect -5141 120858 -763 120948
rect -5128 119854 -5072 120858
rect -5186 117858 -802 117948
rect -5186 116775 -5096 117858
rect -5158 114858 -614 114948
rect -5158 113650 -5068 114858
rect -5192 111858 -768 111948
rect -5192 110633 -5102 111858
rect -5124 108858 -802 108948
rect -5124 107622 -5034 108858
rect -836 104588 -746 105948
rect -5164 104498 -746 104588
rect -5164 104490 -768 104498
rect -892 101548 -802 102948
rect -5175 101458 -802 101548
rect -892 101259 -802 101458
rect -892 98429 -802 99948
rect -5209 98339 -802 98429
rect -892 98077 -802 98339
rect -881 95396 -791 96948
rect -5181 95306 -791 95396
rect -881 95009 -791 95306
rect -870 92316 -780 93948
rect -5232 92226 -780 92316
rect -870 91913 -780 92226
rect -853 89209 -763 90948
rect -5192 89119 -763 89209
rect -853 89016 -763 89119
rect -836 86198 -746 87948
rect -5129 86108 -746 86198
rect -836 85977 -746 86108
rect -796 83153 -706 84948
rect -5221 83063 -706 83153
rect -796 82721 -706 83063
rect -881 80022 -791 81948
rect -5203 79932 -791 80022
rect -881 79527 -791 79932
rect -858 76949 -768 78948
rect -5209 76859 -768 76949
rect -858 76391 -768 76859
rect -5164 73773 -5074 74058
rect -790 73773 -700 75948
rect -5164 73683 -700 73773
rect -790 73477 -700 73683
rect -830 70796 -740 72948
rect -5152 70706 -740 70796
rect -830 70581 -740 70706
rect -5169 67654 -5079 67774
rect -892 67654 -802 69948
rect -5169 67564 -802 67654
rect -892 67370 -802 67564
rect -608 64618 -552 66924
rect -5226 64562 -552 64618
rect -5209 63858 -643 63948
rect -5209 61354 -5119 63858
rect -5243 60858 -700 60948
rect -5243 58378 -5153 60858
rect -5215 57858 -774 57948
rect -5215 55224 -5125 57858
rect -5243 54858 -774 54948
rect -5243 52316 -5153 54858
rect -322 49346 -266 52178
rect -5147 49290 -266 49346
rect -5226 48858 -489 48948
rect -5226 45970 -5136 48858
rect -3541 45858 -802 45948
rect -3541 43182 -3451 45858
rect -5188 43126 -3343 43182
rect -3541 42491 -3451 43126
rect -2360 42948 -2304 43190
rect -2459 42858 -802 42948
rect -2360 40054 -2304 42858
rect -5257 39998 -2304 40054
rect -751 38442 -661 39948
rect -1991 38386 -497 38442
rect -1991 37018 -1935 38386
rect -751 38281 -661 38386
rect -5131 36962 -1935 37018
rect -463 35565 -373 36948
rect -2435 35509 -373 35565
rect -2435 33982 -2379 35509
rect -463 35254 -373 35509
rect -5144 33926 -2379 33982
rect -772 32850 -716 34558
rect -3299 32794 -716 32850
rect -3299 30854 -3243 32794
rect -5175 30798 -3243 30854
rect -720 29741 -630 30948
rect -2905 29685 -584 29741
rect -2905 27818 -2849 29685
rect -720 29385 -584 29685
rect -720 29261 -630 29385
rect -5175 27762 -2849 27818
rect -757 26901 -667 27948
rect -2592 26845 -628 26901
rect -2592 24782 -2536 26845
rect -757 26590 -667 26845
rect -5188 24726 -2536 24782
rect -764 23911 -674 24948
rect -5244 23855 -459 23911
rect -5244 21598 -5188 23855
rect -764 23519 -674 23855
rect -4016 21858 -736 21948
rect -4016 18618 -3926 21858
rect 38313 19214 38563 19226
rect 19851 19189 20101 19202
rect 19851 18979 19874 19189
rect 20084 18979 20101 19189
rect 29084 19062 29304 19071
rect 13790 18930 14040 18950
rect 19851 18944 20101 18979
rect 25909 19007 26226 19029
rect 13650 18925 14040 18930
rect 7470 18887 7720 18911
rect 5317 18785 5567 18810
rect 4518 18780 5567 18785
rect -5180 18510 -3805 18618
rect 4518 18570 5333 18780
rect 5543 18570 5567 18780
rect 7470 18677 7487 18887
rect 7697 18677 7720 18887
rect 7470 18653 7720 18677
rect 10692 18831 10942 18858
rect 4518 18565 5567 18570
rect -5180 18496 -3926 18510
rect 2316 18440 2566 18467
rect 1499 18435 2566 18440
rect 1499 18225 2333 18435
rect 2543 18225 2566 18435
rect 1499 18220 2566 18225
rect -6199 17947 -5999 17956
rect -6199 17738 -5999 17747
rect 1499 16557 1719 18220
rect 2316 18209 2566 18220
rect 4518 16431 4738 18565
rect 5317 18552 5567 18565
rect 7482 16457 7702 18653
rect 10692 18621 10716 18831
rect 10926 18621 10942 18831
rect 10692 18600 10942 18621
rect 13650 18715 13806 18925
rect 14016 18715 14040 18925
rect 13650 18692 14040 18715
rect 16900 18812 17150 18825
rect 10711 16526 10931 18600
rect 13650 16450 13870 18692
rect 16900 18602 16916 18812
rect 17126 18602 17150 18812
rect 16900 18567 17150 18602
rect 16911 16695 17131 18567
rect 16747 16475 17131 16695
rect 19869 16482 20089 18944
rect 25909 18797 25948 19007
rect 26158 18797 26226 19007
rect 29075 18842 29084 19052
rect 29304 18842 29313 19052
rect 35298 19051 35585 19066
rect 32333 18987 32543 18991
rect 32124 18982 32548 18987
rect 25909 18763 26226 18797
rect 22872 18654 23189 18673
rect 22872 18444 22902 18654
rect 23112 18444 23189 18654
rect 22872 18407 23189 18444
rect 22897 16457 23117 18407
rect 25943 16450 26163 18763
rect 29084 16482 29304 18842
rect 32124 18772 32333 18982
rect 32543 18772 32548 18982
rect 35298 18841 35333 19051
rect 35543 18841 35585 19051
rect 38313 19004 38333 19214
rect 38543 19004 38563 19214
rect 56594 19158 56844 19179
rect 38313 18968 38563 19004
rect 47318 19126 47568 19145
rect 35298 18828 35585 18841
rect 32124 18767 32548 18772
rect 32124 18763 32543 18767
rect 32124 16526 32344 18763
rect 35328 17249 35548 18828
rect 35196 17029 35548 17249
rect 35196 16482 35416 17029
rect 38328 16513 38548 18968
rect 44320 18919 44570 18936
rect 41318 18868 41568 18892
rect 41318 18658 41333 18868
rect 41543 18658 41568 18868
rect 44320 18709 44333 18919
rect 44543 18709 44570 18919
rect 47318 18916 47333 19126
rect 47543 18916 47568 19126
rect 53520 19038 53770 19065
rect 47318 18887 47568 18916
rect 50500 19007 50750 19023
rect 44320 18678 44570 18709
rect 41318 18634 41568 18658
rect 41328 16457 41548 18634
rect 44328 16425 44548 18678
rect 47328 17633 47548 18887
rect 50500 18797 50521 19007
rect 50731 18797 50750 19007
rect 53520 18828 53542 19038
rect 53752 18828 53770 19038
rect 56594 18948 56620 19158
rect 56830 18948 56844 19158
rect 174366 19131 174586 19136
rect 75052 19026 75347 19045
rect 108901 19028 109121 19033
rect 68555 18953 68765 18957
rect 56594 18921 56844 18948
rect 68550 18948 69258 18953
rect 53520 18807 53770 18828
rect 50500 18765 50750 18797
rect 47328 17413 47734 17633
rect 47514 16507 47734 17413
rect 50516 16475 50736 18765
rect 53537 17810 53757 18807
rect 53537 17590 53889 17810
rect 53669 16507 53889 17590
rect 56615 16444 56835 18921
rect 59609 18867 59859 18886
rect 65737 18877 66011 18893
rect 59609 18862 60001 18867
rect 59609 18652 59635 18862
rect 59845 18652 60001 18862
rect 59609 18628 60001 18652
rect 59781 16494 60001 18628
rect 62620 18791 62870 18803
rect 62620 18786 62997 18791
rect 62620 18576 62637 18786
rect 62847 18576 62997 18786
rect 65737 18667 65747 18877
rect 65957 18667 66011 18877
rect 68550 18738 68555 18948
rect 68765 18738 69258 18948
rect 75052 18816 75083 19026
rect 75293 18816 75347 19026
rect 96453 18871 96673 18876
rect 90412 18833 90632 18838
rect 75052 18783 75347 18816
rect 68550 18733 69258 18738
rect 68555 18729 68765 18733
rect 65737 18611 66011 18667
rect 62620 18545 62997 18576
rect 62777 16469 62997 18545
rect 65947 16499 66003 18611
rect 69038 16506 69258 18733
rect 71928 18520 72148 18525
rect 71924 18310 71933 18520
rect 72143 18310 72152 18520
rect 71928 17006 72148 18310
rect 71928 16786 72278 17006
rect 72058 16506 72278 16786
rect 75078 16417 75298 18783
rect 81190 18706 81410 18711
rect 81186 18496 81195 18706
rect 81405 18496 81414 18706
rect 90408 18623 90417 18833
rect 90627 18623 90636 18833
rect 93556 18789 93776 18794
rect 78103 18082 78313 18086
rect 78098 18077 78318 18082
rect 78098 17867 78103 18077
rect 78313 17867 78318 18077
rect 78098 17154 78318 17867
rect 78098 16934 78453 17154
rect 78233 16493 78453 16934
rect 81190 16478 81410 18496
rect 87335 18310 87555 18315
rect 87331 18100 87340 18310
rect 87550 18100 87559 18310
rect 84274 17980 84494 17985
rect 84270 17770 84279 17980
rect 84489 17770 84498 17980
rect 84274 16493 84494 17770
rect 87335 16380 87555 18100
rect 90412 16440 90632 18623
rect 93552 18579 93561 18789
rect 93771 18579 93780 18789
rect 96449 18661 96458 18871
rect 96668 18661 96677 18871
rect 108897 18818 108906 19028
rect 109116 18818 109125 19028
rect 157843 18993 158063 18998
rect 114953 18980 115173 18985
rect 111948 18931 112168 18936
rect 105675 18751 105895 18756
rect 102711 18736 102931 18741
rect 93556 16448 93776 18579
rect 96453 17027 96673 18661
rect 102707 18526 102716 18736
rect 102926 18526 102935 18736
rect 105671 18541 105680 18751
rect 105890 18541 105899 18751
rect 99602 18502 99812 18506
rect 99597 18497 99817 18502
rect 99597 18287 99602 18497
rect 99812 18287 99817 18497
rect 96453 16807 96815 17027
rect 96595 16478 96815 16807
rect 99597 16515 99817 18287
rect 102711 16410 102931 18526
rect 105675 16997 105895 18541
rect 105675 16777 106015 16997
rect 105795 16463 106015 16777
rect 108901 16455 109121 18818
rect 111944 18721 111953 18931
rect 112163 18721 112172 18931
rect 114949 18770 114958 18980
rect 115168 18770 115177 18980
rect 117961 18973 118202 18992
rect 111948 16515 112168 18721
rect 114953 16453 115173 18770
rect 117961 18763 117973 18973
rect 118183 18763 118202 18973
rect 127241 18938 127461 18943
rect 117961 18747 118202 18763
rect 121128 18860 121383 18878
rect 117968 17905 118188 18747
rect 121128 18650 121155 18860
rect 121365 18650 121383 18860
rect 124118 18852 124338 18861
rect 124114 18842 124118 18847
rect 121128 18614 121383 18650
rect 124109 18632 124118 18842
rect 124338 18842 124342 18847
rect 124338 18632 124347 18842
rect 127237 18728 127246 18938
rect 127456 18728 127465 18938
rect 133412 18867 133632 18876
rect 133408 18857 133412 18862
rect 130250 18809 130470 18814
rect 117968 17685 118369 17905
rect 118149 16483 118369 17685
rect 121150 16461 121370 18614
rect 124118 16552 124338 18632
rect 127241 16461 127461 18728
rect 130246 18599 130255 18809
rect 130465 18599 130474 18809
rect 133403 18647 133412 18857
rect 133632 18857 133636 18862
rect 133632 18647 133641 18857
rect 154792 18854 155012 18859
rect 145578 18839 145798 18844
rect 148754 18839 148974 18844
rect 142599 18664 142819 18669
rect 130250 16476 130470 18599
rect 133412 16461 133632 18647
rect 139552 18596 139772 18601
rect 139548 18386 139557 18596
rect 139767 18386 139776 18596
rect 142595 18454 142604 18664
rect 142814 18454 142823 18664
rect 145574 18629 145583 18839
rect 145793 18629 145802 18839
rect 148750 18629 148759 18839
rect 148969 18629 148978 18839
rect 151772 18770 151992 18775
rect 136467 18237 136687 18242
rect 136463 18027 136472 18237
rect 136682 18027 136691 18237
rect 136467 16400 136687 18027
rect 139552 16484 139772 18386
rect 142599 16468 142819 18454
rect 145578 16947 145798 18629
rect 145578 16727 145919 16947
rect 145699 16453 145919 16727
rect 148754 16407 148974 18629
rect 151768 18560 151777 18770
rect 151987 18560 151996 18770
rect 154788 18644 154797 18854
rect 155007 18644 155016 18854
rect 157839 18783 157848 18993
rect 158058 18783 158067 18993
rect 174362 18921 174371 19131
rect 174581 18921 174590 19131
rect 305385 19095 305605 19100
rect 290333 18956 290543 18960
rect 290328 18951 293619 18956
rect 229658 18935 229878 18940
rect 151772 16372 151992 18560
rect 154792 17614 155012 18644
rect 154792 17394 155166 17614
rect 154946 16464 155166 17394
rect 157843 17038 158063 18783
rect 160886 18754 161106 18759
rect 160882 18544 160891 18754
rect 161101 18544 161110 18754
rect 160886 17192 161106 18544
rect 173066 18485 173336 18534
rect 163243 18460 163453 18464
rect 163238 18455 164319 18460
rect 163238 18245 163243 18455
rect 163453 18245 164319 18455
rect 163238 18240 164319 18245
rect 163243 18236 163453 18240
rect 164099 17689 164319 18240
rect 173066 18275 173087 18485
rect 173297 18275 173336 18485
rect 173066 18238 173336 18275
rect 165933 18175 166143 18179
rect 165928 18170 167323 18175
rect 165928 17960 165933 18170
rect 166143 17960 167323 18170
rect 165928 17955 167323 17960
rect 165933 17951 166143 17955
rect 164053 17333 164319 17689
rect 157843 16818 158225 17038
rect 160886 16972 161245 17192
rect 158005 16495 158225 16818
rect 161025 16541 161245 16972
rect 164053 16441 164273 17333
rect 167103 16441 167323 17955
rect 173082 17607 173302 18238
rect 168868 17422 169078 17426
rect 168863 17417 170482 17422
rect 168863 17207 168868 17417
rect 169078 17207 170482 17417
rect 173082 17387 173510 17607
rect 168863 17202 170482 17207
rect 168868 17198 169078 17202
rect 170262 16503 170482 17202
rect 173290 16464 173510 17387
rect 174366 17560 174586 18921
rect 176311 18813 176564 18823
rect 176311 18808 179212 18813
rect 176311 18598 176333 18808
rect 176543 18598 179212 18808
rect 229654 18725 229663 18935
rect 229873 18725 229882 18935
rect 290328 18741 290333 18951
rect 290543 18741 293619 18951
rect 305381 18885 305390 19095
rect 305600 18885 305609 19095
rect 290328 18736 293619 18741
rect 290333 18732 290543 18736
rect 176311 18593 179212 18598
rect 176311 18578 176564 18593
rect 174366 17340 176668 17560
rect 176448 16457 176668 17340
rect 178992 17291 179212 18593
rect 215333 18564 215543 18568
rect 215328 18559 219617 18564
rect 206333 18456 206543 18460
rect 206328 18451 208700 18456
rect 206328 18241 206333 18451
rect 206543 18241 208700 18451
rect 215328 18349 215333 18559
rect 215543 18349 219617 18559
rect 227194 18424 227414 18429
rect 215328 18344 219617 18349
rect 215333 18340 215543 18344
rect 206328 18236 208700 18241
rect 206333 18232 206543 18236
rect 185333 18037 185543 18041
rect 185328 18032 188126 18037
rect 182473 17855 182693 17860
rect 182469 17645 182478 17855
rect 182688 17645 182697 17855
rect 185328 17822 185333 18032
rect 185543 17822 188126 18032
rect 200915 17952 201135 17957
rect 196793 17925 197013 17930
rect 185328 17817 188126 17822
rect 185333 17813 185543 17817
rect 178992 17071 179704 17291
rect 179484 16495 179704 17071
rect 182473 16480 182693 17645
rect 184015 17153 184225 17157
rect 184010 17148 185875 17153
rect 184010 16938 184015 17148
rect 184225 16938 185875 17148
rect 184010 16933 185875 16938
rect 184015 16929 184225 16933
rect 185655 16457 185875 16933
rect 187906 16884 188126 17817
rect 196789 17715 196798 17925
rect 197008 17715 197017 17925
rect 200911 17742 200920 17952
rect 201130 17742 201139 17952
rect 206999 17747 207219 17752
rect 188333 17660 188543 17664
rect 188328 17655 191876 17660
rect 188328 17445 188333 17655
rect 188543 17445 191876 17655
rect 188328 17440 191876 17445
rect 188333 17436 188543 17440
rect 187906 16664 188841 16884
rect 188621 16449 188841 16664
rect 191656 16487 191876 17440
rect 193470 17020 193680 17024
rect 196793 17020 197013 17715
rect 193465 17015 195050 17020
rect 193465 16805 193470 17015
rect 193680 16805 195050 17015
rect 193465 16800 195050 16805
rect 196793 16800 198137 17020
rect 193470 16796 193680 16800
rect 194830 16452 195050 16800
rect 197917 16381 198137 16800
rect 200915 16470 201135 17742
rect 206995 17537 207004 17747
rect 207214 17537 207223 17747
rect 202008 16895 202218 16899
rect 202003 16890 204257 16895
rect 202003 16680 202008 16890
rect 202218 16680 204257 16890
rect 202003 16675 204257 16680
rect 202008 16671 202218 16675
rect 204037 16515 204257 16675
rect 206999 16523 207219 17537
rect 208480 17091 208700 18236
rect 213155 18094 213375 18099
rect 213151 17884 213160 18094
rect 213370 17884 213379 18094
rect 208480 16871 210431 17091
rect 210211 16506 210431 16871
rect 213155 16434 213375 17884
rect 213909 17270 214119 17274
rect 213904 17265 216497 17270
rect 213904 17055 213909 17265
rect 214119 17055 216497 17265
rect 213904 17050 216497 17055
rect 213909 17046 214119 17050
rect 216277 16372 216497 17050
rect 219397 16435 219617 18344
rect 227190 18214 227199 18424
rect 227409 18214 227418 18424
rect 221333 17712 221543 17716
rect 221328 17707 225720 17712
rect 221328 17497 221333 17707
rect 221543 17497 225720 17707
rect 221328 17492 225720 17497
rect 221333 17488 221543 17492
rect 220693 17229 220903 17233
rect 220688 17224 222682 17229
rect 220688 17014 220693 17224
rect 220903 17014 222682 17224
rect 220688 17009 222682 17014
rect 220693 17005 220903 17009
rect 222462 16426 222682 17009
rect 225500 16498 225720 17492
rect 227194 17524 227414 18214
rect 227194 17304 228839 17524
rect 228619 16480 228839 17304
rect 229658 17435 229878 18725
rect 254333 18701 254543 18705
rect 254328 18696 257537 18701
rect 233333 18690 233543 18694
rect 233328 18685 237602 18690
rect 233328 18475 233333 18685
rect 233543 18681 237602 18685
rect 233543 18475 237949 18681
rect 242333 18571 242543 18575
rect 242328 18566 245088 18571
rect 241672 18530 241892 18535
rect 233328 18470 237949 18475
rect 233333 18466 233543 18470
rect 237356 18461 237949 18470
rect 234650 18299 235040 18304
rect 234646 18089 234655 18299
rect 234865 18089 235040 18299
rect 234650 18084 235040 18089
rect 229658 17215 231877 17435
rect 231657 16542 231877 17215
rect 234820 16507 235040 18084
rect 237729 17961 237949 18461
rect 241668 18320 241677 18530
rect 241887 18320 241896 18530
rect 242328 18356 242333 18566
rect 242543 18356 245088 18566
rect 253925 18505 254145 18510
rect 242328 18351 245088 18356
rect 242333 18347 242543 18351
rect 240916 18011 241136 18016
rect 237706 17778 237949 17961
rect 240912 17801 240921 18011
rect 241131 17801 241140 18011
rect 237706 16426 237926 17778
rect 240916 16485 241136 17801
rect 241672 17215 241892 18320
rect 241672 16995 244150 17215
rect 243930 16321 244150 16995
rect 244868 16987 245088 18351
rect 253921 18295 253930 18505
rect 254140 18295 254149 18505
rect 254328 18486 254333 18696
rect 254543 18486 257537 18696
rect 279676 18694 279896 18699
rect 269032 18556 269252 18561
rect 254328 18481 257537 18486
rect 254333 18477 254543 18481
rect 249644 17861 249924 17882
rect 249644 17856 253347 17861
rect 249644 17646 249672 17856
rect 249882 17646 253347 17856
rect 249644 17641 253347 17646
rect 249644 17623 249924 17641
rect 248716 17078 248926 17082
rect 248711 17073 250269 17078
rect 244868 16767 247273 16987
rect 248711 16863 248716 17073
rect 248926 16863 250269 17073
rect 248711 16858 250269 16863
rect 248716 16854 248926 16858
rect 247053 16521 247273 16767
rect 250049 16421 250269 16858
rect 253127 16521 253347 17641
rect 253925 17355 254145 18295
rect 257317 17358 257537 18481
rect 269028 18346 269037 18556
rect 269247 18346 269256 18556
rect 279672 18484 279681 18694
rect 279891 18484 279900 18694
rect 261049 18126 261259 18130
rect 261044 18121 265648 18126
rect 261044 17911 261049 18121
rect 261259 17911 265648 18121
rect 265875 17964 266085 17968
rect 261044 17906 265648 17911
rect 261049 17902 261259 17906
rect 259367 17358 259587 17386
rect 253925 17135 256417 17355
rect 257317 17138 259608 17358
rect 260058 17247 260268 17251
rect 260053 17242 262607 17247
rect 256197 16439 256417 17135
rect 259367 16507 259587 17138
rect 260053 17032 260058 17242
rect 260268 17032 262607 17242
rect 260053 17027 262607 17032
rect 260058 17023 260268 17027
rect 262387 16480 262607 17027
rect 265428 16438 265648 17906
rect 265870 17959 267379 17964
rect 265870 17749 265875 17959
rect 266085 17749 267379 17959
rect 265870 17744 267379 17749
rect 265875 17740 266085 17744
rect 267159 17371 267379 17744
rect 267159 17151 268752 17371
rect 267159 17148 267379 17151
rect 268532 16389 268752 17151
rect 269032 17090 269252 18346
rect 269333 18269 269543 18273
rect 269328 18264 274813 18269
rect 269328 18054 269333 18264
rect 269543 18054 274813 18264
rect 278878 18202 279098 18207
rect 269328 18049 274813 18054
rect 269333 18045 269543 18049
rect 269032 16870 271810 17090
rect 271590 16406 271810 16870
rect 274593 16503 274813 18049
rect 278874 17992 278883 18202
rect 279093 17992 279102 18202
rect 277693 17578 277913 17583
rect 277689 17368 277698 17578
rect 277908 17368 277917 17578
rect 277693 16482 277913 17368
rect 278878 17146 279098 17992
rect 279676 17916 279896 18484
rect 292407 18223 292627 18228
rect 284333 18138 284543 18142
rect 284328 18133 287822 18138
rect 284328 17923 284333 18133
rect 284543 17923 287822 18133
rect 292403 18013 292412 18223
rect 292622 18013 292631 18223
rect 284328 17918 287822 17923
rect 279676 17696 284112 17916
rect 284333 17914 284543 17918
rect 278878 16926 280971 17146
rect 280751 16364 280971 16926
rect 283892 16454 284112 17696
rect 286929 17508 287149 17513
rect 286925 17298 286934 17508
rect 287144 17298 287153 17508
rect 286929 16447 287149 17298
rect 287602 16980 287822 17918
rect 287602 16760 290186 16980
rect 289966 16489 290186 16760
rect 292407 16924 292627 18013
rect 293399 17354 293619 18736
rect 299258 17719 299478 17724
rect 299254 17509 299263 17719
rect 299473 17509 299482 17719
rect 293399 17134 296406 17354
rect 292407 16704 293307 16924
rect 293087 16447 293307 16704
rect 296186 16461 296406 17134
rect 299258 16890 299478 17509
rect 300256 17106 300466 17110
rect 299147 16670 299478 16890
rect 300251 17101 302500 17106
rect 300251 16891 300256 17101
rect 300466 16891 302500 17101
rect 300251 16886 302500 16891
rect 300256 16882 300466 16886
rect 299147 16399 299367 16670
rect 302280 16510 302500 16886
rect 305385 16504 305605 18885
rect 306934 17175 307134 17184
rect 306928 16975 306934 17175
rect 307134 16975 307140 17175
rect 306934 16966 307134 16975
rect 108 15588 308 15597
rect 102 15388 108 15588
rect 308 15388 314 15588
rect 108 15379 308 15388
<< via2 >>
rect 302508 324333 302708 324533
rect 19874 18979 20084 19189
rect 5333 18570 5543 18780
rect 7487 18677 7697 18887
rect 2333 18225 2543 18435
rect -6199 17747 -5999 17947
rect 10716 18621 10926 18831
rect 13806 18715 14016 18925
rect 16916 18602 17126 18812
rect 25948 18797 26158 19007
rect 29084 18842 29304 19062
rect 22902 18444 23112 18654
rect 32333 18772 32543 18982
rect 35333 18841 35543 19051
rect 38333 19004 38543 19214
rect 41333 18658 41543 18868
rect 44333 18709 44543 18919
rect 47333 18916 47543 19126
rect 50521 18797 50731 19007
rect 53542 18828 53752 19038
rect 56620 18948 56830 19158
rect 59635 18652 59845 18862
rect 62637 18576 62847 18786
rect 65747 18667 65957 18877
rect 68555 18738 68765 18948
rect 75083 18816 75293 19026
rect 71933 18310 72143 18520
rect 81195 18496 81405 18706
rect 90417 18623 90627 18833
rect 78103 17867 78313 18077
rect 87340 18100 87550 18310
rect 84279 17770 84489 17980
rect 93561 18579 93771 18789
rect 96458 18661 96668 18871
rect 108906 18818 109116 19028
rect 102716 18526 102926 18736
rect 105680 18541 105890 18751
rect 99602 18287 99812 18497
rect 111953 18721 112163 18931
rect 114958 18770 115168 18980
rect 117973 18763 118183 18973
rect 121155 18650 121365 18860
rect 124118 18632 124338 18852
rect 127246 18728 127456 18938
rect 130255 18599 130465 18809
rect 133412 18647 133632 18867
rect 139557 18386 139767 18596
rect 142604 18454 142814 18664
rect 145583 18629 145793 18839
rect 148759 18629 148969 18839
rect 136472 18027 136682 18237
rect 151777 18560 151987 18770
rect 154797 18644 155007 18854
rect 157848 18783 158058 18993
rect 174371 18921 174581 19131
rect 160891 18544 161101 18754
rect 163243 18245 163453 18455
rect 173087 18275 173297 18485
rect 165933 17960 166143 18170
rect 168868 17207 169078 17417
rect 176333 18598 176543 18808
rect 229663 18725 229873 18935
rect 290333 18741 290543 18951
rect 305390 18885 305600 19095
rect 206333 18241 206543 18451
rect 215333 18349 215543 18559
rect 182478 17645 182688 17855
rect 185333 17822 185543 18032
rect 184015 16938 184225 17148
rect 196798 17715 197008 17925
rect 200920 17742 201130 17952
rect 188333 17445 188543 17655
rect 193470 16805 193680 17015
rect 207004 17537 207214 17747
rect 202008 16680 202218 16890
rect 213160 17884 213370 18094
rect 213909 17055 214119 17265
rect 227199 18214 227409 18424
rect 221333 17497 221543 17707
rect 220693 17014 220903 17224
rect 233333 18475 233543 18685
rect 234655 18089 234865 18299
rect 241677 18320 241887 18530
rect 242333 18356 242543 18566
rect 240921 17801 241131 18011
rect 253930 18295 254140 18505
rect 254333 18486 254543 18696
rect 249672 17646 249882 17856
rect 248716 16863 248926 17073
rect 269037 18346 269247 18556
rect 279681 18484 279891 18694
rect 261049 17911 261259 18121
rect 260058 17032 260268 17242
rect 265875 17749 266085 17959
rect 269333 18054 269543 18264
rect 278883 17992 279093 18202
rect 277698 17368 277908 17578
rect 284333 17923 284543 18133
rect 292412 18013 292622 18223
rect 286934 17298 287144 17508
rect 299263 17509 299473 17719
rect 300256 16891 300466 17101
rect 306934 16975 307134 17175
rect 108 15388 308 15588
<< metal3 >>
rect 302503 324538 302713 324544
rect 302503 324333 302508 324338
rect 302708 324333 302713 324338
rect 302503 324328 302713 324333
rect 38328 19218 38548 19219
rect 19870 19194 20088 19199
rect 19869 19193 20089 19194
rect 19869 18975 19870 19193
rect 20088 18975 20089 19193
rect 29079 19062 29309 19067
rect 25944 19012 26162 19017
rect 19869 18974 20089 18975
rect 25943 19011 26163 19012
rect 19870 18969 20088 18974
rect 13802 18930 14020 18935
rect 13801 18929 14021 18930
rect 7482 18891 7702 18892
rect 5329 18785 5547 18790
rect 5328 18784 5548 18785
rect 5328 18566 5329 18784
rect 5547 18566 5548 18784
rect 7477 18673 7483 18891
rect 7701 18673 7707 18891
rect 10712 18836 10930 18841
rect 10711 18835 10931 18836
rect 7482 18672 7702 18673
rect 10711 18617 10712 18835
rect 10930 18617 10931 18835
rect 13801 18711 13802 18929
rect 14020 18711 14021 18929
rect 16912 18817 17130 18822
rect 13801 18710 14021 18711
rect 16911 18816 17131 18817
rect 13802 18705 14020 18710
rect 10711 18616 10931 18617
rect 10712 18611 10930 18616
rect 16911 18598 16912 18816
rect 17130 18598 17131 18816
rect 25943 18793 25944 19011
rect 26162 18793 26163 19011
rect 29079 18842 29084 19062
rect 29304 18842 29309 19062
rect 35328 19055 35548 19056
rect 32329 18987 32547 18992
rect 29079 18837 29309 18842
rect 32328 18986 32548 18987
rect 25943 18792 26163 18793
rect 25944 18787 26162 18792
rect 32328 18768 32329 18986
rect 32547 18768 32548 18986
rect 35323 18837 35329 19055
rect 35547 18837 35553 19055
rect 38323 19000 38329 19218
rect 38547 19000 38553 19218
rect 56616 19163 56834 19168
rect 56615 19162 56835 19163
rect 47328 19130 47548 19131
rect 38328 18999 38548 19000
rect 44328 18923 44548 18924
rect 41328 18872 41548 18873
rect 35328 18836 35548 18837
rect 32328 18767 32548 18768
rect 32329 18762 32547 18767
rect 22898 18659 23116 18664
rect 16911 18597 17131 18598
rect 22897 18658 23117 18659
rect 16912 18592 17130 18597
rect 5328 18565 5548 18566
rect 5329 18560 5547 18565
rect 22897 18440 22898 18658
rect 23116 18440 23117 18658
rect 41323 18654 41329 18872
rect 41547 18654 41553 18872
rect 44323 18705 44329 18923
rect 44547 18705 44553 18923
rect 47323 18912 47329 19130
rect 47547 18912 47553 19130
rect 53538 19043 53756 19048
rect 53537 19042 53757 19043
rect 50517 19012 50735 19017
rect 50516 19011 50736 19012
rect 47328 18911 47548 18912
rect 50516 18793 50517 19011
rect 50735 18793 50736 19011
rect 53537 18824 53538 19042
rect 53756 18824 53757 19042
rect 56615 18944 56616 19162
rect 56834 18944 56835 19162
rect 174366 19135 174586 19136
rect 71929 19061 72147 19066
rect 71928 19060 72148 19061
rect 68328 18952 68770 18953
rect 56615 18943 56835 18944
rect 56616 18938 56834 18943
rect 65743 18882 65961 18887
rect 65742 18881 65962 18882
rect 59631 18867 59849 18872
rect 53537 18823 53757 18824
rect 59630 18866 59850 18867
rect 53538 18818 53756 18823
rect 50516 18792 50736 18793
rect 50517 18787 50735 18792
rect 44328 18704 44548 18705
rect 41328 18653 41548 18654
rect 59630 18648 59631 18866
rect 59849 18648 59850 18866
rect 62633 18791 62851 18796
rect 59630 18647 59850 18648
rect 62632 18790 62852 18791
rect 59631 18642 59849 18647
rect 62632 18572 62633 18790
rect 62851 18572 62852 18790
rect 65742 18663 65743 18881
rect 65961 18663 65962 18881
rect 68323 18734 68329 18952
rect 68547 18948 68770 18952
rect 68547 18738 68555 18948
rect 68765 18738 68770 18948
rect 68547 18734 68770 18738
rect 68328 18733 68770 18734
rect 71928 18842 71929 19060
rect 72147 18842 72148 19060
rect 75079 19031 75297 19036
rect 108902 19033 109120 19038
rect 108901 19032 109121 19033
rect 65742 18662 65962 18663
rect 65743 18657 65961 18662
rect 62632 18571 62852 18572
rect 62633 18566 62851 18571
rect 2328 18439 2548 18440
rect 22897 18439 23117 18440
rect 71928 18520 72148 18842
rect 75078 19030 75298 19031
rect 75078 18812 75079 19030
rect 75297 18812 75298 19030
rect 81190 18905 81410 18906
rect 75078 18811 75298 18812
rect 75079 18806 75297 18811
rect 81185 18687 81191 18905
rect 81409 18687 81415 18905
rect 96453 18875 96673 18876
rect 90412 18837 90632 18838
rect 2323 18221 2329 18439
rect 2547 18221 2553 18439
rect 22898 18434 23116 18439
rect 71928 18310 71933 18520
rect 72143 18310 72148 18520
rect 81190 18496 81195 18687
rect 81405 18496 81410 18687
rect 90407 18619 90413 18837
rect 90631 18619 90637 18837
rect 93556 18793 93776 18794
rect 90412 18618 90632 18619
rect 93551 18575 93557 18793
rect 93775 18575 93781 18793
rect 96448 18657 96454 18875
rect 96672 18657 96678 18875
rect 108901 18814 108902 19032
rect 109120 18814 109121 19032
rect 157844 18998 158062 19003
rect 157843 18997 158063 18998
rect 114954 18985 115172 18990
rect 114953 18984 115173 18985
rect 111949 18936 112167 18941
rect 108901 18813 109121 18814
rect 111948 18935 112168 18936
rect 108902 18808 109120 18813
rect 105675 18755 105895 18756
rect 102712 18741 102930 18746
rect 102711 18740 102931 18741
rect 96453 18656 96673 18657
rect 93556 18574 93776 18575
rect 102711 18522 102712 18740
rect 102930 18522 102931 18740
rect 105670 18537 105676 18755
rect 105894 18537 105900 18755
rect 111948 18717 111949 18935
rect 112167 18717 112168 18935
rect 114953 18766 114954 18984
rect 115172 18766 115173 18984
rect 117969 18978 118187 18983
rect 114953 18765 115173 18766
rect 117968 18977 118188 18978
rect 114954 18760 115172 18765
rect 117968 18759 117969 18977
rect 118187 18759 118188 18977
rect 127242 18943 127460 18948
rect 127241 18942 127461 18943
rect 121151 18865 121369 18870
rect 117968 18758 118188 18759
rect 121150 18864 121370 18865
rect 117969 18753 118187 18758
rect 111948 18716 112168 18717
rect 111949 18711 112167 18716
rect 121150 18646 121151 18864
rect 121369 18646 121370 18864
rect 121150 18645 121370 18646
rect 124113 18852 124343 18857
rect 121151 18640 121369 18645
rect 124113 18632 124118 18852
rect 124338 18632 124343 18852
rect 127241 18724 127242 18942
rect 127460 18724 127461 18942
rect 133407 18867 133637 18872
rect 130251 18814 130469 18819
rect 127241 18723 127461 18724
rect 130250 18813 130470 18814
rect 127242 18718 127460 18723
rect 124113 18627 124343 18632
rect 130250 18595 130251 18813
rect 130469 18595 130470 18813
rect 133407 18647 133412 18867
rect 133632 18647 133637 18867
rect 154793 18859 155011 18864
rect 154792 18858 155012 18859
rect 145579 18844 145797 18849
rect 148755 18844 148973 18849
rect 145578 18843 145798 18844
rect 142600 18669 142818 18674
rect 133407 18642 133637 18647
rect 142599 18668 142819 18669
rect 139553 18601 139771 18606
rect 130250 18594 130470 18595
rect 139552 18600 139772 18601
rect 130251 18589 130469 18594
rect 105675 18536 105895 18537
rect 102711 18521 102931 18522
rect 102712 18516 102930 18521
rect 99598 18502 99816 18507
rect 81190 18491 81410 18496
rect 99597 18501 99817 18502
rect 84275 18404 84493 18409
rect 84274 18403 84494 18404
rect 71928 18305 72148 18310
rect 78099 18307 78317 18312
rect 78098 18306 78318 18307
rect 2328 18220 2548 18221
rect 78098 18088 78099 18306
rect 78317 18088 78318 18306
rect 78098 18077 78318 18088
rect -6204 17947 -5994 17952
rect -6204 17942 -6199 17947
rect -5999 17942 -5994 17947
rect 78098 17867 78103 18077
rect 78313 17867 78318 18077
rect 78098 17862 78318 17867
rect 84274 18185 84275 18403
rect 84493 18185 84494 18403
rect 87336 18315 87554 18320
rect 84274 17980 84494 18185
rect 87335 18314 87555 18315
rect 87335 18096 87336 18314
rect 87554 18096 87555 18314
rect 99597 18283 99598 18501
rect 99816 18283 99817 18501
rect 139552 18382 139553 18600
rect 139771 18382 139772 18600
rect 142599 18450 142600 18668
rect 142818 18450 142819 18668
rect 145578 18625 145579 18843
rect 145797 18625 145798 18843
rect 145578 18624 145798 18625
rect 148754 18843 148974 18844
rect 148754 18625 148755 18843
rect 148973 18625 148974 18843
rect 151773 18775 151991 18780
rect 148754 18624 148974 18625
rect 151772 18774 151992 18775
rect 145579 18619 145797 18624
rect 148755 18619 148973 18624
rect 151772 18556 151773 18774
rect 151991 18556 151992 18774
rect 154792 18640 154793 18858
rect 155011 18640 155012 18858
rect 157843 18779 157844 18997
rect 158062 18779 158063 18997
rect 174361 18917 174367 19135
rect 174585 18917 174591 19135
rect 305386 19100 305604 19105
rect 305385 19099 305605 19100
rect 290329 18956 290547 18961
rect 290328 18955 290548 18956
rect 229658 18939 229878 18940
rect 174366 18916 174586 18917
rect 176328 18812 176548 18813
rect 157843 18778 158063 18779
rect 157844 18773 158062 18778
rect 160886 18758 161106 18759
rect 154792 18639 155012 18640
rect 154793 18634 155011 18639
rect 151772 18555 151992 18556
rect 151773 18550 151991 18555
rect 160881 18540 160887 18758
rect 161105 18540 161111 18758
rect 176323 18594 176329 18812
rect 176547 18594 176553 18812
rect 229653 18721 229659 18939
rect 229877 18721 229883 18939
rect 290328 18737 290329 18955
rect 290547 18737 290548 18955
rect 305385 18881 305386 19099
rect 305604 18881 305605 19099
rect 305385 18880 305605 18881
rect 305386 18875 305604 18880
rect 290328 18736 290548 18737
rect 290329 18731 290547 18736
rect 229658 18720 229878 18721
rect 254329 18701 254547 18706
rect 254328 18700 254548 18701
rect 233329 18690 233547 18695
rect 233328 18689 233548 18690
rect 176328 18593 176548 18594
rect 215329 18564 215547 18569
rect 215328 18563 215548 18564
rect 160886 18539 161106 18540
rect 173083 18490 173301 18495
rect 173082 18489 173302 18490
rect 163238 18459 163458 18460
rect 142599 18449 142819 18450
rect 142600 18444 142818 18449
rect 139552 18381 139772 18382
rect 139553 18376 139771 18381
rect 99597 18282 99817 18283
rect 99598 18277 99816 18282
rect 136467 18241 136687 18242
rect 163233 18241 163239 18459
rect 163457 18241 163463 18459
rect 173082 18271 173083 18489
rect 173301 18271 173302 18489
rect 206329 18456 206547 18461
rect 173082 18270 173302 18271
rect 206328 18455 206548 18456
rect 173083 18265 173301 18270
rect 87335 18095 87555 18096
rect 87336 18090 87554 18095
rect 136462 18023 136468 18241
rect 136686 18023 136692 18241
rect 163238 18240 163458 18241
rect 206328 18237 206329 18455
rect 206547 18237 206548 18455
rect 215328 18345 215329 18563
rect 215547 18345 215548 18563
rect 233328 18471 233329 18689
rect 233547 18471 233548 18689
rect 242329 18571 242547 18576
rect 242328 18570 242548 18571
rect 241673 18535 241891 18540
rect 233328 18470 233548 18471
rect 241672 18534 241892 18535
rect 233329 18465 233547 18470
rect 227194 18428 227414 18429
rect 215328 18344 215548 18345
rect 215329 18339 215547 18344
rect 206328 18236 206548 18237
rect 206329 18231 206547 18236
rect 227189 18210 227195 18428
rect 227413 18210 227419 18428
rect 241672 18316 241673 18534
rect 241891 18316 241892 18534
rect 242328 18352 242329 18570
rect 242547 18352 242548 18570
rect 253925 18509 254145 18510
rect 242328 18351 242548 18352
rect 242329 18346 242547 18351
rect 241672 18315 241892 18316
rect 241673 18310 241891 18315
rect 234650 18303 234870 18304
rect 227194 18209 227414 18210
rect 165929 18175 166147 18180
rect 165928 18174 166148 18175
rect 136467 18022 136687 18023
rect 84274 17770 84279 17980
rect 84489 17770 84494 17980
rect 165928 17956 165929 18174
rect 166147 17956 166148 18174
rect 213156 18099 213374 18104
rect 213155 18098 213375 18099
rect 185329 18037 185547 18042
rect 165928 17955 166148 17956
rect 185328 18036 185548 18037
rect 165929 17950 166147 17955
rect 182473 17859 182693 17860
rect 84274 17765 84494 17770
rect -6204 17736 -5994 17742
rect 182468 17641 182474 17859
rect 182692 17641 182698 17859
rect 185328 17818 185329 18036
rect 185547 17818 185548 18036
rect 200916 17957 201134 17962
rect 200915 17956 201135 17957
rect 196793 17929 197013 17930
rect 185328 17817 185548 17818
rect 185329 17812 185547 17817
rect 196788 17711 196794 17929
rect 197012 17711 197018 17929
rect 200915 17738 200916 17956
rect 201134 17738 201135 17956
rect 213155 17880 213156 18098
rect 213374 17880 213375 18098
rect 234645 18085 234651 18303
rect 234869 18085 234875 18303
rect 253920 18291 253926 18509
rect 254144 18291 254150 18509
rect 254328 18482 254329 18700
rect 254547 18482 254548 18700
rect 279676 18698 279896 18699
rect 269032 18560 269252 18561
rect 254328 18481 254548 18482
rect 254329 18476 254547 18481
rect 269027 18342 269033 18560
rect 269251 18342 269257 18560
rect 279671 18480 279677 18698
rect 279895 18480 279901 18698
rect 279676 18479 279896 18480
rect 269032 18341 269252 18342
rect 253925 18290 254145 18291
rect 269329 18269 269547 18274
rect 269328 18268 269548 18269
rect 261045 18126 261263 18131
rect 261044 18125 261264 18126
rect 234650 18084 234870 18085
rect 240917 18016 241135 18021
rect 213155 17879 213375 17880
rect 240916 18015 241136 18016
rect 213156 17874 213374 17879
rect 240916 17797 240917 18015
rect 241135 17797 241136 18015
rect 261044 17907 261045 18125
rect 261263 17907 261264 18125
rect 269328 18050 269329 18268
rect 269547 18050 269548 18268
rect 292407 18227 292627 18228
rect 278878 18206 279098 18207
rect 269328 18049 269548 18050
rect 269329 18044 269547 18049
rect 278873 17988 278879 18206
rect 279097 17988 279103 18206
rect 284329 18138 284547 18143
rect 284328 18137 284548 18138
rect 278878 17987 279098 17988
rect 265871 17964 266089 17969
rect 261044 17906 261264 17907
rect 265870 17963 266090 17964
rect 261045 17901 261263 17906
rect 249667 17860 249887 17861
rect 240916 17796 241136 17797
rect 240917 17791 241135 17796
rect 207000 17752 207218 17757
rect 200915 17737 201135 17738
rect 206999 17751 207219 17752
rect 200916 17732 201134 17737
rect 196793 17710 197013 17711
rect 188329 17660 188547 17665
rect 188328 17659 188548 17660
rect 182473 17640 182693 17641
rect 188328 17441 188329 17659
rect 188547 17441 188548 17659
rect 206999 17533 207000 17751
rect 207218 17533 207219 17751
rect 221329 17712 221547 17717
rect 206999 17532 207219 17533
rect 221328 17711 221548 17712
rect 207000 17527 207218 17532
rect 221328 17493 221329 17711
rect 221547 17493 221548 17711
rect 249662 17642 249668 17860
rect 249886 17642 249892 17860
rect 265870 17745 265871 17963
rect 266089 17745 266090 17963
rect 284328 17919 284329 18137
rect 284547 17919 284548 18137
rect 292402 18009 292408 18227
rect 292626 18009 292632 18227
rect 292407 18008 292627 18009
rect 284328 17918 284548 17919
rect 284329 17913 284547 17918
rect 265870 17744 266090 17745
rect 265871 17739 266089 17744
rect 299259 17724 299477 17729
rect 299258 17723 299478 17724
rect 249667 17641 249887 17642
rect 277693 17582 277913 17583
rect 221328 17492 221548 17493
rect 221329 17487 221547 17492
rect 188328 17440 188548 17441
rect 188329 17435 188547 17440
rect 168864 17422 169082 17427
rect 168863 17421 169083 17422
rect 168863 17203 168864 17421
rect 169082 17203 169083 17421
rect 277688 17364 277694 17582
rect 277912 17364 277918 17582
rect 286930 17513 287148 17518
rect 286929 17512 287149 17513
rect 277693 17363 277913 17364
rect 286929 17294 286930 17512
rect 287148 17294 287149 17512
rect 299258 17505 299259 17723
rect 299477 17505 299478 17723
rect 299258 17504 299478 17505
rect 299259 17499 299477 17504
rect 286929 17293 287149 17294
rect 286930 17288 287148 17293
rect 213905 17270 214123 17275
rect 168863 17202 169083 17203
rect 213904 17269 214124 17270
rect 168864 17197 169082 17202
rect 184011 17153 184229 17158
rect 184010 17152 184230 17153
rect 184010 16934 184011 17152
rect 184229 16934 184230 17152
rect 213904 17051 213905 17269
rect 214123 17051 214124 17269
rect 260054 17247 260272 17252
rect 260053 17246 260273 17247
rect 220689 17229 220907 17234
rect 213904 17050 214124 17051
rect 220688 17228 220908 17229
rect 213905 17045 214123 17050
rect 193466 17020 193684 17025
rect 184010 16933 184230 16934
rect 193465 17019 193685 17020
rect 184011 16928 184229 16933
rect 193465 16801 193466 17019
rect 193684 16801 193685 17019
rect 220688 17010 220689 17228
rect 220907 17010 220908 17228
rect 248712 17078 248930 17083
rect 220688 17009 220908 17010
rect 248711 17077 248931 17078
rect 220689 17004 220907 17009
rect 202004 16895 202222 16900
rect 193465 16800 193685 16801
rect 202003 16894 202223 16895
rect 193466 16795 193684 16800
rect 202003 16676 202004 16894
rect 202222 16676 202223 16894
rect 248711 16859 248712 17077
rect 248930 16859 248931 17077
rect 260053 17028 260054 17246
rect 260272 17028 260273 17246
rect 306929 17175 307139 17180
rect 306929 17170 306934 17175
rect 307134 17170 307139 17175
rect 300252 17106 300470 17111
rect 260053 17027 260273 17028
rect 300251 17105 300471 17106
rect 260054 17022 260272 17027
rect 300251 16887 300252 17105
rect 300470 16887 300471 17105
rect 306929 16964 307139 16970
rect 300251 16886 300471 16887
rect 300252 16881 300470 16886
rect 248711 16858 248931 16859
rect 248712 16853 248930 16858
rect 202003 16675 202223 16676
rect 202004 16670 202222 16675
rect 103 15588 313 15593
rect 103 15583 108 15588
rect 308 15583 313 15588
rect 103 15377 313 15383
<< via3 >>
rect 302503 324533 302713 324538
rect 302503 324338 302508 324533
rect 302508 324338 302708 324533
rect 302708 324338 302713 324533
rect 19870 19189 20088 19193
rect 19870 18979 19874 19189
rect 19874 18979 20084 19189
rect 20084 18979 20088 19189
rect 19870 18975 20088 18979
rect 5329 18780 5547 18784
rect 5329 18570 5333 18780
rect 5333 18570 5543 18780
rect 5543 18570 5547 18780
rect 5329 18566 5547 18570
rect 7483 18887 7701 18891
rect 7483 18677 7487 18887
rect 7487 18677 7697 18887
rect 7697 18677 7701 18887
rect 7483 18673 7701 18677
rect 10712 18831 10930 18835
rect 10712 18621 10716 18831
rect 10716 18621 10926 18831
rect 10926 18621 10930 18831
rect 10712 18617 10930 18621
rect 13802 18925 14020 18929
rect 13802 18715 13806 18925
rect 13806 18715 14016 18925
rect 14016 18715 14020 18925
rect 13802 18711 14020 18715
rect 16912 18812 17130 18816
rect 16912 18602 16916 18812
rect 16916 18602 17126 18812
rect 17126 18602 17130 18812
rect 16912 18598 17130 18602
rect 25944 19007 26162 19011
rect 25944 18797 25948 19007
rect 25948 18797 26158 19007
rect 26158 18797 26162 19007
rect 25944 18793 26162 18797
rect 29085 18843 29303 19061
rect 32329 18982 32547 18986
rect 32329 18772 32333 18982
rect 32333 18772 32543 18982
rect 32543 18772 32547 18982
rect 32329 18768 32547 18772
rect 35329 19051 35547 19055
rect 35329 18841 35333 19051
rect 35333 18841 35543 19051
rect 35543 18841 35547 19051
rect 35329 18837 35547 18841
rect 38329 19214 38547 19218
rect 38329 19004 38333 19214
rect 38333 19004 38543 19214
rect 38543 19004 38547 19214
rect 38329 19000 38547 19004
rect 22898 18654 23116 18658
rect 22898 18444 22902 18654
rect 22902 18444 23112 18654
rect 23112 18444 23116 18654
rect 22898 18440 23116 18444
rect 41329 18868 41547 18872
rect 41329 18658 41333 18868
rect 41333 18658 41543 18868
rect 41543 18658 41547 18868
rect 41329 18654 41547 18658
rect 44329 18919 44547 18923
rect 44329 18709 44333 18919
rect 44333 18709 44543 18919
rect 44543 18709 44547 18919
rect 44329 18705 44547 18709
rect 47329 19126 47547 19130
rect 47329 18916 47333 19126
rect 47333 18916 47543 19126
rect 47543 18916 47547 19126
rect 47329 18912 47547 18916
rect 50517 19007 50735 19011
rect 50517 18797 50521 19007
rect 50521 18797 50731 19007
rect 50731 18797 50735 19007
rect 50517 18793 50735 18797
rect 53538 19038 53756 19042
rect 53538 18828 53542 19038
rect 53542 18828 53752 19038
rect 53752 18828 53756 19038
rect 53538 18824 53756 18828
rect 56616 19158 56834 19162
rect 56616 18948 56620 19158
rect 56620 18948 56830 19158
rect 56830 18948 56834 19158
rect 56616 18944 56834 18948
rect 59631 18862 59849 18866
rect 59631 18652 59635 18862
rect 59635 18652 59845 18862
rect 59845 18652 59849 18862
rect 59631 18648 59849 18652
rect 62633 18786 62851 18790
rect 62633 18576 62637 18786
rect 62637 18576 62847 18786
rect 62847 18576 62851 18786
rect 62633 18572 62851 18576
rect 65743 18877 65961 18881
rect 65743 18667 65747 18877
rect 65747 18667 65957 18877
rect 65957 18667 65961 18877
rect 65743 18663 65961 18667
rect 68329 18734 68547 18952
rect 71929 18842 72147 19060
rect 75079 19026 75297 19030
rect 75079 18816 75083 19026
rect 75083 18816 75293 19026
rect 75293 18816 75297 19026
rect 75079 18812 75297 18816
rect 81191 18706 81409 18905
rect 81191 18687 81195 18706
rect 81195 18687 81405 18706
rect 81405 18687 81409 18706
rect 2329 18435 2547 18439
rect 2329 18225 2333 18435
rect 2333 18225 2543 18435
rect 2543 18225 2547 18435
rect 2329 18221 2547 18225
rect 90413 18833 90631 18837
rect 90413 18623 90417 18833
rect 90417 18623 90627 18833
rect 90627 18623 90631 18833
rect 90413 18619 90631 18623
rect 93557 18789 93775 18793
rect 93557 18579 93561 18789
rect 93561 18579 93771 18789
rect 93771 18579 93775 18789
rect 93557 18575 93775 18579
rect 96454 18871 96672 18875
rect 96454 18661 96458 18871
rect 96458 18661 96668 18871
rect 96668 18661 96672 18871
rect 96454 18657 96672 18661
rect 108902 19028 109120 19032
rect 108902 18818 108906 19028
rect 108906 18818 109116 19028
rect 109116 18818 109120 19028
rect 108902 18814 109120 18818
rect 102712 18736 102930 18740
rect 102712 18526 102716 18736
rect 102716 18526 102926 18736
rect 102926 18526 102930 18736
rect 102712 18522 102930 18526
rect 105676 18751 105894 18755
rect 105676 18541 105680 18751
rect 105680 18541 105890 18751
rect 105890 18541 105894 18751
rect 105676 18537 105894 18541
rect 111949 18931 112167 18935
rect 111949 18721 111953 18931
rect 111953 18721 112163 18931
rect 112163 18721 112167 18931
rect 111949 18717 112167 18721
rect 114954 18980 115172 18984
rect 114954 18770 114958 18980
rect 114958 18770 115168 18980
rect 115168 18770 115172 18980
rect 114954 18766 115172 18770
rect 117969 18973 118187 18977
rect 117969 18763 117973 18973
rect 117973 18763 118183 18973
rect 118183 18763 118187 18973
rect 117969 18759 118187 18763
rect 121151 18860 121369 18864
rect 121151 18650 121155 18860
rect 121155 18650 121365 18860
rect 121365 18650 121369 18860
rect 121151 18646 121369 18650
rect 124119 18633 124337 18851
rect 127242 18938 127460 18942
rect 127242 18728 127246 18938
rect 127246 18728 127456 18938
rect 127456 18728 127460 18938
rect 127242 18724 127460 18728
rect 130251 18809 130469 18813
rect 130251 18599 130255 18809
rect 130255 18599 130465 18809
rect 130465 18599 130469 18809
rect 130251 18595 130469 18599
rect 133413 18648 133631 18866
rect 78099 18088 78317 18306
rect -6204 17747 -6199 17942
rect -6199 17747 -5999 17942
rect -5999 17747 -5994 17942
rect 84275 18185 84493 18403
rect 87336 18310 87554 18314
rect 87336 18100 87340 18310
rect 87340 18100 87550 18310
rect 87550 18100 87554 18310
rect 87336 18096 87554 18100
rect 99598 18497 99816 18501
rect 99598 18287 99602 18497
rect 99602 18287 99812 18497
rect 99812 18287 99816 18497
rect 99598 18283 99816 18287
rect 139553 18596 139771 18600
rect 139553 18386 139557 18596
rect 139557 18386 139767 18596
rect 139767 18386 139771 18596
rect 139553 18382 139771 18386
rect 142600 18664 142818 18668
rect 142600 18454 142604 18664
rect 142604 18454 142814 18664
rect 142814 18454 142818 18664
rect 142600 18450 142818 18454
rect 145579 18839 145797 18843
rect 145579 18629 145583 18839
rect 145583 18629 145793 18839
rect 145793 18629 145797 18839
rect 145579 18625 145797 18629
rect 148755 18839 148973 18843
rect 148755 18629 148759 18839
rect 148759 18629 148969 18839
rect 148969 18629 148973 18839
rect 148755 18625 148973 18629
rect 151773 18770 151991 18774
rect 151773 18560 151777 18770
rect 151777 18560 151987 18770
rect 151987 18560 151991 18770
rect 151773 18556 151991 18560
rect 154793 18854 155011 18858
rect 154793 18644 154797 18854
rect 154797 18644 155007 18854
rect 155007 18644 155011 18854
rect 154793 18640 155011 18644
rect 157844 18993 158062 18997
rect 157844 18783 157848 18993
rect 157848 18783 158058 18993
rect 158058 18783 158062 18993
rect 157844 18779 158062 18783
rect 174367 19131 174585 19135
rect 174367 18921 174371 19131
rect 174371 18921 174581 19131
rect 174581 18921 174585 19131
rect 174367 18917 174585 18921
rect 160887 18754 161105 18758
rect 160887 18544 160891 18754
rect 160891 18544 161101 18754
rect 161101 18544 161105 18754
rect 160887 18540 161105 18544
rect 176329 18808 176547 18812
rect 176329 18598 176333 18808
rect 176333 18598 176543 18808
rect 176543 18598 176547 18808
rect 176329 18594 176547 18598
rect 229659 18935 229877 18939
rect 229659 18725 229663 18935
rect 229663 18725 229873 18935
rect 229873 18725 229877 18935
rect 229659 18721 229877 18725
rect 290329 18951 290547 18955
rect 290329 18741 290333 18951
rect 290333 18741 290543 18951
rect 290543 18741 290547 18951
rect 290329 18737 290547 18741
rect 305386 19095 305604 19099
rect 305386 18885 305390 19095
rect 305390 18885 305600 19095
rect 305600 18885 305604 19095
rect 305386 18881 305604 18885
rect 163239 18455 163457 18459
rect 163239 18245 163243 18455
rect 163243 18245 163453 18455
rect 163453 18245 163457 18455
rect 163239 18241 163457 18245
rect 173083 18485 173301 18489
rect 173083 18275 173087 18485
rect 173087 18275 173297 18485
rect 173297 18275 173301 18485
rect 173083 18271 173301 18275
rect 136468 18237 136686 18241
rect 136468 18027 136472 18237
rect 136472 18027 136682 18237
rect 136682 18027 136686 18237
rect 136468 18023 136686 18027
rect 206329 18451 206547 18455
rect 206329 18241 206333 18451
rect 206333 18241 206543 18451
rect 206543 18241 206547 18451
rect 206329 18237 206547 18241
rect 215329 18559 215547 18563
rect 215329 18349 215333 18559
rect 215333 18349 215543 18559
rect 215543 18349 215547 18559
rect 215329 18345 215547 18349
rect 233329 18685 233547 18689
rect 233329 18475 233333 18685
rect 233333 18475 233543 18685
rect 233543 18475 233547 18685
rect 233329 18471 233547 18475
rect 227195 18424 227413 18428
rect 227195 18214 227199 18424
rect 227199 18214 227409 18424
rect 227409 18214 227413 18424
rect 227195 18210 227413 18214
rect 241673 18530 241891 18534
rect 241673 18320 241677 18530
rect 241677 18320 241887 18530
rect 241887 18320 241891 18530
rect 241673 18316 241891 18320
rect 242329 18566 242547 18570
rect 242329 18356 242333 18566
rect 242333 18356 242543 18566
rect 242543 18356 242547 18566
rect 242329 18352 242547 18356
rect 165929 18170 166147 18174
rect 165929 17960 165933 18170
rect 165933 17960 166143 18170
rect 166143 17960 166147 18170
rect 165929 17956 166147 17960
rect -6204 17742 -5994 17747
rect 182474 17855 182692 17859
rect 182474 17645 182478 17855
rect 182478 17645 182688 17855
rect 182688 17645 182692 17855
rect 182474 17641 182692 17645
rect 185329 18032 185547 18036
rect 185329 17822 185333 18032
rect 185333 17822 185543 18032
rect 185543 17822 185547 18032
rect 185329 17818 185547 17822
rect 196794 17925 197012 17929
rect 196794 17715 196798 17925
rect 196798 17715 197008 17925
rect 197008 17715 197012 17925
rect 196794 17711 197012 17715
rect 200916 17952 201134 17956
rect 200916 17742 200920 17952
rect 200920 17742 201130 17952
rect 201130 17742 201134 17952
rect 200916 17738 201134 17742
rect 213156 18094 213374 18098
rect 213156 17884 213160 18094
rect 213160 17884 213370 18094
rect 213370 17884 213374 18094
rect 213156 17880 213374 17884
rect 234651 18299 234869 18303
rect 234651 18089 234655 18299
rect 234655 18089 234865 18299
rect 234865 18089 234869 18299
rect 234651 18085 234869 18089
rect 253926 18505 254144 18509
rect 253926 18295 253930 18505
rect 253930 18295 254140 18505
rect 254140 18295 254144 18505
rect 253926 18291 254144 18295
rect 254329 18696 254547 18700
rect 254329 18486 254333 18696
rect 254333 18486 254543 18696
rect 254543 18486 254547 18696
rect 254329 18482 254547 18486
rect 269033 18556 269251 18560
rect 269033 18346 269037 18556
rect 269037 18346 269247 18556
rect 269247 18346 269251 18556
rect 269033 18342 269251 18346
rect 279677 18694 279895 18698
rect 279677 18484 279681 18694
rect 279681 18484 279891 18694
rect 279891 18484 279895 18694
rect 279677 18480 279895 18484
rect 240917 18011 241135 18015
rect 240917 17801 240921 18011
rect 240921 17801 241131 18011
rect 241131 17801 241135 18011
rect 240917 17797 241135 17801
rect 261045 18121 261263 18125
rect 261045 17911 261049 18121
rect 261049 17911 261259 18121
rect 261259 17911 261263 18121
rect 261045 17907 261263 17911
rect 269329 18264 269547 18268
rect 269329 18054 269333 18264
rect 269333 18054 269543 18264
rect 269543 18054 269547 18264
rect 269329 18050 269547 18054
rect 278879 18202 279097 18206
rect 278879 17992 278883 18202
rect 278883 17992 279093 18202
rect 279093 17992 279097 18202
rect 278879 17988 279097 17992
rect 188329 17655 188547 17659
rect 188329 17445 188333 17655
rect 188333 17445 188543 17655
rect 188543 17445 188547 17655
rect 188329 17441 188547 17445
rect 207000 17747 207218 17751
rect 207000 17537 207004 17747
rect 207004 17537 207214 17747
rect 207214 17537 207218 17747
rect 207000 17533 207218 17537
rect 221329 17707 221547 17711
rect 221329 17497 221333 17707
rect 221333 17497 221543 17707
rect 221543 17497 221547 17707
rect 221329 17493 221547 17497
rect 249668 17856 249886 17860
rect 249668 17646 249672 17856
rect 249672 17646 249882 17856
rect 249882 17646 249886 17856
rect 249668 17642 249886 17646
rect 265871 17959 266089 17963
rect 265871 17749 265875 17959
rect 265875 17749 266085 17959
rect 266085 17749 266089 17959
rect 265871 17745 266089 17749
rect 284329 18133 284547 18137
rect 284329 17923 284333 18133
rect 284333 17923 284543 18133
rect 284543 17923 284547 18133
rect 284329 17919 284547 17923
rect 292408 18223 292626 18227
rect 292408 18013 292412 18223
rect 292412 18013 292622 18223
rect 292622 18013 292626 18223
rect 292408 18009 292626 18013
rect 168864 17417 169082 17421
rect 168864 17207 168868 17417
rect 168868 17207 169078 17417
rect 169078 17207 169082 17417
rect 168864 17203 169082 17207
rect 277694 17578 277912 17582
rect 277694 17368 277698 17578
rect 277698 17368 277908 17578
rect 277908 17368 277912 17578
rect 277694 17364 277912 17368
rect 286930 17508 287148 17512
rect 286930 17298 286934 17508
rect 286934 17298 287144 17508
rect 287144 17298 287148 17508
rect 286930 17294 287148 17298
rect 299259 17719 299477 17723
rect 299259 17509 299263 17719
rect 299263 17509 299473 17719
rect 299473 17509 299477 17719
rect 299259 17505 299477 17509
rect 184011 17148 184229 17152
rect 184011 16938 184015 17148
rect 184015 16938 184225 17148
rect 184225 16938 184229 17148
rect 184011 16934 184229 16938
rect 213905 17265 214123 17269
rect 213905 17055 213909 17265
rect 213909 17055 214119 17265
rect 214119 17055 214123 17265
rect 213905 17051 214123 17055
rect 193466 17015 193684 17019
rect 193466 16805 193470 17015
rect 193470 16805 193680 17015
rect 193680 16805 193684 17015
rect 193466 16801 193684 16805
rect 220689 17224 220907 17228
rect 220689 17014 220693 17224
rect 220693 17014 220903 17224
rect 220903 17014 220907 17224
rect 220689 17010 220907 17014
rect 202004 16890 202222 16894
rect 202004 16680 202008 16890
rect 202008 16680 202218 16890
rect 202218 16680 202222 16890
rect 202004 16676 202222 16680
rect 248712 17073 248930 17077
rect 248712 16863 248716 17073
rect 248716 16863 248926 17073
rect 248926 16863 248930 17073
rect 248712 16859 248930 16863
rect 260054 17242 260272 17246
rect 260054 17032 260058 17242
rect 260058 17032 260268 17242
rect 260268 17032 260272 17242
rect 260054 17028 260272 17032
rect 300252 17101 300470 17105
rect 300252 16891 300256 17101
rect 300256 16891 300466 17101
rect 300466 16891 300470 17101
rect 300252 16887 300470 16891
rect 306929 16975 306934 17170
rect 306934 16975 307134 17170
rect 307134 16975 307139 17170
rect 306929 16970 307139 16975
rect 103 15388 108 15583
rect 108 15388 308 15583
rect 308 15388 313 15583
rect 103 15383 313 15388
<< metal4 >>
rect 2328 18467 2548 19498
rect 5328 18810 5548 19607
rect 7470 18892 7720 18911
rect 8328 18892 8548 19654
rect 7470 18891 8548 18892
rect 5317 18784 5567 18810
rect 5317 18566 5329 18784
rect 5547 18566 5567 18784
rect 7470 18673 7483 18891
rect 7701 18673 8548 18891
rect 7470 18672 8548 18673
rect 10692 18836 10942 18858
rect 11328 18836 11548 19678
rect 10692 18835 11548 18836
rect 7470 18653 7720 18672
rect 10692 18617 10712 18835
rect 10930 18617 11548 18835
rect 13790 18930 14040 18950
rect 14328 18930 14548 19678
rect 13790 18929 14548 18930
rect 13790 18711 13802 18929
rect 14020 18711 14548 18929
rect 13790 18710 14548 18711
rect 16900 18817 17150 18825
rect 17328 18817 17548 19673
rect 19851 19194 20101 19202
rect 20328 19194 20548 19678
rect 19851 19193 20548 19194
rect 19851 18975 19870 19193
rect 20088 18975 20548 19193
rect 19851 18974 20548 18975
rect 19851 18944 20101 18974
rect 16900 18816 17548 18817
rect 13790 18692 14040 18710
rect 10692 18616 11548 18617
rect 10692 18600 10942 18616
rect 16900 18598 16912 18816
rect 17130 18598 17548 18816
rect 16900 18597 17548 18598
rect 22872 18659 23189 18673
rect 23328 18659 23548 19678
rect 25909 19012 26226 19029
rect 26328 19012 26548 19678
rect 29328 19062 29548 19678
rect 25909 19011 26548 19012
rect 25909 18793 25944 19011
rect 26162 18793 26548 19011
rect 29084 19061 29548 19062
rect 29084 18843 29085 19061
rect 29303 18843 29548 19061
rect 29084 18842 29548 18843
rect 32328 18986 32548 19678
rect 35328 19066 35548 19597
rect 38328 19226 38548 19635
rect 38313 19218 38563 19226
rect 25909 18792 26548 18793
rect 25909 18763 26226 18792
rect 32328 18768 32329 18986
rect 32547 18768 32548 18986
rect 35298 19055 35585 19066
rect 35298 18837 35329 19055
rect 35547 18837 35585 19055
rect 38313 19000 38329 19218
rect 38547 19000 38563 19218
rect 38313 18968 38563 19000
rect 41328 18892 41548 19678
rect 44328 18936 44548 19673
rect 47328 19145 47548 19678
rect 47318 19130 47568 19145
rect 44320 18923 44570 18936
rect 35298 18828 35585 18837
rect 41318 18872 41568 18892
rect 32328 18767 32548 18768
rect 35328 18759 35548 18828
rect 22872 18658 23548 18659
rect 16900 18567 17150 18597
rect 5317 18552 5567 18566
rect 2316 18439 2566 18467
rect 2316 18221 2329 18439
rect 2547 18221 2566 18439
rect 22872 18440 22898 18658
rect 23116 18440 23548 18658
rect 41318 18654 41329 18872
rect 41547 18654 41568 18872
rect 44320 18705 44329 18923
rect 44547 18705 44570 18923
rect 47318 18912 47329 19130
rect 47547 18912 47568 19130
rect 47318 18887 47568 18912
rect 50328 19023 50548 19654
rect 53328 19065 53548 19678
rect 56328 19163 56548 19666
rect 56328 19162 56835 19163
rect 53328 19042 53770 19065
rect 50328 19011 50750 19023
rect 50328 18793 50517 19011
rect 50735 18793 50750 19011
rect 53328 18824 53538 19042
rect 53756 18824 53770 19042
rect 56328 18944 56616 19162
rect 56834 18944 56835 19162
rect 56328 18943 56835 18944
rect 53328 18823 53770 18824
rect 53520 18807 53770 18823
rect 59328 18867 59548 19678
rect 59328 18866 59850 18867
rect 50328 18792 50750 18793
rect 50500 18765 50750 18792
rect 44320 18678 44570 18705
rect 41318 18634 41568 18654
rect 59328 18648 59631 18866
rect 59849 18648 59850 18866
rect 59328 18647 59850 18648
rect 62328 18791 62548 19678
rect 65328 18882 65548 19645
rect 68328 18952 68548 19638
rect 65328 18881 65962 18882
rect 62328 18790 62852 18791
rect 62328 18572 62633 18790
rect 62851 18572 62852 18790
rect 65328 18663 65743 18881
rect 65961 18663 65962 18881
rect 68328 18734 68329 18952
rect 68547 18734 68548 18952
rect 71328 19061 71548 19631
rect 71328 19060 72148 19061
rect 71328 18842 71929 19060
rect 72147 18842 72148 19060
rect 71328 18841 72148 18842
rect 74328 19031 74548 19676
rect 74328 19030 75298 19031
rect 74328 18812 75079 19030
rect 75297 18812 75298 19030
rect 74328 18811 75298 18812
rect 68328 18733 68548 18734
rect 65328 18662 65962 18663
rect 62328 18571 62852 18572
rect 22872 18439 23548 18440
rect 22872 18407 23189 18439
rect 2316 18209 2566 18221
rect 77328 18307 77548 19678
rect 80328 18906 80548 19677
rect 80328 18905 81410 18906
rect 80328 18687 81191 18905
rect 81409 18687 81410 18905
rect 80328 18686 81410 18687
rect 83328 18404 83548 19662
rect 83328 18403 84494 18404
rect 77328 18306 78318 18307
rect 77328 18088 78099 18306
rect 78317 18088 78318 18306
rect 83328 18185 84275 18403
rect 84493 18185 84494 18403
rect 83328 18184 84494 18185
rect 86328 18315 86548 19678
rect 89328 18838 89548 19632
rect 89328 18837 90632 18838
rect 89328 18619 90413 18837
rect 90631 18619 90632 18837
rect 89328 18618 90632 18619
rect 92328 18794 92548 19624
rect 95328 18876 95548 19632
rect 95328 18875 96673 18876
rect 92328 18793 93776 18794
rect 92328 18575 93557 18793
rect 93775 18575 93776 18793
rect 95328 18657 96454 18875
rect 96672 18657 96673 18875
rect 95328 18656 96673 18657
rect 92328 18574 93776 18575
rect 98328 18502 98548 19639
rect 101328 18741 101548 19610
rect 104328 18756 104548 19632
rect 107328 19033 107548 19624
rect 107328 19032 109121 19033
rect 107328 18814 108902 19032
rect 109120 18814 109121 19032
rect 107328 18813 109121 18814
rect 110328 18936 110548 19647
rect 113328 18985 113548 19658
rect 113328 18984 115173 18985
rect 110328 18935 112168 18936
rect 104328 18755 105895 18756
rect 101328 18740 102931 18741
rect 101328 18522 102712 18740
rect 102930 18522 102931 18740
rect 104328 18537 105676 18755
rect 105894 18537 105895 18755
rect 110328 18717 111949 18935
rect 112167 18717 112168 18935
rect 113328 18766 114954 18984
rect 115172 18766 115173 18984
rect 113328 18765 115173 18766
rect 116328 18978 116548 19613
rect 116328 18977 118188 18978
rect 116328 18759 117969 18977
rect 118187 18759 118188 18977
rect 116328 18758 118188 18759
rect 119328 18865 119548 19678
rect 119328 18864 121370 18865
rect 110328 18716 112168 18717
rect 119328 18646 121151 18864
rect 121369 18646 121370 18864
rect 119328 18645 121370 18646
rect 122328 18852 122548 19659
rect 125328 18943 125548 19678
rect 125328 18942 127461 18943
rect 122328 18851 124338 18852
rect 122328 18633 124119 18851
rect 124337 18633 124338 18851
rect 125328 18724 127242 18942
rect 127460 18724 127461 18942
rect 125328 18723 127461 18724
rect 128328 18814 128548 19644
rect 131328 18867 131548 19675
rect 131328 18866 133632 18867
rect 128328 18813 130470 18814
rect 122328 18632 124338 18633
rect 128328 18595 130251 18813
rect 130469 18595 130470 18813
rect 131328 18648 133413 18866
rect 133631 18648 133632 18866
rect 131328 18647 133632 18648
rect 128328 18594 130470 18595
rect 104328 18536 105895 18537
rect 101328 18521 102931 18522
rect 98328 18501 99817 18502
rect 86328 18314 87555 18315
rect 86328 18096 87336 18314
rect 87554 18096 87555 18314
rect 98328 18283 99598 18501
rect 99816 18283 99817 18501
rect 98328 18282 99817 18283
rect 86328 18095 87555 18096
rect 134328 18242 134548 19659
rect 137328 18601 137548 19614
rect 140328 18669 140548 19678
rect 143328 18844 143548 19675
rect 146328 18844 146548 19667
rect 143328 18843 145798 18844
rect 140328 18668 142819 18669
rect 137328 18600 139772 18601
rect 137328 18382 139553 18600
rect 139771 18382 139772 18600
rect 140328 18450 142600 18668
rect 142818 18450 142819 18668
rect 143328 18625 145579 18843
rect 145797 18625 145798 18843
rect 143328 18624 145798 18625
rect 146328 18843 148974 18844
rect 146328 18625 148755 18843
rect 148973 18625 148974 18843
rect 146328 18624 148974 18625
rect 149328 18775 149548 19658
rect 152328 18859 152548 19658
rect 155328 18998 155548 19658
rect 155328 18997 158063 18998
rect 152328 18858 155012 18859
rect 149328 18774 151992 18775
rect 149328 18556 151773 18774
rect 151991 18556 151992 18774
rect 152328 18640 154793 18858
rect 155011 18640 155012 18858
rect 155328 18779 157844 18997
rect 158062 18779 158063 18997
rect 155328 18778 158063 18779
rect 152328 18639 155012 18640
rect 158328 18759 158548 19678
rect 161328 18890 161548 19666
rect 164328 19028 164548 19666
rect 167328 19136 167548 19658
rect 158328 18758 161153 18759
rect 149328 18555 151992 18556
rect 158328 18540 160887 18758
rect 161105 18540 161153 18758
rect 161328 18670 163556 18890
rect 164328 18808 166148 19028
rect 167328 18916 169083 19136
rect 158328 18539 161153 18540
rect 140328 18449 142819 18450
rect 163238 18459 163458 18670
rect 137328 18381 139772 18382
rect 134328 18241 136687 18242
rect 77328 18087 78318 18088
rect 134328 18023 136468 18241
rect 136686 18023 136687 18241
rect 163238 18241 163239 18459
rect 163457 18241 163458 18459
rect 163238 18240 163458 18241
rect 134328 18022 136687 18023
rect 165928 18174 166148 18808
rect 165928 17956 165929 18174
rect 166147 17956 166148 18174
rect 165928 17955 166148 17956
rect -6095 17942 -5993 17943
rect -5994 17742 -5993 17942
rect -6095 17741 -5993 17742
rect 168863 17421 169083 18916
rect 170328 18490 170548 19643
rect 173328 19136 173548 19678
rect 173328 19135 174586 19136
rect 173328 18917 174367 19135
rect 174585 18917 174586 19135
rect 173328 18916 174586 18917
rect 176328 18812 176548 19628
rect 176328 18594 176329 18812
rect 176547 18594 176548 18812
rect 176328 18593 176548 18594
rect 170328 18489 173302 18490
rect 170328 18271 173083 18489
rect 173301 18271 173302 18489
rect 170328 18270 173302 18271
rect 179328 17860 179548 19678
rect 182328 18782 182548 19658
rect 182328 18562 184230 18782
rect 179328 17859 182693 17860
rect 179328 17641 182474 17859
rect 182692 17641 182693 17859
rect 179328 17640 182693 17641
rect 168863 17203 168864 17421
rect 169082 17203 169083 17421
rect 168863 17202 169083 17203
rect 184010 17152 184230 18562
rect 185328 18036 185548 19678
rect 185328 17818 185329 18036
rect 185547 17818 185548 18036
rect 185328 17817 185548 17818
rect 188328 17659 188548 19658
rect 191328 18626 191548 19634
rect 191328 18406 193685 18626
rect 188328 17441 188329 17659
rect 188547 17441 188548 17659
rect 188328 17440 188548 17441
rect 184010 16934 184011 17152
rect 184229 16934 184230 17152
rect 184010 16933 184230 16934
rect 193465 17019 193685 18406
rect 194328 17930 194548 19625
rect 197328 17957 197548 19661
rect 200328 18804 200548 19625
rect 200328 18584 202223 18804
rect 197328 17956 201135 17957
rect 194328 17929 197013 17930
rect 194328 17711 196794 17929
rect 197012 17711 197013 17929
rect 197328 17738 200916 17956
rect 201134 17738 201135 17956
rect 197328 17737 201135 17738
rect 194328 17710 197013 17711
rect 193465 16801 193466 17019
rect 193684 16801 193685 17019
rect 193465 16800 193685 16801
rect 202003 16894 202223 18584
rect 203328 17752 203548 19670
rect 206328 18455 206548 19678
rect 206328 18237 206329 18455
rect 206547 18237 206548 18455
rect 206328 18236 206548 18237
rect 209328 18099 209548 19652
rect 212328 18885 212548 19634
rect 212328 18665 214124 18885
rect 209328 18098 213375 18099
rect 209328 17880 213156 18098
rect 213374 17880 213375 18098
rect 209328 17879 213375 17880
rect 203328 17751 207219 17752
rect 203328 17533 207000 17751
rect 207218 17533 207219 17751
rect 203328 17532 207219 17533
rect 213904 17269 214124 18665
rect 215328 18563 215548 19666
rect 218328 18895 218548 19678
rect 218328 18675 220908 18895
rect 215328 18345 215329 18563
rect 215547 18345 215548 18563
rect 215328 18344 215548 18345
rect 213904 17051 213905 17269
rect 214123 17051 214124 17269
rect 213904 17050 214124 17051
rect 220688 17228 220908 18675
rect 221328 17711 221548 19666
rect 224328 18429 224548 19657
rect 227328 18940 227548 19675
rect 227328 18939 229878 18940
rect 227328 18721 229659 18939
rect 229877 18721 229878 18939
rect 227328 18720 229878 18721
rect 224328 18428 227414 18429
rect 224328 18210 227195 18428
rect 227413 18210 227414 18428
rect 224328 18209 227414 18210
rect 230328 18304 230548 19648
rect 233328 18689 233548 19678
rect 233328 18471 233329 18689
rect 233547 18471 233548 18689
rect 233328 18470 233548 18471
rect 230328 18303 234870 18304
rect 230328 18085 234651 18303
rect 234869 18085 234870 18303
rect 230328 18084 234870 18085
rect 236328 18016 236548 19498
rect 239328 18535 239548 19610
rect 242328 18570 242548 19678
rect 239328 18534 241892 18535
rect 239328 18316 241673 18534
rect 241891 18316 241892 18534
rect 242328 18352 242329 18570
rect 242547 18352 242548 18570
rect 245328 18599 245548 19678
rect 248328 19091 248548 19655
rect 248328 18871 249887 19091
rect 245328 18379 248931 18599
rect 242328 18351 242548 18352
rect 239328 18315 241892 18316
rect 236328 18015 241136 18016
rect 236328 17797 240917 18015
rect 241135 17797 241136 18015
rect 236328 17796 241136 17797
rect 221328 17493 221329 17711
rect 221547 17493 221548 17711
rect 221328 17492 221548 17493
rect 220688 17010 220689 17228
rect 220907 17010 220908 17228
rect 220688 17009 220908 17010
rect 248711 17077 248931 18379
rect 249667 17860 249887 18871
rect 251328 18510 251548 19678
rect 254328 18700 254548 19678
rect 251328 18509 254145 18510
rect 251328 18291 253926 18509
rect 254144 18291 254145 18509
rect 254328 18482 254329 18700
rect 254547 18482 254548 18700
rect 254328 18481 254548 18482
rect 257328 18577 257548 19671
rect 260328 19117 260548 19678
rect 260328 18897 261264 19117
rect 257328 18357 260273 18577
rect 251328 18290 254145 18291
rect 249667 17642 249668 17860
rect 249886 17642 249887 17860
rect 249667 17641 249887 17642
rect 202003 16676 202004 16894
rect 202222 16676 202223 16894
rect 248711 16859 248712 17077
rect 248930 16859 248931 17077
rect 260053 17246 260273 18357
rect 261044 18125 261264 18897
rect 261044 17907 261045 18125
rect 261263 17907 261264 18125
rect 261044 17906 261264 17907
rect 263328 17964 263548 19678
rect 266328 18561 266548 19621
rect 266328 18560 269252 18561
rect 266328 18342 269033 18560
rect 269251 18342 269252 18560
rect 266328 18341 269252 18342
rect 269328 18268 269548 19594
rect 269328 18050 269329 18268
rect 269547 18050 269548 18268
rect 269328 18049 269548 18050
rect 263328 17963 266146 17964
rect 263328 17745 265871 17963
rect 266089 17745 266146 17963
rect 263328 17744 266146 17745
rect 272328 17583 272548 19649
rect 275328 18207 275548 19649
rect 278328 18699 278548 19670
rect 278328 18698 279896 18699
rect 278328 18480 279677 18698
rect 279895 18480 279896 18698
rect 278328 18479 279896 18480
rect 275328 18206 279098 18207
rect 275328 17988 278879 18206
rect 279097 17988 279098 18206
rect 275328 17987 279098 17988
rect 272328 17582 277913 17583
rect 272328 17364 277694 17582
rect 277912 17364 277913 17582
rect 272328 17363 277913 17364
rect 281328 17513 281548 19678
rect 284328 18137 284548 19678
rect 284328 17919 284329 18137
rect 284547 17919 284548 18137
rect 287328 18228 287548 19670
rect 290328 18955 290548 19678
rect 290328 18737 290329 18955
rect 290547 18737 290548 18955
rect 290328 18736 290548 18737
rect 287328 18227 292627 18228
rect 287328 18009 292408 18227
rect 292626 18009 292627 18227
rect 287328 18008 292627 18009
rect 284328 17918 284548 17919
rect 293328 17724 293548 19642
rect 296328 18328 296548 19655
rect 299328 19100 299548 19678
rect 299328 19099 305605 19100
rect 299328 18881 305386 19099
rect 305604 18881 305605 19099
rect 299328 18880 305605 18881
rect 296328 18108 300471 18328
rect 293328 17723 299478 17724
rect 281328 17512 287149 17513
rect 281328 17294 286930 17512
rect 287148 17294 287149 17512
rect 293328 17505 299259 17723
rect 299477 17505 299478 17723
rect 293328 17504 299478 17505
rect 281328 17293 287149 17294
rect 260053 17028 260054 17246
rect 260272 17028 260273 17246
rect 260053 17027 260273 17028
rect 300251 17105 300471 18108
rect 300251 16887 300252 17105
rect 300470 16887 300471 17105
rect 300251 16886 300471 16887
rect 248711 16858 248931 16859
rect 202003 16675 202223 16676
<< via4 >>
rect 302448 324538 302768 324598
rect 302448 324338 302503 324538
rect 302503 324338 302713 324538
rect 302713 324338 302768 324538
rect 302448 324278 302768 324338
rect -6415 17942 -6095 18002
rect -6415 17742 -6204 17942
rect -6204 17742 -6095 17942
rect -6415 17682 -6095 17742
rect 306874 17170 307194 17230
rect 306874 16970 306929 17170
rect 306929 16970 307139 17170
rect 307139 16970 307194 17170
rect 306874 16910 307194 16970
rect 48 15583 368 15643
rect 48 15383 103 15583
rect 103 15383 313 15583
rect 313 15383 368 15583
rect 48 15323 368 15383
<< metal5 >>
rect 302448 324637 302768 324994
rect -5612 324598 304435 324637
rect -5612 324317 302448 324598
rect 302424 324278 302448 324317
rect 302768 324317 304435 324598
rect 302768 324278 302792 324317
rect 302424 324254 302792 324278
rect -6415 18026 -6095 18186
rect -6439 18002 -6071 18026
rect -6439 17682 -6415 18002
rect -6095 17682 -6071 18002
rect -6439 17658 -6071 17682
rect -6415 17375 -6095 17658
rect 306850 17230 307218 17254
rect 306850 16910 306874 17230
rect 307194 16910 307218 17230
rect 306850 16886 307218 16910
rect 306874 16049 307194 16886
rect 24 15643 392 15667
rect 24 15323 48 15643
rect 368 15323 837 15643
rect 24 15299 392 15323
use shift_registerC  shift_registerC_0
timestamp 1654738065
transform 1 0 58 0 1 590
box -1076 -4 307988 16000
use pixel_array100x100  pixel_array100x100_0
timestamp 1654740282
transform 1 0 2108 0 1 317378
box -3000 -298600 300740 5750
use shift_register  shift_register_0
timestamp 1654738065
transform 0 1 -21072 -1 0 323984
box -1076 -4 307988 16000
<< end >>
