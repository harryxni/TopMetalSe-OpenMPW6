magic
tech sky130A
magscale 1 2
timestamp 1655248532
<< viali >>
rect 1593 13481 1627 13515
rect 4629 13481 4663 13515
rect 7665 13481 7699 13515
rect 10793 13481 10827 13515
rect 14105 13481 14139 13515
rect 16865 13481 16899 13515
rect 19993 13481 20027 13515
rect 23029 13481 23063 13515
rect 25697 13481 25731 13515
rect 29009 13481 29043 13515
rect 31585 13481 31619 13515
rect 47593 13481 47627 13515
rect 50353 13481 50387 13515
rect 50997 13481 51031 13515
rect 142905 13481 142939 13515
rect 144745 13481 144779 13515
rect 148320 13481 148354 13515
rect 157625 13481 157659 13515
rect 182741 13481 182775 13515
rect 185777 13481 185811 13515
rect 210341 13481 210375 13515
rect 213377 13481 213411 13515
rect 269392 13481 269426 13515
rect 274281 13481 274315 13515
rect 274925 13481 274959 13515
rect 277869 13481 277903 13515
rect 280905 13481 280939 13515
rect 284585 13481 284619 13515
rect 287161 13481 287195 13515
rect 290105 13481 290139 13515
rect 293233 13481 293267 13515
rect 296269 13481 296303 13515
rect 299305 13481 299339 13515
rect 301421 13481 301455 13515
rect 301789 13481 301823 13515
rect 302157 13481 302191 13515
rect 302985 13481 303019 13515
rect 303353 13481 303387 13515
rect 44281 13413 44315 13447
rect 60473 13413 60507 13447
rect 63049 13413 63083 13447
rect 75377 13413 75411 13447
rect 93961 13413 93995 13447
rect 101137 13413 101171 13447
rect 109417 13413 109451 13447
rect 111257 13413 111291 13447
rect 121285 13413 121319 13447
rect 124137 13413 124171 13447
rect 136649 13413 136683 13447
rect 140329 13413 140363 13447
rect 155785 13413 155819 13447
rect 170413 13413 170447 13447
rect 173081 13413 173115 13447
rect 173817 13413 173851 13447
rect 175841 13413 175875 13447
rect 178141 13413 178175 13447
rect 181545 13413 181579 13447
rect 199853 13413 199887 13447
rect 203901 13413 203935 13447
rect 216413 13413 216447 13447
rect 220185 13413 220219 13447
rect 226625 13413 226659 13447
rect 229661 13413 229695 13447
rect 239965 13413 239999 13447
rect 247141 13413 247175 13447
rect 249533 13413 249567 13447
rect 252845 13413 252879 13447
rect 255421 13413 255455 13447
rect 259469 13413 259503 13447
rect 262689 13413 262723 13447
rect 266001 13413 266035 13447
rect 26341 13345 26375 13379
rect 27261 13345 27295 13379
rect 34713 13345 34747 13379
rect 37565 13345 37599 13379
rect 45569 13345 45603 13379
rect 51641 13345 51675 13379
rect 72709 13345 72743 13379
rect 73629 13345 73663 13379
rect 78505 13345 78539 13379
rect 80253 13345 80287 13379
rect 81541 13345 81575 13379
rect 81633 13345 81667 13379
rect 98009 13345 98043 13379
rect 98193 13345 98227 13379
rect 112269 13345 112303 13379
rect 120273 13345 120307 13379
rect 125701 13345 125735 13379
rect 126713 13345 126747 13379
rect 130301 13345 130335 13379
rect 132601 13345 132635 13379
rect 148057 13345 148091 13379
rect 150909 13345 150943 13379
rect 153485 13345 153519 13379
rect 160937 13345 160971 13379
rect 166641 13345 166675 13379
rect 167561 13345 167595 13379
rect 174277 13345 174311 13379
rect 174369 13345 174403 13379
rect 178969 13345 179003 13379
rect 182097 13345 182131 13379
rect 188537 13345 188571 13379
rect 189825 13345 189859 13379
rect 198749 13345 198783 13379
rect 201141 13345 201175 13379
rect 204729 13345 204763 13379
rect 207857 13345 207891 13379
rect 224325 13345 224359 13379
rect 227085 13345 227119 13379
rect 227177 13345 227211 13379
rect 230489 13345 230523 13379
rect 232237 13345 232271 13379
rect 237205 13345 237239 13379
rect 237297 13345 237331 13379
rect 240793 13345 240827 13379
rect 243369 13345 243403 13379
rect 245117 13345 245151 13379
rect 250177 13345 250211 13379
rect 262045 13345 262079 13379
rect 263241 13345 263275 13379
rect 266553 13345 266587 13379
rect 269129 13345 269163 13379
rect 271705 13345 271739 13379
rect 304457 13345 304491 13379
rect 304917 13345 304951 13379
rect 305377 13345 305411 13379
rect 1777 13277 1811 13311
rect 4813 13277 4847 13311
rect 7849 13277 7883 13311
rect 10977 13277 11011 13311
rect 14289 13277 14323 13311
rect 17049 13277 17083 13311
rect 20177 13277 20211 13311
rect 23213 13277 23247 13311
rect 26065 13277 26099 13311
rect 29837 13277 29871 13311
rect 32413 13277 32447 13311
rect 40141 13277 40175 13311
rect 42533 13277 42567 13311
rect 47777 13277 47811 13311
rect 50537 13277 50571 13311
rect 51365 13277 51399 13311
rect 53021 13277 53055 13311
rect 55597 13277 55631 13311
rect 57897 13277 57931 13311
rect 60657 13277 60691 13311
rect 63233 13277 63267 13311
rect 66177 13277 66211 13311
rect 69305 13277 69339 13311
rect 72525 13277 72559 13311
rect 76205 13277 76239 13311
rect 82461 13277 82495 13311
rect 83105 13277 83139 13311
rect 83933 13277 83967 13311
rect 86509 13277 86543 13311
rect 88809 13277 88843 13311
rect 94145 13277 94179 13311
rect 96905 13277 96939 13311
rect 99389 13277 99423 13311
rect 101965 13277 101999 13311
rect 104265 13277 104299 13311
rect 109601 13277 109635 13311
rect 111441 13277 111475 13311
rect 114845 13277 114879 13311
rect 117421 13277 117455 13311
rect 120181 13277 120215 13311
rect 121469 13277 121503 13311
rect 124321 13277 124355 13311
rect 126621 13277 126655 13311
rect 127541 13277 127575 13311
rect 136833 13277 136867 13311
rect 140513 13277 140547 13311
rect 143089 13277 143123 13311
rect 144929 13277 144963 13311
rect 145757 13277 145791 13311
rect 155969 13277 156003 13311
rect 156429 13277 156463 13311
rect 157809 13277 157843 13311
rect 158637 13277 158671 13311
rect 163513 13277 163547 13311
rect 170597 13277 170631 13311
rect 173265 13277 173299 13311
rect 174185 13277 174219 13311
rect 175657 13277 175691 13311
rect 176393 13277 176427 13311
rect 182005 13277 182039 13311
rect 182925 13277 182959 13311
rect 185961 13277 185995 13311
rect 187341 13277 187375 13311
rect 188445 13277 188479 13311
rect 189549 13277 189583 13311
rect 191849 13277 191883 13311
rect 194425 13277 194459 13311
rect 200037 13277 200071 13311
rect 202153 13277 202187 13311
rect 207673 13277 207707 13311
rect 210525 13277 210559 13311
rect 213561 13277 213595 13311
rect 216597 13277 216631 13311
rect 220369 13277 220403 13311
rect 222945 13277 222979 13311
rect 225889 13277 225923 13311
rect 227913 13277 227947 13311
rect 233065 13277 233099 13311
rect 233893 13277 233927 13311
rect 235089 13277 235123 13311
rect 237113 13277 237147 13311
rect 238217 13277 238251 13311
rect 247325 13277 247359 13311
rect 249993 13277 250027 13311
rect 251097 13277 251131 13311
rect 253673 13277 253707 13311
rect 256249 13277 256283 13311
rect 259653 13277 259687 13311
rect 264253 13277 264287 13311
rect 268577 13277 268611 13311
rect 274465 13277 274499 13311
rect 275109 13277 275143 13311
rect 278053 13277 278087 13311
rect 281089 13277 281123 13311
rect 284769 13277 284803 13311
rect 287345 13277 287379 13311
rect 290289 13277 290323 13311
rect 293417 13277 293451 13311
rect 296453 13277 296487 13311
rect 299489 13277 299523 13311
rect 303721 13277 303755 13311
rect 27537 13209 27571 13243
rect 30113 13209 30147 13243
rect 32689 13209 32723 13243
rect 34989 13209 35023 13243
rect 37841 13209 37875 13243
rect 40417 13209 40451 13243
rect 42809 13209 42843 13243
rect 45477 13209 45511 13243
rect 53297 13209 53331 13243
rect 55873 13209 55907 13243
rect 58173 13209 58207 13243
rect 73905 13209 73939 13243
rect 76481 13209 76515 13243
rect 78781 13209 78815 13243
rect 84209 13209 84243 13243
rect 86785 13209 86819 13243
rect 89085 13209 89119 13243
rect 91845 13209 91879 13243
rect 92029 13209 92063 13243
rect 99665 13209 99699 13243
rect 102241 13209 102275 13243
rect 104541 13209 104575 13243
rect 112545 13209 112579 13243
rect 115121 13209 115155 13243
rect 117697 13209 117731 13243
rect 120089 13209 120123 13243
rect 125517 13209 125551 13243
rect 127817 13209 127851 13243
rect 130577 13209 130611 13243
rect 132877 13209 132911 13243
rect 146033 13209 146067 13243
rect 150081 13209 150115 13243
rect 151185 13209 151219 13243
rect 153761 13209 153795 13243
rect 156521 13209 156555 13243
rect 158913 13209 158947 13243
rect 161213 13209 161247 13243
rect 163789 13209 163823 13243
rect 166549 13209 166583 13243
rect 167377 13209 167411 13243
rect 176669 13209 176703 13243
rect 179245 13209 179279 13243
rect 181913 13209 181947 13243
rect 187433 13209 187467 13243
rect 192125 13209 192159 13243
rect 193873 13209 193907 13243
rect 194701 13209 194735 13243
rect 196449 13209 196483 13243
rect 197829 13209 197863 13243
rect 198657 13209 198691 13243
rect 202429 13209 202463 13243
rect 205005 13209 205039 13243
rect 228189 13209 228223 13243
rect 230765 13209 230799 13243
rect 238493 13209 238527 13243
rect 241069 13209 241103 13243
rect 243645 13209 243679 13243
rect 251373 13209 251407 13243
rect 253949 13209 253983 13243
rect 256525 13209 256559 13243
rect 261861 13209 261895 13243
rect 263057 13209 263091 13243
rect 264529 13209 264563 13243
rect 266829 13209 266863 13243
rect 271981 13209 272015 13243
rect 26157 13141 26191 13175
rect 34161 13141 34195 13175
rect 36461 13141 36495 13175
rect 39313 13141 39347 13175
rect 41889 13141 41923 13175
rect 45017 13141 45051 13175
rect 45385 13141 45419 13175
rect 51457 13141 51491 13175
rect 54769 13141 54803 13175
rect 57345 13141 57379 13175
rect 59645 13141 59679 13175
rect 65993 13141 66027 13175
rect 69121 13141 69155 13175
rect 72065 13141 72099 13175
rect 72433 13141 72467 13175
rect 77953 13141 77987 13175
rect 81081 13141 81115 13175
rect 81449 13141 81483 13175
rect 82277 13141 82311 13175
rect 82921 13141 82955 13175
rect 85681 13141 85715 13175
rect 88257 13141 88291 13175
rect 90557 13141 90591 13175
rect 96721 13141 96755 13175
rect 97549 13141 97583 13175
rect 97917 13141 97951 13175
rect 103713 13141 103747 13175
rect 106013 13141 106047 13175
rect 114017 13141 114051 13175
rect 116593 13141 116627 13175
rect 119169 13141 119203 13175
rect 119721 13141 119755 13175
rect 126161 13141 126195 13175
rect 126529 13141 126563 13175
rect 129289 13141 129323 13175
rect 132049 13141 132083 13175
rect 134349 13141 134383 13175
rect 147505 13141 147539 13175
rect 152657 13141 152691 13175
rect 155233 13141 155267 13175
rect 160385 13141 160419 13175
rect 162685 13141 162719 13175
rect 165261 13141 165295 13175
rect 166089 13141 166123 13175
rect 166457 13141 166491 13175
rect 180717 13141 180751 13175
rect 187985 13141 188019 13175
rect 188353 13141 188387 13175
rect 191297 13141 191331 13175
rect 198197 13141 198231 13175
rect 198565 13141 198599 13175
rect 200497 13141 200531 13175
rect 200865 13141 200899 13175
rect 200957 13141 200991 13175
rect 206477 13141 206511 13175
rect 207305 13141 207339 13175
rect 207765 13141 207799 13175
rect 222761 13141 222795 13175
rect 223681 13141 223715 13175
rect 224049 13141 224083 13175
rect 224141 13141 224175 13175
rect 225705 13141 225739 13175
rect 226993 13141 227027 13175
rect 233157 13141 233191 13175
rect 233709 13141 233743 13175
rect 234905 13141 234939 13175
rect 236745 13141 236779 13175
rect 242541 13141 242575 13175
rect 249901 13141 249935 13175
rect 257997 13141 258031 13175
rect 263149 13141 263183 13175
rect 270877 13141 270911 13175
rect 273453 13141 273487 13175
rect 295901 13141 295935 13175
rect 26065 12937 26099 12971
rect 27445 12937 27479 12971
rect 33885 12937 33919 12971
rect 34805 12937 34839 12971
rect 35541 12937 35575 12971
rect 36645 12937 36679 12971
rect 42533 12937 42567 12971
rect 43453 12937 43487 12971
rect 44557 12937 44591 12971
rect 52009 12937 52043 12971
rect 53573 12937 53607 12971
rect 53941 12937 53975 12971
rect 58541 12937 58575 12971
rect 72157 12937 72191 12971
rect 89545 12937 89579 12971
rect 91109 12937 91143 12971
rect 112269 12937 112303 12971
rect 118249 12937 118283 12971
rect 118709 12937 118743 12971
rect 126713 12937 126747 12971
rect 128093 12937 128127 12971
rect 128737 12937 128771 12971
rect 129197 12937 129231 12971
rect 130301 12937 130335 12971
rect 133521 12937 133555 12971
rect 134349 12937 134383 12971
rect 145481 12937 145515 12971
rect 151461 12937 151495 12971
rect 152749 12937 152783 12971
rect 153117 12937 153151 12971
rect 153485 12937 153519 12971
rect 153853 12937 153887 12971
rect 154221 12937 154255 12971
rect 154957 12937 154991 12971
rect 156061 12937 156095 12971
rect 156429 12937 156463 12971
rect 156797 12937 156831 12971
rect 157165 12937 157199 12971
rect 163605 12937 163639 12971
rect 164433 12937 164467 12971
rect 167837 12937 167871 12971
rect 175013 12937 175047 12971
rect 175657 12937 175691 12971
rect 180809 12937 180843 12971
rect 192309 12937 192343 12971
rect 195989 12937 196023 12971
rect 206569 12937 206603 12971
rect 252385 12937 252419 12971
rect 264621 12937 264655 12971
rect 302617 12937 302651 12971
rect 304457 12937 304491 12971
rect 29009 12869 29043 12903
rect 36553 12869 36587 12903
rect 37381 12869 37415 12903
rect 38485 12869 38519 12903
rect 39773 12869 39807 12903
rect 58633 12869 58667 12903
rect 77861 12869 77895 12903
rect 78597 12869 78631 12903
rect 99481 12869 99515 12903
rect 104633 12869 104667 12903
rect 104725 12869 104759 12903
rect 112361 12869 112395 12903
rect 114017 12869 114051 12903
rect 115673 12869 115707 12903
rect 133613 12869 133647 12903
rect 145941 12869 145975 12903
rect 159281 12869 159315 12903
rect 164525 12869 164559 12903
rect 181637 12869 181671 12903
rect 189549 12869 189583 12903
rect 190929 12869 190963 12903
rect 193321 12869 193355 12903
rect 195897 12869 195931 12903
rect 231041 12869 231075 12903
rect 238769 12869 238803 12903
rect 240977 12869 241011 12903
rect 245301 12869 245335 12903
rect 251373 12869 251407 12903
rect 252477 12869 252511 12903
rect 261769 12869 261803 12903
rect 263241 12869 263275 12903
rect 263425 12869 263459 12903
rect 265541 12869 265575 12903
rect 271797 12869 271831 12903
rect 272901 12869 272935 12903
rect 305009 12869 305043 12903
rect 305469 12869 305503 12903
rect 26249 12801 26283 12835
rect 27813 12801 27847 12835
rect 34713 12801 34747 12835
rect 35725 12801 35759 12835
rect 38393 12801 38427 12835
rect 41705 12801 41739 12835
rect 42441 12801 42475 12835
rect 44741 12801 44775 12835
rect 52193 12801 52227 12835
rect 52929 12801 52963 12835
rect 54033 12801 54067 12835
rect 54769 12801 54803 12835
rect 57069 12801 57103 12835
rect 72341 12801 72375 12835
rect 75101 12801 75135 12835
rect 75561 12801 75595 12835
rect 77769 12801 77803 12835
rect 78505 12801 78539 12835
rect 79333 12801 79367 12835
rect 79793 12801 79827 12835
rect 86233 12801 86267 12835
rect 90465 12801 90499 12835
rect 91293 12801 91327 12835
rect 98561 12801 98595 12835
rect 106105 12801 106139 12835
rect 113097 12801 113131 12835
rect 113833 12801 113867 12835
rect 114661 12801 114695 12835
rect 118893 12801 118927 12835
rect 126897 12801 126931 12835
rect 127449 12801 127483 12835
rect 128277 12801 128311 12835
rect 129105 12801 129139 12835
rect 130209 12801 130243 12835
rect 130853 12801 130887 12835
rect 134533 12801 134567 12835
rect 135361 12801 135395 12835
rect 142997 12801 143031 12835
rect 145849 12801 145883 12835
rect 147045 12801 147079 12835
rect 149897 12801 149931 12835
rect 154865 12801 154899 12835
rect 159189 12801 159223 12835
rect 160017 12801 160051 12835
rect 161213 12801 161247 12835
rect 161857 12801 161891 12835
rect 165353 12801 165387 12835
rect 166549 12801 166583 12835
rect 167377 12801 167411 12835
rect 168021 12801 168055 12835
rect 175197 12801 175231 12835
rect 175841 12801 175875 12835
rect 176393 12801 176427 12835
rect 178601 12801 178635 12835
rect 180993 12801 181027 12835
rect 181545 12801 181579 12835
rect 182189 12801 182223 12835
rect 188077 12801 188111 12835
rect 188629 12801 188663 12835
rect 189365 12801 189399 12835
rect 191021 12801 191055 12835
rect 192217 12801 192251 12835
rect 195069 12801 195103 12835
rect 197369 12801 197403 12835
rect 197461 12801 197495 12835
rect 198381 12801 198415 12835
rect 200497 12801 200531 12835
rect 201325 12801 201359 12835
rect 204821 12801 204855 12835
rect 207489 12801 207523 12835
rect 226717 12801 226751 12835
rect 227361 12801 227395 12835
rect 227913 12801 227947 12835
rect 230305 12801 230339 12835
rect 230765 12801 230799 12835
rect 233065 12801 233099 12835
rect 237021 12801 237055 12835
rect 237665 12801 237699 12835
rect 238493 12801 238527 12835
rect 240701 12801 240735 12835
rect 243829 12801 243863 12835
rect 244565 12801 244599 12835
rect 244749 12801 244783 12835
rect 245209 12801 245243 12835
rect 250361 12801 250395 12835
rect 251557 12801 251591 12835
rect 256249 12801 256283 12835
rect 257077 12801 257111 12835
rect 262505 12801 262539 12835
rect 264161 12801 264195 12835
rect 264805 12801 264839 12835
rect 265265 12801 265299 12835
rect 267841 12801 267875 12835
rect 269129 12801 269163 12835
rect 271705 12801 271739 12835
rect 302801 12801 302835 12835
rect 304641 12801 304675 12835
rect 27905 12733 27939 12767
rect 28089 12733 28123 12767
rect 29101 12733 29135 12767
rect 29285 12733 29319 12767
rect 29837 12733 29871 12767
rect 30113 12733 30147 12767
rect 32137 12733 32171 12767
rect 32413 12733 32447 12767
rect 34897 12733 34931 12767
rect 37565 12733 37599 12767
rect 38577 12733 38611 12767
rect 39497 12733 39531 12767
rect 43545 12733 43579 12767
rect 43729 12733 43763 12767
rect 54125 12733 54159 12767
rect 55045 12733 55079 12767
rect 58725 12733 58759 12767
rect 75837 12733 75871 12767
rect 80069 12733 80103 12767
rect 84025 12733 84059 12767
rect 84301 12733 84335 12767
rect 86509 12733 86543 12767
rect 89637 12733 89671 12767
rect 89821 12733 89855 12767
rect 99205 12733 99239 12767
rect 101413 12733 101447 12767
rect 101689 12733 101723 12767
rect 104817 12733 104851 12767
rect 112545 12733 112579 12767
rect 113189 12733 113223 12767
rect 115765 12733 115799 12767
rect 115857 12733 115891 12767
rect 116501 12733 116535 12767
rect 116777 12733 116811 12767
rect 129381 12733 129415 12767
rect 131129 12733 131163 12767
rect 132601 12733 132635 12767
rect 133797 12733 133831 12767
rect 143273 12733 143307 12767
rect 146125 12733 146159 12767
rect 147505 12733 147539 12767
rect 147781 12733 147815 12767
rect 149253 12733 149287 12767
rect 151553 12733 151587 12767
rect 151737 12733 151771 12767
rect 155049 12733 155083 12767
rect 159465 12733 159499 12767
rect 162133 12733 162167 12767
rect 164617 12733 164651 12767
rect 176669 12733 176703 12767
rect 178877 12733 178911 12767
rect 191205 12733 191239 12767
rect 192401 12733 192435 12767
rect 193045 12733 193079 12767
rect 196173 12733 196207 12767
rect 197645 12733 197679 12767
rect 198105 12733 198139 12767
rect 200589 12733 200623 12767
rect 202613 12733 202647 12767
rect 202889 12733 202923 12767
rect 205097 12733 205131 12767
rect 228189 12733 228223 12767
rect 233157 12733 233191 12767
rect 252569 12733 252603 12767
rect 253673 12733 253707 12767
rect 253949 12733 253983 12767
rect 255421 12733 255455 12767
rect 256341 12733 256375 12767
rect 256433 12733 256467 12767
rect 267933 12733 267967 12767
rect 268025 12733 268059 12767
rect 269405 12733 269439 12767
rect 271981 12733 272015 12767
rect 272993 12733 273027 12767
rect 273085 12733 273119 12767
rect 74917 12665 74951 12699
rect 79149 12665 79183 12699
rect 81541 12665 81575 12699
rect 100953 12665 100987 12699
rect 105921 12665 105955 12699
rect 135545 12665 135579 12699
rect 152381 12665 152415 12699
rect 154497 12665 154531 12699
rect 158821 12665 158855 12699
rect 160201 12665 160235 12699
rect 167193 12665 167227 12699
rect 187893 12665 187927 12699
rect 207305 12665 207339 12699
rect 227177 12665 227211 12699
rect 237481 12665 237515 12699
rect 250177 12665 250211 12699
rect 255881 12665 255915 12699
rect 262689 12665 262723 12699
rect 28641 12597 28675 12631
rect 31585 12597 31619 12631
rect 34345 12597 34379 12631
rect 38025 12597 38059 12631
rect 41245 12597 41279 12631
rect 41797 12597 41831 12631
rect 43085 12597 43119 12631
rect 53021 12597 53055 12631
rect 56517 12597 56551 12631
rect 57161 12597 57195 12631
rect 58173 12597 58207 12631
rect 77309 12597 77343 12631
rect 85773 12597 85807 12631
rect 87981 12597 88015 12631
rect 89177 12597 89211 12631
rect 90557 12597 90591 12631
rect 98377 12597 98411 12631
rect 103161 12597 103195 12631
rect 104265 12597 104299 12631
rect 111901 12597 111935 12631
rect 114753 12597 114787 12631
rect 115305 12597 115339 12631
rect 127541 12597 127575 12631
rect 133153 12597 133187 12631
rect 146861 12597 146895 12631
rect 149989 12597 150023 12631
rect 151093 12597 151127 12631
rect 161305 12597 161339 12631
rect 164065 12597 164099 12631
rect 165445 12597 165479 12631
rect 166641 12597 166675 12631
rect 178141 12597 178175 12631
rect 180349 12597 180383 12631
rect 182281 12597 182315 12631
rect 188721 12597 188755 12631
rect 190561 12597 190595 12631
rect 191849 12597 191883 12631
rect 195529 12597 195563 12631
rect 197001 12597 197035 12631
rect 198197 12597 198231 12631
rect 201141 12597 201175 12631
rect 204361 12597 204395 12631
rect 226533 12597 226567 12631
rect 229661 12597 229695 12631
rect 230121 12597 230155 12631
rect 232513 12597 232547 12631
rect 236837 12597 236871 12631
rect 240241 12597 240275 12631
rect 242449 12597 242483 12631
rect 243921 12597 243955 12631
rect 252017 12597 252051 12631
rect 257169 12597 257203 12631
rect 261861 12597 261895 12631
rect 263977 12597 264011 12631
rect 267013 12597 267047 12631
rect 267473 12597 267507 12631
rect 270877 12597 270911 12631
rect 271337 12597 271371 12631
rect 272533 12597 272567 12631
rect 31309 12393 31343 12427
rect 33977 12393 34011 12427
rect 34805 12393 34839 12427
rect 37197 12393 37231 12427
rect 38485 12393 38519 12427
rect 39221 12393 39255 12427
rect 43177 12393 43211 12427
rect 43821 12393 43855 12427
rect 54125 12393 54159 12427
rect 54677 12393 54711 12427
rect 57345 12393 57379 12427
rect 57989 12393 58023 12427
rect 75193 12393 75227 12427
rect 79333 12393 79367 12427
rect 80253 12393 80287 12427
rect 85589 12393 85623 12427
rect 86417 12393 86451 12427
rect 88901 12393 88935 12427
rect 90189 12393 90223 12427
rect 99113 12393 99147 12427
rect 99849 12393 99883 12427
rect 103897 12393 103931 12427
rect 105185 12393 105219 12427
rect 113097 12393 113131 12427
rect 113741 12393 113775 12427
rect 118433 12393 118467 12427
rect 127725 12393 127759 12427
rect 130853 12393 130887 12427
rect 132693 12393 132727 12427
rect 147321 12393 147355 12427
rect 152565 12393 152599 12427
rect 154129 12393 154163 12427
rect 165353 12393 165387 12427
rect 175933 12393 175967 12427
rect 181361 12393 181395 12427
rect 188537 12393 188571 12427
rect 190193 12393 190227 12427
rect 201693 12393 201727 12427
rect 206477 12393 206511 12427
rect 227808 12393 227842 12427
rect 232237 12393 232271 12427
rect 239965 12393 239999 12427
rect 243553 12393 243587 12427
rect 244197 12393 244231 12427
rect 251097 12393 251131 12427
rect 256893 12393 256927 12427
rect 262505 12393 262539 12427
rect 264621 12393 264655 12427
rect 271061 12393 271095 12427
rect 305469 12393 305503 12427
rect 77493 12325 77527 12359
rect 89453 12325 89487 12359
rect 148425 12325 148459 12359
rect 153301 12325 153335 12359
rect 160017 12325 160051 12359
rect 166089 12325 166123 12359
rect 180901 12325 180935 12359
rect 192585 12325 192619 12359
rect 201141 12325 201175 12359
rect 229753 12325 229787 12359
rect 238769 12325 238803 12359
rect 242357 12325 242391 12359
rect 252109 12325 252143 12359
rect 254317 12325 254351 12359
rect 256341 12325 256375 12359
rect 264069 12325 264103 12359
rect 271705 12325 271739 12359
rect 27721 12257 27755 12291
rect 28733 12257 28767 12291
rect 28917 12257 28951 12291
rect 29561 12257 29595 12291
rect 31769 12257 31803 12291
rect 40877 12257 40911 12291
rect 52377 12257 52411 12291
rect 55689 12257 55723 12291
rect 56701 12257 56735 12291
rect 76757 12257 76791 12291
rect 76941 12257 76975 12291
rect 78137 12257 78171 12291
rect 84485 12257 84519 12291
rect 84669 12257 84703 12291
rect 87061 12257 87095 12291
rect 88165 12257 88199 12291
rect 100953 12257 100987 12291
rect 103161 12257 103195 12291
rect 104541 12257 104575 12291
rect 114385 12257 114419 12291
rect 117789 12257 117823 12291
rect 131865 12257 131899 12291
rect 152105 12257 152139 12291
rect 152197 12257 152231 12291
rect 153945 12257 153979 12291
rect 161305 12257 161339 12291
rect 161489 12257 161523 12291
rect 162501 12257 162535 12291
rect 162685 12257 162719 12291
rect 163605 12257 163639 12291
rect 177037 12257 177071 12291
rect 177129 12257 177163 12291
rect 190837 12257 190871 12291
rect 193689 12257 193723 12291
rect 197553 12257 197587 12291
rect 203533 12257 203567 12291
rect 204729 12257 204763 12291
rect 231593 12257 231627 12291
rect 239321 12257 239355 12291
rect 241437 12257 241471 12291
rect 242817 12257 242851 12291
rect 242909 12257 242943 12291
rect 252569 12257 252603 12291
rect 255329 12257 255363 12291
rect 265725 12257 265759 12291
rect 265909 12257 265943 12291
rect 268761 12257 268795 12291
rect 272257 12257 272291 12291
rect 27445 12189 27479 12223
rect 28641 12189 28675 12223
rect 34161 12189 34195 12223
rect 34713 12189 34747 12223
rect 35357 12189 35391 12223
rect 36369 12189 36403 12223
rect 37105 12189 37139 12223
rect 38669 12189 38703 12223
rect 39129 12189 39163 12223
rect 40601 12189 40635 12223
rect 41429 12189 41463 12223
rect 43729 12189 43763 12223
rect 54585 12189 54619 12223
rect 56609 12189 56643 12223
rect 57529 12189 57563 12223
rect 58173 12189 58207 12223
rect 75377 12189 75411 12223
rect 76665 12189 76699 12223
rect 77953 12189 77987 12223
rect 79241 12189 79275 12223
rect 80161 12189 80195 12223
rect 84393 12189 84427 12223
rect 85497 12189 85531 12223
rect 86877 12189 86911 12223
rect 87981 12189 88015 12223
rect 88809 12189 88843 12223
rect 89637 12189 89671 12223
rect 90097 12189 90131 12223
rect 99297 12189 99331 12223
rect 99757 12189 99791 12223
rect 102977 12189 103011 12223
rect 103805 12189 103839 12223
rect 104449 12189 104483 12223
rect 105093 12189 105127 12223
rect 113281 12189 113315 12223
rect 113925 12189 113959 12223
rect 117605 12189 117639 12223
rect 118341 12189 118375 12223
rect 127909 12189 127943 12223
rect 128645 12189 128679 12223
rect 129105 12189 129139 12223
rect 131681 12189 131715 12223
rect 132601 12189 132635 12223
rect 137753 12189 137787 12223
rect 147505 12189 147539 12223
rect 148333 12189 148367 12223
rect 149437 12189 149471 12223
rect 152473 12189 152507 12223
rect 154313 12189 154347 12223
rect 160201 12189 160235 12223
rect 161213 12189 161247 12223
rect 176117 12189 176151 12223
rect 176945 12189 176979 12223
rect 179153 12189 179187 12223
rect 181545 12189 181579 12223
rect 188721 12189 188755 12223
rect 189549 12189 189583 12223
rect 190377 12189 190411 12223
rect 194425 12189 194459 12223
rect 196449 12189 196483 12223
rect 196725 12189 196759 12223
rect 197461 12189 197495 12223
rect 201049 12189 201083 12223
rect 201877 12189 201911 12223
rect 203257 12189 203291 12223
rect 227545 12189 227579 12223
rect 229937 12189 229971 12223
rect 232145 12189 232179 12223
rect 238033 12189 238067 12223
rect 239137 12189 239171 12223
rect 239229 12189 239263 12223
rect 240149 12189 240183 12223
rect 241253 12189 241287 12223
rect 243737 12189 243771 12223
rect 244381 12189 244415 12223
rect 251281 12189 251315 12223
rect 251925 12189 251959 12223
rect 255145 12189 255179 12223
rect 256249 12189 256283 12223
rect 257077 12189 257111 12223
rect 262689 12189 262723 12223
rect 263977 12189 264011 12223
rect 264805 12189 264839 12223
rect 266553 12189 266587 12223
rect 270969 12189 271003 12223
rect 272073 12189 272107 12223
rect 29837 12121 29871 12155
rect 32045 12121 32079 12155
rect 35449 12121 35483 12155
rect 41705 12121 41739 12155
rect 52653 12121 52687 12155
rect 55505 12121 55539 12155
rect 100769 12121 100803 12155
rect 100861 12121 100895 12155
rect 101965 12121 101999 12155
rect 102149 12121 102183 12155
rect 114661 12121 114695 12155
rect 117513 12121 117547 12155
rect 129381 12121 129415 12155
rect 138029 12121 138063 12155
rect 145849 12121 145883 12155
rect 146217 12121 146251 12155
rect 153669 12121 153703 12155
rect 163881 12121 163915 12155
rect 165905 12121 165939 12155
rect 177957 12121 177991 12155
rect 179429 12121 179463 12155
rect 191113 12121 191147 12155
rect 193413 12121 193447 12155
rect 194701 12121 194735 12155
rect 205005 12121 205039 12155
rect 249073 12121 249107 12155
rect 249257 12121 249291 12155
rect 252845 12121 252879 12155
rect 265633 12121 265667 12155
rect 266829 12121 266863 12155
rect 269037 12121 269071 12155
rect 27077 12053 27111 12087
rect 27537 12053 27571 12087
rect 28273 12053 28307 12087
rect 33517 12053 33551 12087
rect 36461 12053 36495 12087
rect 40233 12053 40267 12087
rect 40693 12053 40727 12087
rect 56057 12053 56091 12087
rect 56149 12053 56183 12087
rect 56517 12053 56551 12087
rect 76297 12053 76331 12087
rect 77861 12053 77895 12087
rect 84025 12053 84059 12087
rect 86785 12053 86819 12087
rect 87613 12053 87647 12087
rect 88073 12053 88107 12087
rect 100401 12053 100435 12087
rect 102609 12053 102643 12087
rect 103069 12053 103103 12087
rect 116133 12053 116167 12087
rect 117145 12053 117179 12087
rect 128461 12053 128495 12087
rect 131313 12053 131347 12087
rect 131773 12053 131807 12087
rect 150725 12053 150759 12087
rect 151645 12053 151679 12087
rect 152013 12053 152047 12087
rect 153761 12053 153795 12087
rect 160845 12053 160879 12087
rect 162041 12053 162075 12087
rect 162409 12053 162443 12087
rect 176577 12053 176611 12087
rect 178049 12053 178083 12087
rect 189641 12053 189675 12087
rect 193045 12053 193079 12087
rect 193505 12053 193539 12087
rect 196817 12053 196851 12087
rect 197001 12053 197035 12087
rect 197369 12053 197403 12087
rect 202889 12053 202923 12087
rect 203349 12053 203383 12087
rect 229293 12053 229327 12087
rect 230949 12053 230983 12087
rect 231317 12053 231351 12087
rect 231409 12053 231443 12087
rect 238217 12053 238251 12087
rect 240885 12053 240919 12087
rect 241345 12053 241379 12087
rect 242725 12053 242759 12087
rect 254777 12053 254811 12087
rect 255237 12053 255271 12087
rect 265265 12053 265299 12087
rect 268301 12053 268335 12087
rect 270509 12053 270543 12087
rect 272165 12053 272199 12087
rect 27813 11849 27847 11883
rect 32597 11849 32631 11883
rect 33793 11849 33827 11883
rect 34437 11849 34471 11883
rect 34989 11849 35023 11883
rect 38393 11849 38427 11883
rect 39037 11849 39071 11883
rect 39681 11849 39715 11883
rect 40141 11849 40175 11883
rect 41153 11849 41187 11883
rect 41705 11849 41739 11883
rect 52837 11849 52871 11883
rect 53665 11849 53699 11883
rect 54401 11849 54435 11883
rect 55321 11849 55355 11883
rect 56517 11849 56551 11883
rect 57161 11849 57195 11883
rect 75561 11849 75595 11883
rect 76021 11849 76055 11883
rect 76941 11849 76975 11883
rect 77861 11849 77895 11883
rect 78505 11849 78539 11883
rect 84393 11849 84427 11883
rect 86049 11849 86083 11883
rect 87153 11849 87187 11883
rect 87889 11849 87923 11883
rect 88901 11849 88935 11883
rect 100217 11849 100251 11883
rect 100953 11849 100987 11883
rect 101873 11849 101907 11883
rect 113833 11849 113867 11883
rect 115029 11849 115063 11883
rect 116225 11849 116259 11883
rect 116961 11849 116995 11883
rect 117605 11849 117639 11883
rect 129381 11849 129415 11883
rect 130485 11849 130519 11883
rect 130945 11849 130979 11883
rect 132417 11849 132451 11883
rect 151093 11849 151127 11883
rect 152013 11849 152047 11883
rect 152749 11849 152783 11883
rect 162317 11849 162351 11883
rect 162961 11849 162995 11883
rect 163513 11849 163547 11883
rect 164249 11849 164283 11883
rect 164893 11849 164927 11883
rect 176485 11849 176519 11883
rect 177589 11849 177623 11883
rect 178049 11849 178083 11883
rect 179153 11849 179187 11883
rect 180073 11849 180107 11883
rect 190837 11849 190871 11883
rect 196265 11849 196299 11883
rect 202889 11849 202923 11883
rect 204085 11849 204119 11883
rect 205189 11849 205223 11883
rect 228281 11849 228315 11883
rect 229477 11849 229511 11883
rect 230397 11849 230431 11883
rect 231593 11849 231627 11883
rect 238769 11849 238803 11883
rect 240333 11849 240367 11883
rect 241069 11849 241103 11883
rect 241805 11849 241839 11883
rect 251833 11849 251867 11883
rect 254133 11849 254167 11883
rect 254961 11849 254995 11883
rect 255605 11849 255639 11883
rect 264989 11849 265023 11883
rect 267381 11849 267415 11883
rect 268209 11849 268243 11883
rect 271429 11849 271463 11883
rect 28825 11781 28859 11815
rect 40049 11781 40083 11815
rect 202337 11781 202371 11815
rect 203993 11781 204027 11815
rect 205281 11781 205315 11815
rect 228373 11781 228407 11815
rect 229569 11781 229603 11815
rect 238677 11781 238711 11815
rect 254041 11781 254075 11815
rect 264437 11781 264471 11815
rect 27997 11713 28031 11747
rect 29653 11713 29687 11747
rect 32505 11713 32539 11747
rect 33701 11713 33735 11747
rect 34345 11713 34379 11747
rect 35173 11713 35207 11747
rect 38577 11713 38611 11747
rect 39221 11713 39255 11747
rect 41061 11713 41095 11747
rect 41889 11713 41923 11747
rect 42901 11713 42935 11747
rect 53021 11713 53055 11747
rect 53849 11713 53883 11747
rect 54309 11713 54343 11747
rect 56425 11713 56459 11747
rect 57069 11713 57103 11747
rect 75929 11713 75963 11747
rect 77125 11713 77159 11747
rect 77769 11713 77803 11747
rect 78689 11713 78723 11747
rect 84577 11713 84611 11747
rect 85221 11713 85255 11747
rect 86141 11713 86175 11747
rect 86969 11713 87003 11747
rect 87797 11713 87831 11747
rect 88809 11713 88843 11747
rect 100401 11713 100435 11747
rect 100861 11713 100895 11747
rect 103161 11713 103195 11747
rect 114017 11713 114051 11747
rect 115121 11713 115155 11747
rect 116409 11713 116443 11747
rect 116869 11713 116903 11747
rect 117513 11713 117547 11747
rect 129289 11713 129323 11747
rect 130853 11713 130887 11747
rect 131681 11713 131715 11747
rect 132601 11713 132635 11747
rect 147781 11713 147815 11747
rect 151277 11713 151311 11747
rect 152197 11713 152231 11747
rect 152657 11713 152691 11747
rect 161121 11713 161155 11747
rect 161765 11713 161799 11747
rect 162225 11713 162259 11747
rect 162869 11713 162903 11747
rect 163697 11713 163731 11747
rect 164157 11713 164191 11747
rect 164801 11713 164835 11747
rect 176669 11713 176703 11747
rect 177957 11713 177991 11747
rect 179245 11713 179279 11747
rect 179981 11713 180015 11747
rect 189641 11713 189675 11747
rect 190101 11713 190135 11747
rect 190745 11713 190779 11747
rect 191849 11713 191883 11747
rect 194057 11713 194091 11747
rect 196449 11713 196483 11747
rect 202245 11713 202279 11747
rect 203073 11713 203107 11747
rect 230305 11713 230339 11747
rect 230949 11713 230983 11747
rect 231041 11713 231075 11747
rect 231777 11713 231811 11747
rect 240241 11713 240275 11747
rect 241253 11713 241287 11747
rect 241713 11713 241747 11747
rect 242541 11713 242575 11747
rect 252017 11713 252051 11747
rect 252385 11713 252419 11747
rect 252753 11713 252787 11747
rect 254869 11713 254903 11747
rect 255513 11713 255547 11747
rect 264345 11713 264379 11747
rect 265173 11713 265207 11747
rect 265633 11713 265667 11747
rect 269129 11713 269163 11747
rect 271337 11713 271371 11747
rect 28917 11645 28951 11679
rect 29101 11645 29135 11679
rect 29929 11645 29963 11679
rect 32689 11645 32723 11679
rect 40233 11645 40267 11679
rect 43085 11645 43119 11679
rect 55413 11645 55447 11679
rect 55597 11645 55631 11679
rect 76205 11645 76239 11679
rect 86325 11645 86359 11679
rect 101965 11645 101999 11679
rect 102057 11645 102091 11679
rect 115305 11645 115339 11679
rect 131037 11645 131071 11679
rect 148333 11645 148367 11679
rect 148609 11645 148643 11679
rect 178141 11645 178175 11679
rect 179337 11645 179371 11679
rect 192125 11645 192159 11679
rect 194333 11645 194367 11679
rect 195805 11645 195839 11679
rect 204269 11645 204303 11679
rect 205465 11645 205499 11679
rect 228465 11645 228499 11679
rect 229753 11645 229787 11679
rect 240425 11645 240459 11679
rect 254225 11645 254259 11679
rect 265909 11645 265943 11679
rect 268301 11645 268335 11679
rect 268393 11645 268427 11679
rect 269405 11645 269439 11679
rect 270877 11645 270911 11679
rect 43453 11577 43487 11611
rect 147597 11577 147631 11611
rect 160937 11577 160971 11611
rect 161581 11577 161615 11611
rect 178785 11577 178819 11611
rect 190193 11577 190227 11611
rect 227913 11577 227947 11611
rect 239873 11577 239907 11611
rect 252937 11577 252971 11611
rect 28457 11509 28491 11543
rect 31401 11509 31435 11543
rect 32137 11509 32171 11543
rect 54953 11509 54987 11543
rect 85037 11509 85071 11543
rect 85681 11509 85715 11543
rect 101505 11509 101539 11543
rect 102977 11509 103011 11543
rect 114661 11509 114695 11543
rect 131865 11509 131899 11543
rect 150081 11509 150115 11543
rect 189457 11509 189491 11543
rect 193597 11509 193631 11543
rect 203625 11509 203659 11543
rect 204821 11509 204855 11543
rect 229109 11509 229143 11543
rect 242357 11509 242391 11543
rect 253673 11509 253707 11543
rect 267841 11509 267875 11543
rect 28825 11305 28859 11339
rect 33609 11305 33643 11339
rect 40325 11305 40359 11339
rect 41061 11305 41095 11339
rect 41613 11305 41647 11339
rect 55321 11305 55355 11339
rect 56241 11305 56275 11339
rect 76481 11305 76515 11339
rect 78229 11305 78263 11339
rect 86233 11305 86267 11339
rect 86969 11305 87003 11339
rect 88257 11305 88291 11339
rect 102885 11305 102919 11339
rect 116041 11305 116075 11339
rect 117145 11305 117179 11339
rect 130485 11305 130519 11339
rect 131221 11305 131255 11339
rect 131773 11305 131807 11339
rect 148057 11305 148091 11339
rect 150817 11305 150851 11339
rect 157349 11305 157383 11339
rect 162041 11305 162075 11339
rect 162685 11305 162719 11339
rect 163605 11305 163639 11339
rect 239965 11305 239999 11339
rect 240885 11305 240919 11339
rect 241437 11305 241471 11339
rect 242173 11305 242207 11339
rect 252569 11305 252603 11339
rect 253121 11305 253155 11339
rect 253765 11305 253799 11339
rect 265541 11305 265575 11339
rect 268025 11305 268059 11339
rect 42257 11237 42291 11271
rect 87613 11237 87647 11271
rect 103529 11237 103563 11271
rect 115397 11237 115431 11271
rect 149897 11237 149931 11271
rect 254409 11237 254443 11271
rect 266829 11237 266863 11271
rect 29653 11169 29687 11203
rect 32321 11169 32355 11203
rect 32505 11169 32539 11203
rect 102333 11169 102367 11203
rect 148517 11169 148551 11203
rect 148701 11169 148735 11203
rect 177589 11169 177623 11203
rect 178233 11169 178267 11203
rect 190285 11169 190319 11203
rect 192033 11169 192067 11203
rect 193781 11169 193815 11203
rect 194977 11169 195011 11203
rect 202889 11169 202923 11203
rect 264989 11169 265023 11203
rect 267473 11169 267507 11203
rect 268577 11169 268611 11203
rect 269405 11169 269439 11203
rect 270601 11169 270635 11203
rect 29009 11101 29043 11135
rect 32229 11101 32263 11135
rect 33517 11101 33551 11135
rect 40509 11101 40543 11135
rect 40969 11101 41003 11135
rect 41797 11101 41831 11135
rect 42441 11101 42475 11135
rect 55505 11101 55539 11135
rect 56425 11101 56459 11135
rect 76665 11101 76699 11135
rect 78413 11101 78447 11135
rect 86417 11101 86451 11135
rect 86877 11101 86911 11135
rect 87797 11101 87831 11135
rect 88441 11101 88475 11135
rect 102149 11101 102183 11135
rect 103069 11101 103103 11135
rect 103713 11101 103747 11135
rect 115305 11101 115339 11135
rect 116225 11101 116259 11135
rect 117329 11101 117363 11135
rect 130669 11101 130703 11135
rect 131129 11101 131163 11135
rect 131957 11101 131991 11135
rect 142077 11101 142111 11135
rect 151001 11101 151035 11135
rect 162225 11101 162259 11135
rect 162869 11101 162903 11135
rect 163513 11101 163547 11135
rect 177497 11101 177531 11135
rect 178141 11101 178175 11135
rect 179153 11101 179187 11135
rect 190193 11101 190227 11135
rect 190837 11101 190871 11135
rect 190929 11101 190963 11135
rect 194793 11101 194827 11135
rect 195805 11101 195839 11135
rect 202337 11101 202371 11135
rect 202797 11101 202831 11135
rect 203441 11101 203475 11135
rect 204913 11101 204947 11135
rect 229385 11101 229419 11135
rect 239873 11101 239907 11135
rect 240793 11101 240827 11135
rect 241621 11101 241655 11135
rect 242081 11101 242115 11135
rect 252477 11101 252511 11135
rect 253305 11101 253339 11135
rect 253949 11101 253983 11135
rect 254593 11101 254627 11135
rect 264897 11101 264931 11135
rect 265725 11101 265759 11135
rect 267197 11101 267231 11135
rect 268209 11101 268243 11135
rect 270417 11101 270451 11135
rect 270509 11101 270543 11135
rect 29929 11033 29963 11067
rect 140421 11033 140455 11067
rect 149621 11033 149655 11067
rect 156061 11033 156095 11067
rect 192309 11033 192343 11067
rect 267289 11033 267323 11067
rect 269221 11033 269255 11067
rect 269313 11033 269347 11067
rect 31401 10965 31435 10999
rect 31861 10965 31895 10999
rect 148425 10965 148459 10999
rect 178969 10965 179003 10999
rect 194425 10965 194459 10999
rect 194885 10965 194919 10999
rect 195621 10965 195655 10999
rect 202153 10965 202187 10999
rect 203533 10965 203567 10999
rect 204729 10965 204763 10999
rect 229201 10965 229235 10999
rect 268853 10965 268887 10999
rect 270049 10965 270083 10999
rect 29653 10761 29687 10795
rect 30665 10761 30699 10795
rect 30757 10761 30791 10795
rect 32137 10761 32171 10795
rect 32781 10761 32815 10795
rect 33425 10761 33459 10795
rect 101689 10761 101723 10795
rect 130485 10761 130519 10795
rect 141985 10761 142019 10795
rect 148885 10761 148919 10795
rect 150725 10761 150759 10795
rect 191849 10761 191883 10795
rect 194241 10761 194275 10795
rect 202889 10761 202923 10795
rect 253673 10761 253707 10795
rect 266553 10761 266587 10795
rect 267749 10761 267783 10795
rect 268393 10761 268427 10795
rect 140697 10693 140731 10727
rect 156153 10693 156187 10727
rect 193505 10693 193539 10727
rect 29837 10625 29871 10659
rect 32321 10625 32355 10659
rect 32965 10625 32999 10659
rect 33609 10625 33643 10659
rect 101873 10625 101907 10659
rect 130393 10625 130427 10659
rect 149069 10625 149103 10659
rect 150633 10625 150667 10659
rect 187249 10625 187283 10659
rect 191297 10625 191331 10659
rect 192033 10625 192067 10659
rect 192677 10625 192711 10659
rect 194149 10625 194183 10659
rect 203073 10625 203107 10659
rect 253857 10625 253891 10659
rect 266001 10625 266035 10659
rect 266461 10625 266495 10659
rect 267105 10625 267139 10659
rect 267933 10625 267967 10659
rect 268577 10625 268611 10659
rect 269129 10625 269163 10659
rect 269221 10625 269255 10659
rect 30849 10557 30883 10591
rect 187525 10557 187559 10591
rect 30297 10489 30331 10523
rect 191113 10489 191147 10523
rect 192861 10489 192895 10523
rect 193689 10489 193723 10523
rect 267197 10489 267231 10523
rect 157625 10421 157659 10455
rect 265817 10421 265851 10455
rect 30941 10217 30975 10251
rect 31677 10217 31711 10251
rect 32873 10217 32907 10251
rect 33609 10217 33643 10251
rect 191849 10217 191883 10251
rect 193137 10217 193171 10251
rect 267749 10217 267783 10251
rect 269037 10217 269071 10251
rect 30297 10149 30331 10183
rect 32321 10149 32355 10183
rect 267105 10149 267139 10183
rect 268485 10149 268519 10183
rect 157809 10081 157843 10115
rect 30481 10013 30515 10047
rect 31125 10013 31159 10047
rect 31585 10013 31619 10047
rect 32229 10013 32263 10047
rect 33057 10013 33091 10047
rect 33517 10013 33551 10047
rect 140421 10013 140455 10047
rect 156061 10013 156095 10047
rect 192033 10013 192067 10047
rect 192677 10013 192711 10047
rect 193321 10013 193355 10047
rect 267289 10013 267323 10047
rect 267933 10013 267967 10047
rect 268393 10013 268427 10047
rect 269221 10013 269255 10047
rect 304457 10013 304491 10047
rect 304825 9945 304859 9979
rect 141709 9877 141743 9911
rect 192493 9877 192527 9911
rect 32873 9605 32907 9639
rect 140697 9605 140731 9639
rect 156153 9605 156187 9639
rect 157901 9605 157935 9639
rect 193045 9605 193079 9639
rect 267933 9605 267967 9639
rect 31309 9537 31343 9571
rect 32137 9537 32171 9571
rect 32781 9537 32815 9571
rect 192493 9537 192527 9571
rect 192953 9537 192987 9571
rect 267841 9537 267875 9571
rect 32229 9469 32263 9503
rect 31125 9401 31159 9435
rect 192309 9401 192343 9435
rect 141985 9333 142019 9367
rect 1593 8449 1627 8483
rect 1409 8313 1443 8347
rect 1961 8313 1995 8347
rect 2329 8313 2363 8347
rect 2697 8313 2731 8347
rect 3065 8313 3099 8347
rect 303997 6273 304031 6307
rect 304273 6205 304307 6239
<< metal1 >>
rect 189902 13852 189908 13864
rect 72344 13824 75500 13852
rect 28994 13744 29000 13796
rect 29052 13784 29058 13796
rect 32950 13784 32956 13796
rect 29052 13756 32956 13784
rect 29052 13744 29058 13756
rect 32950 13744 32956 13756
rect 33008 13744 33014 13796
rect 46198 13744 46204 13796
rect 46256 13784 46262 13796
rect 63402 13784 63408 13796
rect 46256 13756 63408 13784
rect 46256 13744 46262 13756
rect 63402 13744 63408 13756
rect 63460 13744 63466 13796
rect 69290 13744 69296 13796
rect 69348 13784 69354 13796
rect 72344 13784 72372 13824
rect 75362 13784 75368 13796
rect 69348 13756 72372 13784
rect 72436 13756 75368 13784
rect 69348 13744 69354 13756
rect 72436 13728 72464 13756
rect 75362 13744 75368 13756
rect 75420 13744 75426 13796
rect 75472 13784 75500 13824
rect 189276 13824 189908 13852
rect 76006 13784 76012 13796
rect 75472 13756 76012 13784
rect 76006 13744 76012 13756
rect 76064 13744 76070 13796
rect 90634 13744 90640 13796
rect 90692 13784 90698 13796
rect 102410 13784 102416 13796
rect 90692 13756 102416 13784
rect 90692 13744 90698 13756
rect 102410 13744 102416 13756
rect 102468 13744 102474 13796
rect 113818 13744 113824 13796
rect 113876 13784 113882 13796
rect 125502 13784 125508 13796
rect 113876 13756 125508 13784
rect 113876 13744 113882 13756
rect 125502 13744 125508 13756
rect 125560 13784 125566 13796
rect 131850 13784 131856 13796
rect 125560 13756 131856 13784
rect 125560 13744 125566 13756
rect 131850 13744 131856 13756
rect 131908 13744 131914 13796
rect 161658 13744 161664 13796
rect 161716 13784 161722 13796
rect 166074 13784 166080 13796
rect 161716 13756 166080 13784
rect 161716 13744 161722 13756
rect 166074 13744 166080 13756
rect 166132 13784 166138 13796
rect 167362 13784 167368 13796
rect 166132 13756 167368 13784
rect 166132 13744 166138 13756
rect 167362 13744 167368 13756
rect 167420 13744 167426 13796
rect 174170 13744 174176 13796
rect 174228 13784 174234 13796
rect 177758 13784 177764 13796
rect 174228 13756 177764 13784
rect 174228 13744 174234 13756
rect 177758 13744 177764 13756
rect 177816 13744 177822 13796
rect 181898 13744 181904 13796
rect 181956 13784 181962 13796
rect 189276 13784 189304 13824
rect 189902 13812 189908 13824
rect 189960 13812 189966 13864
rect 181956 13756 189304 13784
rect 181956 13744 181962 13756
rect 189350 13744 189356 13796
rect 189408 13784 189414 13796
rect 193214 13784 193220 13796
rect 189408 13756 193220 13784
rect 189408 13744 189414 13756
rect 193214 13744 193220 13756
rect 193272 13744 193278 13796
rect 195974 13744 195980 13796
rect 196032 13784 196038 13796
rect 302786 13784 302792 13796
rect 196032 13756 302792 13784
rect 196032 13744 196038 13756
rect 302786 13744 302792 13756
rect 302844 13744 302850 13796
rect 27154 13676 27160 13728
rect 27212 13716 27218 13728
rect 36538 13716 36544 13728
rect 27212 13688 36544 13716
rect 27212 13676 27218 13688
rect 36538 13676 36544 13688
rect 36596 13676 36602 13728
rect 42518 13676 42524 13728
rect 42576 13716 42582 13728
rect 47854 13716 47860 13728
rect 42576 13688 47860 13716
rect 42576 13676 42582 13688
rect 47854 13676 47860 13688
rect 47912 13676 47918 13728
rect 51626 13676 51632 13728
rect 51684 13716 51690 13728
rect 54110 13716 54116 13728
rect 51684 13688 54116 13716
rect 51684 13676 51690 13688
rect 54110 13676 54116 13688
rect 54168 13676 54174 13728
rect 66162 13676 66168 13728
rect 66220 13716 66226 13728
rect 72418 13716 72424 13728
rect 66220 13688 72424 13716
rect 66220 13676 66226 13688
rect 72418 13676 72424 13688
rect 72476 13676 72482 13728
rect 73890 13676 73896 13728
rect 73948 13716 73954 13728
rect 76374 13716 76380 13728
rect 73948 13688 76380 13716
rect 73948 13676 73954 13688
rect 76374 13676 76380 13688
rect 76432 13676 76438 13728
rect 83090 13676 83096 13728
rect 83148 13716 83154 13728
rect 86402 13716 86408 13728
rect 83148 13688 86408 13716
rect 83148 13676 83154 13688
rect 86402 13676 86408 13688
rect 86460 13676 86466 13728
rect 91830 13676 91836 13728
rect 91888 13716 91894 13728
rect 101950 13716 101956 13728
rect 91888 13688 101956 13716
rect 91888 13676 91894 13688
rect 101950 13676 101956 13688
rect 102008 13676 102014 13728
rect 114646 13676 114652 13728
rect 114704 13716 114710 13728
rect 127434 13716 127440 13728
rect 114704 13688 127440 13716
rect 114704 13676 114710 13688
rect 127434 13676 127440 13688
rect 127492 13676 127498 13728
rect 127526 13676 127532 13728
rect 127584 13716 127590 13728
rect 129734 13716 129740 13728
rect 127584 13688 129740 13716
rect 127584 13676 127590 13688
rect 129734 13676 129740 13688
rect 129792 13676 129798 13728
rect 133598 13676 133604 13728
rect 133656 13716 133662 13728
rect 136818 13716 136824 13728
rect 133656 13688 136824 13716
rect 133656 13676 133662 13688
rect 136818 13676 136824 13688
rect 136876 13676 136882 13728
rect 148134 13676 148140 13728
rect 148192 13716 148198 13728
rect 150434 13716 150440 13728
rect 148192 13688 150440 13716
rect 148192 13676 148198 13688
rect 150434 13676 150440 13688
rect 150492 13676 150498 13728
rect 157150 13676 157156 13728
rect 157208 13716 157214 13728
rect 301406 13716 301412 13728
rect 157208 13688 301412 13716
rect 157208 13676 157214 13688
rect 301406 13676 301412 13688
rect 301464 13676 301470 13728
rect 1104 13626 305808 13648
rect 1104 13574 39049 13626
rect 39101 13574 39113 13626
rect 39165 13574 39177 13626
rect 39229 13574 39241 13626
rect 39293 13574 39305 13626
rect 39357 13574 115247 13626
rect 115299 13574 115311 13626
rect 115363 13574 115375 13626
rect 115427 13574 115439 13626
rect 115491 13574 115503 13626
rect 115555 13574 191445 13626
rect 191497 13574 191509 13626
rect 191561 13574 191573 13626
rect 191625 13574 191637 13626
rect 191689 13574 191701 13626
rect 191753 13574 267643 13626
rect 267695 13574 267707 13626
rect 267759 13574 267771 13626
rect 267823 13574 267835 13626
rect 267887 13574 267899 13626
rect 267951 13574 305808 13626
rect 1104 13552 305808 13574
rect 1578 13512 1584 13524
rect 1539 13484 1584 13512
rect 1578 13472 1584 13484
rect 1636 13472 1642 13524
rect 4614 13512 4620 13524
rect 4575 13484 4620 13512
rect 4614 13472 4620 13484
rect 4672 13472 4678 13524
rect 7650 13512 7656 13524
rect 7611 13484 7656 13512
rect 7650 13472 7656 13484
rect 7708 13472 7714 13524
rect 10778 13512 10784 13524
rect 10739 13484 10784 13512
rect 10778 13472 10784 13484
rect 10836 13472 10842 13524
rect 13814 13472 13820 13524
rect 13872 13512 13878 13524
rect 14093 13515 14151 13521
rect 14093 13512 14105 13515
rect 13872 13484 14105 13512
rect 13872 13472 13878 13484
rect 14093 13481 14105 13484
rect 14139 13481 14151 13515
rect 16850 13512 16856 13524
rect 16811 13484 16856 13512
rect 14093 13475 14151 13481
rect 16850 13472 16856 13484
rect 16908 13472 16914 13524
rect 19978 13512 19984 13524
rect 19939 13484 19984 13512
rect 19978 13472 19984 13484
rect 20036 13472 20042 13524
rect 23014 13512 23020 13524
rect 22975 13484 23020 13512
rect 23014 13472 23020 13484
rect 23072 13472 23078 13524
rect 25685 13515 25743 13521
rect 25685 13481 25697 13515
rect 25731 13512 25743 13515
rect 27614 13512 27620 13524
rect 25731 13484 27620 13512
rect 25731 13481 25743 13484
rect 25685 13475 25743 13481
rect 27614 13472 27620 13484
rect 27672 13472 27678 13524
rect 27706 13472 27712 13524
rect 27764 13512 27770 13524
rect 28997 13515 29055 13521
rect 28997 13512 29009 13515
rect 27764 13484 29009 13512
rect 27764 13472 27770 13484
rect 28997 13481 29009 13484
rect 29043 13481 29055 13515
rect 28997 13475 29055 13481
rect 30466 13472 30472 13524
rect 30524 13512 30530 13524
rect 31573 13515 31631 13521
rect 31573 13512 31585 13515
rect 30524 13484 31585 13512
rect 30524 13472 30530 13484
rect 31573 13481 31585 13484
rect 31619 13481 31631 13515
rect 31573 13475 31631 13481
rect 36538 13472 36544 13524
rect 36596 13512 36602 13524
rect 46198 13512 46204 13524
rect 36596 13484 46204 13512
rect 36596 13472 36602 13484
rect 46198 13472 46204 13484
rect 46256 13472 46262 13524
rect 47578 13512 47584 13524
rect 47539 13484 47584 13512
rect 47578 13472 47584 13484
rect 47636 13472 47642 13524
rect 50341 13515 50399 13521
rect 50341 13481 50353 13515
rect 50387 13512 50399 13515
rect 50522 13512 50528 13524
rect 50387 13484 50528 13512
rect 50387 13481 50399 13484
rect 50341 13475 50399 13481
rect 50522 13472 50528 13484
rect 50580 13472 50586 13524
rect 50985 13515 51043 13521
rect 50985 13481 50997 13515
rect 51031 13512 51043 13515
rect 53006 13512 53012 13524
rect 51031 13484 53012 13512
rect 51031 13481 51043 13484
rect 50985 13475 51043 13481
rect 53006 13472 53012 13484
rect 53064 13472 53070 13524
rect 55582 13472 55588 13524
rect 55640 13512 55646 13524
rect 57882 13512 57888 13524
rect 55640 13484 57888 13512
rect 55640 13472 55646 13484
rect 57882 13472 57888 13484
rect 57940 13512 57946 13524
rect 61746 13512 61752 13524
rect 57940 13484 61752 13512
rect 57940 13472 57946 13484
rect 61746 13472 61752 13484
rect 61804 13472 61810 13524
rect 63402 13472 63408 13524
rect 63460 13512 63466 13524
rect 142890 13512 142896 13524
rect 63460 13484 142154 13512
rect 142851 13484 142896 13512
rect 63460 13472 63466 13484
rect 27154 13444 27160 13456
rect 6886 13416 27160 13444
rect 6886 13376 6914 13416
rect 27154 13404 27160 13416
rect 27212 13404 27218 13456
rect 44174 13404 44180 13456
rect 44232 13404 44238 13456
rect 44269 13447 44327 13453
rect 44269 13413 44281 13447
rect 44315 13413 44327 13447
rect 44269 13407 44327 13413
rect 26329 13379 26387 13385
rect 1780 13348 6914 13376
rect 10980 13348 26096 13376
rect 1780 13317 1808 13348
rect 1765 13311 1823 13317
rect 1765 13277 1777 13311
rect 1811 13277 1823 13311
rect 4798 13308 4804 13320
rect 4759 13280 4804 13308
rect 1765 13271 1823 13277
rect 4798 13268 4804 13280
rect 4856 13268 4862 13320
rect 10980 13317 11008 13348
rect 7837 13311 7895 13317
rect 7837 13277 7849 13311
rect 7883 13277 7895 13311
rect 7837 13271 7895 13277
rect 10965 13311 11023 13317
rect 10965 13277 10977 13311
rect 11011 13277 11023 13311
rect 14274 13308 14280 13320
rect 14235 13280 14280 13308
rect 10965 13271 11023 13277
rect 7852 13240 7880 13271
rect 14274 13268 14280 13280
rect 14332 13268 14338 13320
rect 17034 13308 17040 13320
rect 16995 13280 17040 13308
rect 17034 13268 17040 13280
rect 17092 13268 17098 13320
rect 20162 13308 20168 13320
rect 20123 13280 20168 13308
rect 20162 13268 20168 13280
rect 20220 13268 20226 13320
rect 23198 13308 23204 13320
rect 23159 13280 23204 13308
rect 23198 13268 23204 13280
rect 23256 13268 23262 13320
rect 26068 13317 26096 13348
rect 26329 13345 26341 13379
rect 26375 13376 26387 13379
rect 26970 13376 26976 13388
rect 26375 13348 26976 13376
rect 26375 13345 26387 13348
rect 26329 13339 26387 13345
rect 26970 13336 26976 13348
rect 27028 13336 27034 13388
rect 27249 13379 27307 13385
rect 27249 13345 27261 13379
rect 27295 13376 27307 13379
rect 34701 13379 34759 13385
rect 34701 13376 34713 13379
rect 27295 13348 34713 13376
rect 27295 13345 27307 13348
rect 27249 13339 27307 13345
rect 34701 13345 34713 13348
rect 34747 13376 34759 13379
rect 37553 13379 37611 13385
rect 34747 13348 37044 13376
rect 34747 13345 34759 13348
rect 34701 13339 34759 13345
rect 26053 13311 26111 13317
rect 26053 13277 26065 13311
rect 26099 13277 26111 13311
rect 29822 13308 29828 13320
rect 29783 13280 29828 13308
rect 26053 13271 26111 13277
rect 26068 13240 26096 13271
rect 29822 13268 29828 13280
rect 29880 13268 29886 13320
rect 32398 13308 32404 13320
rect 32359 13280 32404 13308
rect 32398 13268 32404 13280
rect 32456 13268 32462 13320
rect 33778 13268 33784 13320
rect 33836 13268 33842 13320
rect 37016 13308 37044 13348
rect 37553 13345 37565 13379
rect 37599 13376 37611 13379
rect 44192 13376 44220 13404
rect 37599 13348 44220 13376
rect 37599 13345 37611 13348
rect 37553 13339 37611 13345
rect 44284 13320 44312 13407
rect 44358 13404 44364 13456
rect 44416 13444 44422 13456
rect 44416 13416 51856 13444
rect 44416 13404 44422 13416
rect 45554 13336 45560 13388
rect 45612 13376 45618 13388
rect 51626 13376 51632 13388
rect 45612 13348 45657 13376
rect 51587 13348 51632 13376
rect 45612 13336 45618 13348
rect 51626 13336 51632 13348
rect 51684 13336 51690 13388
rect 51828 13376 51856 13416
rect 59814 13404 59820 13456
rect 59872 13444 59878 13456
rect 60461 13447 60519 13453
rect 60461 13444 60473 13447
rect 59872 13416 60473 13444
rect 59872 13404 59878 13416
rect 60461 13413 60473 13416
rect 60507 13413 60519 13447
rect 63034 13444 63040 13456
rect 62995 13416 63040 13444
rect 60461 13407 60519 13413
rect 63034 13404 63040 13416
rect 63092 13404 63098 13456
rect 75362 13444 75368 13456
rect 63144 13416 73660 13444
rect 75323 13416 75368 13444
rect 63144 13376 63172 13416
rect 72694 13376 72700 13388
rect 51828 13348 63172 13376
rect 64846 13348 69428 13376
rect 72655 13348 72700 13376
rect 37016 13280 37596 13308
rect 27522 13240 27528 13252
rect 7852 13212 22094 13240
rect 26068 13212 27384 13240
rect 27483 13212 27528 13240
rect 22066 13172 22094 13212
rect 26145 13175 26203 13181
rect 26145 13172 26157 13175
rect 22066 13144 26157 13172
rect 26145 13141 26157 13144
rect 26191 13172 26203 13175
rect 27246 13172 27252 13184
rect 26191 13144 27252 13172
rect 26191 13141 26203 13144
rect 26145 13135 26203 13141
rect 27246 13132 27252 13144
rect 27304 13132 27310 13184
rect 27356 13172 27384 13212
rect 27522 13200 27528 13212
rect 27580 13200 27586 13252
rect 30101 13243 30159 13249
rect 28750 13212 29224 13240
rect 27706 13172 27712 13184
rect 27356 13144 27712 13172
rect 27706 13132 27712 13144
rect 27764 13132 27770 13184
rect 29196 13172 29224 13212
rect 30101 13209 30113 13243
rect 30147 13240 30159 13243
rect 30190 13240 30196 13252
rect 30147 13212 30196 13240
rect 30147 13209 30159 13212
rect 30101 13203 30159 13209
rect 30190 13200 30196 13212
rect 30248 13200 30254 13252
rect 32674 13240 32680 13252
rect 31326 13212 31754 13240
rect 32635 13212 32680 13240
rect 30466 13172 30472 13184
rect 29196 13144 30472 13172
rect 30466 13132 30472 13144
rect 30524 13132 30530 13184
rect 31726 13172 31754 13212
rect 32674 13200 32680 13212
rect 32732 13200 32738 13252
rect 34514 13200 34520 13252
rect 34572 13240 34578 13252
rect 34977 13243 35035 13249
rect 34977 13240 34989 13243
rect 34572 13212 34989 13240
rect 34572 13200 34578 13212
rect 34977 13209 34989 13212
rect 35023 13209 35035 13243
rect 34977 13203 35035 13209
rect 35986 13200 35992 13252
rect 36044 13200 36050 13252
rect 33594 13172 33600 13184
rect 31726 13144 33600 13172
rect 33594 13132 33600 13144
rect 33652 13132 33658 13184
rect 34146 13172 34152 13184
rect 34107 13144 34152 13172
rect 34146 13132 34152 13144
rect 34204 13132 34210 13184
rect 34330 13132 34336 13184
rect 34388 13172 34394 13184
rect 36449 13175 36507 13181
rect 36449 13172 36461 13175
rect 34388 13144 36461 13172
rect 34388 13132 34394 13144
rect 36449 13141 36461 13144
rect 36495 13172 36507 13175
rect 37458 13172 37464 13184
rect 36495 13144 37464 13172
rect 36495 13141 36507 13144
rect 36449 13135 36507 13141
rect 37458 13132 37464 13144
rect 37516 13132 37522 13184
rect 37568 13172 37596 13280
rect 38930 13268 38936 13320
rect 38988 13268 38994 13320
rect 40129 13311 40187 13317
rect 40129 13308 40141 13311
rect 39132 13280 40141 13308
rect 37826 13240 37832 13252
rect 37787 13212 37832 13240
rect 37826 13200 37832 13212
rect 37884 13200 37890 13252
rect 39132 13172 39160 13280
rect 40129 13277 40141 13280
rect 40175 13277 40187 13311
rect 42518 13308 42524 13320
rect 42479 13280 42524 13308
rect 40129 13271 40187 13277
rect 39298 13172 39304 13184
rect 37568 13144 39160 13172
rect 39259 13144 39304 13172
rect 39298 13132 39304 13144
rect 39356 13172 39362 13184
rect 39942 13172 39948 13184
rect 39356 13144 39948 13172
rect 39356 13132 39362 13144
rect 39942 13132 39948 13144
rect 40000 13132 40006 13184
rect 40144 13172 40172 13271
rect 42518 13268 42524 13280
rect 42576 13268 42582 13320
rect 44266 13268 44272 13320
rect 44324 13308 44330 13320
rect 47765 13311 47823 13317
rect 47765 13308 47777 13311
rect 44324 13280 47777 13308
rect 44324 13268 44330 13280
rect 47765 13277 47777 13280
rect 47811 13277 47823 13311
rect 47765 13271 47823 13277
rect 50525 13311 50583 13317
rect 50525 13277 50537 13311
rect 50571 13308 50583 13311
rect 51350 13308 51356 13320
rect 50571 13280 51356 13308
rect 50571 13277 50583 13280
rect 50525 13271 50583 13277
rect 40402 13240 40408 13252
rect 40363 13212 40408 13240
rect 40402 13200 40408 13212
rect 40460 13200 40466 13252
rect 41414 13200 41420 13252
rect 41472 13200 41478 13252
rect 42536 13240 42564 13268
rect 41800 13212 42564 13240
rect 42797 13243 42855 13249
rect 41800 13172 41828 13212
rect 42797 13209 42809 13243
rect 42843 13240 42855 13243
rect 42886 13240 42892 13252
rect 42843 13212 42892 13240
rect 42843 13209 42855 13212
rect 42797 13203 42855 13209
rect 42886 13200 42892 13212
rect 42944 13200 42950 13252
rect 43254 13200 43260 13252
rect 43312 13200 43318 13252
rect 45465 13243 45523 13249
rect 45465 13240 45477 13243
rect 44468 13212 45477 13240
rect 40144 13144 41828 13172
rect 41877 13175 41935 13181
rect 41877 13141 41889 13175
rect 41923 13172 41935 13175
rect 42426 13172 42432 13184
rect 41923 13144 42432 13172
rect 41923 13141 41935 13144
rect 41877 13135 41935 13141
rect 42426 13132 42432 13144
rect 42484 13172 42490 13184
rect 44468 13172 44496 13212
rect 45465 13209 45477 13212
rect 45511 13209 45523 13243
rect 45465 13203 45523 13209
rect 45002 13172 45008 13184
rect 42484 13144 44496 13172
rect 44963 13144 45008 13172
rect 42484 13132 42490 13144
rect 45002 13132 45008 13144
rect 45060 13132 45066 13184
rect 45370 13172 45376 13184
rect 45331 13144 45376 13172
rect 45370 13132 45376 13144
rect 45428 13132 45434 13184
rect 47780 13172 47808 13271
rect 51350 13268 51356 13280
rect 51408 13268 51414 13320
rect 53009 13311 53067 13317
rect 53009 13277 53021 13311
rect 53055 13277 53067 13311
rect 53009 13271 53067 13277
rect 47854 13200 47860 13252
rect 47912 13240 47918 13252
rect 53024 13240 53052 13271
rect 54386 13268 54392 13320
rect 54444 13268 54450 13320
rect 54754 13268 54760 13320
rect 54812 13308 54818 13320
rect 55582 13308 55588 13320
rect 54812 13280 55588 13308
rect 54812 13268 54818 13280
rect 55582 13268 55588 13280
rect 55640 13268 55646 13320
rect 57882 13308 57888 13320
rect 57843 13280 57888 13308
rect 57882 13268 57888 13280
rect 57940 13268 57946 13320
rect 60642 13308 60648 13320
rect 60603 13280 60648 13308
rect 60642 13268 60648 13280
rect 60700 13268 60706 13320
rect 63221 13311 63279 13317
rect 63221 13308 63233 13311
rect 61580 13280 63233 13308
rect 53282 13240 53288 13252
rect 47912 13212 53052 13240
rect 53243 13212 53288 13240
rect 47912 13200 47918 13212
rect 51445 13175 51503 13181
rect 51445 13172 51457 13175
rect 47780 13144 51457 13172
rect 51445 13141 51457 13144
rect 51491 13141 51503 13175
rect 53024 13172 53052 13212
rect 53282 13200 53288 13212
rect 53340 13200 53346 13252
rect 55858 13240 55864 13252
rect 54588 13212 54984 13240
rect 55819 13212 55864 13240
rect 54588 13172 54616 13212
rect 53024 13144 54616 13172
rect 51445 13135 51503 13141
rect 54662 13132 54668 13184
rect 54720 13172 54726 13184
rect 54757 13175 54815 13181
rect 54757 13172 54769 13175
rect 54720 13144 54769 13172
rect 54720 13132 54726 13144
rect 54757 13141 54769 13144
rect 54803 13141 54815 13175
rect 54956 13172 54984 13212
rect 55858 13200 55864 13212
rect 55916 13200 55922 13252
rect 56594 13200 56600 13252
rect 56652 13200 56658 13252
rect 57164 13212 57468 13240
rect 57164 13172 57192 13212
rect 57330 13172 57336 13184
rect 54956 13144 57192 13172
rect 57291 13144 57336 13172
rect 54757 13135 54815 13141
rect 57330 13132 57336 13144
rect 57388 13132 57394 13184
rect 57440 13172 57468 13212
rect 57698 13200 57704 13252
rect 57756 13240 57762 13252
rect 58161 13243 58219 13249
rect 58161 13240 58173 13243
rect 57756 13212 58173 13240
rect 57756 13200 57762 13212
rect 58161 13209 58173 13212
rect 58207 13209 58219 13243
rect 58161 13203 58219 13209
rect 58618 13200 58624 13252
rect 58676 13200 58682 13252
rect 61470 13240 61476 13252
rect 59464 13212 61476 13240
rect 59464 13172 59492 13212
rect 61470 13200 61476 13212
rect 61528 13200 61534 13252
rect 59630 13172 59636 13184
rect 57440 13144 59492 13172
rect 59591 13144 59636 13172
rect 59630 13132 59636 13144
rect 59688 13172 59694 13184
rect 61580 13172 61608 13280
rect 63221 13277 63233 13280
rect 63267 13308 63279 13311
rect 64846 13308 64874 13348
rect 66162 13308 66168 13320
rect 63267 13304 63356 13308
rect 63420 13304 64874 13308
rect 63267 13280 64874 13304
rect 66123 13280 66168 13308
rect 63267 13277 63279 13280
rect 63221 13271 63279 13277
rect 63328 13276 63448 13280
rect 66162 13268 66168 13280
rect 66220 13268 66226 13320
rect 69290 13308 69296 13320
rect 69251 13280 69296 13308
rect 69290 13268 69296 13280
rect 69348 13268 69354 13320
rect 69400 13308 69428 13348
rect 72694 13336 72700 13348
rect 72752 13336 72758 13388
rect 73632 13385 73660 13416
rect 75362 13404 75368 13416
rect 75420 13444 75426 13456
rect 75638 13444 75644 13456
rect 75420 13416 75644 13444
rect 75420 13404 75426 13416
rect 75638 13404 75644 13416
rect 75696 13404 75702 13456
rect 80026 13416 82492 13444
rect 73617 13379 73675 13385
rect 73617 13345 73629 13379
rect 73663 13376 73675 13379
rect 78493 13379 78551 13385
rect 78493 13376 78505 13379
rect 73663 13348 78505 13376
rect 73663 13345 73675 13348
rect 73617 13339 73675 13345
rect 78493 13345 78505 13348
rect 78539 13376 78551 13379
rect 80026 13376 80054 13416
rect 80238 13376 80244 13388
rect 78539 13348 80054 13376
rect 80151 13348 80244 13376
rect 78539 13345 78551 13348
rect 78493 13339 78551 13345
rect 80238 13336 80244 13348
rect 80296 13376 80302 13388
rect 81529 13379 81587 13385
rect 81529 13376 81541 13379
rect 80296 13348 81541 13376
rect 80296 13336 80302 13348
rect 81529 13345 81541 13348
rect 81575 13345 81587 13379
rect 81529 13339 81587 13345
rect 81618 13336 81624 13388
rect 81676 13376 81682 13388
rect 82464 13376 82492 13416
rect 93854 13404 93860 13456
rect 93912 13444 93918 13456
rect 93949 13447 94007 13453
rect 93949 13444 93961 13447
rect 93912 13416 93961 13444
rect 93912 13404 93918 13416
rect 93949 13413 93961 13416
rect 93995 13413 94007 13447
rect 93949 13407 94007 13413
rect 94516 13416 99374 13444
rect 94516 13376 94544 13416
rect 97997 13379 98055 13385
rect 97997 13376 98009 13379
rect 81676 13348 81721 13376
rect 82464 13348 94544 13376
rect 94608 13348 98009 13376
rect 81676 13336 81682 13348
rect 72513 13311 72571 13317
rect 72513 13308 72525 13311
rect 69400 13280 72525 13308
rect 72513 13277 72525 13280
rect 72559 13277 72571 13311
rect 72513 13271 72571 13277
rect 76193 13311 76251 13317
rect 76193 13277 76205 13311
rect 76239 13277 76251 13311
rect 78398 13308 78404 13320
rect 77602 13280 78404 13308
rect 76193 13271 76251 13277
rect 61746 13200 61752 13252
rect 61804 13240 61810 13252
rect 61804 13212 73844 13240
rect 61804 13200 61810 13212
rect 59688 13144 61608 13172
rect 59688 13132 59694 13144
rect 61654 13132 61660 13184
rect 61712 13172 61718 13184
rect 65886 13172 65892 13184
rect 61712 13144 65892 13172
rect 61712 13132 61718 13144
rect 65886 13132 65892 13144
rect 65944 13132 65950 13184
rect 65978 13132 65984 13184
rect 66036 13172 66042 13184
rect 69106 13172 69112 13184
rect 66036 13144 66081 13172
rect 69067 13144 69112 13172
rect 66036 13132 66042 13144
rect 69106 13132 69112 13144
rect 69164 13132 69170 13184
rect 72053 13175 72111 13181
rect 72053 13141 72065 13175
rect 72099 13172 72111 13175
rect 72326 13172 72332 13184
rect 72099 13144 72332 13172
rect 72099 13141 72111 13144
rect 72053 13135 72111 13141
rect 72326 13132 72332 13144
rect 72384 13132 72390 13184
rect 72418 13132 72424 13184
rect 72476 13172 72482 13184
rect 73816 13172 73844 13212
rect 73890 13200 73896 13252
rect 73948 13240 73954 13252
rect 75178 13240 75184 13252
rect 73948 13212 73993 13240
rect 75118 13212 75184 13240
rect 73948 13200 73954 13212
rect 75178 13200 75184 13212
rect 75236 13200 75242 13252
rect 76208 13172 76236 13271
rect 78398 13268 78404 13280
rect 78456 13268 78462 13320
rect 81434 13268 81440 13320
rect 81492 13268 81498 13320
rect 82449 13311 82507 13317
rect 82449 13277 82461 13311
rect 82495 13277 82507 13311
rect 83090 13308 83096 13320
rect 83051 13280 83096 13308
rect 82449 13271 82507 13277
rect 76466 13240 76472 13252
rect 76427 13212 76472 13240
rect 76466 13200 76472 13212
rect 76524 13200 76530 13252
rect 78766 13240 78772 13252
rect 77864 13212 78168 13240
rect 78727 13212 78772 13240
rect 77864 13172 77892 13212
rect 72476 13144 72521 13172
rect 73816 13144 77892 13172
rect 72476 13132 72482 13144
rect 77938 13132 77944 13184
rect 77996 13172 78002 13184
rect 78140 13172 78168 13212
rect 78766 13200 78772 13212
rect 78824 13200 78830 13252
rect 79318 13200 79324 13252
rect 79376 13200 79382 13252
rect 80054 13200 80060 13252
rect 80112 13240 80118 13252
rect 81452 13240 81480 13268
rect 82464 13240 82492 13271
rect 83090 13268 83096 13280
rect 83148 13268 83154 13320
rect 83918 13308 83924 13320
rect 83879 13280 83924 13308
rect 83918 13268 83924 13280
rect 83976 13268 83982 13320
rect 86497 13311 86555 13317
rect 86497 13308 86509 13311
rect 85592 13280 86509 13308
rect 83826 13240 83832 13252
rect 80112 13212 81112 13240
rect 81452 13212 82308 13240
rect 82464 13212 83832 13240
rect 80112 13200 80118 13212
rect 80790 13172 80796 13184
rect 77996 13144 78041 13172
rect 78140 13144 80796 13172
rect 77996 13132 78002 13144
rect 80790 13132 80796 13144
rect 80848 13132 80854 13184
rect 81084 13181 81112 13212
rect 81069 13175 81127 13181
rect 81069 13141 81081 13175
rect 81115 13141 81127 13175
rect 81434 13172 81440 13184
rect 81395 13144 81440 13172
rect 81069 13135 81127 13141
rect 81434 13132 81440 13144
rect 81492 13132 81498 13184
rect 82280 13181 82308 13212
rect 83826 13200 83832 13212
rect 83884 13200 83890 13252
rect 84197 13243 84255 13249
rect 84197 13209 84209 13243
rect 84243 13240 84255 13243
rect 84470 13240 84476 13252
rect 84243 13212 84476 13240
rect 84243 13209 84255 13212
rect 84197 13203 84255 13209
rect 84470 13200 84476 13212
rect 84528 13200 84534 13252
rect 85482 13240 85488 13252
rect 85422 13212 85488 13240
rect 85482 13200 85488 13212
rect 85540 13200 85546 13252
rect 82265 13175 82323 13181
rect 82265 13141 82277 13175
rect 82311 13141 82323 13175
rect 82906 13172 82912 13184
rect 82867 13144 82912 13172
rect 82265 13135 82323 13141
rect 82906 13132 82912 13144
rect 82964 13132 82970 13184
rect 83918 13132 83924 13184
rect 83976 13172 83982 13184
rect 85592 13172 85620 13280
rect 86497 13277 86509 13280
rect 86543 13277 86555 13311
rect 86497 13271 86555 13277
rect 83976 13144 85620 13172
rect 85669 13175 85727 13181
rect 83976 13132 83982 13144
rect 85669 13141 85681 13175
rect 85715 13172 85727 13175
rect 86034 13172 86040 13184
rect 85715 13144 86040 13172
rect 85715 13141 85727 13144
rect 85669 13135 85727 13141
rect 86034 13132 86040 13144
rect 86092 13132 86098 13184
rect 86512 13172 86540 13271
rect 87874 13268 87880 13320
rect 87932 13268 87938 13320
rect 88797 13311 88855 13317
rect 88797 13308 88809 13311
rect 88076 13280 88809 13308
rect 86770 13240 86776 13252
rect 86731 13212 86776 13240
rect 86770 13200 86776 13212
rect 86828 13200 86834 13252
rect 88076 13172 88104 13280
rect 88797 13277 88809 13280
rect 88843 13277 88855 13311
rect 94133 13311 94191 13317
rect 94133 13308 94145 13311
rect 88797 13271 88855 13277
rect 93136 13280 94145 13308
rect 88242 13172 88248 13184
rect 86512 13144 88104 13172
rect 88203 13144 88248 13172
rect 88242 13132 88248 13144
rect 88300 13132 88306 13184
rect 88812 13172 88840 13271
rect 89070 13240 89076 13252
rect 89031 13212 89076 13240
rect 89070 13200 89076 13212
rect 89128 13200 89134 13252
rect 89530 13200 89536 13252
rect 89588 13200 89594 13252
rect 91646 13240 91652 13252
rect 90468 13212 91652 13240
rect 90468 13172 90496 13212
rect 91646 13200 91652 13212
rect 91704 13200 91710 13252
rect 91830 13240 91836 13252
rect 91791 13212 91836 13240
rect 91830 13200 91836 13212
rect 91888 13200 91894 13252
rect 92014 13240 92020 13252
rect 91975 13212 92020 13240
rect 92014 13200 92020 13212
rect 92072 13200 92078 13252
rect 88812 13144 90496 13172
rect 90542 13132 90548 13184
rect 90600 13172 90606 13184
rect 93136 13172 93164 13280
rect 94133 13277 94145 13280
rect 94179 13308 94191 13311
rect 94608 13308 94636 13348
rect 97997 13345 98009 13348
rect 98043 13345 98055 13379
rect 97997 13339 98055 13345
rect 98181 13379 98239 13385
rect 98181 13345 98193 13379
rect 98227 13376 98239 13379
rect 99098 13376 99104 13388
rect 98227 13348 99104 13376
rect 98227 13345 98239 13348
rect 98181 13339 98239 13345
rect 99098 13336 99104 13348
rect 99156 13336 99162 13388
rect 99346 13376 99374 13416
rect 100754 13404 100760 13456
rect 100812 13444 100818 13456
rect 101125 13447 101183 13453
rect 101125 13444 101137 13447
rect 100812 13416 101137 13444
rect 100812 13404 100818 13416
rect 101125 13413 101137 13416
rect 101171 13413 101183 13447
rect 101125 13407 101183 13413
rect 109034 13404 109040 13456
rect 109092 13444 109098 13456
rect 109405 13447 109463 13453
rect 109405 13444 109417 13447
rect 109092 13416 109417 13444
rect 109092 13404 109098 13416
rect 109405 13413 109417 13416
rect 109451 13413 109463 13447
rect 109405 13407 109463 13413
rect 111245 13447 111303 13453
rect 111245 13413 111257 13447
rect 111291 13444 111303 13447
rect 111702 13444 111708 13456
rect 111291 13416 111708 13444
rect 111291 13413 111303 13416
rect 111245 13407 111303 13413
rect 111702 13404 111708 13416
rect 111760 13404 111766 13456
rect 118878 13404 118884 13456
rect 118936 13444 118942 13456
rect 121270 13444 121276 13456
rect 118936 13416 120304 13444
rect 121231 13416 121276 13444
rect 118936 13404 118942 13416
rect 112257 13379 112315 13385
rect 112257 13376 112269 13379
rect 99346 13348 112269 13376
rect 112257 13345 112269 13348
rect 112303 13376 112315 13379
rect 112303 13348 114876 13376
rect 112303 13345 112315 13348
rect 112257 13339 112315 13345
rect 114848 13320 114876 13348
rect 118234 13336 118240 13388
rect 118292 13376 118298 13388
rect 120276 13385 120304 13416
rect 121270 13404 121276 13416
rect 121328 13404 121334 13456
rect 124122 13444 124128 13456
rect 124083 13416 124128 13444
rect 124122 13404 124128 13416
rect 124180 13404 124186 13456
rect 127526 13444 127532 13456
rect 126716 13416 127532 13444
rect 126716 13385 126744 13416
rect 127526 13404 127532 13416
rect 127584 13404 127590 13456
rect 136634 13444 136640 13456
rect 136595 13416 136640 13444
rect 136634 13404 136640 13416
rect 136692 13404 136698 13456
rect 139578 13404 139584 13456
rect 139636 13444 139642 13456
rect 140317 13447 140375 13453
rect 140317 13444 140329 13447
rect 139636 13416 140329 13444
rect 139636 13404 139642 13416
rect 140317 13413 140329 13416
rect 140363 13413 140375 13447
rect 142126 13444 142154 13484
rect 142890 13472 142896 13484
rect 142948 13472 142954 13524
rect 144733 13515 144791 13521
rect 144733 13481 144745 13515
rect 144779 13512 144791 13515
rect 145742 13512 145748 13524
rect 144779 13484 145748 13512
rect 144779 13481 144791 13484
rect 144733 13475 144791 13481
rect 145742 13472 145748 13484
rect 145800 13472 145806 13524
rect 148134 13512 148140 13524
rect 145852 13484 148140 13512
rect 145852 13444 145880 13484
rect 148134 13472 148140 13484
rect 148192 13472 148198 13524
rect 148308 13515 148366 13521
rect 148308 13481 148320 13515
rect 148354 13512 148366 13515
rect 150802 13512 150808 13524
rect 148354 13484 150808 13512
rect 148354 13481 148366 13484
rect 148308 13475 148366 13481
rect 150802 13472 150808 13484
rect 150860 13472 150866 13524
rect 157242 13512 157248 13524
rect 152200 13484 157248 13512
rect 142126 13416 145880 13444
rect 140317 13407 140375 13413
rect 120261 13379 120319 13385
rect 118292 13348 120212 13376
rect 118292 13336 118298 13348
rect 94179 13280 94636 13308
rect 96893 13311 96951 13317
rect 94179 13277 94191 13280
rect 94133 13271 94191 13277
rect 96893 13277 96905 13311
rect 96939 13308 96951 13311
rect 99377 13311 99435 13317
rect 96939 13280 97948 13308
rect 96939 13277 96951 13280
rect 96893 13271 96951 13277
rect 96706 13172 96712 13184
rect 90600 13144 93164 13172
rect 96667 13144 96712 13172
rect 90600 13132 90606 13144
rect 96706 13132 96712 13144
rect 96764 13132 96770 13184
rect 97534 13172 97540 13184
rect 97495 13144 97540 13172
rect 97534 13132 97540 13144
rect 97592 13132 97598 13184
rect 97920 13181 97948 13280
rect 99377 13277 99389 13311
rect 99423 13277 99435 13311
rect 99377 13271 99435 13277
rect 97994 13200 98000 13252
rect 98052 13240 98058 13252
rect 99190 13240 99196 13252
rect 98052 13212 99196 13240
rect 98052 13200 98058 13212
rect 99190 13200 99196 13212
rect 99248 13240 99254 13252
rect 99392 13240 99420 13271
rect 101398 13268 101404 13320
rect 101456 13308 101462 13320
rect 101953 13311 102011 13317
rect 101953 13308 101965 13311
rect 101456 13280 101965 13308
rect 101456 13268 101462 13280
rect 101953 13277 101965 13280
rect 101999 13277 102011 13311
rect 101953 13271 102011 13277
rect 99650 13240 99656 13252
rect 99248 13212 99420 13240
rect 99611 13212 99656 13240
rect 99248 13200 99254 13212
rect 99650 13200 99656 13212
rect 99708 13200 99714 13252
rect 100938 13240 100944 13252
rect 100878 13212 100944 13240
rect 100938 13200 100944 13212
rect 100996 13200 101002 13252
rect 97905 13175 97963 13181
rect 97905 13141 97917 13175
rect 97951 13172 97963 13175
rect 101030 13172 101036 13184
rect 97951 13144 101036 13172
rect 97951 13141 97963 13144
rect 97905 13135 97963 13141
rect 101030 13132 101036 13144
rect 101088 13132 101094 13184
rect 101968 13172 101996 13271
rect 103330 13268 103336 13320
rect 103388 13268 103394 13320
rect 104250 13308 104256 13320
rect 103532 13280 104256 13308
rect 102226 13240 102232 13252
rect 102187 13212 102232 13240
rect 102226 13200 102232 13212
rect 102284 13200 102290 13252
rect 103532 13172 103560 13280
rect 104250 13268 104256 13280
rect 104308 13268 104314 13320
rect 109586 13308 109592 13320
rect 109547 13280 109592 13308
rect 109586 13268 109592 13280
rect 109644 13268 109650 13320
rect 111426 13308 111432 13320
rect 111387 13280 111432 13308
rect 111426 13268 111432 13280
rect 111484 13268 111490 13320
rect 114830 13308 114836 13320
rect 114791 13280 114836 13308
rect 114830 13268 114836 13280
rect 114888 13268 114894 13320
rect 117406 13308 117412 13320
rect 117367 13280 117412 13308
rect 117406 13268 117412 13280
rect 117464 13268 117470 13320
rect 118786 13268 118792 13320
rect 118844 13268 118850 13320
rect 120184 13317 120212 13348
rect 120261 13345 120273 13379
rect 120307 13345 120319 13379
rect 120261 13339 120319 13345
rect 125689 13379 125747 13385
rect 125689 13345 125701 13379
rect 125735 13376 125747 13379
rect 126701 13379 126759 13385
rect 126701 13376 126713 13379
rect 125735 13348 126713 13376
rect 125735 13345 125747 13348
rect 125689 13339 125747 13345
rect 126701 13345 126713 13348
rect 126747 13345 126759 13379
rect 130286 13376 130292 13388
rect 126701 13339 126759 13345
rect 127544 13348 130292 13376
rect 127544 13320 127572 13348
rect 130286 13336 130292 13348
rect 130344 13376 130350 13388
rect 132589 13379 132647 13385
rect 132589 13376 132601 13379
rect 130344 13348 132601 13376
rect 130344 13336 130350 13348
rect 132589 13345 132601 13348
rect 132635 13376 132647 13379
rect 142062 13376 142068 13388
rect 132635 13348 142068 13376
rect 132635 13345 132647 13348
rect 132589 13339 132647 13345
rect 142062 13336 142068 13348
rect 142120 13336 142126 13388
rect 148045 13379 148103 13385
rect 144932 13348 147674 13376
rect 120169 13311 120227 13317
rect 120169 13277 120181 13311
rect 120215 13308 120227 13311
rect 121457 13311 121515 13317
rect 121457 13308 121469 13311
rect 120215 13280 121469 13308
rect 120215 13277 120227 13280
rect 120169 13271 120227 13277
rect 121457 13277 121469 13280
rect 121503 13277 121515 13311
rect 124309 13311 124367 13317
rect 124309 13308 124321 13311
rect 121457 13271 121515 13277
rect 122806 13280 124321 13308
rect 104066 13200 104072 13252
rect 104124 13240 104130 13252
rect 104529 13243 104587 13249
rect 104529 13240 104541 13243
rect 104124 13212 104541 13240
rect 104124 13200 104130 13212
rect 104529 13209 104541 13212
rect 104575 13209 104587 13243
rect 104529 13203 104587 13209
rect 104986 13200 104992 13252
rect 105044 13200 105050 13252
rect 112530 13240 112536 13252
rect 112491 13212 112536 13240
rect 112530 13200 112536 13212
rect 112588 13200 112594 13252
rect 114186 13240 114192 13252
rect 113758 13212 114192 13240
rect 114186 13200 114192 13212
rect 114244 13200 114250 13252
rect 115106 13240 115112 13252
rect 115067 13212 115112 13240
rect 115106 13200 115112 13212
rect 115164 13200 115170 13252
rect 116946 13240 116952 13252
rect 116334 13212 116952 13240
rect 116946 13200 116952 13212
rect 117004 13200 117010 13252
rect 117682 13240 117688 13252
rect 117643 13212 117688 13240
rect 117682 13200 117688 13212
rect 117740 13200 117746 13252
rect 120077 13243 120135 13249
rect 120077 13240 120089 13243
rect 119172 13212 120089 13240
rect 101968 13144 103560 13172
rect 103698 13132 103704 13184
rect 103756 13172 103762 13184
rect 104434 13172 104440 13184
rect 103756 13144 104440 13172
rect 103756 13132 103762 13144
rect 104434 13132 104440 13144
rect 104492 13132 104498 13184
rect 104618 13132 104624 13184
rect 104676 13172 104682 13184
rect 106001 13175 106059 13181
rect 106001 13172 106013 13175
rect 104676 13144 106013 13172
rect 104676 13132 104682 13144
rect 106001 13141 106013 13144
rect 106047 13172 106059 13175
rect 109586 13172 109592 13184
rect 106047 13144 109592 13172
rect 106047 13141 106059 13144
rect 106001 13135 106059 13141
rect 109586 13132 109592 13144
rect 109644 13132 109650 13184
rect 114005 13175 114063 13181
rect 114005 13141 114017 13175
rect 114051 13172 114063 13175
rect 114554 13172 114560 13184
rect 114051 13144 114560 13172
rect 114051 13141 114063 13144
rect 114005 13135 114063 13141
rect 114554 13132 114560 13144
rect 114612 13172 114618 13184
rect 114922 13172 114928 13184
rect 114612 13144 114928 13172
rect 114612 13132 114618 13144
rect 114922 13132 114928 13144
rect 114980 13132 114986 13184
rect 115750 13132 115756 13184
rect 115808 13172 115814 13184
rect 116581 13175 116639 13181
rect 116581 13172 116593 13175
rect 115808 13144 116593 13172
rect 115808 13132 115814 13144
rect 116581 13141 116593 13144
rect 116627 13172 116639 13175
rect 118050 13172 118056 13184
rect 116627 13144 118056 13172
rect 116627 13141 116639 13144
rect 116581 13135 116639 13141
rect 118050 13132 118056 13144
rect 118108 13132 118114 13184
rect 119172 13181 119200 13212
rect 120077 13209 120089 13212
rect 120123 13240 120135 13243
rect 122806 13240 122834 13280
rect 124309 13277 124321 13280
rect 124355 13308 124367 13311
rect 126609 13311 126667 13317
rect 126609 13308 126621 13311
rect 124355 13280 126621 13308
rect 124355 13277 124367 13280
rect 124309 13271 124367 13277
rect 126609 13277 126621 13280
rect 126655 13277 126667 13311
rect 127526 13308 127532 13320
rect 127487 13280 127532 13308
rect 126609 13271 126667 13277
rect 127526 13268 127532 13280
rect 127584 13268 127590 13320
rect 129366 13308 129372 13320
rect 128938 13280 129372 13308
rect 129366 13268 129372 13280
rect 129424 13268 129430 13320
rect 136818 13308 136824 13320
rect 136779 13280 136824 13308
rect 136818 13268 136824 13280
rect 136876 13268 136882 13320
rect 140501 13311 140559 13317
rect 140501 13277 140513 13311
rect 140547 13277 140559 13311
rect 143074 13308 143080 13320
rect 143035 13280 143080 13308
rect 140501 13271 140559 13277
rect 125502 13240 125508 13252
rect 120123 13212 122834 13240
rect 125463 13212 125508 13240
rect 120123 13209 120135 13212
rect 120077 13203 120135 13209
rect 125502 13200 125508 13212
rect 125560 13200 125566 13252
rect 127802 13240 127808 13252
rect 127763 13212 127808 13240
rect 127802 13200 127808 13212
rect 127860 13200 127866 13252
rect 130565 13243 130623 13249
rect 130565 13240 130577 13243
rect 129108 13212 130577 13240
rect 119157 13175 119215 13181
rect 119157 13141 119169 13175
rect 119203 13141 119215 13175
rect 119706 13172 119712 13184
rect 119667 13144 119712 13172
rect 119157 13135 119215 13141
rect 119706 13132 119712 13144
rect 119764 13132 119770 13184
rect 126146 13172 126152 13184
rect 126107 13144 126152 13172
rect 126146 13132 126152 13144
rect 126204 13132 126210 13184
rect 126514 13172 126520 13184
rect 126475 13144 126520 13172
rect 126514 13132 126520 13144
rect 126572 13132 126578 13184
rect 128078 13132 128084 13184
rect 128136 13172 128142 13184
rect 129108 13172 129136 13212
rect 130565 13209 130577 13212
rect 130611 13209 130623 13243
rect 130565 13203 130623 13209
rect 131206 13200 131212 13252
rect 131264 13200 131270 13252
rect 132862 13240 132868 13252
rect 132823 13212 132868 13240
rect 132862 13200 132868 13212
rect 132920 13200 132926 13252
rect 133322 13200 133328 13252
rect 133380 13200 133386 13252
rect 140516 13240 140544 13271
rect 143074 13268 143080 13280
rect 143132 13268 143138 13320
rect 144932 13317 144960 13348
rect 144917 13311 144975 13317
rect 144917 13277 144929 13311
rect 144963 13277 144975 13311
rect 145742 13308 145748 13320
rect 145703 13280 145748 13308
rect 144917 13271 144975 13277
rect 145742 13268 145748 13280
rect 145800 13268 145806 13320
rect 147646 13308 147674 13348
rect 148045 13345 148057 13379
rect 148091 13376 148103 13379
rect 150897 13379 150955 13385
rect 150897 13376 150909 13379
rect 148091 13348 150909 13376
rect 148091 13345 148103 13348
rect 148045 13339 148103 13345
rect 150897 13345 150909 13348
rect 150943 13376 150955 13379
rect 152200 13376 152228 13484
rect 157242 13472 157248 13484
rect 157300 13472 157306 13524
rect 157613 13515 157671 13521
rect 157613 13481 157625 13515
rect 157659 13512 157671 13515
rect 157978 13512 157984 13524
rect 157659 13484 157984 13512
rect 157659 13481 157671 13484
rect 157613 13475 157671 13481
rect 157978 13472 157984 13484
rect 158036 13472 158042 13524
rect 159450 13472 159456 13524
rect 159508 13512 159514 13524
rect 161566 13512 161572 13524
rect 159508 13484 161572 13512
rect 159508 13472 159514 13484
rect 161566 13472 161572 13484
rect 161624 13512 161630 13524
rect 162670 13512 162676 13524
rect 161624 13484 162676 13512
rect 161624 13472 161630 13484
rect 162670 13472 162676 13484
rect 162728 13472 162734 13524
rect 163498 13472 163504 13524
rect 163556 13512 163562 13524
rect 176378 13512 176384 13524
rect 163556 13484 176384 13512
rect 163556 13472 163562 13484
rect 176378 13472 176384 13484
rect 176436 13472 176442 13524
rect 182726 13512 182732 13524
rect 176488 13484 182588 13512
rect 182687 13484 182732 13512
rect 154942 13404 154948 13456
rect 155000 13444 155006 13456
rect 155773 13447 155831 13453
rect 155773 13444 155785 13447
rect 155000 13416 155785 13444
rect 155000 13404 155006 13416
rect 155773 13413 155785 13416
rect 155819 13413 155831 13447
rect 155773 13407 155831 13413
rect 166442 13404 166448 13456
rect 166500 13444 166506 13456
rect 170398 13444 170404 13456
rect 166500 13416 170260 13444
rect 170359 13416 170404 13444
rect 166500 13404 166506 13416
rect 150943 13348 152228 13376
rect 153473 13379 153531 13385
rect 150943 13345 150955 13348
rect 150897 13339 150955 13345
rect 153473 13345 153485 13379
rect 153519 13376 153531 13379
rect 160922 13376 160928 13388
rect 153519 13348 158668 13376
rect 160835 13348 160928 13376
rect 153519 13345 153531 13348
rect 153473 13339 153531 13345
rect 158640 13320 158668 13348
rect 160922 13336 160928 13348
rect 160980 13376 160986 13388
rect 160980 13348 165108 13376
rect 160980 13336 160986 13348
rect 165080 13324 165108 13348
rect 165246 13336 165252 13388
rect 165304 13376 165310 13388
rect 166629 13379 166687 13385
rect 166629 13376 166641 13379
rect 165304 13348 166641 13376
rect 165304 13336 165310 13348
rect 166629 13345 166641 13348
rect 166675 13376 166687 13379
rect 167549 13379 167607 13385
rect 167549 13376 167561 13379
rect 166675 13348 167561 13376
rect 166675 13345 166687 13348
rect 166629 13339 166687 13345
rect 167549 13345 167561 13348
rect 167595 13345 167607 13379
rect 167549 13339 167607 13345
rect 147646 13280 148088 13308
rect 145926 13240 145932 13252
rect 134352 13212 145932 13240
rect 128136 13144 129136 13172
rect 128136 13132 128142 13144
rect 129182 13132 129188 13184
rect 129240 13172 129246 13184
rect 129277 13175 129335 13181
rect 129277 13172 129289 13175
rect 129240 13144 129289 13172
rect 129240 13132 129246 13144
rect 129277 13141 129289 13144
rect 129323 13141 129335 13175
rect 129277 13135 129335 13141
rect 131574 13132 131580 13184
rect 131632 13172 131638 13184
rect 132037 13175 132095 13181
rect 132037 13172 132049 13175
rect 131632 13144 132049 13172
rect 131632 13132 131638 13144
rect 132037 13141 132049 13144
rect 132083 13172 132095 13175
rect 133690 13172 133696 13184
rect 132083 13144 133696 13172
rect 132083 13141 132095 13144
rect 132037 13135 132095 13141
rect 133690 13132 133696 13144
rect 133748 13132 133754 13184
rect 134150 13132 134156 13184
rect 134208 13172 134214 13184
rect 134352 13181 134380 13212
rect 145926 13200 145932 13212
rect 145984 13200 145990 13252
rect 146018 13200 146024 13252
rect 146076 13240 146082 13252
rect 147582 13240 147588 13252
rect 146076 13212 146121 13240
rect 147246 13212 147588 13240
rect 146076 13200 146082 13212
rect 147582 13200 147588 13212
rect 147640 13200 147646 13252
rect 134337 13175 134395 13181
rect 134337 13172 134349 13175
rect 134208 13144 134349 13172
rect 134208 13132 134214 13144
rect 134337 13141 134349 13144
rect 134383 13141 134395 13175
rect 134337 13135 134395 13141
rect 145834 13132 145840 13184
rect 145892 13172 145898 13184
rect 147490 13172 147496 13184
rect 145892 13144 147496 13172
rect 145892 13132 145898 13144
rect 147490 13132 147496 13144
rect 147548 13132 147554 13184
rect 148060 13172 148088 13280
rect 155218 13268 155224 13320
rect 155276 13308 155282 13320
rect 155862 13308 155868 13320
rect 155276 13280 155868 13308
rect 155276 13268 155282 13280
rect 155862 13268 155868 13280
rect 155920 13308 155926 13320
rect 155957 13311 156015 13317
rect 155957 13308 155969 13311
rect 155920 13280 155969 13308
rect 155920 13268 155926 13280
rect 155957 13277 155969 13280
rect 156003 13277 156015 13311
rect 156414 13308 156420 13320
rect 156375 13280 156420 13308
rect 155957 13271 156015 13277
rect 156414 13268 156420 13280
rect 156472 13268 156478 13320
rect 157794 13308 157800 13320
rect 157755 13280 157800 13308
rect 157794 13268 157800 13280
rect 157852 13268 157858 13320
rect 158622 13308 158628 13320
rect 158583 13280 158628 13308
rect 158622 13268 158628 13280
rect 158680 13268 158686 13320
rect 162670 13268 162676 13320
rect 162728 13308 162734 13320
rect 163498 13308 163504 13320
rect 162728 13280 163360 13308
rect 163459 13280 163504 13308
rect 162728 13268 162734 13280
rect 150069 13243 150127 13249
rect 149546 13212 150020 13240
rect 149238 13172 149244 13184
rect 148060 13144 149244 13172
rect 149238 13132 149244 13144
rect 149296 13132 149302 13184
rect 149992 13172 150020 13212
rect 150069 13209 150081 13243
rect 150115 13240 150127 13243
rect 150434 13240 150440 13252
rect 150115 13212 150440 13240
rect 150115 13209 150127 13212
rect 150069 13203 150127 13209
rect 150434 13200 150440 13212
rect 150492 13200 150498 13252
rect 151078 13200 151084 13252
rect 151136 13240 151142 13252
rect 151173 13243 151231 13249
rect 151173 13240 151185 13243
rect 151136 13212 151185 13240
rect 151136 13200 151142 13212
rect 151173 13209 151185 13212
rect 151219 13209 151231 13243
rect 152458 13240 152464 13252
rect 152398 13212 152464 13240
rect 151173 13203 151231 13209
rect 152458 13200 152464 13212
rect 152516 13200 152522 13252
rect 153746 13240 153752 13252
rect 152568 13212 152872 13240
rect 153707 13212 153752 13240
rect 152568 13172 152596 13212
rect 149992 13144 152596 13172
rect 152642 13132 152648 13184
rect 152700 13172 152706 13184
rect 152844 13172 152872 13212
rect 153746 13200 153752 13212
rect 153804 13200 153810 13252
rect 154206 13200 154212 13252
rect 154264 13200 154270 13252
rect 156509 13243 156567 13249
rect 156509 13240 156521 13243
rect 155052 13212 156521 13240
rect 155052 13172 155080 13212
rect 156509 13209 156521 13212
rect 156555 13209 156567 13243
rect 156509 13203 156567 13209
rect 156598 13200 156604 13252
rect 156656 13240 156662 13252
rect 158898 13240 158904 13252
rect 156656 13212 157334 13240
rect 158859 13212 158904 13240
rect 156656 13200 156662 13212
rect 155218 13172 155224 13184
rect 152700 13144 152745 13172
rect 152844 13144 155080 13172
rect 155179 13144 155224 13172
rect 152700 13132 152706 13144
rect 155218 13132 155224 13144
rect 155276 13132 155282 13184
rect 157306 13172 157334 13212
rect 158898 13200 158904 13212
rect 158956 13200 158962 13252
rect 161198 13240 161204 13252
rect 160126 13212 160692 13240
rect 161159 13212 161204 13240
rect 159542 13172 159548 13184
rect 157306 13144 159548 13172
rect 159542 13132 159548 13144
rect 159600 13132 159606 13184
rect 160370 13172 160376 13184
rect 160331 13144 160376 13172
rect 160370 13132 160376 13144
rect 160428 13132 160434 13184
rect 160664 13172 160692 13212
rect 161198 13200 161204 13212
rect 161256 13200 161262 13252
rect 162762 13240 162768 13252
rect 162426 13212 162768 13240
rect 162762 13200 162768 13212
rect 162820 13200 162826 13252
rect 162026 13172 162032 13184
rect 160664 13144 162032 13172
rect 162026 13132 162032 13144
rect 162084 13132 162090 13184
rect 162486 13132 162492 13184
rect 162544 13172 162550 13184
rect 162673 13175 162731 13181
rect 162673 13172 162685 13175
rect 162544 13144 162685 13172
rect 162544 13132 162550 13144
rect 162673 13141 162685 13144
rect 162719 13141 162731 13175
rect 163332 13172 163360 13280
rect 163498 13268 163504 13280
rect 163556 13268 163562 13320
rect 164878 13268 164884 13320
rect 164936 13268 164942 13320
rect 165080 13308 165200 13324
rect 170232 13308 170260 13416
rect 170398 13404 170404 13416
rect 170456 13404 170462 13456
rect 173066 13444 173072 13456
rect 173027 13416 173072 13444
rect 173066 13404 173072 13416
rect 173124 13404 173130 13456
rect 173802 13444 173808 13456
rect 173763 13416 173808 13444
rect 173802 13404 173808 13416
rect 173860 13404 173866 13456
rect 175829 13447 175887 13453
rect 175829 13444 175841 13447
rect 174372 13416 175841 13444
rect 174372 13385 174400 13416
rect 175829 13413 175841 13416
rect 175875 13444 175887 13447
rect 175918 13444 175924 13456
rect 175875 13416 175924 13444
rect 175875 13413 175887 13416
rect 175829 13407 175887 13413
rect 175918 13404 175924 13416
rect 175976 13404 175982 13456
rect 176010 13404 176016 13456
rect 176068 13444 176074 13456
rect 176488 13444 176516 13484
rect 176068 13416 176516 13444
rect 176068 13404 176074 13416
rect 177758 13404 177764 13456
rect 177816 13444 177822 13456
rect 178129 13447 178187 13453
rect 178129 13444 178141 13447
rect 177816 13416 178141 13444
rect 177816 13404 177822 13416
rect 178129 13413 178141 13416
rect 178175 13413 178187 13447
rect 178129 13407 178187 13413
rect 180426 13404 180432 13456
rect 180484 13444 180490 13456
rect 181533 13447 181591 13453
rect 181533 13444 181545 13447
rect 180484 13416 181545 13444
rect 180484 13404 180490 13416
rect 181533 13413 181545 13416
rect 181579 13413 181591 13447
rect 181533 13407 181591 13413
rect 174265 13379 174323 13385
rect 174265 13376 174277 13379
rect 170600 13348 174277 13376
rect 170600 13317 170628 13348
rect 174265 13345 174277 13348
rect 174311 13345 174323 13379
rect 174265 13339 174323 13345
rect 174357 13379 174415 13385
rect 174357 13345 174369 13379
rect 174403 13345 174415 13379
rect 178957 13379 179015 13385
rect 178957 13376 178969 13379
rect 174357 13339 174415 13345
rect 174464 13348 175964 13376
rect 170585 13311 170643 13317
rect 170585 13308 170597 13311
rect 165080 13296 170168 13308
rect 165172 13280 170168 13296
rect 170232 13280 170597 13308
rect 163774 13240 163780 13252
rect 163735 13212 163780 13240
rect 163774 13200 163780 13212
rect 163832 13200 163838 13252
rect 165154 13240 165160 13252
rect 165080 13212 165160 13240
rect 164602 13172 164608 13184
rect 163332 13144 164608 13172
rect 162673 13135 162731 13141
rect 164602 13132 164608 13144
rect 164660 13172 164666 13184
rect 165080 13172 165108 13212
rect 165154 13200 165160 13212
rect 165212 13200 165218 13252
rect 166537 13243 166595 13249
rect 166537 13240 166549 13243
rect 165264 13212 166549 13240
rect 165264 13184 165292 13212
rect 166537 13209 166549 13212
rect 166583 13209 166595 13243
rect 167362 13240 167368 13252
rect 167275 13212 167368 13240
rect 166537 13203 166595 13209
rect 167362 13200 167368 13212
rect 167420 13200 167426 13252
rect 170140 13240 170168 13280
rect 170585 13277 170597 13280
rect 170631 13277 170643 13311
rect 170585 13271 170643 13277
rect 173253 13311 173311 13317
rect 173253 13277 173265 13311
rect 173299 13308 173311 13311
rect 174170 13308 174176 13320
rect 173299 13280 174176 13308
rect 173299 13277 173311 13280
rect 173253 13271 173311 13277
rect 174170 13268 174176 13280
rect 174228 13268 174234 13320
rect 174464 13240 174492 13348
rect 175645 13311 175703 13317
rect 175645 13308 175657 13311
rect 170140 13212 174492 13240
rect 174556 13280 175657 13308
rect 165246 13172 165252 13184
rect 164660 13144 165108 13172
rect 165207 13144 165252 13172
rect 164660 13132 164666 13144
rect 165246 13132 165252 13144
rect 165304 13132 165310 13184
rect 165338 13132 165344 13184
rect 165396 13172 165402 13184
rect 166077 13175 166135 13181
rect 166077 13172 166089 13175
rect 165396 13144 166089 13172
rect 165396 13132 165402 13144
rect 166077 13141 166089 13144
rect 166123 13141 166135 13175
rect 166442 13172 166448 13184
rect 166403 13144 166448 13172
rect 166077 13135 166135 13141
rect 166442 13132 166448 13144
rect 166500 13132 166506 13184
rect 167380 13172 167408 13200
rect 174556 13172 174584 13280
rect 175645 13277 175657 13280
rect 175691 13308 175703 13311
rect 175826 13308 175832 13320
rect 175691 13280 175832 13308
rect 175691 13277 175703 13280
rect 175645 13271 175703 13277
rect 175826 13268 175832 13280
rect 175884 13268 175890 13320
rect 175936 13304 175964 13348
rect 176120 13348 178969 13376
rect 176120 13304 176148 13348
rect 178957 13345 178969 13348
rect 179003 13376 179015 13379
rect 181898 13376 181904 13388
rect 179003 13348 181904 13376
rect 179003 13345 179015 13348
rect 178957 13339 179015 13345
rect 181898 13336 181904 13348
rect 181956 13336 181962 13388
rect 182082 13336 182088 13388
rect 182140 13376 182146 13388
rect 182560 13376 182588 13484
rect 182726 13472 182732 13484
rect 182784 13472 182790 13524
rect 185762 13512 185768 13524
rect 185723 13484 185768 13512
rect 185762 13472 185768 13484
rect 185820 13472 185826 13524
rect 189350 13512 189356 13524
rect 185872 13484 189356 13512
rect 185872 13376 185900 13484
rect 189350 13472 189356 13484
rect 189408 13472 189414 13524
rect 189460 13484 190868 13512
rect 188798 13404 188804 13456
rect 188856 13444 188862 13456
rect 189460 13444 189488 13484
rect 188856 13416 189488 13444
rect 188856 13404 188862 13416
rect 189534 13404 189540 13456
rect 189592 13444 189598 13456
rect 190840 13444 190868 13484
rect 190914 13472 190920 13524
rect 190972 13512 190978 13524
rect 193490 13512 193496 13524
rect 190972 13484 193496 13512
rect 190972 13472 190978 13484
rect 193490 13472 193496 13484
rect 193548 13472 193554 13524
rect 207106 13512 207112 13524
rect 197372 13484 207112 13512
rect 191834 13444 191840 13456
rect 189592 13416 189672 13444
rect 190840 13416 191840 13444
rect 189592 13404 189598 13416
rect 188522 13376 188528 13388
rect 182140 13348 182185 13376
rect 182560 13348 185900 13376
rect 185964 13348 187464 13376
rect 188483 13348 188528 13376
rect 182140 13336 182146 13348
rect 176378 13308 176384 13320
rect 175936 13276 176148 13304
rect 176339 13280 176384 13308
rect 176378 13268 176384 13280
rect 176436 13268 176442 13320
rect 180610 13268 180616 13320
rect 180668 13308 180674 13320
rect 185964 13317 185992 13348
rect 181993 13311 182051 13317
rect 181993 13308 182005 13311
rect 180668 13280 182005 13308
rect 180668 13268 180674 13280
rect 181993 13277 182005 13280
rect 182039 13308 182051 13311
rect 182913 13311 182971 13317
rect 182913 13308 182925 13311
rect 182039 13280 182925 13308
rect 182039 13277 182051 13280
rect 181993 13271 182051 13277
rect 182913 13277 182925 13280
rect 182959 13277 182971 13311
rect 182913 13271 182971 13277
rect 185949 13311 186007 13317
rect 185949 13277 185961 13311
rect 185995 13277 186007 13311
rect 185949 13271 186007 13277
rect 187329 13311 187387 13317
rect 187329 13277 187341 13311
rect 187375 13277 187387 13311
rect 187436 13308 187464 13348
rect 188522 13336 188528 13348
rect 188580 13336 188586 13388
rect 189644 13376 189672 13416
rect 191834 13404 191840 13416
rect 191892 13404 191898 13456
rect 197372 13444 197400 13484
rect 207106 13472 207112 13484
rect 207164 13472 207170 13524
rect 210326 13512 210332 13524
rect 207216 13484 207980 13512
rect 210287 13484 210332 13512
rect 195716 13416 197400 13444
rect 199841 13447 199899 13453
rect 189813 13379 189871 13385
rect 189813 13376 189825 13379
rect 189644 13348 189825 13376
rect 189813 13345 189825 13348
rect 189859 13345 189871 13379
rect 189813 13339 189871 13345
rect 189902 13336 189908 13388
rect 189960 13376 189966 13388
rect 195716 13376 195744 13416
rect 199841 13413 199853 13447
rect 199887 13444 199899 13447
rect 201954 13444 201960 13456
rect 199887 13416 201960 13444
rect 199887 13413 199899 13416
rect 199841 13407 199899 13413
rect 201954 13404 201960 13416
rect 202012 13404 202018 13456
rect 203426 13404 203432 13456
rect 203484 13444 203490 13456
rect 203889 13447 203947 13453
rect 203889 13444 203901 13447
rect 203484 13416 203901 13444
rect 203484 13404 203490 13416
rect 203889 13413 203901 13416
rect 203935 13413 203947 13447
rect 203889 13407 203947 13413
rect 206002 13404 206008 13456
rect 206060 13444 206066 13456
rect 207216 13444 207244 13484
rect 206060 13416 207244 13444
rect 206060 13404 206066 13416
rect 207750 13404 207756 13456
rect 207808 13444 207814 13456
rect 207808 13416 207888 13444
rect 207808 13404 207814 13416
rect 189960 13348 195744 13376
rect 189960 13336 189966 13348
rect 197630 13336 197636 13388
rect 197688 13376 197694 13388
rect 198737 13379 198795 13385
rect 198737 13376 198749 13379
rect 197688 13348 198749 13376
rect 197688 13336 197694 13348
rect 198737 13345 198749 13348
rect 198783 13345 198795 13379
rect 198737 13339 198795 13345
rect 201129 13379 201187 13385
rect 201129 13345 201141 13379
rect 201175 13376 201187 13379
rect 202046 13376 202052 13388
rect 201175 13348 202052 13376
rect 201175 13345 201187 13348
rect 201129 13339 201187 13345
rect 202046 13336 202052 13348
rect 202104 13336 202110 13388
rect 207860 13385 207888 13416
rect 204717 13379 204775 13385
rect 204717 13376 204729 13379
rect 202156 13348 204729 13376
rect 202156 13320 202184 13348
rect 204717 13345 204729 13348
rect 204763 13376 204775 13379
rect 207845 13379 207903 13385
rect 204763 13348 207796 13376
rect 204763 13345 204775 13348
rect 204717 13339 204775 13345
rect 188433 13311 188491 13317
rect 188433 13308 188445 13311
rect 187436 13280 188445 13308
rect 187329 13271 187387 13277
rect 188433 13277 188445 13280
rect 188479 13277 188491 13311
rect 189534 13308 189540 13320
rect 189495 13280 189540 13308
rect 188433 13271 188491 13277
rect 175734 13200 175740 13252
rect 175792 13240 175798 13252
rect 176657 13243 176715 13249
rect 176657 13240 176669 13243
rect 175792 13212 176669 13240
rect 175792 13200 175798 13212
rect 176657 13209 176669 13212
rect 176703 13209 176715 13243
rect 176657 13203 176715 13209
rect 177666 13200 177672 13252
rect 177724 13200 177730 13252
rect 179233 13243 179291 13249
rect 179233 13240 179245 13243
rect 177960 13212 179245 13240
rect 167380 13144 174584 13172
rect 174998 13132 175004 13184
rect 175056 13172 175062 13184
rect 177960 13172 177988 13212
rect 179233 13209 179245 13212
rect 179279 13209 179291 13243
rect 179233 13203 179291 13209
rect 179966 13200 179972 13252
rect 180024 13200 180030 13252
rect 180886 13200 180892 13252
rect 180944 13240 180950 13252
rect 181901 13243 181959 13249
rect 181901 13240 181913 13243
rect 180944 13212 181913 13240
rect 180944 13200 180950 13212
rect 181901 13209 181913 13212
rect 181947 13240 181959 13243
rect 185964 13240 185992 13271
rect 181947 13212 185992 13240
rect 181947 13209 181959 13212
rect 181901 13203 181959 13209
rect 180702 13172 180708 13184
rect 175056 13144 177988 13172
rect 180663 13144 180708 13172
rect 175056 13132 175062 13144
rect 180702 13132 180708 13144
rect 180760 13132 180766 13184
rect 187344 13172 187372 13271
rect 189534 13268 189540 13280
rect 189592 13268 189598 13320
rect 191837 13311 191895 13317
rect 191837 13277 191849 13311
rect 191883 13277 191895 13311
rect 191837 13271 191895 13277
rect 194413 13311 194471 13317
rect 194413 13277 194425 13311
rect 194459 13277 194471 13311
rect 194413 13271 194471 13277
rect 200025 13311 200083 13317
rect 200025 13277 200037 13311
rect 200071 13308 200083 13311
rect 201494 13308 201500 13320
rect 200071 13280 201500 13308
rect 200071 13277 200083 13280
rect 200025 13271 200083 13277
rect 187421 13243 187479 13249
rect 187421 13209 187433 13243
rect 187467 13240 187479 13243
rect 191852 13240 191880 13271
rect 187467 13212 190302 13240
rect 191208 13212 191880 13240
rect 187467 13209 187479 13212
rect 187421 13203 187479 13209
rect 187786 13172 187792 13184
rect 187344 13144 187792 13172
rect 187786 13132 187792 13144
rect 187844 13132 187850 13184
rect 187970 13172 187976 13184
rect 187931 13144 187976 13172
rect 187970 13132 187976 13144
rect 188028 13132 188034 13184
rect 188338 13172 188344 13184
rect 188299 13144 188344 13172
rect 188338 13132 188344 13144
rect 188396 13132 188402 13184
rect 189534 13132 189540 13184
rect 189592 13172 189598 13184
rect 191208 13172 191236 13212
rect 189592 13144 191236 13172
rect 191285 13175 191343 13181
rect 189592 13132 189598 13144
rect 191285 13141 191297 13175
rect 191331 13172 191343 13175
rect 191374 13172 191380 13184
rect 191331 13144 191380 13172
rect 191331 13141 191343 13144
rect 191285 13135 191343 13141
rect 191374 13132 191380 13144
rect 191432 13132 191438 13184
rect 191852 13172 191880 13212
rect 192113 13243 192171 13249
rect 192113 13209 192125 13243
rect 192159 13240 192171 13243
rect 192386 13240 192392 13252
rect 192159 13212 192392 13240
rect 192159 13209 192171 13212
rect 192113 13203 192171 13209
rect 192386 13200 192392 13212
rect 192444 13200 192450 13252
rect 193398 13240 193404 13252
rect 193338 13212 193404 13240
rect 193398 13200 193404 13212
rect 193456 13200 193462 13252
rect 193861 13243 193919 13249
rect 193861 13209 193873 13243
rect 193907 13240 193919 13243
rect 193950 13240 193956 13252
rect 193907 13212 193956 13240
rect 193907 13209 193919 13212
rect 193861 13203 193919 13209
rect 193950 13200 193956 13212
rect 194008 13200 194014 13252
rect 194428 13172 194456 13271
rect 201494 13268 201500 13280
rect 201552 13268 201558 13320
rect 202138 13308 202144 13320
rect 202099 13280 202144 13308
rect 202138 13268 202144 13280
rect 202196 13268 202202 13320
rect 207198 13308 207204 13320
rect 206296 13280 207204 13308
rect 194594 13200 194600 13252
rect 194652 13240 194658 13252
rect 194689 13243 194747 13249
rect 194689 13240 194701 13243
rect 194652 13212 194701 13240
rect 194652 13200 194658 13212
rect 194689 13209 194701 13212
rect 194735 13209 194747 13243
rect 194689 13203 194747 13209
rect 194778 13200 194784 13252
rect 194836 13240 194842 13252
rect 196434 13240 196440 13252
rect 194836 13212 195178 13240
rect 196347 13212 196440 13240
rect 194836 13200 194842 13212
rect 196434 13200 196440 13212
rect 196492 13240 196498 13252
rect 197354 13240 197360 13252
rect 196492 13212 197360 13240
rect 196492 13200 196498 13212
rect 197354 13200 197360 13212
rect 197412 13200 197418 13252
rect 197817 13243 197875 13249
rect 197817 13209 197829 13243
rect 197863 13240 197875 13243
rect 198645 13243 198703 13249
rect 197863 13212 198596 13240
rect 197863 13209 197875 13212
rect 197817 13203 197875 13209
rect 198568 13184 198596 13212
rect 198645 13209 198657 13243
rect 198691 13240 198703 13243
rect 202414 13240 202420 13252
rect 198691 13212 202184 13240
rect 202375 13212 202420 13240
rect 198691 13209 198703 13212
rect 198645 13203 198703 13209
rect 197722 13172 197728 13184
rect 191852 13144 197728 13172
rect 197722 13132 197728 13144
rect 197780 13132 197786 13184
rect 197906 13132 197912 13184
rect 197964 13172 197970 13184
rect 198185 13175 198243 13181
rect 198185 13172 198197 13175
rect 197964 13144 198197 13172
rect 197964 13132 197970 13144
rect 198185 13141 198197 13144
rect 198231 13141 198243 13175
rect 198550 13172 198556 13184
rect 198511 13144 198556 13172
rect 198185 13135 198243 13141
rect 198550 13132 198556 13144
rect 198608 13132 198614 13184
rect 200482 13172 200488 13184
rect 200443 13144 200488 13172
rect 200482 13132 200488 13144
rect 200540 13132 200546 13184
rect 200850 13172 200856 13184
rect 200811 13144 200856 13172
rect 200850 13132 200856 13144
rect 200908 13132 200914 13184
rect 200945 13175 201003 13181
rect 200945 13141 200957 13175
rect 200991 13172 201003 13175
rect 201310 13172 201316 13184
rect 200991 13144 201316 13172
rect 200991 13141 201003 13144
rect 200945 13135 201003 13141
rect 201310 13132 201316 13144
rect 201368 13132 201374 13184
rect 202156 13172 202184 13212
rect 202414 13200 202420 13212
rect 202472 13200 202478 13252
rect 203150 13200 203156 13252
rect 203208 13200 203214 13252
rect 203812 13212 204024 13240
rect 203812 13172 203840 13212
rect 202156 13144 203840 13172
rect 203996 13172 204024 13212
rect 204254 13200 204260 13252
rect 204312 13240 204318 13252
rect 204993 13243 205051 13249
rect 204993 13240 205005 13243
rect 204312 13212 205005 13240
rect 204312 13200 204318 13212
rect 204993 13209 205005 13212
rect 205039 13209 205051 13243
rect 204993 13203 205051 13209
rect 205450 13200 205456 13252
rect 205508 13200 205514 13252
rect 205634 13172 205640 13184
rect 203996 13144 205640 13172
rect 205634 13132 205640 13144
rect 205692 13132 205698 13184
rect 205726 13132 205732 13184
rect 205784 13172 205790 13184
rect 206296 13172 206324 13280
rect 207198 13268 207204 13280
rect 207256 13268 207262 13320
rect 207661 13311 207719 13317
rect 207661 13308 207673 13311
rect 207584 13280 207673 13308
rect 207584 13252 207612 13280
rect 207661 13277 207673 13280
rect 207707 13277 207719 13311
rect 207661 13271 207719 13277
rect 206370 13200 206376 13252
rect 206428 13240 206434 13252
rect 206428 13212 206876 13240
rect 206428 13200 206434 13212
rect 206465 13175 206523 13181
rect 206465 13172 206477 13175
rect 205784 13144 206477 13172
rect 205784 13132 205790 13144
rect 206465 13141 206477 13144
rect 206511 13141 206523 13175
rect 206848 13172 206876 13212
rect 207566 13200 207572 13252
rect 207624 13200 207630 13252
rect 207768 13240 207796 13348
rect 207845 13345 207857 13379
rect 207891 13345 207903 13379
rect 207952 13376 207980 13484
rect 210326 13472 210332 13484
rect 210384 13472 210390 13524
rect 213362 13512 213368 13524
rect 213323 13484 213368 13512
rect 213362 13472 213368 13484
rect 213420 13472 213426 13524
rect 268930 13512 268936 13524
rect 213472 13484 268936 13512
rect 208026 13404 208032 13456
rect 208084 13444 208090 13456
rect 213270 13444 213276 13456
rect 208084 13416 213276 13444
rect 208084 13404 208090 13416
rect 213270 13404 213276 13416
rect 213328 13404 213334 13456
rect 213472 13376 213500 13484
rect 268930 13472 268936 13484
rect 268988 13472 268994 13524
rect 269380 13515 269438 13521
rect 269380 13481 269392 13515
rect 269426 13512 269438 13515
rect 269574 13512 269580 13524
rect 269426 13484 269580 13512
rect 269426 13481 269438 13484
rect 269380 13475 269438 13481
rect 269574 13472 269580 13484
rect 269632 13472 269638 13524
rect 271782 13472 271788 13524
rect 271840 13512 271846 13524
rect 274269 13515 274327 13521
rect 274269 13512 274281 13515
rect 271840 13484 274281 13512
rect 271840 13472 271846 13484
rect 274269 13481 274281 13484
rect 274315 13481 274327 13515
rect 274910 13512 274916 13524
rect 274871 13484 274916 13512
rect 274269 13475 274327 13481
rect 274910 13472 274916 13484
rect 274968 13472 274974 13524
rect 277854 13512 277860 13524
rect 277815 13484 277860 13512
rect 277854 13472 277860 13484
rect 277912 13472 277918 13524
rect 280890 13512 280896 13524
rect 280851 13484 280896 13512
rect 280890 13472 280896 13484
rect 280948 13472 280954 13524
rect 284294 13472 284300 13524
rect 284352 13512 284358 13524
rect 284573 13515 284631 13521
rect 284573 13512 284585 13515
rect 284352 13484 284585 13512
rect 284352 13472 284358 13484
rect 284573 13481 284585 13484
rect 284619 13481 284631 13515
rect 284573 13475 284631 13481
rect 287054 13472 287060 13524
rect 287112 13512 287118 13524
rect 287149 13515 287207 13521
rect 287149 13512 287161 13515
rect 287112 13484 287161 13512
rect 287112 13472 287118 13484
rect 287149 13481 287161 13484
rect 287195 13481 287207 13515
rect 290090 13512 290096 13524
rect 290051 13484 290096 13512
rect 287149 13475 287207 13481
rect 290090 13472 290096 13484
rect 290148 13472 290154 13524
rect 293218 13512 293224 13524
rect 293179 13484 293224 13512
rect 293218 13472 293224 13484
rect 293276 13472 293282 13524
rect 296254 13512 296260 13524
rect 296215 13484 296260 13512
rect 296254 13472 296260 13484
rect 296312 13472 296318 13524
rect 299290 13512 299296 13524
rect 299251 13484 299296 13512
rect 299290 13472 299296 13484
rect 299348 13472 299354 13524
rect 301406 13512 301412 13524
rect 301367 13484 301412 13512
rect 301406 13472 301412 13484
rect 301464 13512 301470 13524
rect 301777 13515 301835 13521
rect 301777 13512 301789 13515
rect 301464 13484 301789 13512
rect 301464 13472 301470 13484
rect 301777 13481 301789 13484
rect 301823 13512 301835 13515
rect 302145 13515 302203 13521
rect 302145 13512 302157 13515
rect 301823 13484 302157 13512
rect 301823 13481 301835 13484
rect 301777 13475 301835 13481
rect 302145 13481 302157 13484
rect 302191 13512 302203 13515
rect 302973 13515 303031 13521
rect 302973 13512 302985 13515
rect 302191 13484 302985 13512
rect 302191 13481 302203 13484
rect 302145 13475 302203 13481
rect 302973 13481 302985 13484
rect 303019 13512 303031 13515
rect 303341 13515 303399 13521
rect 303341 13512 303353 13515
rect 303019 13484 303353 13512
rect 303019 13481 303031 13484
rect 302973 13475 303031 13481
rect 303341 13481 303353 13484
rect 303387 13481 303399 13515
rect 303341 13475 303399 13481
rect 216398 13444 216404 13456
rect 216359 13416 216404 13444
rect 216398 13404 216404 13416
rect 216456 13404 216462 13456
rect 219434 13404 219440 13456
rect 219492 13444 219498 13456
rect 220173 13447 220231 13453
rect 220173 13444 220185 13447
rect 219492 13416 220185 13444
rect 219492 13404 219498 13416
rect 220173 13413 220185 13416
rect 220219 13413 220231 13447
rect 224126 13444 224132 13456
rect 220173 13407 220231 13413
rect 220280 13416 224132 13444
rect 207952 13348 213500 13376
rect 207845 13339 207903 13345
rect 207934 13268 207940 13320
rect 207992 13308 207998 13320
rect 210513 13311 210571 13317
rect 210513 13308 210525 13311
rect 207992 13280 210525 13308
rect 207992 13268 207998 13280
rect 210513 13277 210525 13280
rect 210559 13277 210571 13311
rect 213546 13308 213552 13320
rect 213507 13280 213552 13308
rect 210513 13271 210571 13277
rect 213546 13268 213552 13280
rect 213604 13268 213610 13320
rect 216582 13308 216588 13320
rect 216495 13280 216588 13308
rect 216582 13268 216588 13280
rect 216640 13308 216646 13320
rect 220280 13308 220308 13416
rect 224126 13404 224132 13416
rect 224184 13404 224190 13456
rect 226426 13444 226432 13456
rect 224328 13416 226432 13444
rect 224034 13376 224040 13388
rect 220372 13348 224040 13376
rect 220372 13317 220400 13348
rect 224034 13336 224040 13348
rect 224092 13336 224098 13388
rect 224328 13385 224356 13416
rect 226426 13404 226432 13416
rect 226484 13404 226490 13456
rect 226610 13404 226616 13456
rect 226668 13444 226674 13456
rect 226668 13416 226713 13444
rect 226668 13404 226674 13416
rect 226886 13404 226892 13456
rect 226944 13444 226950 13456
rect 227898 13444 227904 13456
rect 226944 13416 227904 13444
rect 226944 13404 226950 13416
rect 227898 13404 227904 13416
rect 227956 13404 227962 13456
rect 229186 13404 229192 13456
rect 229244 13444 229250 13456
rect 229649 13447 229707 13453
rect 229649 13444 229661 13447
rect 229244 13416 229661 13444
rect 229244 13404 229250 13416
rect 229649 13413 229661 13416
rect 229695 13413 229707 13447
rect 229649 13407 229707 13413
rect 231780 13416 238340 13444
rect 224313 13379 224371 13385
rect 224313 13345 224325 13379
rect 224359 13345 224371 13379
rect 224313 13339 224371 13345
rect 224402 13336 224408 13388
rect 224460 13376 224466 13388
rect 227070 13376 227076 13388
rect 224460 13348 227076 13376
rect 224460 13336 224466 13348
rect 227070 13336 227076 13348
rect 227128 13336 227134 13388
rect 227162 13336 227168 13388
rect 227220 13376 227226 13388
rect 230477 13379 230535 13385
rect 230477 13376 230489 13379
rect 227220 13348 227265 13376
rect 227824 13348 230489 13376
rect 227220 13336 227226 13348
rect 216640 13280 220308 13308
rect 220357 13311 220415 13317
rect 216640 13268 216646 13280
rect 220357 13277 220369 13311
rect 220403 13277 220415 13311
rect 220357 13271 220415 13277
rect 222933 13311 222991 13317
rect 222933 13277 222945 13311
rect 222979 13308 222991 13311
rect 225877 13311 225935 13317
rect 225616 13308 225736 13310
rect 222979 13280 224356 13308
rect 222979 13277 222991 13280
rect 222933 13271 222991 13277
rect 224218 13240 224224 13252
rect 207768 13212 224224 13240
rect 224218 13200 224224 13212
rect 224276 13200 224282 13252
rect 207293 13175 207351 13181
rect 207293 13172 207305 13175
rect 206848 13144 207305 13172
rect 206465 13135 206523 13141
rect 207293 13141 207305 13144
rect 207339 13141 207351 13175
rect 207293 13135 207351 13141
rect 207382 13132 207388 13184
rect 207440 13172 207446 13184
rect 207753 13175 207811 13181
rect 207753 13172 207765 13175
rect 207440 13144 207765 13172
rect 207440 13132 207446 13144
rect 207753 13141 207765 13144
rect 207799 13172 207811 13175
rect 213546 13172 213552 13184
rect 207799 13144 213552 13172
rect 207799 13141 207811 13144
rect 207753 13135 207811 13141
rect 213546 13132 213552 13144
rect 213604 13132 213610 13184
rect 222746 13172 222752 13184
rect 222707 13144 222752 13172
rect 222746 13132 222752 13144
rect 222804 13132 222810 13184
rect 223666 13172 223672 13184
rect 223627 13144 223672 13172
rect 223666 13132 223672 13144
rect 223724 13132 223730 13184
rect 224034 13172 224040 13184
rect 223995 13144 224040 13172
rect 224034 13132 224040 13144
rect 224092 13132 224098 13184
rect 224126 13132 224132 13184
rect 224184 13172 224190 13184
rect 224328 13172 224356 13280
rect 225432 13282 225828 13308
rect 225432 13280 225644 13282
rect 225708 13280 225828 13282
rect 224402 13200 224408 13252
rect 224460 13240 224466 13252
rect 225432 13240 225460 13280
rect 224460 13212 225460 13240
rect 225800 13240 225828 13280
rect 225877 13277 225889 13311
rect 225923 13308 225935 13311
rect 227714 13308 227720 13320
rect 225923 13280 227720 13308
rect 225923 13277 225935 13280
rect 225877 13271 225935 13277
rect 227714 13268 227720 13280
rect 227772 13268 227778 13320
rect 227824 13240 227852 13348
rect 230477 13345 230489 13348
rect 230523 13376 230535 13379
rect 231780 13376 231808 13416
rect 230523 13348 231808 13376
rect 230523 13345 230535 13348
rect 230477 13339 230535 13345
rect 231946 13336 231952 13388
rect 232004 13376 232010 13388
rect 232225 13379 232283 13385
rect 232225 13376 232237 13379
rect 232004 13348 232237 13376
rect 232004 13336 232010 13348
rect 232225 13345 232237 13348
rect 232271 13345 232283 13379
rect 233142 13376 233148 13388
rect 232225 13339 232283 13345
rect 232700 13348 233148 13376
rect 227901 13311 227959 13317
rect 227901 13277 227913 13311
rect 227947 13277 227959 13311
rect 230382 13308 230388 13320
rect 229310 13280 230388 13308
rect 227901 13271 227959 13277
rect 225800 13212 227852 13240
rect 224460 13200 224466 13212
rect 227916 13184 227944 13271
rect 230382 13268 230388 13280
rect 230440 13268 230446 13320
rect 231854 13268 231860 13320
rect 231912 13268 231918 13320
rect 232038 13268 232044 13320
rect 232096 13308 232102 13320
rect 232700 13308 232728 13348
rect 233142 13336 233148 13348
rect 233200 13336 233206 13388
rect 233326 13336 233332 13388
rect 233384 13376 233390 13388
rect 237193 13379 237251 13385
rect 237193 13376 237205 13379
rect 233384 13348 237205 13376
rect 233384 13336 233390 13348
rect 233050 13308 233056 13320
rect 232096 13280 232728 13308
rect 233011 13280 233056 13308
rect 232096 13268 232102 13280
rect 233050 13268 233056 13280
rect 233108 13268 233114 13320
rect 233881 13311 233939 13317
rect 233160 13284 233740 13308
rect 233160 13280 233832 13284
rect 228082 13200 228088 13252
rect 228140 13240 228146 13252
rect 228177 13243 228235 13249
rect 228177 13240 228189 13243
rect 228140 13212 228189 13240
rect 228140 13200 228146 13212
rect 228177 13209 228189 13212
rect 228223 13209 228235 13243
rect 230750 13240 230756 13252
rect 230711 13212 230756 13240
rect 228177 13203 228235 13209
rect 230750 13200 230756 13212
rect 230808 13200 230814 13252
rect 233160 13240 233188 13280
rect 233712 13256 233832 13280
rect 233881 13277 233893 13311
rect 233927 13308 233939 13311
rect 233988 13308 234016 13348
rect 237193 13345 237205 13348
rect 237239 13345 237251 13379
rect 237193 13339 237251 13345
rect 237285 13379 237343 13385
rect 237285 13345 237297 13379
rect 237331 13376 237343 13379
rect 237926 13376 237932 13388
rect 237331 13348 237932 13376
rect 237331 13345 237343 13348
rect 237285 13339 237343 13345
rect 237926 13336 237932 13348
rect 237984 13336 237990 13388
rect 238110 13376 238116 13388
rect 238036 13348 238116 13376
rect 233927 13280 234016 13308
rect 235077 13311 235135 13317
rect 233927 13277 233939 13280
rect 233881 13271 233939 13277
rect 235077 13277 235089 13311
rect 235123 13308 235135 13311
rect 237101 13311 237159 13317
rect 237101 13308 237113 13311
rect 235123 13280 237113 13308
rect 235123 13277 235135 13280
rect 235077 13271 235135 13277
rect 237101 13277 237113 13280
rect 237147 13308 237159 13311
rect 238036 13308 238064 13348
rect 238110 13336 238116 13348
rect 238168 13336 238174 13388
rect 238312 13376 238340 13416
rect 239490 13404 239496 13456
rect 239548 13444 239554 13456
rect 239953 13447 240011 13453
rect 239953 13444 239965 13447
rect 239548 13416 239965 13444
rect 239548 13404 239554 13416
rect 239953 13413 239965 13416
rect 239999 13413 240011 13447
rect 239953 13407 240011 13413
rect 244642 13404 244648 13456
rect 244700 13444 244706 13456
rect 245378 13444 245384 13456
rect 244700 13416 245384 13444
rect 244700 13404 244706 13416
rect 245378 13404 245384 13416
rect 245436 13404 245442 13456
rect 247126 13444 247132 13456
rect 247087 13416 247132 13444
rect 247126 13404 247132 13416
rect 247184 13404 247190 13456
rect 249521 13447 249579 13453
rect 249521 13413 249533 13447
rect 249567 13444 249579 13447
rect 251082 13444 251088 13456
rect 249567 13416 251088 13444
rect 249567 13413 249579 13416
rect 249521 13407 249579 13413
rect 251082 13404 251088 13416
rect 251140 13404 251146 13456
rect 252462 13404 252468 13456
rect 252520 13444 252526 13456
rect 252833 13447 252891 13453
rect 252833 13444 252845 13447
rect 252520 13416 252845 13444
rect 252520 13404 252526 13416
rect 252833 13413 252845 13416
rect 252879 13413 252891 13447
rect 252833 13407 252891 13413
rect 254946 13404 254952 13456
rect 255004 13444 255010 13456
rect 255409 13447 255467 13453
rect 255409 13444 255421 13447
rect 255004 13416 255421 13444
rect 255004 13404 255010 13416
rect 255409 13413 255421 13416
rect 255455 13413 255467 13447
rect 259454 13444 259460 13456
rect 259415 13416 259460 13444
rect 255409 13407 255467 13413
rect 259454 13404 259460 13416
rect 259512 13404 259518 13456
rect 262677 13447 262735 13453
rect 262677 13413 262689 13447
rect 262723 13444 262735 13447
rect 263502 13444 263508 13456
rect 262723 13416 263508 13444
rect 262723 13413 262735 13416
rect 262677 13407 262735 13413
rect 263502 13404 263508 13416
rect 263560 13404 263566 13456
rect 265526 13404 265532 13456
rect 265584 13444 265590 13456
rect 265989 13447 266047 13453
rect 265989 13444 266001 13447
rect 265584 13416 266001 13444
rect 265584 13404 265590 13416
rect 265989 13413 266001 13416
rect 266035 13413 266047 13447
rect 265989 13407 266047 13413
rect 270402 13404 270408 13456
rect 270460 13444 270466 13456
rect 270460 13416 271828 13444
rect 270460 13404 270466 13416
rect 240781 13379 240839 13385
rect 240781 13376 240793 13379
rect 238312 13348 240793 13376
rect 240781 13345 240793 13348
rect 240827 13376 240839 13379
rect 243357 13379 243415 13385
rect 243357 13376 243369 13379
rect 240827 13348 243369 13376
rect 240827 13345 240839 13348
rect 240781 13339 240839 13345
rect 243357 13345 243369 13348
rect 243403 13345 243415 13379
rect 243357 13339 243415 13345
rect 244090 13336 244096 13388
rect 244148 13376 244154 13388
rect 245105 13379 245163 13385
rect 245105 13376 245117 13379
rect 244148 13348 245117 13376
rect 244148 13336 244154 13348
rect 245105 13345 245117 13348
rect 245151 13345 245163 13379
rect 245105 13339 245163 13345
rect 250165 13379 250223 13385
rect 250165 13345 250177 13379
rect 250211 13376 250223 13379
rect 250990 13376 250996 13388
rect 250211 13348 250996 13376
rect 250211 13345 250223 13348
rect 250165 13339 250223 13345
rect 238202 13308 238208 13320
rect 237147 13280 238064 13308
rect 238163 13280 238208 13308
rect 237147 13277 237159 13280
rect 237101 13271 237159 13277
rect 238202 13268 238208 13280
rect 238260 13268 238266 13320
rect 239766 13308 239772 13320
rect 239614 13280 239772 13308
rect 239766 13268 239772 13280
rect 239824 13268 239830 13320
rect 245120 13308 245148 13339
rect 250990 13336 250996 13348
rect 251048 13336 251054 13388
rect 262033 13379 262091 13385
rect 251100 13348 259776 13376
rect 251100 13320 251128 13348
rect 247313 13311 247371 13317
rect 247313 13308 247325 13311
rect 245120 13280 247325 13308
rect 247313 13277 247325 13280
rect 247359 13308 247371 13311
rect 249981 13311 250039 13317
rect 249981 13308 249993 13311
rect 247359 13280 249993 13308
rect 247359 13277 247371 13280
rect 247313 13271 247371 13277
rect 249981 13277 249993 13280
rect 250027 13277 250039 13311
rect 251082 13308 251088 13320
rect 251043 13280 251088 13308
rect 249981 13271 250039 13277
rect 251082 13268 251088 13280
rect 251140 13268 251146 13320
rect 253661 13311 253719 13317
rect 253661 13308 253673 13311
rect 252940 13280 253673 13308
rect 232056 13212 233188 13240
rect 233804 13240 233832 13256
rect 233804 13212 238432 13240
rect 225414 13172 225420 13184
rect 224184 13144 224229 13172
rect 224328 13144 225420 13172
rect 224184 13132 224190 13144
rect 225414 13132 225420 13144
rect 225472 13132 225478 13184
rect 225690 13172 225696 13184
rect 225651 13144 225696 13172
rect 225690 13132 225696 13144
rect 225748 13132 225754 13184
rect 226981 13175 227039 13181
rect 226981 13141 226993 13175
rect 227027 13172 227039 13175
rect 227070 13172 227076 13184
rect 227027 13144 227076 13172
rect 227027 13141 227039 13144
rect 226981 13135 227039 13141
rect 227070 13132 227076 13144
rect 227128 13172 227134 13184
rect 227622 13172 227628 13184
rect 227128 13144 227628 13172
rect 227128 13132 227134 13144
rect 227622 13132 227628 13144
rect 227680 13132 227686 13184
rect 227898 13172 227904 13184
rect 227811 13144 227904 13172
rect 227898 13132 227904 13144
rect 227956 13172 227962 13184
rect 232056 13172 232084 13212
rect 227956 13144 232084 13172
rect 227956 13132 227962 13144
rect 232130 13132 232136 13184
rect 232188 13172 232194 13184
rect 233145 13175 233203 13181
rect 233145 13172 233157 13175
rect 232188 13144 233157 13172
rect 232188 13132 232194 13144
rect 233145 13141 233157 13144
rect 233191 13141 233203 13175
rect 233145 13135 233203 13141
rect 233234 13132 233240 13184
rect 233292 13172 233298 13184
rect 233697 13175 233755 13181
rect 233697 13172 233709 13175
rect 233292 13144 233709 13172
rect 233292 13132 233298 13144
rect 233697 13141 233709 13144
rect 233743 13141 233755 13175
rect 234890 13172 234896 13184
rect 234851 13144 234896 13172
rect 233697 13135 233755 13141
rect 234890 13132 234896 13144
rect 234948 13132 234954 13184
rect 236733 13175 236791 13181
rect 236733 13141 236745 13175
rect 236779 13172 236791 13175
rect 237006 13172 237012 13184
rect 236779 13144 237012 13172
rect 236779 13141 236791 13144
rect 236733 13135 236791 13141
rect 237006 13132 237012 13144
rect 237064 13132 237070 13184
rect 238404 13172 238432 13212
rect 238478 13200 238484 13252
rect 238536 13240 238542 13252
rect 241054 13240 241060 13252
rect 238536 13212 238581 13240
rect 239784 13212 240088 13240
rect 241015 13212 241060 13240
rect 238536 13200 238542 13212
rect 239784 13172 239812 13212
rect 238404 13144 239812 13172
rect 240060 13172 240088 13212
rect 241054 13200 241060 13212
rect 241112 13200 241118 13252
rect 241790 13200 241796 13252
rect 241848 13200 241854 13252
rect 243630 13240 243636 13252
rect 242360 13212 242664 13240
rect 243591 13212 243636 13240
rect 242360 13172 242388 13212
rect 242526 13172 242532 13184
rect 240060 13144 242388 13172
rect 242487 13144 242532 13172
rect 242526 13132 242532 13144
rect 242584 13132 242590 13184
rect 242636 13172 242664 13212
rect 243630 13200 243636 13212
rect 243688 13200 243694 13252
rect 244918 13240 244924 13252
rect 244858 13212 244924 13240
rect 244918 13200 244924 13212
rect 244976 13200 244982 13252
rect 249720 13212 251312 13240
rect 249720 13172 249748 13212
rect 242636 13144 249748 13172
rect 249889 13175 249947 13181
rect 249889 13141 249901 13175
rect 249935 13172 249947 13175
rect 251174 13172 251180 13184
rect 249935 13144 251180 13172
rect 249935 13141 249947 13144
rect 249889 13135 249947 13141
rect 251174 13132 251180 13144
rect 251232 13132 251238 13184
rect 251284 13172 251312 13212
rect 251358 13200 251364 13252
rect 251416 13240 251422 13252
rect 251416 13212 251461 13240
rect 251416 13200 251422 13212
rect 252370 13200 252376 13252
rect 252428 13200 252434 13252
rect 252940 13172 252968 13280
rect 253661 13277 253673 13280
rect 253707 13277 253719 13311
rect 256234 13308 256240 13320
rect 253661 13271 253719 13277
rect 255240 13280 256240 13308
rect 253014 13200 253020 13252
rect 253072 13240 253078 13252
rect 253937 13243 253995 13249
rect 253937 13240 253949 13243
rect 253072 13212 253949 13240
rect 253072 13200 253078 13212
rect 253937 13209 253949 13212
rect 253983 13209 253995 13243
rect 253937 13203 253995 13209
rect 254946 13200 254952 13252
rect 255004 13200 255010 13252
rect 253474 13172 253480 13184
rect 251284 13144 253480 13172
rect 253474 13132 253480 13144
rect 253532 13172 253538 13184
rect 255240 13172 255268 13280
rect 256234 13268 256240 13280
rect 256292 13268 256298 13320
rect 259641 13311 259699 13317
rect 259641 13308 259653 13311
rect 257816 13280 259653 13308
rect 255314 13200 255320 13252
rect 255372 13240 255378 13252
rect 256513 13243 256571 13249
rect 256513 13240 256525 13243
rect 255372 13212 256525 13240
rect 255372 13200 255378 13212
rect 256513 13209 256525 13212
rect 256559 13209 256571 13243
rect 256513 13203 256571 13209
rect 256970 13200 256976 13252
rect 257028 13200 257034 13252
rect 253532 13144 255268 13172
rect 253532 13132 253538 13144
rect 256326 13132 256332 13184
rect 256384 13172 256390 13184
rect 257816 13172 257844 13280
rect 259641 13277 259653 13280
rect 259687 13277 259699 13311
rect 259748 13308 259776 13348
rect 262033 13345 262045 13379
rect 262079 13376 262091 13379
rect 263229 13379 263287 13385
rect 263229 13376 263241 13379
rect 262079 13348 263241 13376
rect 262079 13345 262091 13348
rect 262033 13339 262091 13345
rect 263229 13345 263241 13348
rect 263275 13376 263287 13379
rect 264146 13376 264152 13388
rect 263275 13348 264152 13376
rect 263275 13345 263287 13348
rect 263229 13339 263287 13345
rect 264146 13336 264152 13348
rect 264204 13336 264210 13388
rect 266541 13379 266599 13385
rect 266541 13376 266553 13379
rect 264256 13348 266553 13376
rect 264256 13317 264284 13348
rect 266541 13345 266553 13348
rect 266587 13376 266599 13379
rect 269117 13379 269175 13385
rect 269117 13376 269129 13379
rect 266587 13348 269129 13376
rect 266587 13345 266599 13348
rect 266541 13339 266599 13345
rect 269117 13345 269129 13348
rect 269163 13376 269175 13379
rect 271693 13379 271751 13385
rect 271693 13376 271705 13379
rect 269163 13348 271705 13376
rect 269163 13345 269175 13348
rect 269117 13339 269175 13345
rect 271693 13345 271705 13348
rect 271739 13345 271751 13379
rect 271800 13376 271828 13416
rect 272978 13404 272984 13456
rect 273036 13444 273042 13456
rect 273036 13416 278084 13444
rect 273036 13404 273042 13416
rect 271800 13348 273116 13376
rect 271693 13339 271751 13345
rect 264241 13311 264299 13317
rect 264241 13308 264253 13311
rect 259748 13280 264253 13308
rect 259641 13271 259699 13277
rect 264241 13277 264253 13280
rect 264287 13277 264299 13311
rect 264241 13271 264299 13277
rect 268565 13311 268623 13317
rect 268565 13277 268577 13311
rect 268611 13308 268623 13311
rect 268930 13308 268936 13320
rect 268611 13280 268936 13308
rect 268611 13277 268623 13280
rect 268565 13271 268623 13277
rect 268930 13268 268936 13280
rect 268988 13268 268994 13320
rect 273088 13294 273116 13348
rect 273162 13336 273168 13388
rect 273220 13376 273226 13388
rect 273220 13348 277992 13376
rect 273220 13336 273226 13348
rect 273254 13268 273260 13320
rect 273312 13308 273318 13320
rect 274453 13311 274511 13317
rect 274453 13308 274465 13311
rect 273312 13280 274465 13308
rect 273312 13268 273318 13280
rect 274453 13277 274465 13280
rect 274499 13277 274511 13311
rect 275094 13308 275100 13320
rect 275055 13280 275100 13308
rect 274453 13271 274511 13277
rect 275094 13268 275100 13280
rect 275152 13268 275158 13320
rect 261846 13240 261852 13252
rect 261807 13212 261852 13240
rect 261846 13200 261852 13212
rect 261904 13200 261910 13252
rect 263045 13243 263103 13249
rect 263045 13209 263057 13243
rect 263091 13240 263103 13243
rect 263410 13240 263416 13252
rect 263091 13212 263416 13240
rect 263091 13209 263103 13212
rect 263045 13203 263103 13209
rect 263410 13200 263416 13212
rect 263468 13200 263474 13252
rect 263502 13200 263508 13252
rect 263560 13240 263566 13252
rect 264422 13240 264428 13252
rect 263560 13212 264428 13240
rect 263560 13200 263566 13212
rect 264422 13200 264428 13212
rect 264480 13200 264486 13252
rect 264517 13243 264575 13249
rect 264517 13209 264529 13243
rect 264563 13240 264575 13243
rect 264606 13240 264612 13252
rect 264563 13212 264612 13240
rect 264563 13209 264575 13212
rect 264517 13203 264575 13209
rect 264606 13200 264612 13212
rect 264664 13200 264670 13252
rect 264974 13200 264980 13252
rect 265032 13200 265038 13252
rect 266817 13243 266875 13249
rect 265912 13212 266768 13240
rect 256384 13144 257844 13172
rect 256384 13132 256390 13144
rect 257982 13132 257988 13184
rect 258040 13172 258046 13184
rect 262950 13172 262956 13184
rect 258040 13144 262956 13172
rect 258040 13132 258046 13144
rect 262950 13132 262956 13144
rect 263008 13172 263014 13184
rect 263137 13175 263195 13181
rect 263137 13172 263149 13175
rect 263008 13144 263149 13172
rect 263008 13132 263014 13144
rect 263137 13141 263149 13144
rect 263183 13141 263195 13175
rect 263137 13135 263195 13141
rect 263318 13132 263324 13184
rect 263376 13172 263382 13184
rect 265912 13172 265940 13212
rect 263376 13144 265940 13172
rect 266740 13172 266768 13212
rect 266817 13209 266829 13243
rect 266863 13240 266875 13243
rect 266906 13240 266912 13252
rect 266863 13212 266912 13240
rect 266863 13209 266875 13212
rect 266817 13203 266875 13209
rect 266906 13200 266912 13212
rect 266964 13200 266970 13252
rect 268042 13212 268516 13240
rect 267642 13172 267648 13184
rect 266740 13144 267648 13172
rect 263376 13132 263382 13144
rect 267642 13132 267648 13144
rect 267700 13132 267706 13184
rect 268488 13172 268516 13212
rect 268746 13200 268752 13252
rect 268804 13240 268810 13252
rect 268804 13212 269882 13240
rect 268804 13200 268810 13212
rect 270678 13200 270684 13252
rect 270736 13240 270742 13252
rect 270736 13212 270908 13240
rect 270736 13200 270742 13212
rect 270770 13172 270776 13184
rect 268488 13144 270776 13172
rect 270770 13132 270776 13144
rect 270828 13132 270834 13184
rect 270880 13181 270908 13212
rect 270954 13200 270960 13252
rect 271012 13240 271018 13252
rect 271969 13243 272027 13249
rect 271969 13240 271981 13243
rect 271012 13212 271981 13240
rect 271012 13200 271018 13212
rect 271969 13209 271981 13212
rect 272015 13209 272027 13243
rect 277964 13240 277992 13348
rect 278056 13317 278084 13416
rect 303356 13376 303384 13475
rect 304445 13379 304503 13385
rect 304445 13376 304457 13379
rect 278148 13348 293448 13376
rect 303356 13348 304457 13376
rect 278041 13311 278099 13317
rect 278041 13277 278053 13311
rect 278087 13277 278099 13311
rect 278041 13271 278099 13277
rect 278148 13240 278176 13348
rect 281074 13308 281080 13320
rect 281035 13280 281080 13308
rect 281074 13268 281080 13280
rect 281132 13268 281138 13320
rect 284754 13308 284760 13320
rect 284715 13280 284760 13308
rect 284754 13268 284760 13280
rect 284812 13268 284818 13320
rect 287333 13311 287391 13317
rect 287333 13308 287345 13311
rect 287026 13280 287345 13308
rect 287026 13240 287054 13280
rect 287333 13277 287345 13280
rect 287379 13277 287391 13311
rect 290274 13308 290280 13320
rect 290235 13280 290280 13308
rect 287333 13271 287391 13277
rect 290274 13268 290280 13280
rect 290332 13268 290338 13320
rect 293420 13317 293448 13348
rect 304445 13345 304457 13348
rect 304491 13376 304503 13379
rect 304905 13379 304963 13385
rect 304905 13376 304917 13379
rect 304491 13348 304917 13376
rect 304491 13345 304503 13348
rect 304445 13339 304503 13345
rect 304905 13345 304917 13348
rect 304951 13376 304963 13379
rect 304994 13376 305000 13388
rect 304951 13348 305000 13376
rect 304951 13345 304963 13348
rect 304905 13339 304963 13345
rect 304994 13336 305000 13348
rect 305052 13376 305058 13388
rect 305365 13379 305423 13385
rect 305365 13376 305377 13379
rect 305052 13348 305377 13376
rect 305052 13336 305058 13348
rect 305365 13345 305377 13348
rect 305411 13345 305423 13379
rect 305365 13339 305423 13345
rect 293405 13311 293463 13317
rect 293405 13277 293417 13311
rect 293451 13277 293463 13311
rect 296441 13311 296499 13317
rect 296441 13308 296453 13311
rect 293405 13271 293463 13277
rect 295904 13280 296453 13308
rect 277964 13212 278176 13240
rect 282886 13212 287054 13240
rect 271969 13203 272027 13209
rect 270865 13175 270923 13181
rect 270865 13141 270877 13175
rect 270911 13172 270923 13175
rect 271782 13172 271788 13184
rect 270911 13144 271788 13172
rect 270911 13141 270923 13144
rect 270865 13135 270923 13141
rect 271782 13132 271788 13144
rect 271840 13132 271846 13184
rect 272886 13132 272892 13184
rect 272944 13172 272950 13184
rect 273441 13175 273499 13181
rect 273441 13172 273453 13175
rect 272944 13144 273453 13172
rect 272944 13132 272950 13144
rect 273441 13141 273453 13144
rect 273487 13172 273499 13175
rect 282886 13172 282914 13212
rect 295904 13184 295932 13280
rect 296441 13277 296453 13280
rect 296487 13277 296499 13311
rect 299474 13308 299480 13320
rect 299435 13280 299480 13308
rect 296441 13271 296499 13277
rect 299474 13268 299480 13280
rect 299532 13268 299538 13320
rect 303522 13268 303528 13320
rect 303580 13308 303586 13320
rect 303709 13311 303767 13317
rect 303709 13308 303721 13311
rect 303580 13280 303721 13308
rect 303580 13268 303586 13280
rect 303709 13277 303721 13280
rect 303755 13277 303767 13311
rect 303709 13271 303767 13277
rect 295886 13172 295892 13184
rect 273487 13144 282914 13172
rect 295847 13144 295892 13172
rect 273487 13141 273499 13144
rect 273441 13135 273499 13141
rect 295886 13132 295892 13144
rect 295944 13132 295950 13184
rect 1104 13082 305808 13104
rect 1104 13030 77148 13082
rect 77200 13030 77212 13082
rect 77264 13030 77276 13082
rect 77328 13030 77340 13082
rect 77392 13030 77404 13082
rect 77456 13030 153346 13082
rect 153398 13030 153410 13082
rect 153462 13030 153474 13082
rect 153526 13030 153538 13082
rect 153590 13030 153602 13082
rect 153654 13030 229544 13082
rect 229596 13030 229608 13082
rect 229660 13030 229672 13082
rect 229724 13030 229736 13082
rect 229788 13030 229800 13082
rect 229852 13030 305808 13082
rect 1104 13008 305808 13030
rect 26050 12968 26056 12980
rect 26011 12940 26056 12968
rect 26050 12928 26056 12940
rect 26108 12928 26114 12980
rect 27433 12971 27491 12977
rect 27433 12937 27445 12971
rect 27479 12937 27491 12971
rect 32214 12968 32220 12980
rect 27433 12931 27491 12937
rect 27632 12940 32220 12968
rect 20162 12860 20168 12912
rect 20220 12900 20226 12912
rect 20220 12872 22094 12900
rect 20220 12860 20226 12872
rect 22066 12628 22094 12872
rect 27338 12860 27344 12912
rect 27396 12900 27402 12912
rect 27448 12900 27476 12931
rect 27396 12872 27476 12900
rect 27396 12860 27402 12872
rect 26237 12835 26295 12841
rect 26237 12801 26249 12835
rect 26283 12832 26295 12835
rect 27632 12832 27660 12940
rect 32214 12928 32220 12940
rect 32272 12968 32278 12980
rect 33873 12971 33931 12977
rect 33873 12968 33885 12971
rect 32272 12940 33885 12968
rect 32272 12928 32278 12940
rect 33873 12937 33885 12940
rect 33919 12937 33931 12971
rect 33873 12931 33931 12937
rect 34146 12928 34152 12980
rect 34204 12968 34210 12980
rect 34793 12971 34851 12977
rect 34793 12968 34805 12971
rect 34204 12940 34805 12968
rect 34204 12928 34210 12940
rect 34793 12937 34805 12940
rect 34839 12937 34851 12971
rect 35526 12968 35532 12980
rect 35487 12940 35532 12968
rect 34793 12931 34851 12937
rect 35526 12928 35532 12940
rect 35584 12928 35590 12980
rect 36633 12971 36691 12977
rect 36633 12968 36645 12971
rect 35636 12940 36645 12968
rect 28994 12900 29000 12912
rect 26283 12804 27660 12832
rect 27724 12872 29000 12900
rect 26283 12801 26295 12804
rect 26237 12795 26295 12801
rect 23198 12724 23204 12776
rect 23256 12764 23262 12776
rect 27724 12764 27752 12872
rect 28994 12860 29000 12872
rect 29052 12860 29058 12912
rect 30374 12900 30380 12912
rect 29104 12872 30380 12900
rect 27801 12835 27859 12841
rect 27801 12801 27813 12835
rect 27847 12832 27859 12835
rect 27982 12832 27988 12844
rect 27847 12804 27988 12832
rect 27847 12801 27859 12804
rect 27801 12795 27859 12801
rect 27982 12792 27988 12804
rect 28040 12792 28046 12844
rect 23256 12736 27752 12764
rect 27893 12767 27951 12773
rect 23256 12724 23262 12736
rect 27893 12733 27905 12767
rect 27939 12733 27951 12767
rect 28074 12764 28080 12776
rect 28035 12736 28080 12764
rect 27893 12727 27951 12733
rect 27154 12656 27160 12708
rect 27212 12696 27218 12708
rect 27908 12696 27936 12727
rect 28074 12724 28080 12736
rect 28132 12724 28138 12776
rect 29104 12773 29132 12872
rect 30374 12860 30380 12872
rect 30432 12860 30438 12912
rect 31570 12900 31576 12912
rect 31326 12872 31576 12900
rect 31570 12860 31576 12872
rect 31628 12860 31634 12912
rect 34422 12900 34428 12912
rect 33626 12872 34428 12900
rect 34422 12860 34428 12872
rect 34480 12860 34486 12912
rect 35636 12900 35664 12940
rect 36633 12937 36645 12940
rect 36679 12937 36691 12971
rect 42521 12971 42579 12977
rect 36633 12931 36691 12937
rect 37384 12940 41414 12968
rect 37384 12909 37412 12940
rect 34532 12872 35664 12900
rect 36541 12903 36599 12909
rect 33686 12792 33692 12844
rect 33744 12832 33750 12844
rect 34532 12832 34560 12872
rect 36541 12869 36553 12903
rect 36587 12900 36599 12903
rect 37369 12903 37427 12909
rect 37369 12900 37381 12903
rect 36587 12872 37381 12900
rect 36587 12869 36599 12872
rect 36541 12863 36599 12869
rect 37369 12869 37381 12872
rect 37415 12869 37427 12903
rect 37369 12863 37427 12869
rect 37458 12860 37464 12912
rect 37516 12900 37522 12912
rect 38473 12903 38531 12909
rect 38473 12900 38485 12903
rect 37516 12872 38485 12900
rect 37516 12860 37522 12872
rect 38473 12869 38485 12872
rect 38519 12869 38531 12903
rect 38473 12863 38531 12869
rect 39666 12860 39672 12912
rect 39724 12900 39730 12912
rect 39761 12903 39819 12909
rect 39761 12900 39773 12903
rect 39724 12872 39773 12900
rect 39724 12860 39730 12872
rect 39761 12869 39773 12872
rect 39807 12869 39819 12903
rect 41046 12900 41052 12912
rect 40986 12872 41052 12900
rect 39761 12863 39819 12869
rect 41046 12860 41052 12872
rect 41104 12860 41110 12912
rect 41386 12900 41414 12940
rect 42521 12937 42533 12971
rect 42567 12968 42579 12971
rect 43254 12968 43260 12980
rect 42567 12940 43260 12968
rect 42567 12937 42579 12940
rect 42521 12931 42579 12937
rect 43254 12928 43260 12940
rect 43312 12928 43318 12980
rect 43441 12971 43499 12977
rect 43441 12937 43453 12971
rect 43487 12968 43499 12971
rect 44266 12968 44272 12980
rect 43487 12940 44272 12968
rect 43487 12937 43499 12940
rect 43441 12931 43499 12937
rect 44266 12928 44272 12940
rect 44324 12928 44330 12980
rect 44542 12968 44548 12980
rect 44503 12940 44548 12968
rect 44542 12928 44548 12940
rect 44600 12928 44606 12980
rect 51997 12971 52055 12977
rect 51997 12937 52009 12971
rect 52043 12968 52055 12971
rect 53282 12968 53288 12980
rect 52043 12940 53288 12968
rect 52043 12937 52055 12940
rect 51997 12931 52055 12937
rect 53282 12928 53288 12940
rect 53340 12928 53346 12980
rect 53561 12971 53619 12977
rect 53561 12937 53573 12971
rect 53607 12937 53619 12971
rect 53561 12931 53619 12937
rect 53929 12971 53987 12977
rect 53929 12937 53941 12971
rect 53975 12968 53987 12971
rect 54662 12968 54668 12980
rect 53975 12940 54668 12968
rect 53975 12937 53987 12940
rect 53929 12931 53987 12937
rect 42978 12900 42984 12912
rect 41386 12872 42984 12900
rect 42978 12860 42984 12872
rect 43036 12860 43042 12912
rect 53576 12900 53604 12931
rect 54662 12928 54668 12940
rect 54720 12928 54726 12980
rect 55858 12928 55864 12980
rect 55916 12968 55922 12980
rect 57974 12968 57980 12980
rect 55916 12940 57980 12968
rect 55916 12928 55922 12940
rect 57974 12928 57980 12940
rect 58032 12928 58038 12980
rect 58529 12971 58587 12977
rect 58529 12937 58541 12971
rect 58575 12968 58587 12971
rect 59630 12968 59636 12980
rect 58575 12940 59636 12968
rect 58575 12937 58587 12940
rect 58529 12931 58587 12937
rect 59630 12928 59636 12940
rect 59688 12928 59694 12980
rect 72142 12968 72148 12980
rect 72103 12940 72148 12968
rect 72142 12928 72148 12940
rect 72200 12928 72206 12980
rect 72326 12928 72332 12980
rect 72384 12968 72390 12980
rect 74718 12968 74724 12980
rect 72384 12940 74724 12968
rect 72384 12928 72390 12940
rect 74718 12928 74724 12940
rect 74776 12928 74782 12980
rect 83918 12968 83924 12980
rect 75564 12940 83924 12968
rect 52196 12872 53604 12900
rect 33744 12804 34560 12832
rect 34701 12835 34759 12841
rect 33744 12792 33750 12804
rect 34701 12801 34713 12835
rect 34747 12801 34759 12835
rect 34701 12795 34759 12801
rect 35713 12835 35771 12841
rect 35713 12801 35725 12835
rect 35759 12832 35771 12835
rect 38381 12835 38439 12841
rect 38381 12832 38393 12835
rect 35759 12804 38393 12832
rect 35759 12801 35771 12804
rect 35713 12795 35771 12801
rect 38381 12801 38393 12804
rect 38427 12832 38439 12835
rect 39298 12832 39304 12844
rect 38427 12804 39304 12832
rect 38427 12801 38439 12804
rect 38381 12795 38439 12801
rect 29089 12767 29147 12773
rect 29089 12764 29101 12767
rect 28276 12736 29101 12764
rect 27212 12668 27936 12696
rect 27212 12656 27218 12668
rect 28276 12628 28304 12736
rect 29089 12733 29101 12736
rect 29135 12733 29147 12767
rect 29089 12727 29147 12733
rect 29273 12767 29331 12773
rect 29273 12733 29285 12767
rect 29319 12764 29331 12767
rect 29638 12764 29644 12776
rect 29319 12736 29644 12764
rect 29319 12733 29331 12736
rect 29273 12727 29331 12733
rect 29638 12724 29644 12736
rect 29696 12724 29702 12776
rect 29822 12764 29828 12776
rect 29735 12736 29828 12764
rect 29822 12724 29828 12736
rect 29880 12724 29886 12776
rect 30098 12764 30104 12776
rect 30059 12736 30104 12764
rect 30098 12724 30104 12736
rect 30156 12724 30162 12776
rect 32125 12767 32183 12773
rect 32125 12733 32137 12767
rect 32171 12733 32183 12767
rect 32125 12727 32183 12733
rect 32401 12767 32459 12773
rect 32401 12733 32413 12767
rect 32447 12764 32459 12767
rect 33042 12764 33048 12776
rect 32447 12736 33048 12764
rect 32447 12733 32459 12736
rect 32401 12727 32459 12733
rect 22066 12600 28304 12628
rect 28629 12631 28687 12637
rect 28629 12597 28641 12631
rect 28675 12628 28687 12631
rect 28902 12628 28908 12640
rect 28675 12600 28908 12628
rect 28675 12597 28687 12600
rect 28629 12591 28687 12597
rect 28902 12588 28908 12600
rect 28960 12588 28966 12640
rect 29840 12628 29868 12724
rect 32140 12696 32168 12727
rect 33042 12724 33048 12736
rect 33100 12724 33106 12776
rect 33410 12724 33416 12776
rect 33468 12764 33474 12776
rect 34330 12764 34336 12776
rect 33468 12736 34336 12764
rect 33468 12724 33474 12736
rect 34330 12724 34336 12736
rect 34388 12764 34394 12776
rect 34716 12764 34744 12795
rect 39298 12792 39304 12804
rect 39356 12792 39362 12844
rect 41506 12792 41512 12844
rect 41564 12832 41570 12844
rect 41693 12835 41751 12841
rect 41693 12832 41705 12835
rect 41564 12804 41705 12832
rect 41564 12792 41570 12804
rect 41693 12801 41705 12804
rect 41739 12832 41751 12835
rect 42429 12835 42487 12841
rect 42429 12832 42441 12835
rect 41739 12804 42441 12832
rect 41739 12801 41751 12804
rect 41693 12795 41751 12801
rect 42429 12801 42441 12804
rect 42475 12801 42487 12835
rect 44729 12835 44787 12841
rect 44729 12832 44741 12835
rect 42429 12795 42487 12801
rect 43548 12804 44741 12832
rect 34388 12736 34744 12764
rect 34388 12724 34394 12736
rect 34882 12724 34888 12776
rect 34940 12764 34946 12776
rect 34940 12736 34985 12764
rect 34940 12724 34946 12736
rect 35342 12724 35348 12776
rect 35400 12764 35406 12776
rect 37553 12767 37611 12773
rect 37553 12764 37565 12767
rect 35400 12736 37565 12764
rect 35400 12724 35406 12736
rect 37553 12733 37565 12736
rect 37599 12733 37611 12767
rect 37553 12727 37611 12733
rect 38565 12767 38623 12773
rect 38565 12733 38577 12767
rect 38611 12764 38623 12767
rect 39390 12764 39396 12776
rect 38611 12736 39396 12764
rect 38611 12733 38623 12736
rect 38565 12727 38623 12733
rect 39390 12724 39396 12736
rect 39448 12724 39454 12776
rect 39485 12767 39543 12773
rect 39485 12733 39497 12767
rect 39531 12733 39543 12767
rect 39485 12727 39543 12733
rect 39500 12696 39528 12727
rect 40954 12724 40960 12776
rect 41012 12764 41018 12776
rect 43070 12764 43076 12776
rect 41012 12736 43076 12764
rect 41012 12724 41018 12736
rect 43070 12724 43076 12736
rect 43128 12724 43134 12776
rect 43162 12724 43168 12776
rect 43220 12764 43226 12776
rect 43548 12773 43576 12804
rect 44729 12801 44741 12804
rect 44775 12832 44787 12835
rect 45370 12832 45376 12844
rect 44775 12804 45376 12832
rect 44775 12801 44787 12804
rect 44729 12795 44787 12801
rect 45370 12792 45376 12804
rect 45428 12792 45434 12844
rect 52196 12841 52224 12872
rect 55490 12860 55496 12912
rect 55548 12860 55554 12912
rect 57330 12860 57336 12912
rect 57388 12900 57394 12912
rect 58621 12903 58679 12909
rect 58621 12900 58633 12903
rect 57388 12872 58633 12900
rect 57388 12860 57394 12872
rect 58621 12869 58633 12872
rect 58667 12900 58679 12903
rect 60642 12900 60648 12912
rect 58667 12872 60648 12900
rect 58667 12869 58679 12872
rect 58621 12863 58679 12869
rect 60642 12860 60648 12872
rect 60700 12860 60706 12912
rect 65886 12860 65892 12912
rect 65944 12900 65950 12912
rect 75564 12900 75592 12940
rect 77849 12903 77907 12909
rect 77849 12900 77861 12903
rect 65944 12872 75592 12900
rect 77050 12872 77861 12900
rect 65944 12860 65950 12872
rect 52181 12835 52239 12841
rect 52181 12801 52193 12835
rect 52227 12801 52239 12835
rect 52181 12795 52239 12801
rect 52917 12835 52975 12841
rect 52917 12801 52929 12835
rect 52963 12832 52975 12835
rect 53742 12832 53748 12844
rect 52963 12804 53748 12832
rect 52963 12801 52975 12804
rect 52917 12795 52975 12801
rect 53742 12792 53748 12804
rect 53800 12792 53806 12844
rect 54018 12838 54024 12844
rect 53944 12832 54024 12838
rect 53852 12804 54024 12832
rect 43533 12767 43591 12773
rect 43533 12764 43545 12767
rect 43220 12736 43545 12764
rect 43220 12724 43226 12736
rect 43533 12733 43545 12736
rect 43579 12733 43591 12767
rect 43533 12727 43591 12733
rect 43717 12767 43775 12773
rect 43717 12733 43729 12767
rect 43763 12764 43775 12767
rect 43806 12764 43812 12776
rect 43763 12736 43812 12764
rect 43763 12733 43775 12736
rect 43717 12727 43775 12733
rect 43806 12724 43812 12736
rect 43864 12764 43870 12776
rect 45462 12764 45468 12776
rect 43864 12736 45468 12764
rect 43864 12724 43870 12736
rect 45462 12724 45468 12736
rect 45520 12724 45526 12776
rect 51350 12724 51356 12776
rect 51408 12764 51414 12776
rect 53852 12764 53880 12804
rect 54018 12792 54024 12804
rect 54076 12792 54082 12844
rect 54754 12836 54760 12844
rect 54680 12832 54760 12836
rect 54667 12804 54760 12832
rect 54110 12764 54116 12776
rect 51408 12736 53880 12764
rect 54071 12736 54116 12764
rect 51408 12724 51414 12736
rect 54110 12724 54116 12736
rect 54168 12724 54174 12776
rect 54680 12696 54708 12804
rect 54754 12792 54760 12804
rect 54812 12792 54818 12844
rect 57057 12835 57115 12841
rect 57057 12801 57069 12835
rect 57103 12832 57115 12835
rect 57422 12832 57428 12844
rect 57103 12804 57428 12832
rect 57103 12801 57115 12804
rect 57057 12795 57115 12801
rect 57422 12792 57428 12804
rect 57480 12792 57486 12844
rect 72329 12835 72387 12841
rect 72329 12801 72341 12835
rect 72375 12832 72387 12835
rect 74810 12832 74816 12844
rect 72375 12804 74816 12832
rect 72375 12801 72387 12804
rect 72329 12795 72387 12801
rect 74810 12792 74816 12804
rect 74868 12792 74874 12844
rect 75089 12835 75147 12841
rect 75089 12801 75101 12835
rect 75135 12832 75147 12835
rect 75454 12832 75460 12844
rect 75135 12804 75460 12832
rect 75135 12801 75147 12804
rect 75089 12795 75147 12801
rect 75454 12792 75460 12804
rect 75512 12792 75518 12844
rect 75564 12841 75592 12872
rect 77849 12869 77861 12872
rect 77895 12869 77907 12903
rect 77849 12863 77907 12869
rect 78398 12860 78404 12912
rect 78456 12900 78462 12912
rect 78585 12903 78643 12909
rect 78585 12900 78597 12903
rect 78456 12872 78597 12900
rect 78456 12860 78462 12872
rect 78585 12869 78597 12872
rect 78631 12869 78643 12903
rect 78585 12863 78643 12869
rect 75549 12835 75607 12841
rect 75549 12801 75561 12835
rect 75595 12801 75607 12835
rect 75549 12795 75607 12801
rect 77757 12835 77815 12841
rect 77757 12801 77769 12835
rect 77803 12832 77815 12835
rect 78493 12835 78551 12841
rect 78493 12832 78505 12835
rect 77803 12804 78505 12832
rect 77803 12801 77815 12804
rect 77757 12795 77815 12801
rect 78493 12801 78505 12804
rect 78539 12832 78551 12835
rect 79321 12835 79379 12841
rect 78539 12804 78628 12832
rect 78539 12801 78551 12804
rect 78493 12795 78551 12801
rect 78600 12776 78628 12804
rect 79321 12801 79333 12835
rect 79367 12832 79379 12835
rect 79686 12832 79692 12844
rect 79367 12804 79692 12832
rect 79367 12801 79379 12804
rect 79321 12795 79379 12801
rect 79686 12792 79692 12804
rect 79744 12792 79750 12844
rect 79796 12841 79824 12940
rect 83918 12928 83924 12940
rect 83976 12928 83982 12980
rect 86494 12968 86500 12980
rect 84672 12940 86500 12968
rect 80514 12860 80520 12912
rect 80572 12860 80578 12912
rect 82906 12860 82912 12912
rect 82964 12900 82970 12912
rect 84672 12900 84700 12940
rect 86494 12928 86500 12940
rect 86552 12928 86558 12980
rect 87138 12968 87144 12980
rect 86880 12940 87144 12968
rect 86880 12900 86908 12940
rect 87138 12928 87144 12940
rect 87196 12928 87202 12980
rect 89533 12971 89591 12977
rect 89533 12937 89545 12971
rect 89579 12968 89591 12971
rect 89579 12940 89714 12968
rect 89579 12937 89591 12940
rect 89533 12931 89591 12937
rect 89686 12900 89714 12940
rect 90450 12928 90456 12980
rect 90508 12968 90514 12980
rect 91097 12971 91155 12977
rect 91097 12968 91109 12971
rect 90508 12940 91109 12968
rect 90508 12928 90514 12940
rect 91097 12937 91109 12940
rect 91143 12937 91155 12971
rect 91097 12931 91155 12937
rect 91646 12928 91652 12980
rect 91704 12968 91710 12980
rect 97994 12968 98000 12980
rect 91704 12940 98000 12968
rect 91704 12928 91710 12940
rect 97994 12928 98000 12940
rect 98052 12928 98058 12980
rect 99346 12940 108344 12968
rect 90542 12900 90548 12912
rect 82964 12872 84700 12900
rect 85514 12872 86908 12900
rect 87722 12872 89576 12900
rect 89686 12872 90548 12900
rect 82964 12860 82970 12872
rect 79781 12835 79839 12841
rect 79781 12801 79793 12835
rect 79827 12801 79839 12835
rect 86221 12835 86279 12841
rect 86221 12832 86233 12835
rect 79781 12795 79839 12801
rect 85500 12804 86233 12832
rect 55030 12764 55036 12776
rect 54991 12736 55036 12764
rect 55030 12724 55036 12736
rect 55088 12724 55094 12776
rect 58713 12767 58771 12773
rect 58713 12733 58725 12767
rect 58759 12733 58771 12767
rect 75825 12767 75883 12773
rect 75825 12764 75837 12767
rect 58713 12727 58771 12733
rect 74920 12736 75837 12764
rect 58728 12696 58756 12727
rect 74920 12705 74948 12736
rect 75825 12733 75837 12736
rect 75871 12733 75883 12767
rect 75825 12727 75883 12733
rect 78582 12724 78588 12776
rect 78640 12724 78646 12776
rect 80057 12767 80115 12773
rect 80057 12764 80069 12767
rect 79152 12736 80069 12764
rect 31128 12668 32168 12696
rect 31128 12628 31156 12668
rect 29840 12600 31156 12628
rect 31386 12588 31392 12640
rect 31444 12628 31450 12640
rect 31573 12631 31631 12637
rect 31573 12628 31585 12631
rect 31444 12600 31585 12628
rect 31444 12588 31450 12600
rect 31573 12597 31585 12600
rect 31619 12597 31631 12631
rect 32140 12628 32168 12668
rect 33428 12668 39528 12696
rect 32398 12628 32404 12640
rect 32140 12600 32404 12628
rect 31573 12591 31631 12597
rect 32398 12588 32404 12600
rect 32456 12628 32462 12640
rect 33428 12628 33456 12668
rect 32456 12600 33456 12628
rect 32456 12588 32462 12600
rect 34146 12588 34152 12640
rect 34204 12628 34210 12640
rect 34333 12631 34391 12637
rect 34333 12628 34345 12631
rect 34204 12600 34345 12628
rect 34204 12588 34210 12600
rect 34333 12597 34345 12600
rect 34379 12597 34391 12631
rect 38010 12628 38016 12640
rect 37971 12600 38016 12628
rect 34333 12591 34391 12597
rect 38010 12588 38016 12600
rect 38068 12588 38074 12640
rect 39500 12628 39528 12668
rect 40788 12668 54708 12696
rect 56336 12668 58756 12696
rect 74905 12699 74963 12705
rect 40788 12628 40816 12668
rect 56336 12640 56364 12668
rect 41230 12628 41236 12640
rect 39500 12600 40816 12628
rect 41191 12600 41236 12628
rect 41230 12588 41236 12600
rect 41288 12588 41294 12640
rect 41782 12628 41788 12640
rect 41743 12600 41788 12628
rect 41782 12588 41788 12600
rect 41840 12588 41846 12640
rect 42794 12588 42800 12640
rect 42852 12628 42858 12640
rect 43073 12631 43131 12637
rect 43073 12628 43085 12631
rect 42852 12600 43085 12628
rect 42852 12588 42858 12600
rect 43073 12597 43085 12600
rect 43119 12597 43131 12631
rect 43073 12591 43131 12597
rect 43254 12588 43260 12640
rect 43312 12628 43318 12640
rect 43806 12628 43812 12640
rect 43312 12600 43812 12628
rect 43312 12588 43318 12600
rect 43806 12588 43812 12600
rect 43864 12588 43870 12640
rect 53009 12631 53067 12637
rect 53009 12597 53021 12631
rect 53055 12628 53067 12631
rect 53098 12628 53104 12640
rect 53055 12600 53104 12628
rect 53055 12597 53067 12600
rect 53009 12591 53067 12597
rect 53098 12588 53104 12600
rect 53156 12588 53162 12640
rect 54110 12588 54116 12640
rect 54168 12628 54174 12640
rect 55582 12628 55588 12640
rect 54168 12600 55588 12628
rect 54168 12588 54174 12600
rect 55582 12588 55588 12600
rect 55640 12628 55646 12640
rect 56318 12628 56324 12640
rect 55640 12600 56324 12628
rect 55640 12588 55646 12600
rect 56318 12588 56324 12600
rect 56376 12588 56382 12640
rect 56502 12628 56508 12640
rect 56463 12600 56508 12628
rect 56502 12588 56508 12600
rect 56560 12588 56566 12640
rect 57164 12637 57192 12668
rect 74905 12665 74917 12699
rect 74951 12665 74963 12699
rect 77846 12696 77852 12708
rect 74905 12659 74963 12665
rect 76852 12668 77852 12696
rect 57149 12631 57207 12637
rect 57149 12597 57161 12631
rect 57195 12597 57207 12631
rect 57149 12591 57207 12597
rect 57238 12588 57244 12640
rect 57296 12628 57302 12640
rect 58161 12631 58219 12637
rect 58161 12628 58173 12631
rect 57296 12600 58173 12628
rect 57296 12588 57302 12600
rect 58161 12597 58173 12600
rect 58207 12597 58219 12631
rect 58161 12591 58219 12597
rect 72694 12588 72700 12640
rect 72752 12628 72758 12640
rect 74994 12628 75000 12640
rect 72752 12600 75000 12628
rect 72752 12588 72758 12600
rect 74994 12588 75000 12600
rect 75052 12588 75058 12640
rect 75178 12588 75184 12640
rect 75236 12628 75242 12640
rect 76852 12628 76880 12668
rect 77846 12656 77852 12668
rect 77904 12656 77910 12708
rect 78122 12656 78128 12708
rect 78180 12696 78186 12708
rect 79152 12705 79180 12736
rect 80057 12733 80069 12736
rect 80103 12733 80115 12767
rect 80057 12727 80115 12733
rect 80790 12724 80796 12776
rect 80848 12764 80854 12776
rect 84013 12767 84071 12773
rect 84013 12764 84025 12767
rect 80848 12736 84025 12764
rect 80848 12724 80854 12736
rect 84013 12733 84025 12736
rect 84059 12733 84071 12767
rect 84013 12727 84071 12733
rect 84289 12767 84347 12773
rect 84289 12733 84301 12767
rect 84335 12764 84347 12767
rect 84838 12764 84844 12776
rect 84335 12736 84844 12764
rect 84335 12733 84347 12736
rect 84289 12727 84347 12733
rect 79137 12699 79195 12705
rect 78180 12668 78720 12696
rect 78180 12656 78186 12668
rect 75236 12600 76880 12628
rect 75236 12588 75242 12600
rect 77202 12588 77208 12640
rect 77260 12628 77266 12640
rect 77297 12631 77355 12637
rect 77297 12628 77309 12631
rect 77260 12600 77309 12628
rect 77260 12588 77266 12600
rect 77297 12597 77309 12600
rect 77343 12597 77355 12631
rect 78692 12628 78720 12668
rect 79137 12665 79149 12699
rect 79183 12665 79195 12699
rect 79137 12659 79195 12665
rect 81434 12656 81440 12708
rect 81492 12696 81498 12708
rect 81529 12699 81587 12705
rect 81529 12696 81541 12699
rect 81492 12668 81541 12696
rect 81492 12656 81498 12668
rect 81529 12665 81541 12668
rect 81575 12665 81587 12699
rect 81529 12659 81587 12665
rect 81618 12628 81624 12640
rect 78692 12600 81624 12628
rect 77297 12591 77355 12597
rect 81618 12588 81624 12600
rect 81676 12588 81682 12640
rect 84028 12628 84056 12727
rect 84838 12724 84844 12736
rect 84896 12724 84902 12776
rect 85500 12764 85528 12804
rect 85316 12736 85528 12764
rect 85316 12628 85344 12736
rect 85758 12628 85764 12640
rect 84028 12600 85344 12628
rect 85719 12600 85764 12628
rect 85758 12588 85764 12600
rect 85816 12588 85822 12640
rect 86144 12628 86172 12804
rect 86221 12801 86233 12804
rect 86267 12801 86279 12835
rect 89548 12832 89576 12872
rect 90542 12860 90548 12872
rect 90600 12860 90606 12912
rect 90726 12860 90732 12912
rect 90784 12900 90790 12912
rect 99346 12900 99374 12940
rect 99466 12900 99472 12912
rect 90784 12872 99374 12900
rect 99427 12872 99472 12900
rect 90784 12860 90790 12872
rect 99466 12860 99472 12872
rect 99524 12860 99530 12912
rect 99926 12860 99932 12912
rect 99984 12860 99990 12912
rect 104618 12900 104624 12912
rect 104579 12872 104624 12900
rect 104618 12860 104624 12872
rect 104676 12860 104682 12912
rect 104710 12860 104716 12912
rect 104768 12900 104774 12912
rect 104768 12872 106136 12900
rect 104768 12860 104774 12872
rect 90174 12832 90180 12844
rect 89548 12804 90180 12832
rect 86221 12795 86279 12801
rect 90174 12792 90180 12804
rect 90232 12792 90238 12844
rect 90450 12832 90456 12844
rect 90363 12804 90456 12832
rect 90450 12792 90456 12804
rect 90508 12832 90514 12844
rect 90634 12832 90640 12844
rect 90508 12804 90640 12832
rect 90508 12792 90514 12804
rect 90634 12792 90640 12804
rect 90692 12792 90698 12844
rect 91281 12835 91339 12841
rect 91281 12801 91293 12835
rect 91327 12801 91339 12835
rect 91281 12795 91339 12801
rect 98549 12835 98607 12841
rect 98549 12801 98561 12835
rect 98595 12801 98607 12835
rect 105170 12832 105176 12844
rect 102810 12804 105176 12832
rect 98549 12795 98607 12801
rect 86494 12764 86500 12776
rect 86455 12736 86500 12764
rect 86494 12724 86500 12736
rect 86552 12724 86558 12776
rect 88242 12724 88248 12776
rect 88300 12764 88306 12776
rect 89625 12767 89683 12773
rect 89625 12764 89637 12767
rect 88300 12736 89637 12764
rect 88300 12724 88306 12736
rect 89625 12733 89637 12736
rect 89671 12764 89683 12767
rect 89714 12764 89720 12776
rect 89671 12736 89720 12764
rect 89671 12733 89683 12736
rect 89625 12727 89683 12733
rect 89714 12724 89720 12736
rect 89772 12724 89778 12776
rect 89809 12767 89867 12773
rect 89809 12733 89821 12767
rect 89855 12764 89867 12767
rect 89855 12736 89944 12764
rect 89855 12733 89867 12736
rect 89809 12727 89867 12733
rect 89916 12640 89944 12736
rect 90082 12724 90088 12776
rect 90140 12764 90146 12776
rect 91296 12764 91324 12795
rect 90140 12736 91324 12764
rect 90140 12724 90146 12736
rect 98564 12696 98592 12795
rect 105170 12792 105176 12804
rect 105228 12792 105234 12844
rect 106108 12841 106136 12872
rect 106093 12835 106151 12841
rect 106093 12801 106105 12835
rect 106139 12801 106151 12835
rect 106093 12795 106151 12801
rect 99190 12764 99196 12776
rect 99103 12736 99196 12764
rect 99190 12724 99196 12736
rect 99248 12764 99254 12776
rect 101398 12764 101404 12776
rect 99248 12736 101404 12764
rect 99248 12724 99254 12736
rect 101398 12724 101404 12736
rect 101456 12724 101462 12776
rect 101674 12764 101680 12776
rect 101635 12736 101680 12764
rect 101674 12724 101680 12736
rect 101732 12724 101738 12776
rect 104805 12767 104863 12773
rect 104805 12733 104817 12767
rect 104851 12733 104863 12767
rect 104805 12727 104863 12733
rect 100941 12699 100999 12705
rect 98564 12668 99328 12696
rect 87782 12628 87788 12640
rect 86144 12600 87788 12628
rect 87782 12588 87788 12600
rect 87840 12588 87846 12640
rect 87966 12628 87972 12640
rect 87927 12600 87972 12628
rect 87966 12588 87972 12600
rect 88024 12588 88030 12640
rect 88426 12588 88432 12640
rect 88484 12628 88490 12640
rect 89165 12631 89223 12637
rect 89165 12628 89177 12631
rect 88484 12600 89177 12628
rect 88484 12588 88490 12600
rect 89165 12597 89177 12600
rect 89211 12597 89223 12631
rect 89898 12628 89904 12640
rect 89811 12600 89904 12628
rect 89165 12591 89223 12597
rect 89898 12588 89904 12600
rect 89956 12628 89962 12640
rect 90545 12631 90603 12637
rect 90545 12628 90557 12631
rect 89956 12600 90557 12628
rect 89956 12588 89962 12600
rect 90545 12597 90557 12600
rect 90591 12597 90603 12631
rect 90545 12591 90603 12597
rect 98365 12631 98423 12637
rect 98365 12597 98377 12631
rect 98411 12628 98423 12631
rect 99190 12628 99196 12640
rect 98411 12600 99196 12628
rect 98411 12597 98423 12600
rect 98365 12591 98423 12597
rect 99190 12588 99196 12600
rect 99248 12588 99254 12640
rect 99300 12628 99328 12668
rect 100941 12665 100953 12699
rect 100987 12696 100999 12699
rect 101030 12696 101036 12708
rect 100987 12668 101036 12696
rect 100987 12665 100999 12668
rect 100941 12659 100999 12665
rect 101030 12656 101036 12668
rect 101088 12656 101094 12708
rect 103238 12656 103244 12708
rect 103296 12696 103302 12708
rect 104820 12696 104848 12727
rect 105906 12696 105912 12708
rect 103296 12668 104848 12696
rect 105867 12668 105912 12696
rect 103296 12656 103302 12668
rect 105906 12656 105912 12668
rect 105964 12656 105970 12708
rect 108316 12696 108344 12940
rect 111426 12928 111432 12980
rect 111484 12968 111490 12980
rect 112257 12971 112315 12977
rect 112257 12968 112269 12971
rect 111484 12940 112269 12968
rect 111484 12928 111490 12940
rect 112257 12937 112269 12940
rect 112303 12968 112315 12971
rect 114554 12968 114560 12980
rect 112303 12940 114560 12968
rect 112303 12937 112315 12940
rect 112257 12931 112315 12937
rect 114554 12928 114560 12940
rect 114612 12928 114618 12980
rect 114738 12928 114744 12980
rect 114796 12968 114802 12980
rect 117406 12968 117412 12980
rect 114796 12940 117412 12968
rect 114796 12928 114802 12940
rect 117406 12928 117412 12940
rect 117464 12928 117470 12980
rect 118234 12968 118240 12980
rect 118195 12940 118240 12968
rect 118234 12928 118240 12940
rect 118292 12928 118298 12980
rect 118694 12968 118700 12980
rect 118655 12940 118700 12968
rect 118694 12928 118700 12940
rect 118752 12928 118758 12980
rect 126701 12971 126759 12977
rect 126701 12937 126713 12971
rect 126747 12968 126759 12971
rect 126882 12968 126888 12980
rect 126747 12940 126888 12968
rect 126747 12937 126759 12940
rect 126701 12931 126759 12937
rect 126882 12928 126888 12940
rect 126940 12928 126946 12980
rect 128078 12968 128084 12980
rect 128039 12940 128084 12968
rect 128078 12928 128084 12940
rect 128136 12928 128142 12980
rect 128630 12928 128636 12980
rect 128688 12968 128694 12980
rect 128725 12971 128783 12977
rect 128725 12968 128737 12971
rect 128688 12940 128737 12968
rect 128688 12928 128694 12940
rect 128725 12937 128737 12940
rect 128771 12937 128783 12971
rect 129182 12968 129188 12980
rect 129143 12940 129188 12968
rect 128725 12931 128783 12937
rect 129182 12928 129188 12940
rect 129240 12928 129246 12980
rect 130289 12971 130347 12977
rect 130289 12937 130301 12971
rect 130335 12968 130347 12971
rect 133322 12968 133328 12980
rect 130335 12940 133328 12968
rect 130335 12937 130347 12940
rect 130289 12931 130347 12937
rect 133322 12928 133328 12940
rect 133380 12928 133386 12980
rect 133509 12971 133567 12977
rect 133509 12937 133521 12971
rect 133555 12968 133567 12971
rect 133555 12940 133828 12968
rect 133555 12937 133567 12940
rect 133509 12931 133567 12937
rect 109586 12860 109592 12912
rect 109644 12900 109650 12912
rect 112349 12903 112407 12909
rect 112349 12900 112361 12903
rect 109644 12872 112361 12900
rect 109644 12860 109650 12872
rect 112349 12869 112361 12872
rect 112395 12869 112407 12903
rect 114005 12903 114063 12909
rect 114005 12900 114017 12903
rect 112349 12863 112407 12869
rect 112548 12872 114017 12900
rect 112548 12773 112576 12872
rect 114005 12869 114017 12872
rect 114051 12900 114063 12903
rect 115661 12903 115719 12909
rect 114051 12872 115612 12900
rect 114051 12869 114063 12872
rect 114005 12863 114063 12869
rect 113082 12832 113088 12844
rect 113043 12804 113088 12832
rect 113082 12792 113088 12804
rect 113140 12792 113146 12844
rect 113818 12832 113824 12844
rect 113779 12804 113824 12832
rect 113818 12792 113824 12804
rect 113876 12792 113882 12844
rect 114646 12792 114652 12844
rect 114704 12832 114710 12844
rect 115584 12832 115612 12872
rect 115661 12869 115673 12903
rect 115707 12900 115719 12903
rect 115750 12900 115756 12912
rect 115707 12872 115756 12900
rect 115707 12869 115719 12872
rect 115661 12863 115719 12869
rect 115750 12860 115756 12872
rect 115808 12860 115814 12912
rect 117314 12860 117320 12912
rect 117372 12860 117378 12912
rect 126514 12860 126520 12912
rect 126572 12900 126578 12912
rect 129200 12900 129228 12928
rect 132402 12900 132408 12912
rect 126572 12872 129228 12900
rect 132342 12872 132408 12900
rect 126572 12860 126578 12872
rect 114704 12804 114749 12832
rect 115584 12804 115888 12832
rect 114704 12792 114710 12804
rect 115860 12776 115888 12804
rect 118050 12792 118056 12844
rect 118108 12832 118114 12844
rect 126900 12841 126928 12872
rect 132402 12860 132408 12872
rect 132460 12860 132466 12912
rect 133598 12900 133604 12912
rect 133559 12872 133604 12900
rect 133598 12860 133604 12872
rect 133656 12860 133662 12912
rect 133800 12900 133828 12940
rect 133874 12928 133880 12980
rect 133932 12968 133938 12980
rect 134337 12971 134395 12977
rect 134337 12968 134349 12971
rect 133932 12940 134349 12968
rect 133932 12928 133938 12940
rect 134337 12937 134349 12940
rect 134383 12937 134395 12971
rect 134337 12931 134395 12937
rect 145469 12971 145527 12977
rect 145469 12937 145481 12971
rect 145515 12968 145527 12971
rect 147674 12968 147680 12980
rect 145515 12940 147680 12968
rect 145515 12937 145527 12940
rect 145469 12931 145527 12937
rect 147674 12928 147680 12940
rect 147732 12928 147738 12980
rect 151449 12971 151507 12977
rect 148152 12940 149836 12968
rect 134150 12900 134156 12912
rect 133800 12872 134156 12900
rect 134150 12860 134156 12872
rect 134208 12860 134214 12912
rect 143074 12860 143080 12912
rect 143132 12900 143138 12912
rect 145926 12900 145932 12912
rect 143132 12872 145788 12900
rect 145887 12872 145932 12900
rect 143132 12860 143138 12872
rect 118881 12835 118939 12841
rect 118881 12832 118893 12835
rect 118108 12804 118893 12832
rect 118108 12792 118114 12804
rect 118881 12801 118893 12804
rect 118927 12801 118939 12835
rect 118881 12795 118939 12801
rect 126885 12835 126943 12841
rect 126885 12801 126897 12835
rect 126931 12801 126943 12835
rect 127434 12832 127440 12844
rect 127395 12804 127440 12832
rect 126885 12795 126943 12801
rect 127434 12792 127440 12804
rect 127492 12832 127498 12844
rect 128265 12835 128323 12841
rect 127492 12804 128216 12832
rect 127492 12792 127498 12804
rect 112533 12767 112591 12773
rect 112533 12733 112545 12767
rect 112579 12733 112591 12767
rect 112533 12727 112591 12733
rect 113177 12767 113235 12773
rect 113177 12733 113189 12767
rect 113223 12764 113235 12767
rect 113910 12764 113916 12776
rect 113223 12736 113916 12764
rect 113223 12733 113235 12736
rect 113177 12727 113235 12733
rect 113910 12724 113916 12736
rect 113968 12724 113974 12776
rect 114738 12724 114744 12776
rect 114796 12724 114802 12776
rect 115658 12724 115664 12776
rect 115716 12764 115722 12776
rect 115753 12767 115811 12773
rect 115753 12764 115765 12767
rect 115716 12736 115765 12764
rect 115716 12724 115722 12736
rect 115753 12733 115765 12736
rect 115799 12733 115811 12767
rect 115753 12727 115811 12733
rect 115842 12724 115848 12776
rect 115900 12764 115906 12776
rect 116489 12767 116547 12773
rect 115900 12736 115945 12764
rect 115900 12724 115906 12736
rect 116489 12733 116501 12767
rect 116535 12733 116547 12767
rect 116762 12764 116768 12776
rect 116723 12736 116768 12764
rect 116489 12727 116547 12733
rect 114756 12696 114784 12724
rect 108316 12668 114784 12696
rect 114830 12656 114836 12708
rect 114888 12696 114894 12708
rect 116504 12696 116532 12727
rect 116762 12724 116768 12736
rect 116820 12724 116826 12776
rect 127526 12764 127532 12776
rect 117792 12736 127532 12764
rect 114888 12668 116532 12696
rect 114888 12656 114894 12668
rect 100754 12628 100760 12640
rect 99300 12600 100760 12628
rect 100754 12588 100760 12600
rect 100812 12588 100818 12640
rect 103054 12588 103060 12640
rect 103112 12628 103118 12640
rect 103149 12631 103207 12637
rect 103149 12628 103161 12631
rect 103112 12600 103161 12628
rect 103112 12588 103118 12600
rect 103149 12597 103161 12600
rect 103195 12597 103207 12631
rect 103149 12591 103207 12597
rect 103606 12588 103612 12640
rect 103664 12628 103670 12640
rect 104253 12631 104311 12637
rect 104253 12628 104265 12631
rect 103664 12600 104265 12628
rect 103664 12588 103670 12600
rect 104253 12597 104265 12600
rect 104299 12597 104311 12631
rect 111886 12628 111892 12640
rect 111847 12600 111892 12628
rect 104253 12591 104311 12597
rect 111886 12588 111892 12600
rect 111944 12588 111950 12640
rect 113082 12588 113088 12640
rect 113140 12628 113146 12640
rect 114738 12628 114744 12640
rect 113140 12600 114744 12628
rect 113140 12588 113146 12600
rect 114738 12588 114744 12600
rect 114796 12588 114802 12640
rect 115293 12631 115351 12637
rect 115293 12597 115305 12631
rect 115339 12628 115351 12631
rect 115842 12628 115848 12640
rect 115339 12600 115848 12628
rect 115339 12597 115351 12600
rect 115293 12591 115351 12597
rect 115842 12588 115848 12600
rect 115900 12588 115906 12640
rect 116504 12628 116532 12668
rect 117792 12628 117820 12736
rect 127526 12724 127532 12736
rect 127584 12724 127590 12776
rect 116504 12600 117820 12628
rect 127529 12631 127587 12637
rect 127529 12597 127541 12631
rect 127575 12628 127587 12631
rect 128078 12628 128084 12640
rect 127575 12600 128084 12628
rect 127575 12597 127587 12600
rect 127529 12591 127587 12597
rect 128078 12588 128084 12600
rect 128136 12588 128142 12640
rect 128188 12628 128216 12804
rect 128265 12801 128277 12835
rect 128311 12801 128323 12835
rect 129090 12832 129096 12844
rect 129051 12804 129096 12832
rect 128265 12795 128323 12801
rect 128280 12696 128308 12795
rect 129090 12792 129096 12804
rect 129148 12792 129154 12844
rect 130197 12835 130255 12841
rect 130197 12832 130209 12835
rect 129200 12804 130209 12832
rect 128354 12724 128360 12776
rect 128412 12764 128418 12776
rect 129200 12764 129228 12804
rect 130197 12801 130209 12804
rect 130243 12801 130255 12835
rect 130197 12795 130255 12801
rect 130286 12792 130292 12844
rect 130344 12832 130350 12844
rect 130841 12835 130899 12841
rect 130841 12832 130853 12835
rect 130344 12804 130853 12832
rect 130344 12792 130350 12804
rect 130841 12801 130853 12804
rect 130887 12801 130899 12835
rect 130841 12795 130899 12801
rect 128412 12736 129228 12764
rect 129369 12767 129427 12773
rect 128412 12724 128418 12736
rect 129369 12733 129381 12767
rect 129415 12764 129427 12767
rect 129734 12764 129740 12776
rect 129415 12736 129740 12764
rect 129415 12733 129427 12736
rect 129369 12727 129427 12733
rect 129734 12724 129740 12736
rect 129792 12724 129798 12776
rect 131114 12764 131120 12776
rect 131075 12736 131120 12764
rect 131114 12724 131120 12736
rect 131172 12724 131178 12776
rect 132586 12724 132592 12776
rect 132644 12764 132650 12776
rect 133616 12764 133644 12860
rect 133690 12792 133696 12844
rect 133748 12836 133754 12844
rect 133748 12832 133828 12836
rect 134521 12835 134579 12841
rect 134521 12832 134533 12835
rect 133748 12808 134533 12832
rect 133748 12792 133754 12808
rect 133800 12804 134533 12808
rect 134521 12801 134533 12804
rect 134567 12801 134579 12835
rect 134521 12795 134579 12801
rect 135349 12835 135407 12841
rect 135349 12801 135361 12835
rect 135395 12832 135407 12835
rect 142985 12835 143043 12841
rect 142985 12832 142997 12835
rect 135395 12804 142997 12832
rect 135395 12801 135407 12804
rect 135349 12795 135407 12801
rect 142985 12801 142997 12804
rect 143031 12832 143043 12835
rect 145760 12832 145788 12872
rect 145926 12860 145932 12872
rect 145984 12860 145990 12912
rect 148152 12900 148180 12940
rect 146036 12872 148180 12900
rect 149808 12900 149836 12940
rect 151449 12937 151461 12971
rect 151495 12968 151507 12971
rect 152642 12968 152648 12980
rect 151495 12940 152648 12968
rect 151495 12937 151507 12940
rect 151449 12931 151507 12937
rect 152642 12928 152648 12940
rect 152700 12928 152706 12980
rect 152737 12971 152795 12977
rect 152737 12937 152749 12971
rect 152783 12968 152795 12971
rect 152826 12968 152832 12980
rect 152783 12940 152832 12968
rect 152783 12937 152795 12940
rect 152737 12931 152795 12937
rect 152826 12928 152832 12940
rect 152884 12968 152890 12980
rect 153105 12971 153163 12977
rect 153105 12968 153117 12971
rect 152884 12940 153117 12968
rect 152884 12928 152890 12940
rect 153105 12937 153117 12940
rect 153151 12968 153163 12971
rect 153473 12971 153531 12977
rect 153473 12968 153485 12971
rect 153151 12940 153485 12968
rect 153151 12937 153163 12940
rect 153105 12931 153163 12937
rect 153473 12937 153485 12940
rect 153519 12968 153531 12971
rect 153841 12971 153899 12977
rect 153841 12968 153853 12971
rect 153519 12940 153853 12968
rect 153519 12937 153531 12940
rect 153473 12931 153531 12937
rect 153841 12937 153853 12940
rect 153887 12968 153899 12971
rect 154209 12971 154267 12977
rect 154209 12968 154221 12971
rect 153887 12940 154221 12968
rect 153887 12937 153899 12940
rect 153841 12931 153899 12937
rect 154209 12937 154221 12940
rect 154255 12968 154267 12971
rect 154945 12971 155003 12977
rect 154945 12968 154957 12971
rect 154255 12940 154957 12968
rect 154255 12937 154267 12940
rect 154209 12931 154267 12937
rect 154945 12937 154957 12940
rect 154991 12968 155003 12971
rect 156049 12971 156107 12977
rect 156049 12968 156061 12971
rect 154991 12940 156061 12968
rect 154991 12937 155003 12940
rect 154945 12931 155003 12937
rect 156049 12937 156061 12940
rect 156095 12968 156107 12971
rect 156417 12971 156475 12977
rect 156417 12968 156429 12971
rect 156095 12940 156429 12968
rect 156095 12937 156107 12940
rect 156049 12931 156107 12937
rect 156417 12937 156429 12940
rect 156463 12968 156475 12971
rect 156785 12971 156843 12977
rect 156785 12968 156797 12971
rect 156463 12940 156797 12968
rect 156463 12937 156475 12940
rect 156417 12931 156475 12937
rect 156785 12937 156797 12940
rect 156831 12968 156843 12971
rect 157150 12968 157156 12980
rect 156831 12940 157156 12968
rect 156831 12937 156843 12940
rect 156785 12931 156843 12937
rect 157150 12928 157156 12940
rect 157208 12928 157214 12980
rect 158622 12928 158628 12980
rect 158680 12968 158686 12980
rect 163498 12968 163504 12980
rect 158680 12940 163504 12968
rect 158680 12928 158686 12940
rect 156598 12900 156604 12912
rect 149808 12872 156604 12900
rect 145834 12832 145840 12844
rect 143031 12804 145696 12832
rect 145747 12804 145840 12832
rect 143031 12801 143043 12804
rect 142985 12795 143043 12801
rect 132644 12736 133644 12764
rect 133785 12767 133843 12773
rect 132644 12724 132650 12736
rect 133785 12733 133797 12767
rect 133831 12733 133843 12767
rect 143258 12764 143264 12776
rect 143219 12736 143264 12764
rect 133785 12727 133843 12733
rect 130286 12696 130292 12708
rect 128280 12668 130292 12696
rect 130286 12656 130292 12668
rect 130344 12656 130350 12708
rect 133690 12696 133696 12708
rect 132466 12668 133696 12696
rect 132466 12628 132494 12668
rect 133690 12656 133696 12668
rect 133748 12656 133754 12708
rect 133138 12628 133144 12640
rect 128188 12600 132494 12628
rect 133099 12600 133144 12628
rect 133138 12588 133144 12600
rect 133196 12588 133202 12640
rect 133230 12588 133236 12640
rect 133288 12628 133294 12640
rect 133800 12628 133828 12727
rect 143258 12724 143264 12736
rect 143316 12724 143322 12776
rect 145668 12764 145696 12804
rect 145834 12792 145840 12804
rect 145892 12792 145898 12844
rect 146036 12832 146064 12872
rect 156598 12860 156604 12872
rect 156656 12860 156662 12912
rect 159269 12903 159327 12909
rect 159269 12900 159281 12903
rect 157306 12872 159281 12900
rect 145944 12804 146064 12832
rect 147033 12835 147091 12841
rect 145944 12764 145972 12804
rect 147033 12801 147045 12835
rect 147079 12832 147091 12835
rect 147306 12832 147312 12844
rect 147079 12804 147312 12832
rect 147079 12801 147091 12804
rect 147033 12795 147091 12801
rect 147306 12792 147312 12804
rect 147364 12792 147370 12844
rect 148902 12804 149008 12832
rect 148980 12776 149008 12804
rect 149330 12792 149336 12844
rect 149388 12832 149394 12844
rect 149885 12835 149943 12841
rect 149885 12832 149897 12835
rect 149388 12804 149897 12832
rect 149388 12792 149394 12804
rect 149885 12801 149897 12804
rect 149931 12832 149943 12835
rect 149931 12804 150388 12832
rect 149931 12801 149943 12804
rect 149885 12795 149943 12801
rect 145668 12736 145972 12764
rect 146113 12767 146171 12773
rect 146113 12733 146125 12767
rect 146159 12764 146171 12767
rect 147398 12764 147404 12776
rect 146159 12736 147404 12764
rect 146159 12733 146171 12736
rect 146113 12727 146171 12733
rect 147398 12724 147404 12736
rect 147456 12724 147462 12776
rect 147493 12767 147551 12773
rect 147493 12733 147505 12767
rect 147539 12733 147551 12767
rect 147766 12764 147772 12776
rect 147727 12736 147772 12764
rect 147493 12727 147551 12733
rect 133874 12656 133880 12708
rect 133932 12696 133938 12708
rect 135533 12699 135591 12705
rect 135533 12696 135545 12699
rect 133932 12668 135545 12696
rect 133932 12656 133938 12668
rect 135533 12665 135545 12668
rect 135579 12665 135591 12699
rect 135533 12659 135591 12665
rect 145742 12656 145748 12708
rect 145800 12696 145806 12708
rect 147508 12696 147536 12727
rect 147766 12724 147772 12736
rect 147824 12724 147830 12776
rect 148962 12724 148968 12776
rect 149020 12724 149026 12776
rect 149238 12764 149244 12776
rect 149199 12736 149244 12764
rect 149238 12724 149244 12736
rect 149296 12724 149302 12776
rect 150360 12708 150388 12804
rect 150434 12792 150440 12844
rect 150492 12832 150498 12844
rect 154853 12835 154911 12841
rect 154853 12832 154865 12835
rect 150492 12804 154865 12832
rect 150492 12792 150498 12804
rect 154853 12801 154865 12804
rect 154899 12801 154911 12835
rect 154853 12795 154911 12801
rect 155862 12792 155868 12844
rect 155920 12832 155926 12844
rect 157306 12832 157334 12872
rect 159269 12869 159281 12872
rect 159315 12869 159327 12903
rect 160370 12900 160376 12912
rect 159269 12863 159327 12869
rect 159928 12872 160376 12900
rect 155920 12804 157334 12832
rect 155920 12792 155926 12804
rect 157794 12792 157800 12844
rect 157852 12832 157858 12844
rect 159177 12835 159235 12841
rect 159177 12832 159189 12835
rect 157852 12804 159189 12832
rect 157852 12792 157858 12804
rect 159177 12801 159189 12804
rect 159223 12832 159235 12835
rect 159928 12832 159956 12872
rect 160370 12860 160376 12872
rect 160428 12860 160434 12912
rect 161124 12872 161796 12900
rect 159223 12804 159956 12832
rect 160005 12835 160063 12841
rect 159223 12801 159235 12804
rect 159177 12795 159235 12801
rect 160005 12801 160017 12835
rect 160051 12832 160063 12835
rect 161124 12832 161152 12872
rect 160051 12804 161152 12832
rect 161201 12835 161259 12841
rect 160051 12801 160063 12804
rect 160005 12795 160063 12801
rect 161201 12801 161213 12835
rect 161247 12832 161259 12835
rect 161658 12832 161664 12844
rect 161247 12804 161664 12832
rect 161247 12801 161259 12804
rect 161201 12795 161259 12801
rect 161658 12792 161664 12804
rect 161716 12792 161722 12844
rect 151538 12764 151544 12776
rect 151499 12736 151544 12764
rect 151538 12724 151544 12736
rect 151596 12724 151602 12776
rect 151725 12767 151783 12773
rect 151725 12733 151737 12767
rect 151771 12733 151783 12767
rect 151725 12727 151783 12733
rect 145800 12668 147536 12696
rect 145800 12656 145806 12668
rect 150342 12656 150348 12708
rect 150400 12696 150406 12708
rect 151630 12696 151636 12708
rect 150400 12668 151636 12696
rect 150400 12656 150406 12668
rect 151630 12656 151636 12668
rect 151688 12656 151694 12708
rect 133288 12600 133828 12628
rect 146849 12631 146907 12637
rect 133288 12588 133294 12600
rect 146849 12597 146861 12631
rect 146895 12628 146907 12631
rect 148502 12628 148508 12640
rect 146895 12600 148508 12628
rect 146895 12597 146907 12600
rect 146849 12591 146907 12597
rect 148502 12588 148508 12600
rect 148560 12588 148566 12640
rect 149974 12628 149980 12640
rect 149935 12600 149980 12628
rect 149974 12588 149980 12600
rect 150032 12588 150038 12640
rect 151081 12631 151139 12637
rect 151081 12597 151093 12631
rect 151127 12628 151139 12631
rect 151262 12628 151268 12640
rect 151127 12600 151268 12628
rect 151127 12597 151139 12600
rect 151081 12591 151139 12597
rect 151262 12588 151268 12600
rect 151320 12588 151326 12640
rect 151354 12588 151360 12640
rect 151412 12628 151418 12640
rect 151740 12628 151768 12727
rect 152734 12724 152740 12776
rect 152792 12764 152798 12776
rect 152792 12736 154988 12764
rect 152792 12724 152798 12736
rect 152369 12699 152427 12705
rect 152369 12665 152381 12699
rect 152415 12696 152427 12699
rect 152826 12696 152832 12708
rect 152415 12668 152832 12696
rect 152415 12665 152427 12668
rect 152369 12659 152427 12665
rect 152826 12656 152832 12668
rect 152884 12656 152890 12708
rect 153102 12656 153108 12708
rect 153160 12696 153166 12708
rect 154485 12699 154543 12705
rect 154485 12696 154497 12699
rect 153160 12668 154497 12696
rect 153160 12656 153166 12668
rect 154485 12665 154497 12668
rect 154531 12665 154543 12699
rect 154960 12696 154988 12736
rect 155034 12724 155040 12776
rect 155092 12764 155098 12776
rect 159450 12764 159456 12776
rect 155092 12736 155137 12764
rect 155236 12736 159312 12764
rect 159411 12736 159456 12764
rect 155092 12724 155098 12736
rect 155236 12696 155264 12736
rect 158806 12696 158812 12708
rect 154960 12668 155264 12696
rect 158767 12668 158812 12696
rect 154485 12659 154543 12665
rect 158806 12656 158812 12668
rect 158864 12656 158870 12708
rect 159284 12696 159312 12736
rect 159450 12724 159456 12736
rect 159508 12724 159514 12776
rect 159542 12724 159548 12776
rect 159600 12764 159606 12776
rect 161566 12764 161572 12776
rect 159600 12736 161572 12764
rect 159600 12724 159606 12736
rect 161566 12724 161572 12736
rect 161624 12724 161630 12776
rect 160189 12699 160247 12705
rect 160189 12696 160201 12699
rect 159284 12668 160201 12696
rect 160189 12665 160201 12668
rect 160235 12665 160247 12699
rect 160189 12659 160247 12665
rect 154114 12628 154120 12640
rect 151412 12600 154120 12628
rect 151412 12588 151418 12600
rect 154114 12588 154120 12600
rect 154172 12628 154178 12640
rect 157886 12628 157892 12640
rect 154172 12600 157892 12628
rect 154172 12588 154178 12600
rect 157886 12588 157892 12600
rect 157944 12588 157950 12640
rect 160278 12588 160284 12640
rect 160336 12628 160342 12640
rect 161293 12631 161351 12637
rect 161293 12628 161305 12631
rect 160336 12600 161305 12628
rect 160336 12588 160342 12600
rect 161293 12597 161305 12600
rect 161339 12597 161351 12631
rect 161768 12628 161796 12872
rect 161860 12841 161888 12940
rect 163498 12928 163504 12940
rect 163556 12928 163562 12980
rect 163593 12971 163651 12977
rect 163593 12937 163605 12971
rect 163639 12937 163651 12971
rect 163593 12931 163651 12937
rect 164421 12971 164479 12977
rect 164421 12937 164433 12971
rect 164467 12968 164479 12971
rect 165246 12968 165252 12980
rect 164467 12940 165252 12968
rect 164467 12937 164479 12940
rect 164421 12931 164479 12937
rect 163406 12900 163412 12912
rect 163346 12872 163412 12900
rect 163406 12860 163412 12872
rect 163464 12860 163470 12912
rect 163608 12900 163636 12931
rect 165246 12928 165252 12940
rect 165304 12968 165310 12980
rect 165304 12940 166994 12968
rect 165304 12928 165310 12940
rect 164513 12903 164571 12909
rect 164513 12900 164525 12903
rect 163608 12872 164525 12900
rect 161845 12835 161903 12841
rect 161845 12801 161857 12835
rect 161891 12801 161903 12835
rect 161845 12795 161903 12801
rect 162118 12764 162124 12776
rect 162079 12736 162124 12764
rect 162118 12724 162124 12736
rect 162176 12724 162182 12776
rect 162854 12724 162860 12776
rect 162912 12764 162918 12776
rect 163608 12764 163636 12872
rect 164513 12869 164525 12872
rect 164559 12900 164571 12903
rect 166966 12900 166994 12940
rect 167178 12928 167184 12980
rect 167236 12968 167242 12980
rect 167825 12971 167883 12977
rect 167825 12968 167837 12971
rect 167236 12940 167837 12968
rect 167236 12928 167242 12940
rect 167825 12937 167837 12940
rect 167871 12937 167883 12971
rect 174998 12968 175004 12980
rect 174959 12940 175004 12968
rect 167825 12931 167883 12937
rect 174998 12928 175004 12940
rect 175056 12928 175062 12980
rect 175645 12971 175703 12977
rect 175645 12937 175657 12971
rect 175691 12968 175703 12971
rect 175734 12968 175740 12980
rect 175691 12940 175740 12968
rect 175691 12937 175703 12940
rect 175645 12931 175703 12937
rect 175734 12928 175740 12940
rect 175792 12928 175798 12980
rect 176378 12928 176384 12980
rect 176436 12968 176442 12980
rect 180150 12968 180156 12980
rect 176436 12940 180156 12968
rect 176436 12928 176442 12940
rect 164559 12872 166672 12900
rect 166966 12872 168052 12900
rect 164559 12869 164571 12872
rect 164513 12863 164571 12869
rect 165341 12835 165399 12841
rect 165341 12801 165353 12835
rect 165387 12832 165399 12835
rect 165430 12832 165436 12844
rect 165387 12804 165436 12832
rect 165387 12801 165399 12804
rect 165341 12795 165399 12801
rect 165430 12792 165436 12804
rect 165488 12792 165494 12844
rect 166166 12792 166172 12844
rect 166224 12832 166230 12844
rect 166534 12832 166540 12844
rect 166224 12804 166540 12832
rect 166224 12792 166230 12804
rect 166534 12792 166540 12804
rect 166592 12792 166598 12844
rect 166644 12832 166672 12872
rect 168024 12841 168052 12872
rect 173802 12860 173808 12912
rect 173860 12900 173866 12912
rect 173860 12872 175872 12900
rect 173860 12860 173866 12872
rect 175844 12841 175872 12872
rect 175918 12860 175924 12912
rect 175976 12900 175982 12912
rect 176930 12900 176936 12912
rect 175976 12872 176936 12900
rect 175976 12860 175982 12872
rect 176930 12860 176936 12872
rect 176988 12860 176994 12912
rect 177942 12900 177948 12912
rect 177882 12872 177948 12900
rect 177942 12860 177948 12872
rect 178000 12860 178006 12912
rect 167365 12835 167423 12841
rect 167365 12832 167377 12835
rect 166644 12804 167377 12832
rect 167365 12801 167377 12804
rect 167411 12801 167423 12835
rect 167365 12795 167423 12801
rect 168009 12835 168067 12841
rect 168009 12801 168021 12835
rect 168055 12801 168067 12835
rect 168009 12795 168067 12801
rect 175185 12835 175243 12841
rect 175185 12801 175197 12835
rect 175231 12801 175243 12835
rect 175185 12795 175243 12801
rect 175829 12835 175887 12841
rect 175829 12801 175841 12835
rect 175875 12801 175887 12835
rect 176378 12832 176384 12844
rect 176339 12804 176384 12832
rect 175829 12795 175887 12801
rect 164602 12764 164608 12776
rect 162912 12736 163636 12764
rect 164563 12736 164608 12764
rect 162912 12724 162918 12736
rect 164602 12724 164608 12736
rect 164660 12724 164666 12776
rect 163608 12668 164188 12696
rect 163608 12628 163636 12668
rect 161768 12600 163636 12628
rect 161293 12591 161351 12597
rect 163682 12588 163688 12640
rect 163740 12628 163746 12640
rect 164053 12631 164111 12637
rect 164053 12628 164065 12631
rect 163740 12600 164065 12628
rect 163740 12588 163746 12600
rect 164053 12597 164065 12600
rect 164099 12597 164111 12631
rect 164160 12628 164188 12668
rect 164234 12656 164240 12708
rect 164292 12696 164298 12708
rect 167181 12699 167239 12705
rect 167181 12696 167193 12699
rect 164292 12668 167193 12696
rect 164292 12656 164298 12668
rect 167181 12665 167193 12668
rect 167227 12665 167239 12699
rect 175200 12696 175228 12795
rect 176378 12792 176384 12804
rect 176436 12792 176442 12844
rect 178604 12841 178632 12940
rect 180150 12928 180156 12940
rect 180208 12928 180214 12980
rect 180242 12928 180248 12980
rect 180300 12968 180306 12980
rect 180797 12971 180855 12977
rect 180797 12968 180809 12971
rect 180300 12940 180809 12968
rect 180300 12928 180306 12940
rect 180797 12937 180809 12940
rect 180843 12937 180855 12971
rect 188338 12968 188344 12980
rect 180797 12931 180855 12937
rect 188080 12940 188344 12968
rect 181625 12903 181683 12909
rect 181625 12900 181637 12903
rect 180260 12872 181637 12900
rect 178589 12835 178647 12841
rect 178589 12801 178601 12835
rect 178635 12801 178647 12835
rect 180260 12832 180288 12872
rect 181625 12869 181637 12872
rect 181671 12869 181683 12903
rect 181625 12863 181683 12869
rect 179998 12804 180288 12832
rect 178589 12795 178647 12801
rect 180334 12792 180340 12844
rect 180392 12832 180398 12844
rect 180981 12835 181039 12841
rect 180981 12832 180993 12835
rect 180392 12804 180993 12832
rect 180392 12792 180398 12804
rect 180981 12801 180993 12804
rect 181027 12801 181039 12835
rect 181530 12832 181536 12844
rect 181443 12804 181536 12832
rect 180981 12795 181039 12801
rect 181530 12792 181536 12804
rect 181588 12832 181594 12844
rect 188080 12841 188108 12940
rect 188338 12928 188344 12940
rect 188396 12968 188402 12980
rect 191374 12968 191380 12980
rect 188396 12940 191380 12968
rect 188396 12928 188402 12940
rect 191374 12928 191380 12940
rect 191432 12968 191438 12980
rect 192297 12971 192355 12977
rect 192297 12968 192309 12971
rect 191432 12940 192309 12968
rect 191432 12928 191438 12940
rect 192297 12937 192309 12940
rect 192343 12937 192355 12971
rect 192297 12931 192355 12937
rect 192478 12928 192484 12980
rect 192536 12968 192542 12980
rect 192536 12940 193444 12968
rect 192536 12928 192542 12940
rect 188522 12860 188528 12912
rect 188580 12900 188586 12912
rect 189537 12903 189595 12909
rect 189537 12900 189549 12903
rect 188580 12872 189549 12900
rect 188580 12860 188586 12872
rect 189537 12869 189549 12872
rect 189583 12900 189595 12903
rect 190914 12900 190920 12912
rect 189583 12872 190454 12900
rect 190875 12872 190920 12900
rect 189583 12869 189595 12872
rect 189537 12863 189595 12869
rect 182177 12835 182235 12841
rect 182177 12832 182189 12835
rect 181588 12804 182189 12832
rect 181588 12792 181594 12804
rect 182177 12801 182189 12804
rect 182223 12801 182235 12835
rect 182177 12795 182235 12801
rect 188065 12835 188123 12841
rect 188065 12801 188077 12835
rect 188111 12801 188123 12835
rect 188065 12795 188123 12801
rect 188338 12792 188344 12844
rect 188396 12832 188402 12844
rect 188617 12835 188675 12841
rect 188617 12832 188629 12835
rect 188396 12804 188629 12832
rect 188396 12792 188402 12804
rect 188617 12801 188629 12804
rect 188663 12832 188675 12835
rect 188798 12832 188804 12844
rect 188663 12804 188804 12832
rect 188663 12801 188675 12804
rect 188617 12795 188675 12801
rect 188798 12792 188804 12804
rect 188856 12792 188862 12844
rect 189350 12832 189356 12844
rect 189311 12804 189356 12832
rect 189350 12792 189356 12804
rect 189408 12792 189414 12844
rect 176657 12767 176715 12773
rect 176657 12733 176669 12767
rect 176703 12764 176715 12767
rect 176746 12764 176752 12776
rect 176703 12736 176752 12764
rect 176703 12733 176715 12736
rect 176657 12727 176715 12733
rect 176746 12724 176752 12736
rect 176804 12724 176810 12776
rect 178865 12767 178923 12773
rect 178865 12733 178877 12767
rect 178911 12764 178923 12767
rect 178911 12736 180104 12764
rect 178911 12733 178923 12736
rect 178865 12727 178923 12733
rect 180076 12696 180104 12736
rect 180150 12724 180156 12776
rect 180208 12764 180214 12776
rect 189534 12764 189540 12776
rect 180208 12736 189540 12764
rect 180208 12724 180214 12736
rect 189534 12724 189540 12736
rect 189592 12724 189598 12776
rect 190426 12764 190454 12872
rect 190914 12860 190920 12872
rect 190972 12860 190978 12912
rect 191742 12860 191748 12912
rect 191800 12900 191806 12912
rect 193309 12903 193367 12909
rect 193309 12900 193321 12903
rect 191800 12872 193321 12900
rect 191800 12860 191806 12872
rect 193309 12869 193321 12872
rect 193355 12869 193367 12903
rect 193416 12900 193444 12940
rect 193950 12928 193956 12980
rect 194008 12968 194014 12980
rect 194870 12968 194876 12980
rect 194008 12940 194876 12968
rect 194008 12928 194014 12940
rect 194870 12928 194876 12940
rect 194928 12968 194934 12980
rect 195974 12968 195980 12980
rect 194928 12940 195980 12968
rect 194928 12928 194934 12940
rect 195974 12928 195980 12940
rect 196032 12928 196038 12980
rect 197722 12928 197728 12980
rect 197780 12968 197786 12980
rect 197780 12940 206508 12968
rect 197780 12928 197786 12940
rect 195885 12903 195943 12909
rect 195885 12900 195897 12903
rect 193416 12872 193798 12900
rect 195072 12872 195897 12900
rect 193309 12863 193367 12869
rect 195072 12844 195100 12872
rect 195885 12869 195897 12872
rect 195931 12869 195943 12903
rect 202966 12900 202972 12912
rect 195885 12863 195943 12869
rect 202524 12872 202972 12900
rect 191009 12835 191067 12841
rect 191009 12801 191021 12835
rect 191055 12832 191067 12835
rect 192205 12835 192263 12841
rect 192205 12832 192217 12835
rect 191055 12804 192217 12832
rect 191055 12801 191067 12804
rect 191009 12795 191067 12801
rect 192205 12801 192217 12804
rect 192251 12832 192263 12835
rect 192570 12832 192576 12844
rect 192251 12804 192576 12832
rect 192251 12801 192263 12804
rect 192205 12795 192263 12801
rect 192570 12792 192576 12804
rect 192628 12792 192634 12844
rect 195054 12832 195060 12844
rect 195015 12804 195060 12832
rect 195054 12792 195060 12804
rect 195112 12792 195118 12844
rect 197354 12832 197360 12844
rect 197315 12804 197360 12832
rect 197354 12792 197360 12804
rect 197412 12792 197418 12844
rect 197446 12792 197452 12844
rect 197504 12832 197510 12844
rect 198366 12832 198372 12844
rect 197504 12804 198136 12832
rect 198327 12804 198372 12832
rect 197504 12792 197510 12804
rect 191193 12767 191251 12773
rect 191193 12764 191205 12767
rect 190426 12736 191205 12764
rect 191193 12733 191205 12736
rect 191239 12764 191251 12767
rect 192389 12767 192447 12773
rect 192389 12764 192401 12767
rect 191239 12736 192401 12764
rect 191239 12733 191251 12736
rect 191193 12727 191251 12733
rect 192389 12733 192401 12736
rect 192435 12764 192447 12767
rect 192662 12764 192668 12776
rect 192435 12736 192668 12764
rect 192435 12733 192447 12736
rect 192389 12727 192447 12733
rect 192662 12724 192668 12736
rect 192720 12724 192726 12776
rect 193030 12764 193036 12776
rect 192991 12736 193036 12764
rect 193030 12724 193036 12736
rect 193088 12724 193094 12776
rect 194778 12764 194784 12776
rect 193140 12736 194784 12764
rect 180242 12696 180248 12708
rect 175200 12668 176148 12696
rect 180076 12668 180248 12696
rect 167181 12659 167239 12665
rect 165433 12631 165491 12637
rect 165433 12628 165445 12631
rect 164160 12600 165445 12628
rect 164053 12591 164111 12597
rect 165433 12597 165445 12600
rect 165479 12628 165491 12631
rect 166166 12628 166172 12640
rect 165479 12600 166172 12628
rect 165479 12597 165491 12600
rect 165433 12591 165491 12597
rect 166166 12588 166172 12600
rect 166224 12588 166230 12640
rect 166626 12628 166632 12640
rect 166587 12600 166632 12628
rect 166626 12588 166632 12600
rect 166684 12588 166690 12640
rect 176120 12628 176148 12668
rect 180242 12656 180248 12668
rect 180300 12656 180306 12708
rect 180518 12656 180524 12708
rect 180576 12696 180582 12708
rect 182082 12696 182088 12708
rect 180576 12668 182088 12696
rect 180576 12656 180582 12668
rect 182082 12656 182088 12668
rect 182140 12656 182146 12708
rect 187881 12699 187939 12705
rect 187881 12665 187893 12699
rect 187927 12696 187939 12699
rect 188614 12696 188620 12708
rect 187927 12668 188620 12696
rect 187927 12665 187939 12668
rect 187881 12659 187939 12665
rect 188614 12656 188620 12668
rect 188672 12656 188678 12708
rect 189166 12656 189172 12708
rect 189224 12696 189230 12708
rect 191742 12696 191748 12708
rect 189224 12668 191748 12696
rect 189224 12656 189230 12668
rect 191742 12656 191748 12668
rect 191800 12656 191806 12708
rect 191926 12656 191932 12708
rect 191984 12696 191990 12708
rect 192478 12696 192484 12708
rect 191984 12668 192484 12696
rect 191984 12656 191990 12668
rect 192478 12656 192484 12668
rect 192536 12656 192542 12708
rect 193140 12696 193168 12736
rect 194778 12724 194784 12736
rect 194836 12724 194842 12776
rect 195790 12724 195796 12776
rect 195848 12764 195854 12776
rect 196161 12767 196219 12773
rect 196161 12764 196173 12767
rect 195848 12736 196173 12764
rect 195848 12724 195854 12736
rect 196161 12733 196173 12736
rect 196207 12764 196219 12767
rect 197630 12764 197636 12776
rect 196207 12736 197636 12764
rect 196207 12733 196219 12736
rect 196161 12727 196219 12733
rect 197630 12724 197636 12736
rect 197688 12724 197694 12776
rect 198108 12773 198136 12804
rect 198366 12792 198372 12804
rect 198424 12792 198430 12844
rect 200485 12835 200543 12841
rect 200485 12801 200497 12835
rect 200531 12832 200543 12835
rect 200666 12832 200672 12844
rect 200531 12804 200672 12832
rect 200531 12801 200543 12804
rect 200485 12795 200543 12801
rect 200666 12792 200672 12804
rect 200724 12792 200730 12844
rect 201310 12832 201316 12844
rect 201271 12804 201316 12832
rect 201310 12792 201316 12804
rect 201368 12792 201374 12844
rect 198093 12767 198151 12773
rect 198093 12733 198105 12767
rect 198139 12764 198151 12767
rect 198550 12764 198556 12776
rect 198139 12736 198556 12764
rect 198139 12733 198151 12736
rect 198093 12727 198151 12733
rect 198550 12724 198556 12736
rect 198608 12764 198614 12776
rect 200390 12764 200396 12776
rect 198608 12736 200396 12764
rect 198608 12724 198614 12736
rect 200390 12724 200396 12736
rect 200448 12724 200454 12776
rect 200577 12767 200635 12773
rect 200577 12733 200589 12767
rect 200623 12764 200635 12767
rect 202524 12764 202552 12872
rect 202966 12860 202972 12872
rect 203024 12860 203030 12912
rect 203334 12860 203340 12912
rect 203392 12860 203398 12912
rect 204824 12841 204852 12940
rect 205634 12860 205640 12912
rect 205692 12860 205698 12912
rect 204809 12835 204867 12841
rect 204809 12801 204821 12835
rect 204855 12801 204867 12835
rect 206480 12832 206508 12940
rect 206554 12928 206560 12980
rect 206612 12968 206618 12980
rect 207382 12968 207388 12980
rect 206612 12940 207388 12968
rect 206612 12928 206618 12940
rect 207382 12928 207388 12940
rect 207440 12928 207446 12980
rect 207842 12928 207848 12980
rect 207900 12968 207906 12980
rect 207900 12940 219756 12968
rect 207900 12928 207906 12940
rect 206664 12872 207612 12900
rect 206664 12832 206692 12872
rect 206480 12804 206692 12832
rect 207477 12835 207535 12841
rect 204809 12795 204867 12801
rect 207477 12801 207489 12835
rect 207523 12801 207535 12835
rect 207477 12795 207535 12801
rect 200623 12736 202552 12764
rect 202601 12767 202659 12773
rect 200623 12733 200635 12736
rect 200577 12727 200635 12733
rect 202601 12733 202613 12767
rect 202647 12733 202659 12767
rect 202874 12764 202880 12776
rect 202835 12736 202880 12764
rect 202601 12727 202659 12733
rect 202138 12696 202144 12708
rect 192588 12668 193168 12696
rect 194336 12668 202144 12696
rect 177390 12628 177396 12640
rect 176120 12600 177396 12628
rect 177390 12588 177396 12600
rect 177448 12588 177454 12640
rect 177850 12588 177856 12640
rect 177908 12628 177914 12640
rect 178129 12631 178187 12637
rect 178129 12628 178141 12631
rect 177908 12600 178141 12628
rect 177908 12588 177914 12600
rect 178129 12597 178141 12600
rect 178175 12597 178187 12631
rect 178129 12591 178187 12597
rect 179874 12588 179880 12640
rect 179932 12628 179938 12640
rect 180337 12631 180395 12637
rect 180337 12628 180349 12631
rect 179932 12600 180349 12628
rect 179932 12588 179938 12600
rect 180337 12597 180349 12600
rect 180383 12628 180395 12631
rect 180610 12628 180616 12640
rect 180383 12600 180616 12628
rect 180383 12597 180395 12600
rect 180337 12591 180395 12597
rect 180610 12588 180616 12600
rect 180668 12588 180674 12640
rect 181438 12588 181444 12640
rect 181496 12628 181502 12640
rect 182269 12631 182327 12637
rect 182269 12628 182281 12631
rect 181496 12600 182281 12628
rect 181496 12588 181502 12600
rect 182269 12597 182281 12600
rect 182315 12597 182327 12631
rect 182269 12591 182327 12597
rect 187786 12588 187792 12640
rect 187844 12628 187850 12640
rect 188709 12631 188767 12637
rect 188709 12628 188721 12631
rect 187844 12600 188721 12628
rect 187844 12588 187850 12600
rect 188709 12597 188721 12600
rect 188755 12628 188767 12631
rect 188982 12628 188988 12640
rect 188755 12600 188988 12628
rect 188755 12597 188767 12600
rect 188709 12591 188767 12597
rect 188982 12588 188988 12600
rect 189040 12588 189046 12640
rect 190546 12628 190552 12640
rect 190507 12600 190552 12628
rect 190546 12588 190552 12600
rect 190604 12588 190610 12640
rect 191837 12631 191895 12637
rect 191837 12597 191849 12631
rect 191883 12628 191895 12631
rect 192018 12628 192024 12640
rect 191883 12600 192024 12628
rect 191883 12597 191895 12600
rect 191837 12591 191895 12597
rect 192018 12588 192024 12600
rect 192076 12588 192082 12640
rect 192110 12588 192116 12640
rect 192168 12628 192174 12640
rect 192588 12628 192616 12668
rect 192168 12600 192616 12628
rect 192168 12588 192174 12600
rect 193030 12588 193036 12640
rect 193088 12628 193094 12640
rect 194336 12628 194364 12668
rect 202138 12656 202144 12668
rect 202196 12696 202202 12708
rect 202616 12696 202644 12727
rect 202874 12724 202880 12736
rect 202932 12724 202938 12776
rect 202966 12724 202972 12776
rect 203024 12764 203030 12776
rect 204162 12764 204168 12776
rect 203024 12736 204168 12764
rect 203024 12724 203030 12736
rect 204162 12724 204168 12736
rect 204220 12724 204226 12776
rect 205082 12764 205088 12776
rect 205043 12736 205088 12764
rect 205082 12724 205088 12736
rect 205140 12724 205146 12776
rect 205174 12724 205180 12776
rect 205232 12764 205238 12776
rect 207492 12764 207520 12795
rect 205232 12736 207520 12764
rect 207584 12764 207612 12872
rect 210602 12860 210608 12912
rect 210660 12900 210666 12912
rect 219728 12900 219756 12940
rect 219802 12928 219808 12980
rect 219860 12968 219866 12980
rect 238202 12968 238208 12980
rect 219860 12940 238208 12968
rect 219860 12928 219866 12940
rect 228266 12900 228272 12912
rect 210660 12872 217364 12900
rect 219728 12872 228272 12900
rect 210660 12860 210666 12872
rect 207658 12792 207664 12844
rect 207716 12832 207722 12844
rect 210344 12832 210464 12836
rect 216582 12832 216588 12844
rect 207716 12808 216588 12832
rect 207716 12804 210372 12808
rect 210436 12804 216588 12808
rect 207716 12792 207722 12804
rect 216582 12792 216588 12804
rect 216640 12792 216646 12844
rect 217336 12832 217364 12872
rect 228266 12860 228272 12872
rect 228324 12860 228330 12912
rect 230382 12900 230388 12912
rect 229402 12872 230388 12900
rect 230382 12860 230388 12872
rect 230440 12860 230446 12912
rect 219802 12832 219808 12844
rect 217336 12804 219808 12832
rect 219802 12792 219808 12804
rect 219860 12792 219866 12844
rect 223666 12792 223672 12844
rect 223724 12832 223730 12844
rect 226705 12835 226763 12841
rect 226705 12832 226717 12835
rect 223724 12804 226717 12832
rect 223724 12792 223730 12804
rect 226705 12801 226717 12804
rect 226751 12801 226763 12835
rect 226705 12795 226763 12801
rect 226794 12792 226800 12844
rect 226852 12832 226858 12844
rect 227349 12835 227407 12841
rect 227349 12832 227361 12835
rect 226852 12804 227361 12832
rect 226852 12792 226858 12804
rect 227349 12801 227361 12804
rect 227395 12801 227407 12835
rect 227898 12832 227904 12844
rect 227859 12804 227904 12832
rect 227349 12795 227407 12801
rect 227898 12792 227904 12804
rect 227956 12792 227962 12844
rect 230290 12832 230296 12844
rect 230251 12804 230296 12832
rect 230290 12792 230296 12804
rect 230348 12792 230354 12844
rect 230768 12841 230796 12940
rect 238202 12928 238208 12940
rect 238260 12968 238266 12980
rect 251082 12968 251088 12980
rect 238260 12940 251088 12968
rect 238260 12928 238266 12940
rect 231026 12900 231032 12912
rect 230987 12872 231032 12900
rect 231026 12860 231032 12872
rect 231084 12860 231090 12912
rect 232314 12860 232320 12912
rect 232372 12900 232378 12912
rect 238294 12900 238300 12912
rect 232372 12872 238300 12900
rect 232372 12860 232378 12872
rect 238294 12860 238300 12872
rect 238352 12860 238358 12912
rect 238588 12900 238616 12940
rect 238496 12872 238616 12900
rect 238757 12903 238815 12909
rect 230753 12835 230811 12841
rect 230753 12801 230765 12835
rect 230799 12801 230811 12835
rect 233050 12832 233056 12844
rect 232162 12804 232728 12832
rect 233011 12804 233056 12832
rect 230753 12795 230811 12801
rect 227916 12764 227944 12792
rect 228177 12767 228235 12773
rect 228177 12764 228189 12767
rect 207584 12736 215294 12764
rect 205232 12724 205238 12736
rect 207290 12696 207296 12708
rect 202196 12668 202644 12696
rect 206480 12668 206784 12696
rect 207251 12668 207296 12696
rect 202196 12656 202202 12668
rect 193088 12600 194364 12628
rect 193088 12588 193094 12600
rect 194410 12588 194416 12640
rect 194468 12628 194474 12640
rect 195517 12631 195575 12637
rect 195517 12628 195529 12631
rect 194468 12600 195529 12628
rect 194468 12588 194474 12600
rect 195517 12597 195529 12600
rect 195563 12597 195575 12631
rect 195517 12591 195575 12597
rect 195974 12588 195980 12640
rect 196032 12628 196038 12640
rect 196989 12631 197047 12637
rect 196989 12628 197001 12631
rect 196032 12600 197001 12628
rect 196032 12588 196038 12600
rect 196989 12597 197001 12600
rect 197035 12597 197047 12631
rect 198182 12628 198188 12640
rect 198143 12600 198188 12628
rect 196989 12591 197047 12597
rect 198182 12588 198188 12600
rect 198240 12588 198246 12640
rect 201126 12628 201132 12640
rect 201087 12600 201132 12628
rect 201126 12588 201132 12600
rect 201184 12588 201190 12640
rect 201954 12588 201960 12640
rect 202012 12628 202018 12640
rect 204254 12628 204260 12640
rect 202012 12600 204260 12628
rect 202012 12588 202018 12600
rect 204254 12588 204260 12600
rect 204312 12588 204318 12640
rect 204349 12631 204407 12637
rect 204349 12597 204361 12631
rect 204395 12628 204407 12631
rect 204530 12628 204536 12640
rect 204395 12600 204536 12628
rect 204395 12597 204407 12600
rect 204349 12591 204407 12597
rect 204530 12588 204536 12600
rect 204588 12628 204594 12640
rect 205174 12628 205180 12640
rect 204588 12600 205180 12628
rect 204588 12588 204594 12600
rect 205174 12588 205180 12600
rect 205232 12588 205238 12640
rect 205266 12588 205272 12640
rect 205324 12628 205330 12640
rect 206480 12628 206508 12668
rect 205324 12600 206508 12628
rect 206756 12628 206784 12668
rect 207290 12656 207296 12668
rect 207348 12656 207354 12708
rect 210602 12628 210608 12640
rect 206756 12600 210608 12628
rect 205324 12588 205330 12600
rect 210602 12588 210608 12600
rect 210660 12588 210666 12640
rect 215266 12628 215294 12736
rect 219728 12736 227944 12764
rect 228008 12736 228189 12764
rect 219728 12628 219756 12736
rect 219802 12656 219808 12708
rect 219860 12696 219866 12708
rect 227165 12699 227223 12705
rect 219860 12668 227116 12696
rect 219860 12656 219866 12668
rect 215266 12600 219756 12628
rect 226521 12631 226579 12637
rect 226521 12597 226533 12631
rect 226567 12628 226579 12631
rect 226886 12628 226892 12640
rect 226567 12600 226892 12628
rect 226567 12597 226579 12600
rect 226521 12591 226579 12597
rect 226886 12588 226892 12600
rect 226944 12588 226950 12640
rect 227088 12628 227116 12668
rect 227165 12665 227177 12699
rect 227211 12696 227223 12699
rect 228008 12696 228036 12736
rect 228177 12733 228189 12736
rect 228223 12733 228235 12767
rect 228177 12727 228235 12733
rect 228266 12724 228272 12776
rect 228324 12764 228330 12776
rect 230198 12764 230204 12776
rect 228324 12736 230204 12764
rect 228324 12724 228330 12736
rect 230198 12724 230204 12736
rect 230256 12724 230262 12776
rect 232700 12764 232728 12804
rect 233050 12792 233056 12804
rect 233108 12792 233114 12844
rect 237006 12832 237012 12844
rect 236967 12804 237012 12832
rect 237006 12792 237012 12804
rect 237064 12792 237070 12844
rect 237653 12835 237711 12841
rect 237653 12801 237665 12835
rect 237699 12832 237711 12835
rect 238386 12832 238392 12844
rect 237699 12804 238392 12832
rect 237699 12801 237711 12804
rect 237653 12795 237711 12801
rect 238386 12792 238392 12804
rect 238444 12792 238450 12844
rect 238496 12841 238524 12872
rect 238757 12869 238769 12903
rect 238803 12900 238815 12903
rect 239030 12900 239036 12912
rect 238803 12872 239036 12900
rect 238803 12869 238815 12872
rect 238757 12863 238815 12869
rect 239030 12860 239036 12872
rect 239088 12860 239094 12912
rect 240042 12900 240048 12912
rect 239982 12872 240048 12900
rect 240042 12860 240048 12872
rect 240100 12860 240106 12912
rect 240704 12841 240732 12940
rect 251082 12928 251088 12940
rect 251140 12928 251146 12980
rect 252373 12971 252431 12977
rect 252373 12937 252385 12971
rect 252419 12968 252431 12971
rect 254670 12968 254676 12980
rect 252419 12940 254676 12968
rect 252419 12937 252431 12940
rect 252373 12931 252431 12937
rect 254670 12928 254676 12940
rect 254728 12928 254734 12980
rect 256234 12928 256240 12980
rect 256292 12968 256298 12980
rect 264606 12968 264612 12980
rect 256292 12940 263594 12968
rect 264567 12940 264612 12968
rect 256292 12928 256298 12940
rect 240962 12900 240968 12912
rect 240923 12872 240968 12900
rect 240962 12860 240968 12872
rect 241020 12860 241026 12912
rect 244642 12900 244648 12912
rect 244246 12872 244648 12900
rect 238481 12835 238539 12841
rect 238481 12801 238493 12835
rect 238527 12801 238539 12835
rect 238481 12795 238539 12801
rect 240689 12835 240747 12841
rect 240689 12801 240701 12835
rect 240735 12801 240747 12835
rect 240689 12795 240747 12801
rect 242066 12792 242072 12844
rect 242124 12792 242130 12844
rect 242250 12792 242256 12844
rect 242308 12832 242314 12844
rect 243817 12835 243875 12841
rect 243817 12832 243829 12835
rect 242308 12804 243829 12832
rect 242308 12792 242314 12804
rect 243817 12801 243829 12804
rect 243863 12832 243875 12835
rect 244246 12832 244274 12872
rect 244642 12860 244648 12872
rect 244700 12860 244706 12912
rect 244918 12860 244924 12912
rect 244976 12900 244982 12912
rect 245289 12903 245347 12909
rect 245289 12900 245301 12903
rect 244976 12872 245301 12900
rect 244976 12860 244982 12872
rect 245289 12869 245301 12872
rect 245335 12869 245347 12903
rect 245289 12863 245347 12869
rect 245378 12860 245384 12912
rect 245436 12900 245442 12912
rect 251361 12903 251419 12909
rect 251361 12900 251373 12903
rect 245436 12872 251373 12900
rect 245436 12860 245442 12872
rect 251361 12869 251373 12872
rect 251407 12900 251419 12903
rect 251634 12900 251640 12912
rect 251407 12872 251640 12900
rect 251407 12869 251419 12872
rect 251361 12863 251419 12869
rect 251634 12860 251640 12872
rect 251692 12860 251698 12912
rect 252462 12860 252468 12912
rect 252520 12900 252526 12912
rect 257246 12900 257252 12912
rect 252520 12872 252565 12900
rect 255162 12872 256740 12900
rect 252520 12860 252526 12872
rect 244550 12832 244556 12844
rect 243863 12804 244274 12832
rect 244511 12804 244556 12832
rect 243863 12801 243875 12804
rect 243817 12795 243875 12801
rect 244550 12792 244556 12804
rect 244608 12792 244614 12844
rect 244737 12835 244795 12841
rect 244737 12801 244749 12835
rect 244783 12832 244795 12835
rect 244826 12832 244832 12844
rect 244783 12804 244832 12832
rect 244783 12801 244795 12804
rect 244737 12795 244795 12801
rect 244826 12792 244832 12804
rect 244884 12832 244890 12844
rect 245197 12835 245255 12841
rect 245197 12832 245209 12835
rect 244884 12804 245209 12832
rect 244884 12792 244890 12804
rect 245197 12801 245209 12804
rect 245243 12801 245255 12835
rect 245197 12795 245255 12801
rect 250349 12835 250407 12841
rect 250349 12801 250361 12835
rect 250395 12832 250407 12835
rect 251174 12832 251180 12844
rect 250395 12804 251180 12832
rect 250395 12801 250407 12804
rect 250349 12795 250407 12801
rect 251146 12792 251180 12804
rect 251232 12792 251238 12844
rect 251542 12832 251548 12844
rect 251503 12804 251548 12832
rect 251542 12792 251548 12804
rect 251600 12792 251606 12844
rect 251652 12830 252416 12832
rect 252480 12830 252508 12860
rect 251652 12804 252508 12830
rect 233145 12767 233203 12773
rect 233145 12764 233157 12767
rect 230308 12736 232084 12764
rect 232700 12736 233157 12764
rect 230308 12696 230336 12736
rect 227211 12668 228036 12696
rect 229204 12668 230336 12696
rect 232056 12696 232084 12736
rect 233145 12733 233157 12736
rect 233191 12733 233203 12767
rect 251146 12764 251174 12792
rect 251652 12764 251680 12804
rect 252388 12802 252508 12804
rect 256237 12835 256295 12841
rect 256237 12801 256249 12835
rect 256283 12832 256295 12835
rect 256602 12832 256608 12844
rect 256283 12804 256608 12832
rect 256283 12801 256295 12804
rect 256237 12795 256295 12801
rect 256602 12792 256608 12804
rect 256660 12792 256666 12844
rect 233145 12727 233203 12733
rect 234586 12736 240548 12764
rect 234586 12696 234614 12736
rect 232056 12668 234614 12696
rect 237469 12699 237527 12705
rect 227211 12665 227223 12668
rect 227165 12659 227223 12665
rect 229204 12628 229232 12668
rect 237469 12665 237481 12699
rect 237515 12696 237527 12699
rect 237834 12696 237840 12708
rect 237515 12668 237840 12696
rect 237515 12665 237527 12668
rect 237469 12659 237527 12665
rect 237834 12656 237840 12668
rect 237892 12656 237898 12708
rect 237926 12656 237932 12708
rect 237984 12696 237990 12708
rect 237984 12668 238616 12696
rect 237984 12656 237990 12668
rect 227088 12600 229232 12628
rect 229554 12588 229560 12640
rect 229612 12628 229618 12640
rect 229649 12631 229707 12637
rect 229649 12628 229661 12631
rect 229612 12600 229661 12628
rect 229612 12588 229618 12600
rect 229649 12597 229661 12600
rect 229695 12597 229707 12631
rect 230106 12628 230112 12640
rect 230067 12600 230112 12628
rect 229649 12591 229707 12597
rect 230106 12588 230112 12600
rect 230164 12588 230170 12640
rect 230198 12588 230204 12640
rect 230256 12628 230262 12640
rect 232314 12628 232320 12640
rect 230256 12600 232320 12628
rect 230256 12588 230262 12600
rect 232314 12588 232320 12600
rect 232372 12588 232378 12640
rect 232498 12628 232504 12640
rect 232459 12600 232504 12628
rect 232498 12588 232504 12600
rect 232556 12628 232562 12640
rect 233142 12628 233148 12640
rect 232556 12600 233148 12628
rect 232556 12588 232562 12600
rect 233142 12588 233148 12600
rect 233200 12588 233206 12640
rect 236825 12631 236883 12637
rect 236825 12597 236837 12631
rect 236871 12628 236883 12631
rect 238478 12628 238484 12640
rect 236871 12600 238484 12628
rect 236871 12597 236883 12600
rect 236825 12591 236883 12597
rect 238478 12588 238484 12600
rect 238536 12588 238542 12640
rect 238588 12628 238616 12668
rect 238846 12628 238852 12640
rect 238588 12600 238852 12628
rect 238846 12588 238852 12600
rect 238904 12588 238910 12640
rect 239122 12588 239128 12640
rect 239180 12628 239186 12640
rect 240229 12631 240287 12637
rect 240229 12628 240241 12631
rect 239180 12600 240241 12628
rect 239180 12588 239186 12600
rect 240229 12597 240241 12600
rect 240275 12628 240287 12631
rect 240318 12628 240324 12640
rect 240275 12600 240324 12628
rect 240275 12597 240287 12600
rect 240229 12591 240287 12597
rect 240318 12588 240324 12600
rect 240376 12588 240382 12640
rect 240520 12628 240548 12736
rect 242084 12736 250300 12764
rect 251146 12736 251680 12764
rect 242084 12628 242112 12736
rect 242158 12656 242164 12708
rect 242216 12696 242222 12708
rect 242216 12668 244274 12696
rect 242216 12656 242222 12668
rect 242434 12628 242440 12640
rect 240520 12600 242112 12628
rect 242395 12600 242440 12628
rect 242434 12588 242440 12600
rect 242492 12588 242498 12640
rect 242894 12588 242900 12640
rect 242952 12628 242958 12640
rect 243909 12631 243967 12637
rect 243909 12628 243921 12631
rect 242952 12600 243921 12628
rect 242952 12588 242958 12600
rect 243909 12597 243921 12600
rect 243955 12597 243967 12631
rect 244246 12628 244274 12668
rect 244642 12656 244648 12708
rect 244700 12696 244706 12708
rect 248322 12696 248328 12708
rect 244700 12668 248328 12696
rect 244700 12656 244706 12668
rect 248322 12656 248328 12668
rect 248380 12656 248386 12708
rect 250162 12696 250168 12708
rect 250123 12668 250168 12696
rect 250162 12656 250168 12668
rect 250220 12656 250226 12708
rect 250272 12696 250300 12736
rect 252094 12724 252100 12776
rect 252152 12764 252158 12776
rect 252557 12767 252615 12773
rect 252557 12764 252569 12767
rect 252152 12736 252569 12764
rect 252152 12724 252158 12736
rect 252557 12733 252569 12736
rect 252603 12733 252615 12767
rect 252557 12727 252615 12733
rect 253658 12724 253664 12776
rect 253716 12764 253722 12776
rect 253716 12736 253761 12764
rect 253716 12724 253722 12736
rect 253934 12724 253940 12776
rect 253992 12764 253998 12776
rect 253992 12736 254037 12764
rect 253992 12724 253998 12736
rect 255130 12724 255136 12776
rect 255188 12764 255194 12776
rect 255409 12767 255467 12773
rect 255409 12764 255421 12767
rect 255188 12736 255421 12764
rect 255188 12724 255194 12736
rect 255409 12733 255421 12736
rect 255455 12764 255467 12767
rect 256326 12764 256332 12776
rect 255455 12736 256332 12764
rect 255455 12733 255467 12736
rect 255409 12727 255467 12733
rect 256326 12724 256332 12736
rect 256384 12724 256390 12776
rect 256418 12724 256424 12776
rect 256476 12764 256482 12776
rect 256476 12736 256521 12764
rect 256476 12724 256482 12736
rect 251818 12696 251824 12708
rect 250272 12668 251824 12696
rect 251818 12656 251824 12668
rect 251876 12656 251882 12708
rect 255038 12656 255044 12708
rect 255096 12696 255102 12708
rect 255869 12699 255927 12705
rect 255869 12696 255881 12699
rect 255096 12668 255881 12696
rect 255096 12656 255102 12668
rect 255869 12665 255881 12668
rect 255915 12665 255927 12699
rect 255869 12659 255927 12665
rect 251910 12628 251916 12640
rect 244246 12600 251916 12628
rect 243909 12591 243967 12597
rect 251910 12588 251916 12600
rect 251968 12588 251974 12640
rect 252002 12588 252008 12640
rect 252060 12628 252066 12640
rect 256712 12628 256740 12872
rect 257080 12872 257252 12900
rect 257080 12841 257108 12872
rect 257246 12860 257252 12872
rect 257304 12860 257310 12912
rect 261754 12900 261760 12912
rect 261667 12872 261760 12900
rect 261754 12860 261760 12872
rect 261812 12900 261818 12912
rect 263229 12903 263287 12909
rect 263229 12900 263241 12903
rect 261812 12872 263241 12900
rect 261812 12860 261818 12872
rect 263229 12869 263241 12872
rect 263275 12869 263287 12903
rect 263229 12863 263287 12869
rect 263318 12860 263324 12912
rect 263376 12900 263382 12912
rect 263413 12903 263471 12909
rect 263413 12900 263425 12903
rect 263376 12872 263425 12900
rect 263376 12860 263382 12872
rect 263413 12869 263425 12872
rect 263459 12869 263471 12903
rect 263566 12900 263594 12940
rect 264606 12928 264612 12940
rect 264664 12928 264670 12980
rect 268378 12968 268384 12980
rect 265268 12940 268384 12968
rect 265268 12900 265296 12940
rect 268378 12928 268384 12940
rect 268436 12928 268442 12980
rect 302602 12968 302608 12980
rect 268488 12940 296714 12968
rect 302563 12940 302608 12968
rect 265526 12900 265532 12912
rect 263566 12872 265296 12900
rect 265487 12872 265532 12900
rect 263413 12863 263471 12869
rect 257065 12835 257123 12841
rect 257065 12801 257077 12835
rect 257111 12801 257123 12835
rect 257065 12795 257123 12801
rect 261846 12792 261852 12844
rect 261904 12832 261910 12844
rect 262493 12835 262551 12841
rect 262493 12832 262505 12835
rect 261904 12804 262505 12832
rect 261904 12792 261910 12804
rect 262493 12801 262505 12804
rect 262539 12801 262551 12835
rect 262493 12795 262551 12801
rect 264149 12835 264207 12841
rect 264149 12801 264161 12835
rect 264195 12832 264207 12835
rect 264330 12832 264336 12844
rect 264195 12804 264336 12832
rect 264195 12801 264207 12804
rect 264149 12795 264207 12801
rect 264330 12792 264336 12804
rect 264388 12792 264394 12844
rect 264422 12792 264428 12844
rect 264480 12832 264486 12844
rect 265268 12841 265296 12872
rect 265526 12860 265532 12872
rect 265584 12860 265590 12912
rect 266538 12860 266544 12912
rect 266596 12860 266602 12912
rect 268488 12900 268516 12940
rect 271046 12900 271052 12912
rect 266832 12872 268516 12900
rect 270618 12872 271052 12900
rect 264793 12835 264851 12841
rect 264793 12832 264805 12835
rect 264480 12804 264805 12832
rect 264480 12792 264486 12804
rect 264793 12801 264805 12804
rect 264839 12801 264851 12835
rect 264793 12795 264851 12801
rect 265253 12835 265311 12841
rect 265253 12801 265265 12835
rect 265299 12801 265311 12835
rect 265253 12795 265311 12801
rect 257154 12724 257160 12776
rect 257212 12764 257218 12776
rect 262306 12764 262312 12776
rect 257212 12736 262312 12764
rect 257212 12724 257218 12736
rect 262306 12724 262312 12736
rect 262364 12724 262370 12776
rect 266832 12764 266860 12872
rect 271046 12860 271052 12872
rect 271104 12860 271110 12912
rect 271782 12900 271788 12912
rect 271695 12872 271788 12900
rect 271782 12860 271788 12872
rect 271840 12900 271846 12912
rect 272794 12900 272800 12912
rect 271840 12872 272800 12900
rect 271840 12860 271846 12872
rect 272794 12860 272800 12872
rect 272852 12860 272858 12912
rect 272889 12903 272947 12909
rect 272889 12869 272901 12903
rect 272935 12900 272947 12903
rect 273162 12900 273168 12912
rect 272935 12872 273168 12900
rect 272935 12869 272947 12872
rect 272889 12863 272947 12869
rect 273162 12860 273168 12872
rect 273220 12860 273226 12912
rect 295886 12900 295892 12912
rect 282886 12872 295892 12900
rect 267829 12835 267887 12841
rect 267829 12801 267841 12835
rect 267875 12832 267887 12835
rect 268286 12832 268292 12844
rect 267875 12804 268292 12832
rect 267875 12801 267887 12804
rect 267829 12795 267887 12801
rect 268286 12792 268292 12804
rect 268344 12832 268350 12844
rect 269022 12832 269028 12844
rect 268344 12804 269028 12832
rect 268344 12792 268350 12804
rect 269022 12792 269028 12804
rect 269080 12792 269086 12844
rect 269117 12835 269175 12841
rect 269117 12801 269129 12835
rect 269163 12801 269175 12835
rect 269117 12795 269175 12801
rect 263428 12736 266860 12764
rect 257062 12656 257068 12708
rect 257120 12696 257126 12708
rect 262674 12696 262680 12708
rect 257120 12668 262536 12696
rect 262635 12668 262680 12696
rect 257120 12656 257126 12668
rect 257157 12631 257215 12637
rect 257157 12628 257169 12631
rect 252060 12600 252105 12628
rect 256712 12600 257169 12628
rect 252060 12588 252066 12600
rect 257157 12597 257169 12600
rect 257203 12597 257215 12631
rect 257157 12591 257215 12597
rect 261849 12631 261907 12637
rect 261849 12597 261861 12631
rect 261895 12628 261907 12631
rect 262214 12628 262220 12640
rect 261895 12600 262220 12628
rect 261895 12597 261907 12600
rect 261849 12591 261907 12597
rect 262214 12588 262220 12600
rect 262272 12588 262278 12640
rect 262508 12628 262536 12668
rect 262674 12656 262680 12668
rect 262732 12656 262738 12708
rect 263428 12628 263456 12736
rect 266998 12724 267004 12776
rect 267056 12764 267062 12776
rect 267550 12764 267556 12776
rect 267056 12736 267556 12764
rect 267056 12724 267062 12736
rect 267550 12724 267556 12736
rect 267608 12764 267614 12776
rect 267921 12767 267979 12773
rect 267921 12764 267933 12767
rect 267608 12736 267933 12764
rect 267608 12724 267614 12736
rect 267921 12733 267933 12736
rect 267967 12733 267979 12767
rect 267921 12727 267979 12733
rect 268010 12724 268016 12776
rect 268068 12764 268074 12776
rect 268068 12736 268113 12764
rect 268068 12724 268074 12736
rect 268378 12724 268384 12776
rect 268436 12764 268442 12776
rect 269132 12764 269160 12795
rect 270862 12792 270868 12844
rect 270920 12832 270926 12844
rect 271693 12835 271751 12841
rect 271693 12832 271705 12835
rect 270920 12804 271705 12832
rect 270920 12792 270926 12804
rect 271693 12801 271705 12804
rect 271739 12832 271751 12835
rect 272610 12832 272616 12844
rect 271739 12804 272616 12832
rect 271739 12801 271751 12804
rect 271693 12795 271751 12801
rect 272610 12792 272616 12804
rect 272668 12792 272674 12844
rect 282886 12832 282914 12872
rect 295886 12860 295892 12872
rect 295944 12860 295950 12912
rect 296686 12900 296714 12940
rect 302602 12928 302608 12940
rect 302660 12928 302666 12980
rect 304445 12971 304503 12977
rect 304445 12937 304457 12971
rect 304491 12968 304503 12971
rect 305362 12968 305368 12980
rect 304491 12940 305368 12968
rect 304491 12937 304503 12940
rect 304445 12931 304503 12937
rect 305362 12928 305368 12940
rect 305420 12928 305426 12980
rect 304994 12900 305000 12912
rect 296686 12872 304672 12900
rect 304955 12872 305000 12900
rect 290274 12832 290280 12844
rect 272720 12804 282914 12832
rect 287026 12804 290280 12832
rect 269390 12764 269396 12776
rect 268436 12736 269160 12764
rect 269351 12736 269396 12764
rect 268436 12724 268442 12736
rect 269390 12724 269396 12736
rect 269448 12724 269454 12776
rect 271969 12767 272027 12773
rect 270880 12736 271460 12764
rect 263502 12656 263508 12708
rect 263560 12696 263566 12708
rect 270880 12696 270908 12736
rect 263560 12668 264100 12696
rect 263560 12656 263566 12668
rect 263962 12628 263968 12640
rect 262508 12600 263456 12628
rect 263923 12600 263968 12628
rect 263962 12588 263968 12600
rect 264020 12588 264026 12640
rect 264072 12628 264100 12668
rect 266556 12668 269252 12696
rect 266556 12628 266584 12668
rect 266998 12628 267004 12640
rect 264072 12600 266584 12628
rect 266959 12600 267004 12628
rect 266998 12588 267004 12600
rect 267056 12588 267062 12640
rect 267090 12588 267096 12640
rect 267148 12628 267154 12640
rect 267461 12631 267519 12637
rect 267461 12628 267473 12631
rect 267148 12600 267473 12628
rect 267148 12588 267154 12600
rect 267461 12597 267473 12600
rect 267507 12597 267519 12631
rect 267461 12591 267519 12597
rect 267550 12588 267556 12640
rect 267608 12628 267614 12640
rect 269114 12628 269120 12640
rect 267608 12600 269120 12628
rect 267608 12588 267614 12600
rect 269114 12588 269120 12600
rect 269172 12588 269178 12640
rect 269224 12628 269252 12668
rect 270420 12668 270908 12696
rect 271432 12696 271460 12736
rect 271969 12733 271981 12767
rect 272015 12764 272027 12767
rect 272242 12764 272248 12776
rect 272015 12736 272248 12764
rect 272015 12733 272027 12736
rect 271969 12727 272027 12733
rect 272242 12724 272248 12736
rect 272300 12724 272306 12776
rect 272720 12696 272748 12804
rect 272886 12724 272892 12776
rect 272944 12764 272950 12776
rect 272981 12767 273039 12773
rect 272981 12764 272993 12767
rect 272944 12736 272993 12764
rect 272944 12724 272950 12736
rect 272981 12733 272993 12736
rect 273027 12733 273039 12767
rect 272981 12727 273039 12733
rect 273073 12767 273131 12773
rect 273073 12733 273085 12767
rect 273119 12733 273131 12767
rect 273073 12727 273131 12733
rect 271432 12668 272748 12696
rect 270420 12628 270448 12668
rect 272794 12656 272800 12708
rect 272852 12696 272858 12708
rect 273088 12696 273116 12727
rect 273162 12724 273168 12776
rect 273220 12764 273226 12776
rect 287026 12764 287054 12804
rect 290274 12792 290280 12804
rect 290332 12792 290338 12844
rect 302786 12832 302792 12844
rect 302747 12804 302792 12832
rect 302786 12792 302792 12804
rect 302844 12792 302850 12844
rect 304644 12841 304672 12872
rect 304994 12860 305000 12872
rect 305052 12900 305058 12912
rect 305454 12900 305460 12912
rect 305052 12872 305460 12900
rect 305052 12860 305058 12872
rect 305454 12860 305460 12872
rect 305512 12860 305518 12912
rect 304629 12835 304687 12841
rect 304629 12801 304641 12835
rect 304675 12801 304687 12835
rect 304629 12795 304687 12801
rect 273220 12736 287054 12764
rect 273220 12724 273226 12736
rect 272852 12668 273116 12696
rect 272852 12656 272858 12668
rect 270862 12628 270868 12640
rect 269224 12600 270448 12628
rect 270823 12600 270868 12628
rect 270862 12588 270868 12600
rect 270920 12588 270926 12640
rect 271138 12588 271144 12640
rect 271196 12628 271202 12640
rect 271325 12631 271383 12637
rect 271325 12628 271337 12631
rect 271196 12600 271337 12628
rect 271196 12588 271202 12600
rect 271325 12597 271337 12600
rect 271371 12597 271383 12631
rect 272518 12628 272524 12640
rect 272479 12600 272524 12628
rect 271325 12591 271383 12597
rect 272518 12588 272524 12600
rect 272576 12588 272582 12640
rect 272610 12588 272616 12640
rect 272668 12628 272674 12640
rect 281074 12628 281080 12640
rect 272668 12600 281080 12628
rect 272668 12588 272674 12600
rect 281074 12588 281080 12600
rect 281132 12588 281138 12640
rect 1104 12538 305808 12560
rect 1104 12486 39049 12538
rect 39101 12486 39113 12538
rect 39165 12486 39177 12538
rect 39229 12486 39241 12538
rect 39293 12486 39305 12538
rect 39357 12486 115247 12538
rect 115299 12486 115311 12538
rect 115363 12486 115375 12538
rect 115427 12486 115439 12538
rect 115491 12486 115503 12538
rect 115555 12486 191445 12538
rect 191497 12486 191509 12538
rect 191561 12486 191573 12538
rect 191625 12486 191637 12538
rect 191689 12486 191701 12538
rect 191753 12486 267643 12538
rect 267695 12486 267707 12538
rect 267759 12486 267771 12538
rect 267823 12486 267835 12538
rect 267887 12486 267899 12538
rect 267951 12486 305808 12538
rect 1104 12464 305808 12486
rect 26970 12384 26976 12436
rect 27028 12424 27034 12436
rect 28074 12424 28080 12436
rect 27028 12396 28080 12424
rect 27028 12384 27034 12396
rect 28074 12384 28080 12396
rect 28132 12424 28138 12436
rect 28132 12396 28488 12424
rect 28132 12384 28138 12396
rect 14274 12316 14280 12368
rect 14332 12356 14338 12368
rect 28460 12356 28488 12396
rect 28810 12384 28816 12436
rect 28868 12424 28874 12436
rect 31297 12427 31355 12433
rect 31297 12424 31309 12427
rect 28868 12396 31309 12424
rect 28868 12384 28874 12396
rect 31297 12393 31309 12396
rect 31343 12393 31355 12427
rect 31297 12387 31355 12393
rect 32582 12384 32588 12436
rect 32640 12424 32646 12436
rect 33965 12427 34023 12433
rect 32640 12396 33088 12424
rect 32640 12384 32646 12396
rect 33060 12356 33088 12396
rect 33965 12393 33977 12427
rect 34011 12424 34023 12427
rect 34514 12424 34520 12436
rect 34011 12396 34520 12424
rect 34011 12393 34023 12396
rect 33965 12387 34023 12393
rect 34514 12384 34520 12396
rect 34572 12384 34578 12436
rect 34793 12427 34851 12433
rect 34793 12393 34805 12427
rect 34839 12424 34851 12427
rect 35986 12424 35992 12436
rect 34839 12396 35992 12424
rect 34839 12393 34851 12396
rect 34793 12387 34851 12393
rect 35986 12384 35992 12396
rect 36044 12384 36050 12436
rect 37185 12427 37243 12433
rect 37185 12393 37197 12427
rect 37231 12393 37243 12427
rect 37185 12387 37243 12393
rect 34882 12356 34888 12368
rect 14332 12328 28396 12356
rect 28460 12328 28948 12356
rect 33060 12328 34888 12356
rect 14332 12316 14338 12328
rect 26878 12288 26884 12300
rect 16960 12260 26884 12288
rect 4798 12044 4804 12096
rect 4856 12084 4862 12096
rect 16960 12084 16988 12260
rect 26878 12248 26884 12260
rect 26936 12248 26942 12300
rect 27709 12291 27767 12297
rect 27709 12257 27721 12291
rect 27755 12288 27767 12291
rect 28074 12288 28080 12300
rect 27755 12260 28080 12288
rect 27755 12257 27767 12260
rect 27709 12251 27767 12257
rect 28074 12248 28080 12260
rect 28132 12248 28138 12300
rect 28368 12288 28396 12328
rect 28718 12288 28724 12300
rect 28368 12260 28724 12288
rect 28718 12248 28724 12260
rect 28776 12248 28782 12300
rect 28920 12297 28948 12328
rect 34882 12316 34888 12328
rect 34940 12356 34946 12368
rect 37200 12356 37228 12387
rect 37826 12384 37832 12436
rect 37884 12424 37890 12436
rect 38473 12427 38531 12433
rect 38473 12424 38485 12427
rect 37884 12396 38485 12424
rect 37884 12384 37890 12396
rect 38473 12393 38485 12396
rect 38519 12393 38531 12427
rect 38473 12387 38531 12393
rect 38930 12384 38936 12436
rect 38988 12424 38994 12436
rect 39209 12427 39267 12433
rect 39209 12424 39221 12427
rect 38988 12396 39221 12424
rect 38988 12384 38994 12396
rect 39209 12393 39221 12396
rect 39255 12393 39267 12427
rect 39209 12387 39267 12393
rect 39390 12384 39396 12436
rect 39448 12424 39454 12436
rect 40954 12424 40960 12436
rect 39448 12396 40960 12424
rect 39448 12384 39454 12396
rect 40954 12384 40960 12396
rect 41012 12384 41018 12436
rect 43162 12424 43168 12436
rect 41524 12396 43024 12424
rect 43123 12396 43168 12424
rect 41524 12356 41552 12396
rect 34940 12328 37228 12356
rect 37292 12328 41552 12356
rect 42996 12356 43024 12396
rect 43162 12384 43168 12396
rect 43220 12384 43226 12436
rect 43806 12424 43812 12436
rect 43767 12396 43812 12424
rect 43806 12384 43812 12396
rect 43864 12384 43870 12436
rect 54018 12384 54024 12436
rect 54076 12424 54082 12436
rect 54113 12427 54171 12433
rect 54113 12424 54125 12427
rect 54076 12396 54125 12424
rect 54076 12384 54082 12396
rect 54113 12393 54125 12396
rect 54159 12393 54171 12427
rect 54113 12387 54171 12393
rect 54665 12427 54723 12433
rect 54665 12393 54677 12427
rect 54711 12424 54723 12427
rect 55490 12424 55496 12436
rect 54711 12396 55496 12424
rect 54711 12393 54723 12396
rect 54665 12387 54723 12393
rect 55490 12384 55496 12396
rect 55548 12384 55554 12436
rect 56686 12384 56692 12436
rect 56744 12424 56750 12436
rect 57333 12427 57391 12433
rect 57333 12424 57345 12427
rect 56744 12396 57345 12424
rect 56744 12384 56750 12396
rect 57333 12393 57345 12396
rect 57379 12393 57391 12427
rect 57974 12424 57980 12436
rect 57935 12396 57980 12424
rect 57333 12387 57391 12393
rect 57974 12384 57980 12396
rect 58032 12384 58038 12436
rect 75086 12384 75092 12436
rect 75144 12424 75150 12436
rect 75181 12427 75239 12433
rect 75181 12424 75193 12427
rect 75144 12396 75193 12424
rect 75144 12384 75150 12396
rect 75181 12393 75193 12396
rect 75227 12393 75239 12427
rect 79318 12424 79324 12436
rect 75181 12387 75239 12393
rect 75288 12396 78536 12424
rect 79279 12396 79324 12424
rect 43714 12356 43720 12368
rect 42996 12328 43720 12356
rect 34940 12316 34946 12328
rect 28905 12291 28963 12297
rect 28905 12257 28917 12291
rect 28951 12288 28963 12291
rect 28994 12288 29000 12300
rect 28951 12260 29000 12288
rect 28951 12257 28963 12260
rect 28905 12251 28963 12257
rect 28994 12248 29000 12260
rect 29052 12248 29058 12300
rect 29546 12288 29552 12300
rect 29459 12260 29552 12288
rect 29546 12248 29552 12260
rect 29604 12288 29610 12300
rect 31757 12291 31815 12297
rect 31757 12288 31769 12291
rect 29604 12260 31769 12288
rect 29604 12248 29610 12260
rect 31757 12257 31769 12260
rect 31803 12288 31815 12291
rect 31803 12260 35572 12288
rect 31803 12257 31815 12260
rect 31757 12251 31815 12257
rect 17034 12180 17040 12232
rect 17092 12220 17098 12232
rect 17092 12192 22094 12220
rect 17092 12180 17098 12192
rect 22066 12152 22094 12192
rect 27080 12192 27384 12220
rect 27080 12152 27108 12192
rect 22066 12124 27108 12152
rect 27356 12152 27384 12192
rect 27430 12180 27436 12232
rect 27488 12220 27494 12232
rect 28629 12223 28687 12229
rect 28629 12220 28641 12223
rect 27488 12192 27533 12220
rect 28000 12192 28641 12220
rect 27488 12180 27494 12192
rect 28000 12152 28028 12192
rect 28629 12189 28641 12192
rect 28675 12220 28687 12223
rect 29362 12220 29368 12232
rect 28675 12192 29368 12220
rect 28675 12189 28687 12192
rect 28629 12183 28687 12189
rect 29362 12180 29368 12192
rect 29420 12180 29426 12232
rect 34146 12220 34152 12232
rect 34107 12192 34152 12220
rect 34146 12180 34152 12192
rect 34204 12180 34210 12232
rect 34698 12220 34704 12232
rect 34611 12192 34704 12220
rect 34698 12180 34704 12192
rect 34756 12220 34762 12232
rect 35342 12220 35348 12232
rect 34756 12192 35348 12220
rect 34756 12180 34762 12192
rect 35342 12180 35348 12192
rect 35400 12180 35406 12232
rect 29454 12152 29460 12164
rect 27356 12124 28028 12152
rect 28276 12124 29460 12152
rect 27062 12084 27068 12096
rect 4856 12056 16988 12084
rect 27023 12056 27068 12084
rect 4856 12044 4862 12056
rect 27062 12044 27068 12056
rect 27120 12044 27126 12096
rect 27154 12044 27160 12096
rect 27212 12084 27218 12096
rect 27525 12087 27583 12093
rect 27525 12084 27537 12087
rect 27212 12056 27537 12084
rect 27212 12044 27218 12056
rect 27525 12053 27537 12056
rect 27571 12084 27583 12087
rect 27982 12084 27988 12096
rect 27571 12056 27988 12084
rect 27571 12053 27583 12056
rect 27525 12047 27583 12053
rect 27982 12044 27988 12056
rect 28040 12044 28046 12096
rect 28276 12093 28304 12124
rect 29454 12112 29460 12124
rect 29512 12112 29518 12164
rect 29822 12152 29828 12164
rect 29783 12124 29828 12152
rect 29822 12112 29828 12124
rect 29880 12112 29886 12164
rect 31202 12152 31208 12164
rect 31050 12124 31208 12152
rect 31202 12112 31208 12124
rect 31260 12112 31266 12164
rect 32030 12152 32036 12164
rect 31991 12124 32036 12152
rect 32030 12112 32036 12124
rect 32088 12112 32094 12164
rect 35437 12155 35495 12161
rect 35437 12152 35449 12155
rect 33258 12124 35449 12152
rect 35437 12121 35449 12124
rect 35483 12121 35495 12155
rect 35544 12152 35572 12260
rect 36357 12223 36415 12229
rect 36357 12189 36369 12223
rect 36403 12220 36415 12223
rect 37093 12223 37151 12229
rect 37093 12220 37105 12223
rect 36403 12192 37105 12220
rect 36403 12189 36415 12192
rect 36357 12183 36415 12189
rect 37093 12189 37105 12192
rect 37139 12220 37151 12223
rect 37292 12220 37320 12328
rect 43714 12316 43720 12328
rect 43772 12316 43778 12368
rect 75288 12356 75316 12396
rect 53668 12328 75316 12356
rect 40865 12291 40923 12297
rect 40865 12257 40877 12291
rect 40911 12288 40923 12291
rect 40954 12288 40960 12300
rect 40911 12260 40960 12288
rect 40911 12257 40923 12260
rect 40865 12251 40923 12257
rect 40954 12248 40960 12260
rect 41012 12248 41018 12300
rect 52365 12291 52423 12297
rect 52365 12288 52377 12291
rect 41432 12260 52377 12288
rect 37139 12192 37320 12220
rect 37139 12189 37151 12192
rect 37093 12183 37151 12189
rect 38010 12180 38016 12232
rect 38068 12220 38074 12232
rect 38657 12223 38715 12229
rect 38657 12220 38669 12223
rect 38068 12192 38669 12220
rect 38068 12180 38074 12192
rect 38657 12189 38669 12192
rect 38703 12189 38715 12223
rect 38657 12183 38715 12189
rect 39117 12223 39175 12229
rect 39117 12189 39129 12223
rect 39163 12220 39175 12223
rect 40310 12220 40316 12232
rect 39163 12192 40316 12220
rect 39163 12189 39175 12192
rect 39117 12183 39175 12189
rect 40310 12180 40316 12192
rect 40368 12180 40374 12232
rect 40586 12220 40592 12232
rect 40547 12192 40592 12220
rect 40586 12180 40592 12192
rect 40644 12180 40650 12232
rect 41432 12229 41460 12260
rect 52365 12257 52377 12260
rect 52411 12288 52423 12291
rect 53668 12288 53696 12328
rect 76006 12316 76012 12368
rect 76064 12356 76070 12368
rect 77202 12356 77208 12368
rect 76064 12328 77208 12356
rect 76064 12316 76070 12328
rect 52411 12260 53696 12288
rect 52411 12257 52423 12260
rect 52365 12251 52423 12257
rect 53834 12248 53840 12300
rect 53892 12248 53898 12300
rect 55677 12291 55735 12297
rect 55677 12288 55689 12291
rect 55186 12260 55689 12288
rect 41417 12223 41475 12229
rect 41417 12189 41429 12223
rect 41463 12189 41475 12223
rect 43714 12220 43720 12232
rect 43675 12192 43720 12220
rect 41417 12183 41475 12189
rect 41432 12152 41460 12183
rect 43714 12180 43720 12192
rect 43772 12220 43778 12232
rect 53852 12220 53880 12248
rect 54573 12223 54631 12229
rect 54573 12220 54585 12223
rect 43772 12192 48314 12220
rect 53852 12192 54585 12220
rect 43772 12180 43778 12192
rect 35544 12124 41460 12152
rect 35437 12115 35495 12121
rect 41598 12112 41604 12164
rect 41656 12152 41662 12164
rect 41693 12155 41751 12161
rect 41693 12152 41705 12155
rect 41656 12124 41705 12152
rect 41656 12112 41662 12124
rect 41693 12121 41705 12124
rect 41739 12121 41751 12155
rect 41693 12115 41751 12121
rect 41782 12112 41788 12164
rect 41840 12152 41846 12164
rect 41840 12124 42182 12152
rect 41840 12112 41846 12124
rect 28261 12087 28319 12093
rect 28261 12053 28273 12087
rect 28307 12053 28319 12087
rect 28261 12047 28319 12053
rect 28902 12044 28908 12096
rect 28960 12084 28966 12096
rect 31110 12084 31116 12096
rect 28960 12056 31116 12084
rect 28960 12044 28966 12056
rect 31110 12044 31116 12056
rect 31168 12044 31174 12096
rect 32306 12044 32312 12096
rect 32364 12084 32370 12096
rect 32950 12084 32956 12096
rect 32364 12056 32956 12084
rect 32364 12044 32370 12056
rect 32950 12044 32956 12056
rect 33008 12084 33014 12096
rect 33505 12087 33563 12093
rect 33505 12084 33517 12087
rect 33008 12056 33517 12084
rect 33008 12044 33014 12056
rect 33505 12053 33517 12056
rect 33551 12053 33563 12087
rect 36446 12084 36452 12096
rect 36407 12056 36452 12084
rect 33505 12047 33563 12053
rect 36446 12044 36452 12056
rect 36504 12044 36510 12096
rect 40221 12087 40279 12093
rect 40221 12053 40233 12087
rect 40267 12084 40279 12087
rect 40494 12084 40500 12096
rect 40267 12056 40500 12084
rect 40267 12053 40279 12056
rect 40221 12047 40279 12053
rect 40494 12044 40500 12056
rect 40552 12044 40558 12096
rect 40678 12084 40684 12096
rect 40639 12056 40684 12084
rect 40678 12044 40684 12056
rect 40736 12044 40742 12096
rect 48286 12084 48314 12192
rect 54573 12189 54585 12192
rect 54619 12220 54631 12223
rect 55186 12220 55214 12260
rect 55677 12257 55689 12260
rect 55723 12257 55735 12291
rect 55677 12251 55735 12257
rect 56410 12248 56416 12300
rect 56468 12288 56474 12300
rect 56689 12291 56747 12297
rect 56689 12288 56701 12291
rect 56468 12260 56701 12288
rect 56468 12248 56474 12260
rect 56689 12257 56701 12260
rect 56735 12257 56747 12291
rect 56689 12251 56747 12257
rect 74810 12248 74816 12300
rect 74868 12288 74874 12300
rect 76760 12297 76788 12328
rect 77202 12316 77208 12328
rect 77260 12316 77266 12368
rect 77481 12359 77539 12365
rect 77481 12325 77493 12359
rect 77527 12356 77539 12359
rect 78398 12356 78404 12368
rect 77527 12328 78404 12356
rect 77527 12325 77539 12328
rect 77481 12319 77539 12325
rect 78398 12316 78404 12328
rect 78456 12316 78462 12368
rect 76745 12291 76803 12297
rect 74868 12260 76696 12288
rect 74868 12248 74874 12260
rect 54619 12192 55214 12220
rect 54619 12189 54631 12192
rect 54573 12183 54631 12189
rect 55306 12180 55312 12232
rect 55364 12220 55370 12232
rect 56502 12220 56508 12232
rect 55364 12192 56508 12220
rect 55364 12180 55370 12192
rect 56502 12180 56508 12192
rect 56560 12220 56566 12232
rect 76668 12229 76696 12260
rect 76745 12257 76757 12291
rect 76791 12257 76803 12291
rect 76745 12251 76803 12257
rect 76926 12248 76932 12300
rect 76984 12288 76990 12300
rect 78122 12288 78128 12300
rect 76984 12260 78128 12288
rect 76984 12248 76990 12260
rect 78122 12248 78128 12260
rect 78180 12248 78186 12300
rect 56597 12223 56655 12229
rect 56597 12220 56609 12223
rect 56560 12192 56609 12220
rect 56560 12180 56566 12192
rect 56597 12189 56609 12192
rect 56643 12220 56655 12223
rect 57517 12223 57575 12229
rect 57517 12220 57529 12223
rect 56643 12192 57529 12220
rect 56643 12189 56655 12192
rect 56597 12183 56655 12189
rect 57517 12189 57529 12192
rect 57563 12189 57575 12223
rect 57517 12183 57575 12189
rect 58161 12223 58219 12229
rect 58161 12189 58173 12223
rect 58207 12189 58219 12223
rect 58161 12183 58219 12189
rect 75365 12223 75423 12229
rect 75365 12189 75377 12223
rect 75411 12220 75423 12223
rect 76653 12223 76711 12229
rect 75411 12192 76604 12220
rect 75411 12189 75423 12192
rect 75365 12183 75423 12189
rect 52638 12152 52644 12164
rect 52599 12124 52644 12152
rect 52638 12112 52644 12124
rect 52696 12112 52702 12164
rect 53098 12112 53104 12164
rect 53156 12112 53162 12164
rect 55493 12155 55551 12161
rect 53944 12124 55214 12152
rect 53944 12084 53972 12124
rect 48286 12056 53972 12084
rect 55186 12084 55214 12124
rect 55493 12121 55505 12155
rect 55539 12152 55551 12155
rect 58176 12152 58204 12183
rect 55539 12124 56088 12152
rect 55539 12121 55551 12124
rect 55493 12115 55551 12121
rect 56060 12096 56088 12124
rect 56152 12124 58204 12152
rect 76576 12152 76604 12192
rect 76653 12189 76665 12223
rect 76699 12220 76711 12223
rect 77938 12220 77944 12232
rect 76699 12192 77944 12220
rect 76699 12189 76711 12192
rect 76653 12183 76711 12189
rect 77938 12180 77944 12192
rect 77996 12180 78002 12232
rect 78508 12152 78536 12396
rect 79318 12384 79324 12396
rect 79376 12384 79382 12436
rect 80241 12427 80299 12433
rect 80241 12393 80253 12427
rect 80287 12424 80299 12427
rect 80514 12424 80520 12436
rect 80287 12396 80520 12424
rect 80287 12393 80299 12396
rect 80241 12387 80299 12393
rect 80514 12384 80520 12396
rect 80572 12384 80578 12436
rect 85482 12384 85488 12436
rect 85540 12424 85546 12436
rect 85577 12427 85635 12433
rect 85577 12424 85589 12427
rect 85540 12396 85589 12424
rect 85540 12384 85546 12396
rect 85577 12393 85589 12396
rect 85623 12393 85635 12427
rect 86402 12424 86408 12436
rect 86363 12396 86408 12424
rect 85577 12387 85635 12393
rect 86402 12384 86408 12396
rect 86460 12384 86466 12436
rect 87874 12384 87880 12436
rect 87932 12424 87938 12436
rect 88889 12427 88947 12433
rect 88889 12424 88901 12427
rect 87932 12396 88901 12424
rect 87932 12384 87938 12396
rect 88889 12393 88901 12396
rect 88935 12393 88947 12427
rect 90174 12424 90180 12436
rect 90135 12396 90180 12424
rect 88889 12387 88947 12393
rect 90174 12384 90180 12396
rect 90232 12384 90238 12436
rect 99101 12427 99159 12433
rect 99101 12393 99113 12427
rect 99147 12424 99159 12427
rect 99466 12424 99472 12436
rect 99147 12396 99472 12424
rect 99147 12393 99159 12396
rect 99101 12387 99159 12393
rect 99466 12384 99472 12396
rect 99524 12384 99530 12436
rect 99837 12427 99895 12433
rect 99837 12393 99849 12427
rect 99883 12424 99895 12427
rect 99926 12424 99932 12436
rect 99883 12396 99932 12424
rect 99883 12393 99895 12396
rect 99837 12387 99895 12393
rect 99926 12384 99932 12396
rect 99984 12384 99990 12436
rect 103885 12427 103943 12433
rect 103885 12393 103897 12427
rect 103931 12424 103943 12427
rect 104986 12424 104992 12436
rect 103931 12396 104992 12424
rect 103931 12393 103943 12396
rect 103885 12387 103943 12393
rect 104986 12384 104992 12396
rect 105044 12384 105050 12436
rect 105170 12424 105176 12436
rect 105131 12396 105176 12424
rect 105170 12384 105176 12396
rect 105228 12384 105234 12436
rect 112530 12384 112536 12436
rect 112588 12424 112594 12436
rect 113085 12427 113143 12433
rect 113085 12424 113097 12427
rect 112588 12396 113097 12424
rect 112588 12384 112594 12396
rect 113085 12393 113097 12396
rect 113131 12393 113143 12427
rect 113085 12387 113143 12393
rect 113729 12427 113787 12433
rect 113729 12393 113741 12427
rect 113775 12424 113787 12427
rect 115014 12424 115020 12436
rect 113775 12396 115020 12424
rect 113775 12393 113787 12396
rect 113729 12387 113787 12393
rect 115014 12384 115020 12396
rect 115072 12384 115078 12436
rect 116946 12384 116952 12436
rect 117004 12424 117010 12436
rect 118421 12427 118479 12433
rect 118421 12424 118433 12427
rect 117004 12396 118433 12424
rect 117004 12384 117010 12396
rect 118421 12393 118433 12396
rect 118467 12393 118479 12427
rect 118421 12387 118479 12393
rect 127713 12427 127771 12433
rect 127713 12393 127725 12427
rect 127759 12424 127771 12427
rect 127802 12424 127808 12436
rect 127759 12396 127808 12424
rect 127759 12393 127771 12396
rect 127713 12387 127771 12393
rect 127802 12384 127808 12396
rect 127860 12384 127866 12436
rect 129090 12384 129096 12436
rect 129148 12424 129154 12436
rect 130841 12427 130899 12433
rect 130841 12424 130853 12427
rect 129148 12396 130853 12424
rect 129148 12384 129154 12396
rect 130841 12393 130853 12396
rect 130887 12424 130899 12427
rect 130930 12424 130936 12436
rect 130887 12396 130936 12424
rect 130887 12393 130899 12396
rect 130841 12387 130899 12393
rect 130930 12384 130936 12396
rect 130988 12384 130994 12436
rect 132402 12384 132408 12436
rect 132460 12424 132466 12436
rect 132681 12427 132739 12433
rect 132681 12424 132693 12427
rect 132460 12396 132693 12424
rect 132460 12384 132466 12396
rect 132681 12393 132693 12396
rect 132727 12393 132739 12427
rect 132681 12387 132739 12393
rect 147309 12427 147367 12433
rect 147309 12393 147321 12427
rect 147355 12424 147367 12427
rect 147766 12424 147772 12436
rect 147355 12396 147772 12424
rect 147355 12393 147367 12396
rect 147309 12387 147367 12393
rect 147766 12384 147772 12396
rect 147824 12384 147830 12436
rect 152458 12384 152464 12436
rect 152516 12424 152522 12436
rect 152553 12427 152611 12433
rect 152553 12424 152565 12427
rect 152516 12396 152565 12424
rect 152516 12384 152522 12396
rect 152553 12393 152565 12396
rect 152599 12393 152611 12427
rect 152553 12387 152611 12393
rect 152844 12396 153424 12424
rect 86126 12356 86132 12368
rect 80164 12328 86132 12356
rect 78582 12180 78588 12232
rect 78640 12220 78646 12232
rect 80164 12229 80192 12328
rect 86126 12316 86132 12328
rect 86184 12316 86190 12368
rect 87414 12316 87420 12368
rect 87472 12356 87478 12368
rect 89441 12359 89499 12365
rect 89441 12356 89453 12359
rect 87472 12328 89453 12356
rect 87472 12316 87478 12328
rect 89441 12325 89453 12328
rect 89487 12325 89499 12359
rect 89441 12319 89499 12325
rect 94516 12328 113174 12356
rect 81434 12248 81440 12300
rect 81492 12288 81498 12300
rect 84473 12291 84531 12297
rect 84473 12288 84485 12291
rect 81492 12260 84485 12288
rect 81492 12248 81498 12260
rect 84473 12257 84485 12260
rect 84519 12257 84531 12291
rect 84654 12288 84660 12300
rect 84615 12260 84660 12288
rect 84473 12251 84531 12257
rect 84654 12248 84660 12260
rect 84712 12248 84718 12300
rect 85758 12288 85764 12300
rect 85040 12260 85764 12288
rect 79229 12223 79287 12229
rect 79229 12220 79241 12223
rect 78640 12192 79241 12220
rect 78640 12180 78646 12192
rect 79229 12189 79241 12192
rect 79275 12220 79287 12223
rect 80149 12223 80207 12229
rect 80149 12220 80161 12223
rect 79275 12192 80161 12220
rect 79275 12189 79287 12192
rect 79229 12183 79287 12189
rect 80149 12189 80161 12192
rect 80195 12189 80207 12223
rect 80149 12183 80207 12189
rect 83826 12180 83832 12232
rect 83884 12220 83890 12232
rect 84381 12223 84439 12229
rect 84381 12220 84393 12223
rect 83884 12192 84393 12220
rect 83884 12180 83890 12192
rect 84381 12189 84393 12192
rect 84427 12220 84439 12223
rect 85040 12220 85068 12260
rect 85758 12248 85764 12260
rect 85816 12248 85822 12300
rect 86310 12248 86316 12300
rect 86368 12288 86374 12300
rect 87049 12291 87107 12297
rect 87049 12288 87061 12291
rect 86368 12260 87061 12288
rect 86368 12248 86374 12260
rect 87049 12257 87061 12260
rect 87095 12288 87107 12291
rect 88150 12288 88156 12300
rect 87095 12260 88156 12288
rect 87095 12257 87107 12260
rect 87049 12251 87107 12257
rect 88150 12248 88156 12260
rect 88208 12248 88214 12300
rect 89162 12288 89168 12300
rect 88904 12260 89168 12288
rect 85482 12220 85488 12232
rect 84427 12192 85068 12220
rect 85443 12192 85488 12220
rect 84427 12189 84439 12192
rect 84381 12183 84439 12189
rect 85482 12180 85488 12192
rect 85540 12180 85546 12232
rect 86034 12180 86040 12232
rect 86092 12220 86098 12232
rect 86865 12223 86923 12229
rect 86865 12220 86877 12223
rect 86092 12192 86877 12220
rect 86092 12180 86098 12192
rect 86865 12189 86877 12192
rect 86911 12189 86923 12223
rect 86865 12183 86923 12189
rect 87969 12223 88027 12229
rect 87969 12189 87981 12223
rect 88015 12220 88027 12223
rect 88242 12220 88248 12232
rect 88015 12192 88248 12220
rect 88015 12189 88027 12192
rect 87969 12183 88027 12189
rect 88242 12180 88248 12192
rect 88300 12180 88306 12232
rect 88797 12223 88855 12229
rect 88797 12189 88809 12223
rect 88843 12222 88855 12223
rect 88904 12222 88932 12260
rect 89162 12248 89168 12260
rect 89220 12288 89226 12300
rect 89220 12260 90128 12288
rect 89220 12248 89226 12260
rect 88843 12194 88932 12222
rect 88843 12189 88855 12194
rect 88797 12183 88855 12189
rect 88978 12180 88984 12232
rect 89036 12220 89042 12232
rect 90100 12229 90128 12260
rect 89625 12223 89683 12229
rect 89625 12220 89637 12223
rect 89036 12192 89637 12220
rect 89036 12180 89042 12192
rect 89625 12189 89637 12192
rect 89671 12189 89683 12223
rect 89625 12183 89683 12189
rect 90085 12223 90143 12229
rect 90085 12189 90097 12223
rect 90131 12220 90143 12223
rect 92014 12220 92020 12232
rect 90131 12192 92020 12220
rect 90131 12189 90143 12192
rect 90085 12183 90143 12189
rect 92014 12180 92020 12192
rect 92072 12180 92078 12232
rect 94516 12152 94544 12328
rect 99098 12248 99104 12300
rect 99156 12288 99162 12300
rect 100941 12291 100999 12297
rect 100941 12288 100953 12291
rect 99156 12260 100953 12288
rect 99156 12248 99162 12260
rect 100941 12257 100953 12260
rect 100987 12288 100999 12291
rect 102042 12288 102048 12300
rect 100987 12260 102048 12288
rect 100987 12257 100999 12260
rect 100941 12251 100999 12257
rect 102042 12248 102048 12260
rect 102100 12288 102106 12300
rect 103149 12291 103207 12297
rect 103149 12288 103161 12291
rect 102100 12260 103161 12288
rect 102100 12248 102106 12260
rect 103149 12257 103161 12260
rect 103195 12288 103207 12291
rect 103238 12288 103244 12300
rect 103195 12260 103244 12288
rect 103195 12257 103207 12260
rect 103149 12251 103207 12257
rect 103238 12248 103244 12260
rect 103296 12248 103302 12300
rect 103330 12248 103336 12300
rect 103388 12288 103394 12300
rect 104529 12291 104587 12297
rect 104529 12288 104541 12291
rect 103388 12260 104541 12288
rect 103388 12248 103394 12260
rect 104529 12257 104541 12260
rect 104575 12257 104587 12291
rect 113146 12288 113174 12328
rect 115750 12316 115756 12368
rect 115808 12356 115814 12368
rect 141970 12356 141976 12368
rect 115808 12328 117820 12356
rect 115808 12316 115814 12328
rect 117792 12297 117820 12328
rect 130396 12328 141976 12356
rect 114373 12291 114431 12297
rect 114373 12288 114385 12291
rect 113146 12260 114385 12288
rect 104529 12251 104587 12257
rect 114373 12257 114385 12260
rect 114419 12288 114431 12291
rect 117777 12291 117835 12297
rect 114419 12260 116808 12288
rect 114419 12257 114431 12260
rect 114373 12251 114431 12257
rect 97534 12180 97540 12232
rect 97592 12220 97598 12232
rect 99285 12223 99343 12229
rect 99285 12220 99297 12223
rect 97592 12192 99297 12220
rect 97592 12180 97598 12192
rect 99285 12189 99297 12192
rect 99331 12189 99343 12223
rect 99285 12183 99343 12189
rect 99745 12223 99803 12229
rect 99745 12189 99757 12223
rect 99791 12220 99803 12223
rect 102965 12223 103023 12229
rect 99791 12192 102180 12220
rect 99791 12189 99803 12192
rect 99745 12183 99803 12189
rect 102152 12164 102180 12192
rect 102965 12189 102977 12223
rect 103011 12220 103023 12223
rect 103698 12220 103704 12232
rect 103011 12192 103704 12220
rect 103011 12189 103023 12192
rect 102965 12183 103023 12189
rect 103698 12180 103704 12192
rect 103756 12180 103762 12232
rect 103793 12223 103851 12229
rect 103793 12189 103805 12223
rect 103839 12220 103851 12223
rect 104437 12223 104495 12229
rect 104437 12220 104449 12223
rect 103839 12192 104449 12220
rect 103839 12189 103851 12192
rect 103793 12183 103851 12189
rect 104437 12189 104449 12192
rect 104483 12220 104495 12223
rect 105081 12223 105139 12229
rect 105081 12220 105093 12223
rect 104483 12192 105093 12220
rect 104483 12189 104495 12192
rect 104437 12183 104495 12189
rect 105081 12189 105093 12192
rect 105127 12189 105139 12223
rect 105081 12183 105139 12189
rect 100754 12152 100760 12164
rect 76576 12124 77892 12152
rect 78508 12124 88840 12152
rect 55858 12084 55864 12096
rect 55186 12056 55864 12084
rect 55858 12044 55864 12056
rect 55916 12044 55922 12096
rect 56042 12084 56048 12096
rect 56003 12056 56048 12084
rect 56042 12044 56048 12056
rect 56100 12044 56106 12096
rect 56152 12093 56180 12124
rect 56137 12087 56195 12093
rect 56137 12053 56149 12087
rect 56183 12053 56195 12087
rect 56137 12047 56195 12053
rect 56505 12087 56563 12093
rect 56505 12053 56517 12087
rect 56551 12084 56563 12087
rect 57330 12084 57336 12096
rect 56551 12056 57336 12084
rect 56551 12053 56563 12056
rect 56505 12047 56563 12053
rect 57330 12044 57336 12056
rect 57388 12044 57394 12096
rect 76282 12084 76288 12096
rect 76243 12056 76288 12084
rect 76282 12044 76288 12056
rect 76340 12044 76346 12096
rect 77864 12093 77892 12124
rect 77849 12087 77907 12093
rect 77849 12053 77861 12087
rect 77895 12084 77907 12087
rect 80238 12084 80244 12096
rect 77895 12056 80244 12084
rect 77895 12053 77907 12056
rect 77849 12047 77907 12053
rect 80238 12044 80244 12056
rect 80296 12044 80302 12096
rect 84010 12084 84016 12096
rect 83971 12056 84016 12084
rect 84010 12044 84016 12056
rect 84068 12044 84074 12096
rect 84654 12044 84660 12096
rect 84712 12084 84718 12096
rect 86310 12084 86316 12096
rect 84712 12056 86316 12084
rect 84712 12044 84718 12056
rect 86310 12044 86316 12056
rect 86368 12044 86374 12096
rect 86773 12087 86831 12093
rect 86773 12053 86785 12087
rect 86819 12084 86831 12087
rect 87506 12084 87512 12096
rect 86819 12056 87512 12084
rect 86819 12053 86831 12056
rect 86773 12047 86831 12053
rect 87506 12044 87512 12056
rect 87564 12044 87570 12096
rect 87601 12087 87659 12093
rect 87601 12053 87613 12087
rect 87647 12084 87659 12087
rect 87782 12084 87788 12096
rect 87647 12056 87788 12084
rect 87647 12053 87659 12056
rect 87601 12047 87659 12053
rect 87782 12044 87788 12056
rect 87840 12044 87846 12096
rect 87966 12044 87972 12096
rect 88024 12084 88030 12096
rect 88061 12087 88119 12093
rect 88061 12084 88073 12087
rect 88024 12056 88073 12084
rect 88024 12044 88030 12056
rect 88061 12053 88073 12056
rect 88107 12084 88119 12087
rect 88702 12084 88708 12096
rect 88107 12056 88708 12084
rect 88107 12053 88119 12056
rect 88061 12047 88119 12053
rect 88702 12044 88708 12056
rect 88760 12044 88766 12096
rect 88812 12084 88840 12124
rect 89686 12124 94544 12152
rect 100715 12124 100760 12152
rect 89686 12084 89714 12124
rect 100754 12112 100760 12124
rect 100812 12112 100818 12164
rect 100849 12155 100907 12161
rect 100849 12121 100861 12155
rect 100895 12152 100907 12155
rect 101030 12152 101036 12164
rect 100895 12124 101036 12152
rect 100895 12121 100907 12124
rect 100849 12115 100907 12121
rect 101030 12112 101036 12124
rect 101088 12112 101094 12164
rect 101950 12152 101956 12164
rect 101911 12124 101956 12152
rect 101950 12112 101956 12124
rect 102008 12112 102014 12164
rect 102134 12112 102140 12164
rect 102192 12152 102198 12164
rect 103808 12152 103836 12183
rect 111886 12180 111892 12232
rect 111944 12220 111950 12232
rect 113269 12223 113327 12229
rect 113269 12220 113281 12223
rect 111944 12192 113281 12220
rect 111944 12180 111950 12192
rect 113269 12189 113281 12192
rect 113315 12189 113327 12223
rect 113269 12183 113327 12189
rect 113913 12223 113971 12229
rect 113913 12189 113925 12223
rect 113959 12220 113971 12223
rect 114278 12220 114284 12232
rect 113959 12192 114284 12220
rect 113959 12189 113971 12192
rect 113913 12183 113971 12189
rect 114278 12180 114284 12192
rect 114336 12180 114342 12232
rect 116780 12220 116808 12260
rect 117777 12257 117789 12291
rect 117823 12288 117835 12291
rect 118878 12288 118884 12300
rect 117823 12260 118884 12288
rect 117823 12257 117835 12260
rect 117777 12251 117835 12257
rect 118878 12248 118884 12260
rect 118936 12248 118942 12300
rect 130396 12288 130424 12328
rect 141970 12316 141976 12328
rect 142028 12316 142034 12368
rect 147582 12316 147588 12368
rect 147640 12356 147646 12368
rect 148413 12359 148471 12365
rect 148413 12356 148425 12359
rect 147640 12328 148425 12356
rect 147640 12316 147646 12328
rect 148413 12325 148425 12328
rect 148459 12325 148471 12359
rect 148413 12319 148471 12325
rect 151630 12316 151636 12368
rect 151688 12356 151694 12368
rect 152734 12356 152740 12368
rect 151688 12328 152740 12356
rect 151688 12316 151694 12328
rect 129108 12260 130424 12288
rect 117593 12223 117651 12229
rect 116780 12192 117268 12220
rect 102192 12124 103836 12152
rect 102192 12112 102198 12124
rect 113818 12112 113824 12164
rect 113876 12152 113882 12164
rect 114649 12155 114707 12161
rect 114649 12152 114661 12155
rect 113876 12124 114661 12152
rect 113876 12112 113882 12124
rect 114649 12121 114661 12124
rect 114695 12121 114707 12155
rect 114649 12115 114707 12121
rect 114756 12124 115138 12152
rect 100386 12084 100392 12096
rect 88812 12056 89714 12084
rect 100347 12056 100392 12084
rect 100386 12044 100392 12056
rect 100444 12044 100450 12096
rect 101968 12084 101996 12112
rect 102318 12084 102324 12096
rect 101968 12056 102324 12084
rect 102318 12044 102324 12056
rect 102376 12044 102382 12096
rect 102594 12084 102600 12096
rect 102555 12056 102600 12084
rect 102594 12044 102600 12056
rect 102652 12044 102658 12096
rect 103054 12084 103060 12096
rect 103015 12056 103060 12084
rect 103054 12044 103060 12056
rect 103112 12044 103118 12096
rect 113910 12044 113916 12096
rect 113968 12084 113974 12096
rect 114756 12084 114784 12124
rect 113968 12056 114784 12084
rect 113968 12044 113974 12056
rect 115658 12044 115664 12096
rect 115716 12084 115722 12096
rect 116121 12087 116179 12093
rect 116121 12084 116133 12087
rect 115716 12056 116133 12084
rect 115716 12044 115722 12056
rect 116121 12053 116133 12056
rect 116167 12053 116179 12087
rect 116121 12047 116179 12053
rect 116394 12044 116400 12096
rect 116452 12084 116458 12096
rect 117133 12087 117191 12093
rect 117133 12084 117145 12087
rect 116452 12056 117145 12084
rect 116452 12044 116458 12056
rect 117133 12053 117145 12056
rect 117179 12053 117191 12087
rect 117240 12084 117268 12192
rect 117593 12189 117605 12223
rect 117639 12220 117651 12223
rect 118050 12220 118056 12232
rect 117639 12192 118056 12220
rect 117639 12189 117651 12192
rect 117593 12183 117651 12189
rect 118050 12180 118056 12192
rect 118108 12180 118114 12232
rect 118326 12220 118332 12232
rect 118287 12192 118332 12220
rect 118326 12180 118332 12192
rect 118384 12180 118390 12232
rect 126146 12180 126152 12232
rect 126204 12220 126210 12232
rect 127897 12223 127955 12229
rect 127897 12220 127909 12223
rect 126204 12192 127909 12220
rect 126204 12180 126210 12192
rect 127897 12189 127909 12192
rect 127943 12189 127955 12223
rect 128630 12220 128636 12232
rect 128591 12192 128636 12220
rect 127897 12183 127955 12189
rect 128630 12180 128636 12192
rect 128688 12180 128694 12232
rect 129108 12229 129136 12260
rect 131022 12248 131028 12300
rect 131080 12288 131086 12300
rect 131853 12291 131911 12297
rect 131853 12288 131865 12291
rect 131080 12260 131865 12288
rect 131080 12248 131086 12260
rect 131853 12257 131865 12260
rect 131899 12288 131911 12291
rect 133230 12288 133236 12300
rect 131899 12260 133236 12288
rect 131899 12257 131911 12260
rect 131853 12251 131911 12257
rect 133230 12248 133236 12260
rect 133288 12248 133294 12300
rect 149054 12248 149060 12300
rect 149112 12288 149118 12300
rect 152093 12291 152151 12297
rect 152093 12288 152105 12291
rect 149112 12260 152105 12288
rect 149112 12248 149118 12260
rect 152093 12257 152105 12260
rect 152139 12257 152151 12291
rect 152093 12251 152151 12257
rect 152185 12291 152243 12297
rect 152185 12257 152197 12291
rect 152231 12257 152243 12291
rect 152185 12251 152243 12257
rect 129093 12223 129151 12229
rect 129093 12189 129105 12223
rect 129139 12189 129151 12223
rect 129093 12183 129151 12189
rect 117501 12155 117559 12161
rect 117501 12121 117513 12155
rect 117547 12152 117559 12155
rect 118234 12152 118240 12164
rect 117547 12124 118240 12152
rect 117547 12121 117559 12124
rect 117501 12115 117559 12121
rect 118234 12112 118240 12124
rect 118292 12112 118298 12164
rect 129108 12152 129136 12183
rect 130470 12180 130476 12232
rect 130528 12180 130534 12232
rect 131669 12223 131727 12229
rect 131669 12189 131681 12223
rect 131715 12220 131727 12223
rect 132402 12220 132408 12232
rect 131715 12192 132408 12220
rect 131715 12189 131727 12192
rect 131669 12183 131727 12189
rect 132402 12180 132408 12192
rect 132460 12180 132466 12232
rect 132586 12220 132592 12232
rect 132547 12192 132592 12220
rect 132586 12180 132592 12192
rect 132644 12180 132650 12232
rect 137738 12220 137744 12232
rect 137699 12192 137744 12220
rect 137738 12180 137744 12192
rect 137796 12180 137802 12232
rect 147493 12223 147551 12229
rect 147493 12189 147505 12223
rect 147539 12220 147551 12223
rect 148042 12220 148048 12232
rect 147539 12192 148048 12220
rect 147539 12189 147551 12192
rect 147493 12183 147551 12189
rect 148042 12180 148048 12192
rect 148100 12180 148106 12232
rect 148321 12223 148379 12229
rect 148321 12189 148333 12223
rect 148367 12220 148379 12223
rect 149330 12220 149336 12232
rect 148367 12192 149336 12220
rect 148367 12189 148379 12192
rect 148321 12183 148379 12189
rect 149330 12180 149336 12192
rect 149388 12180 149394 12232
rect 149422 12180 149428 12232
rect 149480 12220 149486 12232
rect 149480 12192 149525 12220
rect 149480 12180 149486 12192
rect 151354 12180 151360 12232
rect 151412 12220 151418 12232
rect 152200 12220 152228 12251
rect 152476 12229 152504 12328
rect 152734 12316 152740 12328
rect 152792 12316 152798 12368
rect 151412 12192 152228 12220
rect 152461 12223 152519 12229
rect 151412 12180 151418 12192
rect 152461 12189 152473 12223
rect 152507 12189 152519 12223
rect 152461 12183 152519 12189
rect 122806 12124 129136 12152
rect 129369 12155 129427 12161
rect 122806 12084 122834 12124
rect 129369 12121 129381 12155
rect 129415 12121 129427 12155
rect 132494 12152 132500 12164
rect 129369 12115 129427 12121
rect 131316 12124 132500 12152
rect 117240 12056 122834 12084
rect 128449 12087 128507 12093
rect 117133 12047 117191 12053
rect 128449 12053 128461 12087
rect 128495 12084 128507 12087
rect 129384 12084 129412 12115
rect 131316 12093 131344 12124
rect 132494 12112 132500 12124
rect 132552 12112 132558 12164
rect 138014 12152 138020 12164
rect 137975 12124 138020 12152
rect 138014 12112 138020 12124
rect 138072 12152 138078 12164
rect 145837 12155 145895 12161
rect 145837 12152 145849 12155
rect 138072 12124 145849 12152
rect 138072 12112 138078 12124
rect 145837 12121 145849 12124
rect 145883 12121 145895 12155
rect 145837 12115 145895 12121
rect 146205 12155 146263 12161
rect 146205 12121 146217 12155
rect 146251 12152 146263 12155
rect 152844 12152 152872 12396
rect 153289 12359 153347 12365
rect 153289 12325 153301 12359
rect 153335 12325 153347 12359
rect 153396 12356 153424 12396
rect 153746 12384 153752 12436
rect 153804 12424 153810 12436
rect 154117 12427 154175 12433
rect 154117 12424 154129 12427
rect 153804 12396 154129 12424
rect 153804 12384 153810 12396
rect 154117 12393 154129 12396
rect 154163 12393 154175 12427
rect 154117 12387 154175 12393
rect 157242 12384 157248 12436
rect 157300 12424 157306 12436
rect 160922 12424 160928 12436
rect 157300 12396 160928 12424
rect 157300 12384 157306 12396
rect 160922 12384 160928 12396
rect 160980 12384 160986 12436
rect 161566 12384 161572 12436
rect 161624 12424 161630 12436
rect 165341 12427 165399 12433
rect 161624 12396 164924 12424
rect 161624 12384 161630 12396
rect 155034 12356 155040 12368
rect 153396 12328 155040 12356
rect 153289 12319 153347 12325
rect 153304 12220 153332 12319
rect 155034 12316 155040 12328
rect 155092 12316 155098 12368
rect 158898 12316 158904 12368
rect 158956 12356 158962 12368
rect 160005 12359 160063 12365
rect 160005 12356 160017 12359
rect 158956 12328 160017 12356
rect 158956 12316 158962 12328
rect 160005 12325 160017 12328
rect 160051 12325 160063 12359
rect 164896 12356 164924 12396
rect 165341 12393 165353 12427
rect 165387 12424 165399 12427
rect 166442 12424 166448 12436
rect 165387 12396 166448 12424
rect 165387 12393 165399 12396
rect 165341 12387 165399 12393
rect 166442 12384 166448 12396
rect 166500 12384 166506 12436
rect 175921 12427 175979 12433
rect 175921 12393 175933 12427
rect 175967 12424 175979 12427
rect 176470 12424 176476 12436
rect 175967 12396 176476 12424
rect 175967 12393 175979 12396
rect 175921 12387 175979 12393
rect 176470 12384 176476 12396
rect 176528 12384 176534 12436
rect 179506 12384 179512 12436
rect 179564 12424 179570 12436
rect 181349 12427 181407 12433
rect 181349 12424 181361 12427
rect 179564 12396 181361 12424
rect 179564 12384 179570 12396
rect 181349 12393 181361 12396
rect 181395 12393 181407 12427
rect 181349 12387 181407 12393
rect 188525 12427 188583 12433
rect 188525 12393 188537 12427
rect 188571 12424 188583 12427
rect 189166 12424 189172 12436
rect 188571 12396 189172 12424
rect 188571 12393 188583 12396
rect 188525 12387 188583 12393
rect 189166 12384 189172 12396
rect 189224 12384 189230 12436
rect 189626 12384 189632 12436
rect 189684 12424 189690 12436
rect 190181 12427 190239 12433
rect 190181 12424 190193 12427
rect 189684 12396 190193 12424
rect 189684 12384 189690 12396
rect 190181 12393 190193 12396
rect 190227 12393 190239 12427
rect 190181 12387 190239 12393
rect 190822 12384 190828 12436
rect 190880 12424 190886 12436
rect 194042 12424 194048 12436
rect 190880 12396 194048 12424
rect 190880 12384 190886 12396
rect 194042 12384 194048 12396
rect 194100 12384 194106 12436
rect 201681 12427 201739 12433
rect 194152 12396 197584 12424
rect 165430 12356 165436 12368
rect 164896 12328 165436 12356
rect 160005 12319 160063 12325
rect 165430 12316 165436 12328
rect 165488 12316 165494 12368
rect 166074 12356 166080 12368
rect 166035 12328 166080 12356
rect 166074 12316 166080 12328
rect 166132 12316 166138 12368
rect 177758 12356 177764 12368
rect 177040 12328 177764 12356
rect 153933 12291 153991 12297
rect 153933 12257 153945 12291
rect 153979 12288 153991 12291
rect 154114 12288 154120 12300
rect 153979 12260 154120 12288
rect 153979 12257 153991 12260
rect 153933 12251 153991 12257
rect 154114 12248 154120 12260
rect 154172 12248 154178 12300
rect 160370 12248 160376 12300
rect 160428 12288 160434 12300
rect 161293 12291 161351 12297
rect 161293 12288 161305 12291
rect 160428 12260 161305 12288
rect 160428 12248 160434 12260
rect 161293 12257 161305 12260
rect 161339 12257 161351 12291
rect 161293 12251 161351 12257
rect 161474 12248 161480 12300
rect 161532 12288 161538 12300
rect 162486 12288 162492 12300
rect 161532 12260 161577 12288
rect 162447 12260 162492 12288
rect 161532 12248 161538 12260
rect 162486 12248 162492 12260
rect 162544 12248 162550 12300
rect 162670 12288 162676 12300
rect 162631 12260 162676 12288
rect 162670 12248 162676 12260
rect 162728 12248 162734 12300
rect 163590 12288 163596 12300
rect 163551 12260 163596 12288
rect 163590 12248 163596 12260
rect 163648 12248 163654 12300
rect 177040 12297 177068 12328
rect 177758 12316 177764 12328
rect 177816 12316 177822 12368
rect 180886 12356 180892 12368
rect 180847 12328 180892 12356
rect 180886 12316 180892 12328
rect 180944 12316 180950 12368
rect 192570 12356 192576 12368
rect 185596 12328 190500 12356
rect 192531 12328 192576 12356
rect 177025 12291 177083 12297
rect 177025 12257 177037 12291
rect 177071 12257 177083 12291
rect 177025 12251 177083 12257
rect 177114 12248 177120 12300
rect 177172 12288 177178 12300
rect 185596 12288 185624 12328
rect 177172 12260 177217 12288
rect 179156 12260 185624 12288
rect 177172 12248 177178 12260
rect 154301 12223 154359 12229
rect 154301 12220 154313 12223
rect 153304 12192 154313 12220
rect 154301 12189 154313 12192
rect 154347 12189 154359 12223
rect 154301 12183 154359 12189
rect 158806 12180 158812 12232
rect 158864 12220 158870 12232
rect 160189 12223 160247 12229
rect 160189 12220 160201 12223
rect 158864 12192 160201 12220
rect 158864 12180 158870 12192
rect 160189 12189 160201 12192
rect 160235 12189 160247 12223
rect 160189 12183 160247 12189
rect 161201 12223 161259 12229
rect 161201 12189 161213 12223
rect 161247 12220 161259 12223
rect 161750 12220 161756 12232
rect 161247 12192 161756 12220
rect 161247 12189 161259 12192
rect 161201 12183 161259 12189
rect 161750 12180 161756 12192
rect 161808 12220 161814 12232
rect 162504 12220 162532 12248
rect 179156 12232 179184 12260
rect 187970 12248 187976 12300
rect 188028 12288 188034 12300
rect 188028 12260 190408 12288
rect 188028 12248 188034 12260
rect 161808 12192 162532 12220
rect 176105 12223 176163 12229
rect 161808 12180 161814 12192
rect 176105 12189 176117 12223
rect 176151 12220 176163 12223
rect 176933 12223 176991 12229
rect 176933 12220 176945 12223
rect 176151 12192 176945 12220
rect 176151 12189 176163 12192
rect 176105 12183 176163 12189
rect 176933 12189 176945 12192
rect 176979 12220 176991 12223
rect 177850 12220 177856 12232
rect 176979 12192 177856 12220
rect 176979 12189 176991 12192
rect 176933 12183 176991 12189
rect 177850 12180 177856 12192
rect 177908 12180 177914 12232
rect 179138 12220 179144 12232
rect 179099 12192 179144 12220
rect 179138 12180 179144 12192
rect 179196 12180 179202 12232
rect 180702 12180 180708 12232
rect 180760 12220 180766 12232
rect 181533 12223 181591 12229
rect 181533 12220 181545 12223
rect 180760 12192 181545 12220
rect 180760 12180 180766 12192
rect 181533 12189 181545 12192
rect 181579 12189 181591 12223
rect 181533 12183 181591 12189
rect 188709 12223 188767 12229
rect 188709 12189 188721 12223
rect 188755 12189 188767 12223
rect 189534 12220 189540 12232
rect 189495 12192 189540 12220
rect 188709 12183 188767 12189
rect 146251 12124 147674 12152
rect 146251 12121 146263 12124
rect 146205 12115 146263 12121
rect 128495 12056 129412 12084
rect 131301 12087 131359 12093
rect 128495 12053 128507 12056
rect 128449 12047 128507 12053
rect 131301 12053 131313 12087
rect 131347 12053 131359 12087
rect 131301 12047 131359 12053
rect 131574 12044 131580 12096
rect 131632 12084 131638 12096
rect 131761 12087 131819 12093
rect 131761 12084 131773 12087
rect 131632 12056 131773 12084
rect 131632 12044 131638 12056
rect 131761 12053 131773 12056
rect 131807 12053 131819 12087
rect 147646 12084 147674 12124
rect 149440 12124 152872 12152
rect 153657 12155 153715 12161
rect 149440 12084 149468 12124
rect 153657 12121 153669 12155
rect 153703 12152 153715 12155
rect 155862 12152 155868 12164
rect 153703 12124 155868 12152
rect 153703 12121 153715 12124
rect 153657 12115 153715 12121
rect 155862 12112 155868 12124
rect 155920 12112 155926 12164
rect 156414 12112 156420 12164
rect 156472 12152 156478 12164
rect 162578 12152 162584 12164
rect 156472 12124 162584 12152
rect 156472 12112 156478 12124
rect 162578 12112 162584 12124
rect 162636 12112 162642 12164
rect 162670 12112 162676 12164
rect 162728 12152 162734 12164
rect 163869 12155 163927 12161
rect 163869 12152 163881 12155
rect 162728 12124 163881 12152
rect 162728 12112 162734 12124
rect 163869 12121 163881 12124
rect 163915 12121 163927 12155
rect 163869 12115 163927 12121
rect 164326 12112 164332 12164
rect 164384 12112 164390 12164
rect 165890 12152 165896 12164
rect 165851 12124 165896 12152
rect 165890 12112 165896 12124
rect 165948 12112 165954 12164
rect 166534 12112 166540 12164
rect 166592 12152 166598 12164
rect 177945 12155 178003 12161
rect 177945 12152 177957 12155
rect 166592 12124 177957 12152
rect 166592 12112 166598 12124
rect 177945 12121 177957 12124
rect 177991 12152 178003 12155
rect 179414 12152 179420 12164
rect 177991 12124 179276 12152
rect 179375 12124 179420 12152
rect 177991 12121 178003 12124
rect 177945 12115 178003 12121
rect 147646 12056 149468 12084
rect 131761 12047 131819 12053
rect 149514 12044 149520 12096
rect 149572 12084 149578 12096
rect 150713 12087 150771 12093
rect 150713 12084 150725 12087
rect 149572 12056 150725 12084
rect 149572 12044 149578 12056
rect 150713 12053 150725 12056
rect 150759 12053 150771 12087
rect 151630 12084 151636 12096
rect 151591 12056 151636 12084
rect 150713 12047 150771 12053
rect 151630 12044 151636 12056
rect 151688 12044 151694 12096
rect 151722 12044 151728 12096
rect 151780 12084 151786 12096
rect 152001 12087 152059 12093
rect 152001 12084 152013 12087
rect 151780 12056 152013 12084
rect 151780 12044 151786 12056
rect 152001 12053 152013 12056
rect 152047 12053 152059 12087
rect 152001 12047 152059 12053
rect 152182 12044 152188 12096
rect 152240 12084 152246 12096
rect 152550 12084 152556 12096
rect 152240 12056 152556 12084
rect 152240 12044 152246 12056
rect 152550 12044 152556 12056
rect 152608 12084 152614 12096
rect 153749 12087 153807 12093
rect 153749 12084 153761 12087
rect 152608 12056 153761 12084
rect 152608 12044 152614 12056
rect 153749 12053 153761 12056
rect 153795 12053 153807 12087
rect 153749 12047 153807 12053
rect 160833 12087 160891 12093
rect 160833 12053 160845 12087
rect 160879 12084 160891 12087
rect 161106 12084 161112 12096
rect 160879 12056 161112 12084
rect 160879 12053 160891 12056
rect 160833 12047 160891 12053
rect 161106 12044 161112 12056
rect 161164 12044 161170 12096
rect 162029 12087 162087 12093
rect 162029 12053 162041 12087
rect 162075 12084 162087 12087
rect 162210 12084 162216 12096
rect 162075 12056 162216 12084
rect 162075 12053 162087 12056
rect 162029 12047 162087 12053
rect 162210 12044 162216 12056
rect 162268 12044 162274 12096
rect 162397 12087 162455 12093
rect 162397 12053 162409 12087
rect 162443 12084 162455 12087
rect 162854 12084 162860 12096
rect 162443 12056 162860 12084
rect 162443 12053 162455 12056
rect 162397 12047 162455 12053
rect 162854 12044 162860 12056
rect 162912 12044 162918 12096
rect 176565 12087 176623 12093
rect 176565 12053 176577 12087
rect 176611 12084 176623 12087
rect 176654 12084 176660 12096
rect 176611 12056 176660 12084
rect 176611 12053 176623 12056
rect 176565 12047 176623 12053
rect 176654 12044 176660 12056
rect 176712 12044 176718 12096
rect 178034 12084 178040 12096
rect 177995 12056 178040 12084
rect 178034 12044 178040 12056
rect 178092 12044 178098 12096
rect 179248 12084 179276 12124
rect 179414 12112 179420 12124
rect 179472 12112 179478 12164
rect 181438 12152 181444 12164
rect 180642 12124 181444 12152
rect 181438 12112 181444 12124
rect 181496 12112 181502 12164
rect 188724 12152 188752 12183
rect 189534 12180 189540 12192
rect 189592 12180 189598 12232
rect 190380 12229 190408 12260
rect 190365 12223 190423 12229
rect 190365 12189 190377 12223
rect 190411 12189 190423 12223
rect 190472 12220 190500 12328
rect 192570 12316 192576 12328
rect 192628 12316 192634 12368
rect 190825 12291 190883 12297
rect 190825 12257 190837 12291
rect 190871 12288 190883 12291
rect 191834 12288 191840 12300
rect 190871 12260 191840 12288
rect 190871 12257 190883 12260
rect 190825 12251 190883 12257
rect 190840 12220 190868 12251
rect 191834 12248 191840 12260
rect 191892 12248 191898 12300
rect 192662 12248 192668 12300
rect 192720 12288 192726 12300
rect 193677 12291 193735 12297
rect 193677 12288 193689 12291
rect 192720 12260 193689 12288
rect 192720 12248 192726 12260
rect 193677 12257 193689 12260
rect 193723 12288 193735 12291
rect 194152 12288 194180 12396
rect 197446 12356 197452 12368
rect 196452 12328 197452 12356
rect 193723 12260 194180 12288
rect 194428 12260 196020 12288
rect 193723 12257 193735 12260
rect 193677 12251 193735 12257
rect 194428 12232 194456 12260
rect 194410 12220 194416 12232
rect 190472 12192 190868 12220
rect 192404 12192 193812 12220
rect 194371 12192 194416 12220
rect 190365 12183 190423 12189
rect 190822 12152 190828 12164
rect 188724 12124 190828 12152
rect 190822 12112 190828 12124
rect 190880 12112 190886 12164
rect 191098 12152 191104 12164
rect 191059 12124 191104 12152
rect 191098 12112 191104 12124
rect 191156 12112 191162 12164
rect 191190 12112 191196 12164
rect 191248 12152 191254 12164
rect 191248 12124 191590 12152
rect 191248 12112 191254 12124
rect 180150 12084 180156 12096
rect 179248 12056 180156 12084
rect 180150 12044 180156 12056
rect 180208 12044 180214 12096
rect 189629 12087 189687 12093
rect 189629 12053 189641 12087
rect 189675 12084 189687 12087
rect 192404 12084 192432 12192
rect 193398 12152 193404 12164
rect 193359 12124 193404 12152
rect 193398 12112 193404 12124
rect 193456 12112 193462 12164
rect 193030 12084 193036 12096
rect 189675 12056 192432 12084
rect 192991 12056 193036 12084
rect 189675 12053 189687 12056
rect 189629 12047 189687 12053
rect 193030 12044 193036 12056
rect 193088 12044 193094 12096
rect 193493 12087 193551 12093
rect 193493 12053 193505 12087
rect 193539 12084 193551 12087
rect 193674 12084 193680 12096
rect 193539 12056 193680 12084
rect 193539 12053 193551 12056
rect 193493 12047 193551 12053
rect 193674 12044 193680 12056
rect 193732 12044 193738 12096
rect 193784 12084 193812 12192
rect 194410 12180 194416 12192
rect 194468 12180 194474 12232
rect 194686 12152 194692 12164
rect 194647 12124 194692 12152
rect 194686 12112 194692 12124
rect 194744 12112 194750 12164
rect 195992 12152 196020 12260
rect 196452 12229 196480 12328
rect 197446 12316 197452 12328
rect 197504 12316 197510 12368
rect 197556 12297 197584 12396
rect 201681 12393 201693 12427
rect 201727 12424 201739 12427
rect 202414 12424 202420 12436
rect 201727 12396 202420 12424
rect 201727 12393 201739 12396
rect 201681 12387 201739 12393
rect 202414 12384 202420 12396
rect 202472 12384 202478 12436
rect 205634 12424 205640 12436
rect 203628 12396 205640 12424
rect 201129 12359 201187 12365
rect 201129 12325 201141 12359
rect 201175 12356 201187 12359
rect 203628 12356 203656 12396
rect 205634 12384 205640 12396
rect 205692 12384 205698 12436
rect 206465 12427 206523 12433
rect 206465 12393 206477 12427
rect 206511 12424 206523 12427
rect 207658 12424 207664 12436
rect 206511 12396 207664 12424
rect 206511 12393 206523 12396
rect 206465 12387 206523 12393
rect 207658 12384 207664 12396
rect 207716 12384 207722 12436
rect 227796 12427 227854 12433
rect 227796 12393 227808 12427
rect 227842 12424 227854 12427
rect 230106 12424 230112 12436
rect 227842 12396 230112 12424
rect 227842 12393 227854 12396
rect 227796 12387 227854 12393
rect 230106 12384 230112 12396
rect 230164 12384 230170 12436
rect 231854 12384 231860 12436
rect 231912 12424 231918 12436
rect 232225 12427 232283 12433
rect 232225 12424 232237 12427
rect 231912 12396 232237 12424
rect 231912 12384 231918 12396
rect 232225 12393 232237 12396
rect 232271 12393 232283 12427
rect 232225 12387 232283 12393
rect 239030 12384 239036 12436
rect 239088 12424 239094 12436
rect 239953 12427 240011 12433
rect 239953 12424 239965 12427
rect 239088 12396 239965 12424
rect 239088 12384 239094 12396
rect 239953 12393 239965 12396
rect 239999 12393 240011 12427
rect 239953 12387 240011 12393
rect 240134 12384 240140 12436
rect 240192 12424 240198 12436
rect 243541 12427 243599 12433
rect 240192 12396 241192 12424
rect 240192 12384 240198 12396
rect 201175 12328 203656 12356
rect 201175 12325 201187 12328
rect 201129 12319 201187 12325
rect 228818 12316 228824 12368
rect 228876 12356 228882 12368
rect 229741 12359 229799 12365
rect 229741 12356 229753 12359
rect 228876 12328 229753 12356
rect 228876 12316 228882 12328
rect 229741 12325 229753 12328
rect 229787 12325 229799 12359
rect 229741 12319 229799 12325
rect 231118 12316 231124 12368
rect 231176 12356 231182 12368
rect 232498 12356 232504 12368
rect 231176 12328 232504 12356
rect 231176 12316 231182 12328
rect 232498 12316 232504 12328
rect 232556 12316 232562 12368
rect 238757 12359 238815 12365
rect 238757 12325 238769 12359
rect 238803 12356 238815 12359
rect 241164 12356 241192 12396
rect 242360 12396 243124 12424
rect 242250 12356 242256 12368
rect 238803 12328 239720 12356
rect 238803 12325 238815 12328
rect 238757 12319 238815 12325
rect 197541 12291 197599 12297
rect 196544 12260 196848 12288
rect 196437 12223 196495 12229
rect 196437 12189 196449 12223
rect 196483 12189 196495 12223
rect 196437 12183 196495 12189
rect 196544 12152 196572 12260
rect 196713 12223 196771 12229
rect 196713 12220 196725 12223
rect 194796 12124 195178 12152
rect 195992 12124 196572 12152
rect 196636 12192 196725 12220
rect 194796 12084 194824 12124
rect 193784 12056 194824 12084
rect 194962 12044 194968 12096
rect 195020 12084 195026 12096
rect 196636 12084 196664 12192
rect 196713 12189 196725 12192
rect 196759 12189 196771 12223
rect 196713 12183 196771 12189
rect 196820 12152 196848 12260
rect 197541 12257 197553 12291
rect 197587 12257 197599 12291
rect 197541 12251 197599 12257
rect 200482 12248 200488 12300
rect 200540 12288 200546 12300
rect 200540 12260 201908 12288
rect 200540 12248 200546 12260
rect 197446 12220 197452 12232
rect 197359 12192 197452 12220
rect 197446 12180 197452 12192
rect 197504 12220 197510 12232
rect 198366 12220 198372 12232
rect 197504 12192 198372 12220
rect 197504 12180 197510 12192
rect 198366 12180 198372 12192
rect 198424 12180 198430 12232
rect 200574 12180 200580 12232
rect 200632 12220 200638 12232
rect 201034 12220 201040 12232
rect 200632 12192 201040 12220
rect 200632 12180 200638 12192
rect 201034 12180 201040 12192
rect 201092 12180 201098 12232
rect 201880 12229 201908 12260
rect 202046 12248 202052 12300
rect 202104 12288 202110 12300
rect 203518 12288 203524 12300
rect 202104 12260 203524 12288
rect 202104 12248 202110 12260
rect 203518 12248 203524 12260
rect 203576 12248 203582 12300
rect 204717 12291 204775 12297
rect 204717 12257 204729 12291
rect 204763 12288 204775 12291
rect 231581 12291 231639 12297
rect 204763 12260 209774 12288
rect 204763 12257 204775 12260
rect 204717 12251 204775 12257
rect 201865 12223 201923 12229
rect 201865 12189 201877 12223
rect 201911 12189 201923 12223
rect 201865 12183 201923 12189
rect 203245 12223 203303 12229
rect 203245 12189 203257 12223
rect 203291 12220 203303 12223
rect 204530 12220 204536 12232
rect 203291 12192 204536 12220
rect 203291 12189 203303 12192
rect 203245 12183 203303 12189
rect 204530 12180 204536 12192
rect 204588 12180 204594 12232
rect 204732 12152 204760 12251
rect 209746 12220 209774 12260
rect 227548 12260 231440 12288
rect 227548 12229 227576 12260
rect 227533 12223 227591 12229
rect 227533 12220 227545 12223
rect 209746 12192 227545 12220
rect 227533 12189 227545 12192
rect 227579 12189 227591 12223
rect 229922 12220 229928 12232
rect 229835 12192 229928 12220
rect 227533 12183 227591 12189
rect 229922 12180 229928 12192
rect 229980 12220 229986 12232
rect 231302 12220 231308 12232
rect 229980 12192 231308 12220
rect 229980 12180 229986 12192
rect 231302 12180 231308 12192
rect 231360 12180 231366 12232
rect 204990 12152 204996 12164
rect 196820 12124 204760 12152
rect 204951 12124 204996 12152
rect 204990 12112 204996 12124
rect 205048 12112 205054 12164
rect 230842 12152 230848 12164
rect 205100 12124 205482 12152
rect 229034 12124 230848 12152
rect 196802 12084 196808 12096
rect 195020 12056 196664 12084
rect 196763 12056 196808 12084
rect 195020 12044 195026 12056
rect 196802 12044 196808 12056
rect 196860 12044 196866 12096
rect 196986 12084 196992 12096
rect 196947 12056 196992 12084
rect 196986 12044 196992 12056
rect 197044 12044 197050 12096
rect 197354 12084 197360 12096
rect 197315 12056 197360 12084
rect 197354 12044 197360 12056
rect 197412 12044 197418 12096
rect 202877 12087 202935 12093
rect 202877 12053 202889 12087
rect 202923 12084 202935 12087
rect 203058 12084 203064 12096
rect 202923 12056 203064 12084
rect 202923 12053 202935 12056
rect 202877 12047 202935 12053
rect 203058 12044 203064 12056
rect 203116 12044 203122 12096
rect 203337 12087 203395 12093
rect 203337 12053 203349 12087
rect 203383 12084 203395 12087
rect 203426 12084 203432 12096
rect 203383 12056 203432 12084
rect 203383 12053 203395 12056
rect 203337 12047 203395 12053
rect 203426 12044 203432 12056
rect 203484 12044 203490 12096
rect 204254 12044 204260 12096
rect 204312 12084 204318 12096
rect 205100 12084 205128 12124
rect 230842 12112 230848 12124
rect 230900 12112 230906 12164
rect 231118 12112 231124 12164
rect 231176 12152 231182 12164
rect 231412 12152 231440 12260
rect 231581 12257 231593 12291
rect 231627 12288 231639 12291
rect 231670 12288 231676 12300
rect 231627 12260 231676 12288
rect 231627 12257 231639 12260
rect 231581 12251 231639 12257
rect 231670 12248 231676 12260
rect 231728 12248 231734 12300
rect 238846 12248 238852 12300
rect 238904 12288 238910 12300
rect 239306 12288 239312 12300
rect 238904 12260 239312 12288
rect 238904 12248 238910 12260
rect 239306 12248 239312 12260
rect 239364 12248 239370 12300
rect 232130 12220 232136 12232
rect 232043 12192 232136 12220
rect 232130 12180 232136 12192
rect 232188 12220 232194 12232
rect 233050 12220 233056 12232
rect 232188 12192 233056 12220
rect 232188 12180 232194 12192
rect 233050 12180 233056 12192
rect 233108 12180 233114 12232
rect 238018 12220 238024 12232
rect 237979 12192 238024 12220
rect 238018 12180 238024 12192
rect 238076 12180 238082 12232
rect 238386 12180 238392 12232
rect 238444 12220 238450 12232
rect 239122 12220 239128 12232
rect 238444 12192 239128 12220
rect 238444 12180 238450 12192
rect 239122 12180 239128 12192
rect 239180 12180 239186 12232
rect 239217 12223 239275 12229
rect 239217 12189 239229 12223
rect 239263 12220 239275 12223
rect 239490 12220 239496 12232
rect 239263 12192 239496 12220
rect 239263 12189 239275 12192
rect 239217 12183 239275 12189
rect 239490 12180 239496 12192
rect 239548 12180 239554 12232
rect 239692 12220 239720 12328
rect 239968 12328 241008 12356
rect 241164 12328 242256 12356
rect 239968 12300 239996 12328
rect 239950 12248 239956 12300
rect 240008 12248 240014 12300
rect 240980 12288 241008 12328
rect 242250 12316 242256 12328
rect 242308 12316 242314 12368
rect 242360 12365 242388 12396
rect 242345 12359 242403 12365
rect 242345 12325 242357 12359
rect 242391 12325 242403 12359
rect 242986 12356 242992 12368
rect 242345 12319 242403 12325
rect 242728 12328 242992 12356
rect 241425 12291 241483 12297
rect 241425 12288 241437 12291
rect 240980 12260 241437 12288
rect 241425 12257 241437 12260
rect 241471 12288 241483 12291
rect 241471 12260 242296 12288
rect 241471 12257 241483 12260
rect 241425 12251 241483 12257
rect 242268 12236 242296 12260
rect 242434 12248 242440 12300
rect 242492 12288 242498 12300
rect 242728 12288 242756 12328
rect 242986 12316 242992 12328
rect 243044 12316 243050 12368
rect 242805 12291 242863 12297
rect 242805 12288 242817 12291
rect 242492 12260 242817 12288
rect 242492 12248 242498 12260
rect 242805 12257 242817 12260
rect 242851 12257 242863 12291
rect 242805 12251 242863 12257
rect 242894 12248 242900 12300
rect 242952 12288 242958 12300
rect 242952 12260 243045 12288
rect 242952 12248 242958 12260
rect 240137 12223 240195 12229
rect 240137 12220 240149 12223
rect 239692 12192 240149 12220
rect 240137 12189 240149 12192
rect 240183 12189 240195 12223
rect 240137 12183 240195 12189
rect 241241 12223 241299 12229
rect 241241 12189 241253 12223
rect 241287 12220 241299 12223
rect 242158 12220 242164 12232
rect 241287 12192 242164 12220
rect 241287 12189 241299 12192
rect 241241 12183 241299 12189
rect 242158 12180 242164 12192
rect 242216 12180 242222 12232
rect 242268 12220 242388 12236
rect 242268 12216 242848 12220
rect 242912 12216 242940 12248
rect 242268 12208 242940 12216
rect 242360 12192 242940 12208
rect 243096 12220 243124 12396
rect 243541 12393 243553 12427
rect 243587 12424 243599 12427
rect 243630 12424 243636 12436
rect 243587 12396 243636 12424
rect 243587 12393 243599 12396
rect 243541 12387 243599 12393
rect 243630 12384 243636 12396
rect 243688 12384 243694 12436
rect 244182 12424 244188 12436
rect 244143 12396 244188 12424
rect 244182 12384 244188 12396
rect 244240 12384 244246 12436
rect 251085 12427 251143 12433
rect 251085 12393 251097 12427
rect 251131 12424 251143 12427
rect 251358 12424 251364 12436
rect 251131 12396 251364 12424
rect 251131 12393 251143 12396
rect 251085 12387 251143 12393
rect 251358 12384 251364 12396
rect 251416 12384 251422 12436
rect 251910 12384 251916 12436
rect 251968 12424 251974 12436
rect 251968 12396 256280 12424
rect 251968 12384 251974 12396
rect 251450 12316 251456 12368
rect 251508 12356 251514 12368
rect 252094 12356 252100 12368
rect 251508 12328 252100 12356
rect 251508 12316 251514 12328
rect 252094 12316 252100 12328
rect 252152 12316 252158 12368
rect 254302 12356 254308 12368
rect 254215 12328 254308 12356
rect 254302 12316 254308 12328
rect 254360 12356 254366 12368
rect 255222 12356 255228 12368
rect 254360 12328 255228 12356
rect 254360 12316 254366 12328
rect 255222 12316 255228 12328
rect 255280 12316 255286 12368
rect 243170 12248 243176 12300
rect 243228 12288 243234 12300
rect 243228 12260 244412 12288
rect 243228 12248 243234 12260
rect 244384 12229 244412 12260
rect 248322 12248 248328 12300
rect 248380 12288 248386 12300
rect 249242 12288 249248 12300
rect 248380 12260 249248 12288
rect 248380 12248 248386 12260
rect 249242 12248 249248 12260
rect 249300 12248 249306 12300
rect 252557 12291 252615 12297
rect 252557 12288 252569 12291
rect 251146 12260 252569 12288
rect 243725 12223 243783 12229
rect 243725 12220 243737 12223
rect 243096 12192 243737 12220
rect 242820 12188 242940 12192
rect 243725 12189 243737 12192
rect 243771 12189 243783 12223
rect 243725 12183 243783 12189
rect 244369 12223 244427 12229
rect 244369 12189 244381 12223
rect 244415 12189 244427 12223
rect 251146 12220 251174 12260
rect 252557 12257 252569 12260
rect 252603 12288 252615 12291
rect 255317 12291 255375 12297
rect 252603 12260 255268 12288
rect 252603 12257 252615 12260
rect 252557 12251 252615 12257
rect 244369 12183 244427 12189
rect 248386 12192 251174 12220
rect 248386 12152 248414 12192
rect 251266 12180 251272 12232
rect 251324 12220 251330 12232
rect 251910 12220 251916 12232
rect 251324 12192 251369 12220
rect 251871 12192 251916 12220
rect 251324 12180 251330 12192
rect 251910 12180 251916 12192
rect 251968 12180 251974 12232
rect 255130 12220 255136 12232
rect 255091 12192 255136 12220
rect 255130 12180 255136 12192
rect 255188 12180 255194 12232
rect 249058 12152 249064 12164
rect 231176 12124 231348 12152
rect 231412 12124 248414 12152
rect 249019 12124 249064 12152
rect 231176 12112 231182 12124
rect 204312 12056 205128 12084
rect 204312 12044 204318 12056
rect 228818 12044 228824 12096
rect 228876 12084 228882 12096
rect 229281 12087 229339 12093
rect 229281 12084 229293 12087
rect 228876 12056 229293 12084
rect 228876 12044 228882 12056
rect 229281 12053 229293 12056
rect 229327 12053 229339 12087
rect 229281 12047 229339 12053
rect 230937 12087 230995 12093
rect 230937 12053 230949 12087
rect 230983 12084 230995 12087
rect 231210 12084 231216 12096
rect 230983 12056 231216 12084
rect 230983 12053 230995 12056
rect 230937 12047 230995 12053
rect 231210 12044 231216 12056
rect 231268 12044 231274 12096
rect 231320 12093 231348 12124
rect 249058 12112 249064 12124
rect 249116 12112 249122 12164
rect 249242 12112 249248 12164
rect 249300 12152 249306 12164
rect 251928 12152 251956 12180
rect 249300 12124 251956 12152
rect 252833 12155 252891 12161
rect 249300 12112 249306 12124
rect 252833 12121 252845 12155
rect 252879 12152 252891 12155
rect 253106 12152 253112 12164
rect 252879 12124 253112 12152
rect 252879 12121 252891 12124
rect 252833 12115 252891 12121
rect 253106 12112 253112 12124
rect 253164 12112 253170 12164
rect 255240 12152 255268 12260
rect 255317 12257 255329 12291
rect 255363 12288 255375 12291
rect 255590 12288 255596 12300
rect 255363 12260 255596 12288
rect 255363 12257 255375 12260
rect 255317 12251 255375 12257
rect 255590 12248 255596 12260
rect 255648 12248 255654 12300
rect 256252 12288 256280 12396
rect 256510 12384 256516 12436
rect 256568 12424 256574 12436
rect 256881 12427 256939 12433
rect 256881 12424 256893 12427
rect 256568 12396 256893 12424
rect 256568 12384 256574 12396
rect 256881 12393 256893 12396
rect 256927 12393 256939 12427
rect 262490 12424 262496 12436
rect 262451 12396 262496 12424
rect 256881 12387 256939 12393
rect 262490 12384 262496 12396
rect 262548 12384 262554 12436
rect 264609 12427 264667 12433
rect 264609 12393 264621 12427
rect 264655 12424 264667 12427
rect 265526 12424 265532 12436
rect 264655 12396 265532 12424
rect 264655 12393 264667 12396
rect 264609 12387 264667 12393
rect 265526 12384 265532 12396
rect 265584 12384 265590 12436
rect 268010 12424 268016 12436
rect 265912 12396 268016 12424
rect 256329 12359 256387 12365
rect 256329 12325 256341 12359
rect 256375 12356 256387 12359
rect 256970 12356 256976 12368
rect 256375 12328 256976 12356
rect 256375 12325 256387 12328
rect 256329 12319 256387 12325
rect 256970 12316 256976 12328
rect 257028 12316 257034 12368
rect 264057 12359 264115 12365
rect 264057 12325 264069 12359
rect 264103 12356 264115 12359
rect 264974 12356 264980 12368
rect 264103 12328 264980 12356
rect 264103 12325 264115 12328
rect 264057 12319 264115 12325
rect 264974 12316 264980 12328
rect 265032 12316 265038 12368
rect 265912 12356 265940 12396
rect 268010 12384 268016 12396
rect 268068 12384 268074 12436
rect 268378 12384 268384 12436
rect 268436 12424 268442 12436
rect 271046 12424 271052 12436
rect 268436 12396 270080 12424
rect 271007 12396 271052 12424
rect 268436 12384 268442 12396
rect 265084 12328 265940 12356
rect 270052 12356 270080 12396
rect 271046 12384 271052 12396
rect 271104 12384 271110 12436
rect 305454 12424 305460 12436
rect 305415 12396 305460 12424
rect 305454 12384 305460 12396
rect 305512 12384 305518 12436
rect 271693 12359 271751 12365
rect 271693 12356 271705 12359
rect 270052 12328 271705 12356
rect 261846 12288 261852 12300
rect 256252 12260 261852 12288
rect 261846 12248 261852 12260
rect 261904 12248 261910 12300
rect 262398 12248 262404 12300
rect 262456 12288 262462 12300
rect 262456 12260 264008 12288
rect 262456 12248 262462 12260
rect 256234 12220 256240 12232
rect 256195 12192 256240 12220
rect 256234 12180 256240 12192
rect 256292 12180 256298 12232
rect 256326 12180 256332 12232
rect 256384 12220 256390 12232
rect 257065 12223 257123 12229
rect 257065 12220 257077 12223
rect 256384 12192 257077 12220
rect 256384 12180 256390 12192
rect 257065 12189 257077 12192
rect 257111 12189 257123 12223
rect 257065 12183 257123 12189
rect 262677 12223 262735 12229
rect 262677 12189 262689 12223
rect 262723 12220 262735 12223
rect 263042 12220 263048 12232
rect 262723 12192 263048 12220
rect 262723 12189 262735 12192
rect 262677 12183 262735 12189
rect 263042 12180 263048 12192
rect 263100 12180 263106 12232
rect 263980 12229 264008 12260
rect 264146 12248 264152 12300
rect 264204 12288 264210 12300
rect 265084 12288 265112 12328
rect 264204 12260 265112 12288
rect 264204 12248 264210 12260
rect 265158 12248 265164 12300
rect 265216 12288 265222 12300
rect 265216 12260 265388 12288
rect 265216 12248 265222 12260
rect 263965 12223 264023 12229
rect 263965 12189 263977 12223
rect 264011 12220 264023 12223
rect 264330 12220 264336 12232
rect 264011 12192 264336 12220
rect 264011 12189 264023 12192
rect 263965 12183 264023 12189
rect 264330 12180 264336 12192
rect 264388 12180 264394 12232
rect 264793 12223 264851 12229
rect 264793 12189 264805 12223
rect 264839 12220 264851 12223
rect 265360 12220 265388 12260
rect 265618 12248 265624 12300
rect 265676 12288 265682 12300
rect 265912 12297 265940 12328
rect 271693 12325 271705 12328
rect 271739 12325 271751 12359
rect 271693 12319 271751 12325
rect 265713 12291 265771 12297
rect 265713 12288 265725 12291
rect 265676 12260 265725 12288
rect 265676 12248 265682 12260
rect 265713 12257 265725 12260
rect 265759 12257 265771 12291
rect 265713 12251 265771 12257
rect 265897 12291 265955 12297
rect 265897 12257 265909 12291
rect 265943 12257 265955 12291
rect 268749 12291 268807 12297
rect 268749 12288 268761 12291
rect 265897 12251 265955 12257
rect 266556 12260 268761 12288
rect 266556 12229 266584 12260
rect 268749 12257 268761 12260
rect 268795 12288 268807 12291
rect 269114 12288 269120 12300
rect 268795 12260 269120 12288
rect 268795 12257 268807 12260
rect 268749 12251 268807 12257
rect 269114 12248 269120 12260
rect 269172 12248 269178 12300
rect 269666 12248 269672 12300
rect 269724 12288 269730 12300
rect 271138 12288 271144 12300
rect 269724 12260 271144 12288
rect 269724 12248 269730 12260
rect 271138 12248 271144 12260
rect 271196 12248 271202 12300
rect 272242 12288 272248 12300
rect 272203 12260 272248 12288
rect 272242 12248 272248 12260
rect 272300 12288 272306 12300
rect 272794 12288 272800 12300
rect 272300 12260 272800 12288
rect 272300 12248 272306 12260
rect 272794 12248 272800 12260
rect 272852 12248 272858 12300
rect 266541 12223 266599 12229
rect 266541 12220 266553 12223
rect 264839 12192 265296 12220
rect 265360 12192 266553 12220
rect 264839 12189 264851 12192
rect 264793 12183 264851 12189
rect 265158 12152 265164 12164
rect 254058 12124 255084 12152
rect 255240 12124 256464 12152
rect 255056 12096 255084 12124
rect 231305 12087 231363 12093
rect 231305 12053 231317 12087
rect 231351 12053 231363 12087
rect 231305 12047 231363 12053
rect 231394 12044 231400 12096
rect 231452 12084 231458 12096
rect 231762 12084 231768 12096
rect 231452 12056 231768 12084
rect 231452 12044 231458 12056
rect 231762 12044 231768 12056
rect 231820 12044 231826 12096
rect 233050 12044 233056 12096
rect 233108 12084 233114 12096
rect 238205 12087 238263 12093
rect 238205 12084 238217 12087
rect 233108 12056 238217 12084
rect 233108 12044 233114 12056
rect 238205 12053 238217 12056
rect 238251 12053 238263 12087
rect 240870 12084 240876 12096
rect 240831 12056 240876 12084
rect 238205 12047 238263 12053
rect 240870 12044 240876 12056
rect 240928 12044 240934 12096
rect 241333 12087 241391 12093
rect 241333 12053 241345 12087
rect 241379 12084 241391 12087
rect 241514 12084 241520 12096
rect 241379 12056 241520 12084
rect 241379 12053 241391 12056
rect 241333 12047 241391 12053
rect 241514 12044 241520 12056
rect 241572 12084 241578 12096
rect 242526 12084 242532 12096
rect 241572 12056 242532 12084
rect 241572 12044 241578 12056
rect 242526 12044 242532 12056
rect 242584 12044 242590 12096
rect 242713 12087 242771 12093
rect 242713 12053 242725 12087
rect 242759 12084 242771 12087
rect 244090 12084 244096 12096
rect 242759 12056 244096 12084
rect 242759 12053 242771 12056
rect 242713 12047 242771 12053
rect 244090 12044 244096 12056
rect 244148 12044 244154 12096
rect 254394 12044 254400 12096
rect 254452 12084 254458 12096
rect 254765 12087 254823 12093
rect 254765 12084 254777 12087
rect 254452 12056 254777 12084
rect 254452 12044 254458 12056
rect 254765 12053 254777 12056
rect 254811 12053 254823 12087
rect 254765 12047 254823 12053
rect 255038 12044 255044 12096
rect 255096 12044 255102 12096
rect 255222 12044 255228 12096
rect 255280 12084 255286 12096
rect 256326 12084 256332 12096
rect 255280 12056 256332 12084
rect 255280 12044 255286 12056
rect 256326 12044 256332 12056
rect 256384 12044 256390 12096
rect 256436 12084 256464 12124
rect 263566 12124 265164 12152
rect 263566 12084 263594 12124
rect 265158 12112 265164 12124
rect 265216 12112 265222 12164
rect 265268 12093 265296 12192
rect 266541 12189 266553 12192
rect 266587 12189 266599 12223
rect 266541 12183 266599 12189
rect 268102 12180 268108 12232
rect 268160 12220 268166 12232
rect 268654 12220 268660 12232
rect 268160 12192 268660 12220
rect 268160 12180 268166 12192
rect 268654 12180 268660 12192
rect 268712 12180 268718 12232
rect 270957 12223 271015 12229
rect 270957 12220 270969 12223
rect 270328 12192 270969 12220
rect 265621 12155 265679 12161
rect 265621 12121 265633 12155
rect 265667 12152 265679 12155
rect 266814 12152 266820 12164
rect 265667 12124 266676 12152
rect 266775 12124 266820 12152
rect 265667 12121 265679 12124
rect 265621 12115 265679 12121
rect 256436 12056 263594 12084
rect 265253 12087 265311 12093
rect 265253 12053 265265 12087
rect 265299 12053 265311 12087
rect 266648 12084 266676 12124
rect 266814 12112 266820 12124
rect 266872 12112 266878 12164
rect 267274 12112 267280 12164
rect 267332 12112 267338 12164
rect 268194 12112 268200 12164
rect 268252 12152 268258 12164
rect 269025 12155 269083 12161
rect 269025 12152 269037 12155
rect 268252 12124 269037 12152
rect 268252 12112 268258 12124
rect 269025 12121 269037 12124
rect 269071 12121 269083 12155
rect 269025 12115 269083 12121
rect 269482 12112 269488 12164
rect 269540 12112 269546 12164
rect 266998 12084 267004 12096
rect 266648 12056 267004 12084
rect 265253 12047 265311 12053
rect 266998 12044 267004 12056
rect 267056 12044 267062 12096
rect 268289 12087 268347 12093
rect 268289 12053 268301 12087
rect 268335 12084 268347 12087
rect 268470 12084 268476 12096
rect 268335 12056 268476 12084
rect 268335 12053 268347 12056
rect 268289 12047 268347 12053
rect 268470 12044 268476 12056
rect 268528 12044 268534 12096
rect 268654 12044 268660 12096
rect 268712 12084 268718 12096
rect 270328 12084 270356 12192
rect 270957 12189 270969 12192
rect 271003 12220 271015 12223
rect 271322 12220 271328 12232
rect 271003 12192 271328 12220
rect 271003 12189 271015 12192
rect 270957 12183 271015 12189
rect 271322 12180 271328 12192
rect 271380 12180 271386 12232
rect 272061 12223 272119 12229
rect 272061 12189 272073 12223
rect 272107 12220 272119 12223
rect 272886 12220 272892 12232
rect 272107 12192 272892 12220
rect 272107 12189 272119 12192
rect 272061 12183 272119 12189
rect 272886 12180 272892 12192
rect 272944 12180 272950 12232
rect 270512 12124 272196 12152
rect 268712 12056 270356 12084
rect 268712 12044 268718 12056
rect 270402 12044 270408 12096
rect 270460 12084 270466 12096
rect 270512 12093 270540 12124
rect 272168 12093 272196 12124
rect 270497 12087 270555 12093
rect 270497 12084 270509 12087
rect 270460 12056 270509 12084
rect 270460 12044 270466 12056
rect 270497 12053 270509 12056
rect 270543 12053 270555 12087
rect 270497 12047 270555 12053
rect 272153 12087 272211 12093
rect 272153 12053 272165 12087
rect 272199 12084 272211 12087
rect 284754 12084 284760 12096
rect 272199 12056 284760 12084
rect 272199 12053 272211 12056
rect 272153 12047 272211 12053
rect 284754 12044 284760 12056
rect 284812 12044 284818 12096
rect 1104 11994 305808 12016
rect 1104 11942 77148 11994
rect 77200 11942 77212 11994
rect 77264 11942 77276 11994
rect 77328 11942 77340 11994
rect 77392 11942 77404 11994
rect 77456 11942 153346 11994
rect 153398 11942 153410 11994
rect 153462 11942 153474 11994
rect 153526 11942 153538 11994
rect 153590 11942 153602 11994
rect 153654 11942 229544 11994
rect 229596 11942 229608 11994
rect 229660 11942 229672 11994
rect 229724 11942 229736 11994
rect 229788 11942 229800 11994
rect 229852 11942 305808 11994
rect 1104 11920 305808 11942
rect 27801 11883 27859 11889
rect 27801 11849 27813 11883
rect 27847 11880 27859 11883
rect 29086 11880 29092 11892
rect 27847 11852 29092 11880
rect 27847 11849 27859 11852
rect 27801 11843 27859 11849
rect 29086 11840 29092 11852
rect 29144 11840 29150 11892
rect 29454 11840 29460 11892
rect 29512 11880 29518 11892
rect 30926 11880 30932 11892
rect 29512 11852 30932 11880
rect 29512 11840 29518 11852
rect 30926 11840 30932 11852
rect 30984 11840 30990 11892
rect 32214 11840 32220 11892
rect 32272 11880 32278 11892
rect 32585 11883 32643 11889
rect 32585 11880 32597 11883
rect 32272 11852 32597 11880
rect 32272 11840 32278 11852
rect 32585 11849 32597 11852
rect 32631 11849 32643 11883
rect 33778 11880 33784 11892
rect 33739 11852 33784 11880
rect 32585 11843 32643 11849
rect 33778 11840 33784 11852
rect 33836 11840 33842 11892
rect 34422 11880 34428 11892
rect 34383 11852 34428 11880
rect 34422 11840 34428 11852
rect 34480 11840 34486 11892
rect 34977 11883 35035 11889
rect 34977 11849 34989 11883
rect 35023 11849 35035 11883
rect 38378 11880 38384 11892
rect 38339 11852 38384 11880
rect 34977 11843 35035 11849
rect 27706 11772 27712 11824
rect 27764 11812 27770 11824
rect 27764 11784 28120 11812
rect 27764 11772 27770 11784
rect 27985 11747 28043 11753
rect 27985 11713 27997 11747
rect 28031 11713 28043 11747
rect 27985 11707 28043 11713
rect 28000 11608 28028 11707
rect 28092 11676 28120 11784
rect 28718 11772 28724 11824
rect 28776 11812 28782 11824
rect 28813 11815 28871 11821
rect 28813 11812 28825 11815
rect 28776 11784 28825 11812
rect 28776 11772 28782 11784
rect 28813 11781 28825 11784
rect 28859 11781 28871 11815
rect 28813 11775 28871 11781
rect 28994 11772 29000 11824
rect 29052 11812 29058 11824
rect 30006 11812 30012 11824
rect 29052 11784 30012 11812
rect 29052 11772 29058 11784
rect 28902 11676 28908 11688
rect 28092 11648 28908 11676
rect 28902 11636 28908 11648
rect 28960 11636 28966 11688
rect 29104 11685 29132 11784
rect 30006 11772 30012 11784
rect 30064 11772 30070 11824
rect 32030 11772 32036 11824
rect 32088 11812 32094 11824
rect 34992 11812 35020 11843
rect 38378 11840 38384 11852
rect 38436 11840 38442 11892
rect 39025 11883 39083 11889
rect 39025 11849 39037 11883
rect 39071 11880 39083 11883
rect 39574 11880 39580 11892
rect 39071 11852 39580 11880
rect 39071 11849 39083 11852
rect 39025 11843 39083 11849
rect 39574 11840 39580 11852
rect 39632 11840 39638 11892
rect 39669 11883 39727 11889
rect 39669 11849 39681 11883
rect 39715 11849 39727 11883
rect 39669 11843 39727 11849
rect 32088 11784 35020 11812
rect 32088 11772 32094 11784
rect 29546 11704 29552 11756
rect 29604 11744 29610 11756
rect 29641 11747 29699 11753
rect 29641 11744 29653 11747
rect 29604 11716 29653 11744
rect 29604 11704 29610 11716
rect 29641 11713 29653 11716
rect 29687 11713 29699 11747
rect 32398 11744 32404 11756
rect 31050 11716 32404 11744
rect 29641 11707 29699 11713
rect 32398 11704 32404 11716
rect 32456 11704 32462 11756
rect 32493 11747 32551 11753
rect 32493 11713 32505 11747
rect 32539 11744 32551 11747
rect 33689 11747 33747 11753
rect 32539 11716 32812 11744
rect 32539 11713 32551 11716
rect 32493 11707 32551 11713
rect 29089 11679 29147 11685
rect 29089 11645 29101 11679
rect 29135 11645 29147 11679
rect 29914 11676 29920 11688
rect 29875 11648 29920 11676
rect 29089 11639 29147 11645
rect 29914 11636 29920 11648
rect 29972 11636 29978 11688
rect 32508 11676 32536 11707
rect 30944 11648 32536 11676
rect 28000 11580 29776 11608
rect 28442 11540 28448 11552
rect 28403 11512 28448 11540
rect 28442 11500 28448 11512
rect 28500 11500 28506 11552
rect 29748 11540 29776 11580
rect 30944 11540 30972 11648
rect 32582 11636 32588 11688
rect 32640 11676 32646 11688
rect 32677 11679 32735 11685
rect 32677 11676 32689 11679
rect 32640 11648 32689 11676
rect 32640 11636 32646 11648
rect 32677 11645 32689 11648
rect 32723 11645 32735 11679
rect 32784 11676 32812 11716
rect 33689 11713 33701 11747
rect 33735 11744 33747 11747
rect 34333 11747 34391 11753
rect 34333 11744 34345 11747
rect 33735 11716 34345 11744
rect 33735 11713 33747 11716
rect 33689 11707 33747 11713
rect 34333 11713 34345 11716
rect 34379 11744 34391 11747
rect 34698 11744 34704 11756
rect 34379 11716 34704 11744
rect 34379 11713 34391 11716
rect 34333 11707 34391 11713
rect 34698 11704 34704 11716
rect 34756 11704 34762 11756
rect 35161 11747 35219 11753
rect 35161 11713 35173 11747
rect 35207 11713 35219 11747
rect 35161 11707 35219 11713
rect 38565 11747 38623 11753
rect 38565 11713 38577 11747
rect 38611 11713 38623 11747
rect 38565 11707 38623 11713
rect 39209 11747 39267 11753
rect 39209 11713 39221 11747
rect 39255 11744 39267 11747
rect 39684 11744 39712 11843
rect 39942 11840 39948 11892
rect 40000 11880 40006 11892
rect 40129 11883 40187 11889
rect 40129 11880 40141 11883
rect 40000 11852 40141 11880
rect 40000 11840 40006 11852
rect 40129 11849 40141 11852
rect 40175 11849 40187 11883
rect 40129 11843 40187 11849
rect 41141 11883 41199 11889
rect 41141 11849 41153 11883
rect 41187 11880 41199 11883
rect 41414 11880 41420 11892
rect 41187 11852 41420 11880
rect 41187 11849 41199 11852
rect 41141 11843 41199 11849
rect 41414 11840 41420 11852
rect 41472 11840 41478 11892
rect 41693 11883 41751 11889
rect 41693 11849 41705 11883
rect 41739 11880 41751 11883
rect 42886 11880 42892 11892
rect 41739 11852 42892 11880
rect 41739 11849 41751 11852
rect 41693 11843 41751 11849
rect 42886 11840 42892 11852
rect 42944 11840 42950 11892
rect 52638 11840 52644 11892
rect 52696 11880 52702 11892
rect 52825 11883 52883 11889
rect 52825 11880 52837 11883
rect 52696 11852 52837 11880
rect 52696 11840 52702 11852
rect 52825 11849 52837 11852
rect 52871 11849 52883 11883
rect 53650 11880 53656 11892
rect 53611 11852 53656 11880
rect 52825 11843 52883 11849
rect 53650 11840 53656 11852
rect 53708 11840 53714 11892
rect 54386 11880 54392 11892
rect 54347 11852 54392 11880
rect 54386 11840 54392 11852
rect 54444 11840 54450 11892
rect 55306 11880 55312 11892
rect 55267 11852 55312 11880
rect 55306 11840 55312 11852
rect 55364 11840 55370 11892
rect 56505 11883 56563 11889
rect 56505 11849 56517 11883
rect 56551 11880 56563 11883
rect 56594 11880 56600 11892
rect 56551 11852 56600 11880
rect 56551 11849 56563 11852
rect 56505 11843 56563 11849
rect 56594 11840 56600 11852
rect 56652 11840 56658 11892
rect 57149 11883 57207 11889
rect 57149 11849 57161 11883
rect 57195 11880 57207 11883
rect 58618 11880 58624 11892
rect 57195 11852 58624 11880
rect 57195 11849 57207 11852
rect 57149 11843 57207 11849
rect 58618 11840 58624 11852
rect 58676 11840 58682 11892
rect 75454 11840 75460 11892
rect 75512 11880 75518 11892
rect 75549 11883 75607 11889
rect 75549 11880 75561 11883
rect 75512 11852 75561 11880
rect 75512 11840 75518 11852
rect 75549 11849 75561 11852
rect 75595 11849 75607 11883
rect 75549 11843 75607 11849
rect 75638 11840 75644 11892
rect 75696 11880 75702 11892
rect 76009 11883 76067 11889
rect 76009 11880 76021 11883
rect 75696 11852 76021 11880
rect 75696 11840 75702 11852
rect 76009 11849 76021 11852
rect 76055 11849 76067 11883
rect 76009 11843 76067 11849
rect 76466 11840 76472 11892
rect 76524 11880 76530 11892
rect 76929 11883 76987 11889
rect 76929 11880 76941 11883
rect 76524 11852 76941 11880
rect 76524 11840 76530 11852
rect 76929 11849 76941 11852
rect 76975 11849 76987 11883
rect 77846 11880 77852 11892
rect 77807 11852 77852 11880
rect 76929 11843 76987 11849
rect 77846 11840 77852 11852
rect 77904 11840 77910 11892
rect 78490 11880 78496 11892
rect 78451 11852 78496 11880
rect 78490 11840 78496 11852
rect 78548 11840 78554 11892
rect 84286 11840 84292 11892
rect 84344 11880 84350 11892
rect 84381 11883 84439 11889
rect 84381 11880 84393 11883
rect 84344 11852 84393 11880
rect 84344 11840 84350 11852
rect 84381 11849 84393 11852
rect 84427 11849 84439 11883
rect 86034 11880 86040 11892
rect 84381 11843 84439 11849
rect 85040 11852 86040 11880
rect 40037 11815 40095 11821
rect 40037 11781 40049 11815
rect 40083 11812 40095 11815
rect 40678 11812 40684 11824
rect 40083 11784 40684 11812
rect 40083 11781 40095 11784
rect 40037 11775 40095 11781
rect 39255 11716 39712 11744
rect 39255 11713 39267 11716
rect 39209 11707 39267 11713
rect 34054 11676 34060 11688
rect 32784 11648 34060 11676
rect 32677 11639 32735 11645
rect 34054 11636 34060 11648
rect 34112 11636 34118 11688
rect 31110 11568 31116 11620
rect 31168 11608 31174 11620
rect 35176 11608 35204 11707
rect 38580 11676 38608 11707
rect 40052 11676 40080 11775
rect 40678 11772 40684 11784
rect 40736 11812 40742 11824
rect 41230 11812 41236 11824
rect 40736 11784 41236 11812
rect 40736 11772 40742 11784
rect 41230 11772 41236 11784
rect 41288 11772 41294 11824
rect 53742 11772 53748 11824
rect 53800 11812 53806 11824
rect 53800 11784 56456 11812
rect 53800 11772 53806 11784
rect 40310 11704 40316 11756
rect 40368 11744 40374 11756
rect 41049 11747 41107 11753
rect 41049 11744 41061 11747
rect 40368 11716 41061 11744
rect 40368 11704 40374 11716
rect 41049 11713 41061 11716
rect 41095 11744 41107 11747
rect 41877 11747 41935 11753
rect 41095 11716 41414 11744
rect 41095 11713 41107 11716
rect 41049 11707 41107 11713
rect 41386 11688 41414 11716
rect 41877 11713 41889 11747
rect 41923 11744 41935 11747
rect 42794 11744 42800 11756
rect 41923 11716 42800 11744
rect 41923 11713 41935 11716
rect 41877 11707 41935 11713
rect 42794 11704 42800 11716
rect 42852 11704 42858 11756
rect 42889 11747 42947 11753
rect 42889 11713 42901 11747
rect 42935 11744 42947 11747
rect 42978 11744 42984 11756
rect 42935 11716 42984 11744
rect 42935 11713 42947 11716
rect 42889 11707 42947 11713
rect 42978 11704 42984 11716
rect 43036 11744 43042 11756
rect 53006 11744 53012 11756
rect 43036 11716 43484 11744
rect 52967 11716 53012 11744
rect 43036 11704 43042 11716
rect 38580 11648 40080 11676
rect 40221 11679 40279 11685
rect 40221 11645 40233 11679
rect 40267 11676 40279 11679
rect 40954 11676 40960 11688
rect 40267 11648 40960 11676
rect 40267 11645 40279 11648
rect 40221 11639 40279 11645
rect 40954 11636 40960 11648
rect 41012 11636 41018 11688
rect 41386 11648 41420 11688
rect 41414 11636 41420 11648
rect 41472 11676 41478 11688
rect 43073 11679 43131 11685
rect 43073 11676 43085 11679
rect 41472 11648 43085 11676
rect 41472 11636 41478 11648
rect 43073 11645 43085 11648
rect 43119 11645 43131 11679
rect 43073 11639 43131 11645
rect 43456 11617 43484 11716
rect 53006 11704 53012 11716
rect 53064 11704 53070 11756
rect 54312 11753 54340 11784
rect 56428 11753 56456 11784
rect 57422 11772 57428 11824
rect 57480 11812 57486 11824
rect 84930 11812 84936 11824
rect 57480 11784 84936 11812
rect 57480 11772 57486 11784
rect 84930 11772 84936 11784
rect 84988 11772 84994 11824
rect 53837 11747 53895 11753
rect 53837 11713 53849 11747
rect 53883 11713 53895 11747
rect 53837 11707 53895 11713
rect 54297 11747 54355 11753
rect 54297 11713 54309 11747
rect 54343 11713 54355 11747
rect 54297 11707 54355 11713
rect 56413 11747 56471 11753
rect 56413 11713 56425 11747
rect 56459 11744 56471 11747
rect 57057 11747 57115 11753
rect 57057 11744 57069 11747
rect 56459 11716 57069 11744
rect 56459 11713 56471 11716
rect 56413 11707 56471 11713
rect 57057 11713 57069 11716
rect 57103 11713 57115 11747
rect 57057 11707 57115 11713
rect 53852 11676 53880 11707
rect 54662 11676 54668 11688
rect 53852 11648 54668 11676
rect 54662 11636 54668 11648
rect 54720 11676 54726 11688
rect 55401 11679 55459 11685
rect 55401 11676 55413 11679
rect 54720 11648 55413 11676
rect 54720 11636 54726 11648
rect 55401 11645 55413 11648
rect 55447 11645 55459 11679
rect 55582 11676 55588 11688
rect 55543 11648 55588 11676
rect 55401 11639 55459 11645
rect 55582 11636 55588 11648
rect 55640 11636 55646 11688
rect 55858 11636 55864 11688
rect 55916 11676 55922 11688
rect 57440 11676 57468 11772
rect 75917 11747 75975 11753
rect 75917 11713 75929 11747
rect 75963 11744 75975 11747
rect 76006 11744 76012 11756
rect 75963 11716 76012 11744
rect 75963 11713 75975 11716
rect 75917 11707 75975 11713
rect 76006 11704 76012 11716
rect 76064 11704 76070 11756
rect 76282 11704 76288 11756
rect 76340 11744 76346 11756
rect 77113 11747 77171 11753
rect 77113 11744 77125 11747
rect 76340 11716 77125 11744
rect 76340 11704 76346 11716
rect 77113 11713 77125 11716
rect 77159 11713 77171 11747
rect 77113 11707 77171 11713
rect 77757 11747 77815 11753
rect 77757 11713 77769 11747
rect 77803 11744 77815 11747
rect 78582 11744 78588 11756
rect 77803 11716 78588 11744
rect 77803 11713 77815 11716
rect 77757 11707 77815 11713
rect 78582 11704 78588 11716
rect 78640 11704 78646 11756
rect 78677 11747 78735 11753
rect 78677 11713 78689 11747
rect 78723 11744 78735 11747
rect 81434 11744 81440 11756
rect 78723 11716 81440 11744
rect 78723 11713 78735 11716
rect 78677 11707 78735 11713
rect 81434 11704 81440 11716
rect 81492 11704 81498 11756
rect 84565 11747 84623 11753
rect 84565 11713 84577 11747
rect 84611 11744 84623 11747
rect 85040 11744 85068 11852
rect 86034 11840 86040 11852
rect 86092 11840 86098 11892
rect 86126 11840 86132 11892
rect 86184 11880 86190 11892
rect 87141 11883 87199 11889
rect 87141 11880 87153 11883
rect 86184 11852 87153 11880
rect 86184 11840 86190 11852
rect 87141 11849 87153 11852
rect 87187 11849 87199 11883
rect 87874 11880 87880 11892
rect 87835 11852 87880 11880
rect 87141 11843 87199 11849
rect 87874 11840 87880 11852
rect 87932 11840 87938 11892
rect 88889 11883 88947 11889
rect 88889 11849 88901 11883
rect 88935 11880 88947 11883
rect 89530 11880 89536 11892
rect 88935 11852 89536 11880
rect 88935 11849 88947 11852
rect 88889 11843 88947 11849
rect 89530 11840 89536 11852
rect 89588 11840 89594 11892
rect 99650 11840 99656 11892
rect 99708 11880 99714 11892
rect 100205 11883 100263 11889
rect 100205 11880 100217 11883
rect 99708 11852 100217 11880
rect 99708 11840 99714 11852
rect 100205 11849 100217 11852
rect 100251 11849 100263 11883
rect 100938 11880 100944 11892
rect 100899 11852 100944 11880
rect 100205 11843 100263 11849
rect 100938 11840 100944 11852
rect 100996 11840 101002 11892
rect 101861 11883 101919 11889
rect 101861 11849 101873 11883
rect 101907 11880 101919 11883
rect 103054 11880 103060 11892
rect 101907 11852 103060 11880
rect 101907 11849 101919 11852
rect 101861 11843 101919 11849
rect 103054 11840 103060 11852
rect 103112 11840 103118 11892
rect 103514 11840 103520 11892
rect 103572 11880 103578 11892
rect 113818 11880 113824 11892
rect 103572 11852 113174 11880
rect 113779 11852 113824 11880
rect 103572 11840 103578 11852
rect 85298 11772 85304 11824
rect 85356 11812 85362 11824
rect 113146 11812 113174 11852
rect 113818 11840 113824 11852
rect 113876 11840 113882 11892
rect 114278 11840 114284 11892
rect 114336 11880 114342 11892
rect 115017 11883 115075 11889
rect 115017 11880 115029 11883
rect 114336 11852 115029 11880
rect 114336 11840 114342 11852
rect 115017 11849 115029 11852
rect 115063 11880 115075 11883
rect 115658 11880 115664 11892
rect 115063 11852 115664 11880
rect 115063 11849 115075 11852
rect 115017 11843 115075 11849
rect 115658 11840 115664 11852
rect 115716 11840 115722 11892
rect 116213 11883 116271 11889
rect 116213 11849 116225 11883
rect 116259 11880 116271 11883
rect 116762 11880 116768 11892
rect 116259 11852 116768 11880
rect 116259 11849 116271 11852
rect 116213 11843 116271 11849
rect 116762 11840 116768 11852
rect 116820 11840 116826 11892
rect 116949 11883 117007 11889
rect 116949 11849 116961 11883
rect 116995 11880 117007 11883
rect 117314 11880 117320 11892
rect 116995 11852 117320 11880
rect 116995 11849 117007 11852
rect 116949 11843 117007 11849
rect 117314 11840 117320 11852
rect 117372 11840 117378 11892
rect 117593 11883 117651 11889
rect 117593 11849 117605 11883
rect 117639 11880 117651 11883
rect 118786 11880 118792 11892
rect 117639 11852 118792 11880
rect 117639 11849 117651 11852
rect 117593 11843 117651 11849
rect 118786 11840 118792 11852
rect 118844 11840 118850 11892
rect 129366 11880 129372 11892
rect 129327 11852 129372 11880
rect 129366 11840 129372 11852
rect 129424 11840 129430 11892
rect 130286 11840 130292 11892
rect 130344 11880 130350 11892
rect 130473 11883 130531 11889
rect 130473 11880 130485 11883
rect 130344 11852 130485 11880
rect 130344 11840 130350 11852
rect 130473 11849 130485 11852
rect 130519 11849 130531 11883
rect 130930 11880 130936 11892
rect 130891 11852 130936 11880
rect 130473 11843 130531 11849
rect 130930 11840 130936 11852
rect 130988 11840 130994 11892
rect 131114 11840 131120 11892
rect 131172 11880 131178 11892
rect 132405 11883 132463 11889
rect 132405 11880 132417 11883
rect 131172 11852 132417 11880
rect 131172 11840 131178 11852
rect 132405 11849 132417 11852
rect 132451 11849 132463 11883
rect 132405 11843 132463 11849
rect 137738 11840 137744 11892
rect 137796 11880 137802 11892
rect 151078 11880 151084 11892
rect 137796 11852 150940 11880
rect 151039 11852 151084 11880
rect 137796 11840 137802 11852
rect 114554 11812 114560 11824
rect 85356 11784 108252 11812
rect 113146 11784 114560 11812
rect 85356 11772 85362 11784
rect 84611 11716 85068 11744
rect 85209 11747 85267 11753
rect 84611 11713 84623 11716
rect 84565 11707 84623 11713
rect 85209 11713 85221 11747
rect 85255 11713 85267 11747
rect 85209 11707 85267 11713
rect 55916 11648 57468 11676
rect 55916 11636 55922 11648
rect 74994 11636 75000 11688
rect 75052 11676 75058 11688
rect 76193 11679 76251 11685
rect 76193 11676 76205 11679
rect 75052 11648 76205 11676
rect 75052 11636 75058 11648
rect 76193 11645 76205 11648
rect 76239 11676 76251 11679
rect 76926 11676 76932 11688
rect 76239 11648 76932 11676
rect 76239 11645 76251 11648
rect 76193 11639 76251 11645
rect 76926 11636 76932 11648
rect 76984 11636 76990 11688
rect 84010 11636 84016 11688
rect 84068 11676 84074 11688
rect 85224 11676 85252 11707
rect 85758 11704 85764 11756
rect 85816 11744 85822 11756
rect 86129 11747 86187 11753
rect 86129 11744 86141 11747
rect 85816 11716 86141 11744
rect 85816 11704 85822 11716
rect 86129 11713 86141 11716
rect 86175 11713 86187 11747
rect 86129 11707 86187 11713
rect 86954 11704 86960 11756
rect 87012 11744 87018 11756
rect 87785 11747 87843 11753
rect 87012 11716 87057 11744
rect 87012 11704 87018 11716
rect 87785 11713 87797 11747
rect 87831 11744 87843 11747
rect 88797 11747 88855 11753
rect 87831 11716 87920 11744
rect 87831 11713 87843 11716
rect 87785 11707 87843 11713
rect 86310 11676 86316 11688
rect 84068 11648 85252 11676
rect 86271 11648 86316 11676
rect 84068 11636 84074 11648
rect 86310 11636 86316 11648
rect 86368 11636 86374 11688
rect 87892 11676 87920 11716
rect 88797 11713 88809 11747
rect 88843 11744 88855 11747
rect 89162 11744 89168 11756
rect 88843 11716 89168 11744
rect 88843 11713 88855 11716
rect 88797 11707 88855 11713
rect 89162 11704 89168 11716
rect 89220 11704 89226 11756
rect 100386 11744 100392 11756
rect 100347 11716 100392 11744
rect 100386 11704 100392 11716
rect 100444 11704 100450 11756
rect 100849 11747 100907 11753
rect 100849 11713 100861 11747
rect 100895 11744 100907 11747
rect 102134 11744 102140 11756
rect 100895 11716 102140 11744
rect 100895 11713 100907 11716
rect 100849 11707 100907 11713
rect 102134 11704 102140 11716
rect 102192 11704 102198 11756
rect 103149 11747 103207 11753
rect 103149 11713 103161 11747
rect 103195 11744 103207 11747
rect 103606 11744 103612 11756
rect 103195 11716 103612 11744
rect 103195 11713 103207 11716
rect 103149 11707 103207 11713
rect 103606 11704 103612 11716
rect 103664 11704 103670 11756
rect 90450 11676 90456 11688
rect 86420 11648 86954 11676
rect 87892 11648 90456 11676
rect 31168 11580 35204 11608
rect 43441 11611 43499 11617
rect 31168 11568 31174 11580
rect 43441 11577 43453 11611
rect 43487 11608 43499 11611
rect 56042 11608 56048 11620
rect 43487 11580 56048 11608
rect 43487 11577 43499 11580
rect 43441 11571 43499 11577
rect 56042 11568 56048 11580
rect 56100 11608 56106 11620
rect 86420 11608 86448 11648
rect 56100 11580 86448 11608
rect 86926 11608 86954 11648
rect 90450 11636 90456 11648
rect 90508 11636 90514 11688
rect 100754 11636 100760 11688
rect 100812 11676 100818 11688
rect 101953 11679 102011 11685
rect 101953 11676 101965 11679
rect 100812 11648 101965 11676
rect 100812 11636 100818 11648
rect 101953 11645 101965 11648
rect 101999 11645 102011 11679
rect 101953 11639 102011 11645
rect 102042 11636 102048 11688
rect 102100 11676 102106 11688
rect 102100 11648 102145 11676
rect 102100 11636 102106 11648
rect 102318 11636 102324 11688
rect 102376 11676 102382 11688
rect 103514 11676 103520 11688
rect 102376 11648 103520 11676
rect 102376 11636 102382 11648
rect 103514 11636 103520 11648
rect 103572 11636 103578 11688
rect 108224 11676 108252 11784
rect 114554 11772 114560 11784
rect 114612 11772 114618 11824
rect 138014 11812 138020 11824
rect 114940 11784 138020 11812
rect 114002 11744 114008 11756
rect 113963 11716 114008 11744
rect 114002 11704 114008 11716
rect 114060 11704 114066 11756
rect 114940 11676 114968 11784
rect 138014 11772 138020 11784
rect 138072 11772 138078 11824
rect 149974 11812 149980 11824
rect 149822 11784 149980 11812
rect 149974 11772 149980 11784
rect 150032 11772 150038 11824
rect 150912 11812 150940 11852
rect 151078 11840 151084 11852
rect 151136 11840 151142 11892
rect 151998 11880 152004 11892
rect 151959 11852 152004 11880
rect 151998 11840 152004 11852
rect 152056 11840 152062 11892
rect 152737 11883 152795 11889
rect 152737 11849 152749 11883
rect 152783 11880 152795 11883
rect 154206 11880 154212 11892
rect 152783 11852 154212 11880
rect 152783 11849 152795 11852
rect 152737 11843 152795 11849
rect 154206 11840 154212 11852
rect 154264 11840 154270 11892
rect 157306 11852 161980 11880
rect 157306 11812 157334 11852
rect 150912 11784 157334 11812
rect 115014 11704 115020 11756
rect 115072 11744 115078 11756
rect 115109 11747 115167 11753
rect 115109 11744 115121 11747
rect 115072 11716 115121 11744
rect 115072 11704 115078 11716
rect 115109 11713 115121 11716
rect 115155 11713 115167 11747
rect 116394 11744 116400 11756
rect 116355 11716 116400 11744
rect 115109 11707 115167 11713
rect 116394 11704 116400 11716
rect 116452 11704 116458 11756
rect 116857 11747 116915 11753
rect 116857 11713 116869 11747
rect 116903 11744 116915 11747
rect 117501 11747 117559 11753
rect 117501 11744 117513 11747
rect 116903 11716 117513 11744
rect 116903 11713 116915 11716
rect 116857 11707 116915 11713
rect 117501 11713 117513 11716
rect 117547 11744 117559 11747
rect 118326 11744 118332 11756
rect 117547 11716 118332 11744
rect 117547 11713 117559 11716
rect 117501 11707 117559 11713
rect 108224 11648 114968 11676
rect 115293 11679 115351 11685
rect 115293 11645 115305 11679
rect 115339 11676 115351 11679
rect 115658 11676 115664 11688
rect 115339 11648 115664 11676
rect 115339 11645 115351 11648
rect 115293 11639 115351 11645
rect 115658 11636 115664 11648
rect 115716 11636 115722 11688
rect 115750 11636 115756 11688
rect 115808 11676 115814 11688
rect 116872 11676 116900 11707
rect 118326 11704 118332 11716
rect 118384 11704 118390 11756
rect 128354 11704 128360 11756
rect 128412 11744 128418 11756
rect 129277 11747 129335 11753
rect 129277 11744 129289 11747
rect 128412 11716 129289 11744
rect 128412 11704 128418 11716
rect 129277 11713 129289 11716
rect 129323 11744 129335 11747
rect 130286 11744 130292 11756
rect 129323 11716 130292 11744
rect 129323 11713 129335 11716
rect 129277 11707 129335 11713
rect 130286 11704 130292 11716
rect 130344 11704 130350 11756
rect 130841 11747 130899 11753
rect 130841 11713 130853 11747
rect 130887 11744 130899 11747
rect 131574 11744 131580 11756
rect 130887 11716 131580 11744
rect 130887 11713 130899 11716
rect 130841 11707 130899 11713
rect 131574 11704 131580 11716
rect 131632 11704 131638 11756
rect 131669 11747 131727 11753
rect 131669 11713 131681 11747
rect 131715 11713 131727 11747
rect 131669 11707 131727 11713
rect 115808 11648 116900 11676
rect 115808 11636 115814 11648
rect 129734 11636 129740 11688
rect 129792 11676 129798 11688
rect 131022 11676 131028 11688
rect 129792 11648 131028 11676
rect 129792 11636 129798 11648
rect 131022 11636 131028 11648
rect 131080 11636 131086 11688
rect 131684 11676 131712 11707
rect 132494 11704 132500 11756
rect 132552 11744 132558 11756
rect 132589 11747 132647 11753
rect 132589 11744 132601 11747
rect 132552 11716 132601 11744
rect 132552 11704 132558 11716
rect 132589 11713 132601 11716
rect 132635 11713 132647 11747
rect 132589 11707 132647 11713
rect 147674 11704 147680 11756
rect 147732 11744 147738 11756
rect 147769 11747 147827 11753
rect 147769 11744 147781 11747
rect 147732 11716 147781 11744
rect 147732 11704 147738 11716
rect 147769 11713 147781 11716
rect 147815 11713 147827 11747
rect 151262 11744 151268 11756
rect 151223 11716 151268 11744
rect 147769 11707 147827 11713
rect 151262 11704 151268 11716
rect 151320 11704 151326 11756
rect 152182 11744 152188 11756
rect 152143 11716 152188 11744
rect 152182 11704 152188 11716
rect 152240 11704 152246 11756
rect 152645 11747 152703 11753
rect 152645 11713 152657 11747
rect 152691 11744 152703 11747
rect 152734 11744 152740 11756
rect 152691 11716 152740 11744
rect 152691 11713 152703 11716
rect 152645 11707 152703 11713
rect 152734 11704 152740 11716
rect 152792 11704 152798 11756
rect 161106 11744 161112 11756
rect 161067 11716 161112 11744
rect 161106 11704 161112 11716
rect 161164 11704 161170 11756
rect 161750 11744 161756 11756
rect 161711 11716 161756 11744
rect 161750 11704 161756 11716
rect 161808 11704 161814 11756
rect 137738 11676 137744 11688
rect 131684 11648 137744 11676
rect 137738 11636 137744 11648
rect 137796 11636 137802 11688
rect 148318 11676 148324 11688
rect 148279 11648 148324 11676
rect 148318 11636 148324 11648
rect 148376 11636 148382 11688
rect 148594 11676 148600 11688
rect 148555 11648 148600 11676
rect 148594 11636 148600 11648
rect 148652 11636 148658 11688
rect 143258 11608 143264 11620
rect 86926 11580 143264 11608
rect 56100 11568 56106 11580
rect 143258 11568 143264 11580
rect 143316 11568 143322 11620
rect 146018 11568 146024 11620
rect 146076 11608 146082 11620
rect 147585 11611 147643 11617
rect 147585 11608 147597 11611
rect 146076 11580 147597 11608
rect 146076 11568 146082 11580
rect 147585 11577 147597 11580
rect 147631 11577 147643 11611
rect 147585 11571 147643 11577
rect 160925 11611 160983 11617
rect 160925 11577 160937 11611
rect 160971 11608 160983 11611
rect 161198 11608 161204 11620
rect 160971 11580 161204 11608
rect 160971 11577 160983 11580
rect 160925 11571 160983 11577
rect 161198 11568 161204 11580
rect 161256 11568 161262 11620
rect 161290 11568 161296 11620
rect 161348 11608 161354 11620
rect 161569 11611 161627 11617
rect 161569 11608 161581 11611
rect 161348 11580 161581 11608
rect 161348 11568 161354 11580
rect 161569 11577 161581 11580
rect 161615 11577 161627 11611
rect 161952 11608 161980 11852
rect 162026 11840 162032 11892
rect 162084 11880 162090 11892
rect 162305 11883 162363 11889
rect 162305 11880 162317 11883
rect 162084 11852 162317 11880
rect 162084 11840 162090 11852
rect 162305 11849 162317 11852
rect 162351 11849 162363 11883
rect 162305 11843 162363 11849
rect 162762 11840 162768 11892
rect 162820 11880 162826 11892
rect 162949 11883 163007 11889
rect 162949 11880 162961 11883
rect 162820 11852 162961 11880
rect 162820 11840 162826 11852
rect 162949 11849 162961 11852
rect 162995 11849 163007 11883
rect 162949 11843 163007 11849
rect 163501 11883 163559 11889
rect 163501 11849 163513 11883
rect 163547 11880 163559 11883
rect 163774 11880 163780 11892
rect 163547 11852 163780 11880
rect 163547 11849 163559 11852
rect 163501 11843 163559 11849
rect 163774 11840 163780 11852
rect 163832 11840 163838 11892
rect 164237 11883 164295 11889
rect 164237 11849 164249 11883
rect 164283 11880 164295 11883
rect 164326 11880 164332 11892
rect 164283 11852 164332 11880
rect 164283 11849 164295 11852
rect 164237 11843 164295 11849
rect 164326 11840 164332 11852
rect 164384 11840 164390 11892
rect 164878 11880 164884 11892
rect 164839 11852 164884 11880
rect 164878 11840 164884 11852
rect 164936 11840 164942 11892
rect 176473 11883 176531 11889
rect 176473 11849 176485 11883
rect 176519 11880 176531 11883
rect 176746 11880 176752 11892
rect 176519 11852 176752 11880
rect 176519 11849 176531 11852
rect 176473 11843 176531 11849
rect 176746 11840 176752 11852
rect 176804 11840 176810 11892
rect 177390 11840 177396 11892
rect 177448 11880 177454 11892
rect 177577 11883 177635 11889
rect 177577 11880 177589 11883
rect 177448 11852 177589 11880
rect 177448 11840 177454 11852
rect 177577 11849 177589 11852
rect 177623 11849 177635 11883
rect 177577 11843 177635 11849
rect 177850 11840 177856 11892
rect 177908 11880 177914 11892
rect 178037 11883 178095 11889
rect 178037 11880 178049 11883
rect 177908 11852 178049 11880
rect 177908 11840 177914 11852
rect 178037 11849 178049 11852
rect 178083 11849 178095 11883
rect 178037 11843 178095 11849
rect 179141 11883 179199 11889
rect 179141 11849 179153 11883
rect 179187 11880 179199 11883
rect 179874 11880 179880 11892
rect 179187 11852 179880 11880
rect 179187 11849 179199 11852
rect 179141 11843 179199 11849
rect 179874 11840 179880 11852
rect 179932 11840 179938 11892
rect 179966 11840 179972 11892
rect 180024 11880 180030 11892
rect 180061 11883 180119 11889
rect 180061 11880 180073 11883
rect 180024 11852 180073 11880
rect 180024 11840 180030 11852
rect 180061 11849 180073 11852
rect 180107 11849 180119 11883
rect 180061 11843 180119 11849
rect 180150 11840 180156 11892
rect 180208 11880 180214 11892
rect 188338 11880 188344 11892
rect 180208 11852 188344 11880
rect 180208 11840 180214 11852
rect 188338 11840 188344 11852
rect 188396 11840 188402 11892
rect 190825 11883 190883 11889
rect 190825 11849 190837 11883
rect 190871 11880 190883 11883
rect 191742 11880 191748 11892
rect 190871 11852 191748 11880
rect 190871 11849 190883 11852
rect 190825 11843 190883 11849
rect 191742 11840 191748 11852
rect 191800 11840 191806 11892
rect 191834 11840 191840 11892
rect 191892 11880 191898 11892
rect 194410 11880 194416 11892
rect 191892 11852 194416 11880
rect 191892 11840 191898 11852
rect 162578 11772 162584 11824
rect 162636 11812 162642 11824
rect 189534 11812 189540 11824
rect 162636 11784 189540 11812
rect 162636 11772 162642 11784
rect 189534 11772 189540 11784
rect 189592 11772 189598 11824
rect 193858 11812 193864 11824
rect 193338 11784 193864 11812
rect 193858 11772 193864 11784
rect 193916 11772 193922 11824
rect 162213 11747 162271 11753
rect 162213 11713 162225 11747
rect 162259 11744 162271 11747
rect 162857 11747 162915 11753
rect 162857 11744 162869 11747
rect 162259 11716 162869 11744
rect 162259 11713 162271 11716
rect 162213 11707 162271 11713
rect 162857 11713 162869 11716
rect 162903 11713 162915 11747
rect 163682 11744 163688 11756
rect 163643 11716 163688 11744
rect 162857 11707 162915 11713
rect 162872 11676 162900 11707
rect 163682 11704 163688 11716
rect 163740 11704 163746 11756
rect 164145 11747 164203 11753
rect 164145 11713 164157 11747
rect 164191 11744 164203 11747
rect 164789 11747 164847 11753
rect 164789 11744 164801 11747
rect 164191 11716 164801 11744
rect 164191 11713 164203 11716
rect 164145 11707 164203 11713
rect 164789 11713 164801 11716
rect 164835 11744 164847 11747
rect 166626 11744 166632 11756
rect 164835 11716 166632 11744
rect 164835 11713 164847 11716
rect 164789 11707 164847 11713
rect 163498 11676 163504 11688
rect 162872 11648 163504 11676
rect 163498 11636 163504 11648
rect 163556 11676 163562 11688
rect 164160 11676 164188 11707
rect 166626 11704 166632 11716
rect 166684 11704 166690 11756
rect 176654 11744 176660 11756
rect 176615 11716 176660 11744
rect 176654 11704 176660 11716
rect 176712 11704 176718 11756
rect 177945 11747 178003 11753
rect 177945 11713 177957 11747
rect 177991 11744 178003 11747
rect 179233 11747 179291 11753
rect 179233 11744 179245 11747
rect 177991 11716 179245 11744
rect 177991 11713 178003 11716
rect 177945 11707 178003 11713
rect 179233 11713 179245 11716
rect 179279 11744 179291 11747
rect 179874 11744 179880 11756
rect 179279 11716 179880 11744
rect 179279 11713 179291 11716
rect 179233 11707 179291 11713
rect 179874 11704 179880 11716
rect 179932 11704 179938 11756
rect 179969 11747 180027 11753
rect 179969 11713 179981 11747
rect 180015 11713 180027 11747
rect 179969 11707 180027 11713
rect 163556 11648 164188 11676
rect 163556 11636 163562 11648
rect 177114 11636 177120 11688
rect 177172 11676 177178 11688
rect 178129 11679 178187 11685
rect 178129 11676 178141 11679
rect 177172 11648 178141 11676
rect 177172 11636 177178 11648
rect 178129 11645 178141 11648
rect 178175 11676 178187 11679
rect 179325 11679 179383 11685
rect 179325 11676 179337 11679
rect 178175 11648 179337 11676
rect 178175 11645 178187 11648
rect 178129 11639 178187 11645
rect 165890 11608 165896 11620
rect 161952 11580 165896 11608
rect 161569 11571 161627 11577
rect 165890 11568 165896 11580
rect 165948 11568 165954 11620
rect 31386 11540 31392 11552
rect 29748 11512 30972 11540
rect 31347 11512 31392 11540
rect 31386 11500 31392 11512
rect 31444 11500 31450 11552
rect 32125 11543 32183 11549
rect 32125 11509 32137 11543
rect 32171 11540 32183 11543
rect 32950 11540 32956 11552
rect 32171 11512 32956 11540
rect 32171 11509 32183 11512
rect 32125 11503 32183 11509
rect 32950 11500 32956 11512
rect 33008 11500 33014 11552
rect 54941 11543 54999 11549
rect 54941 11509 54953 11543
rect 54987 11540 54999 11543
rect 55490 11540 55496 11552
rect 54987 11512 55496 11540
rect 54987 11509 54999 11512
rect 54941 11503 54999 11509
rect 55490 11500 55496 11512
rect 55548 11500 55554 11552
rect 84838 11500 84844 11552
rect 84896 11540 84902 11552
rect 85025 11543 85083 11549
rect 85025 11540 85037 11543
rect 84896 11512 85037 11540
rect 84896 11500 84902 11512
rect 85025 11509 85037 11512
rect 85071 11509 85083 11543
rect 85025 11503 85083 11509
rect 85669 11543 85727 11549
rect 85669 11509 85681 11543
rect 85715 11540 85727 11543
rect 86402 11540 86408 11552
rect 85715 11512 86408 11540
rect 85715 11509 85727 11512
rect 85669 11503 85727 11509
rect 86402 11500 86408 11512
rect 86460 11500 86466 11552
rect 101493 11543 101551 11549
rect 101493 11509 101505 11543
rect 101539 11540 101551 11543
rect 101858 11540 101864 11552
rect 101539 11512 101864 11540
rect 101539 11509 101551 11512
rect 101493 11503 101551 11509
rect 101858 11500 101864 11512
rect 101916 11500 101922 11552
rect 102965 11543 103023 11549
rect 102965 11509 102977 11543
rect 103011 11540 103023 11543
rect 104066 11540 104072 11552
rect 103011 11512 104072 11540
rect 103011 11509 103023 11512
rect 102965 11503 103023 11509
rect 104066 11500 104072 11512
rect 104124 11500 104130 11552
rect 114002 11500 114008 11552
rect 114060 11540 114066 11552
rect 114649 11543 114707 11549
rect 114649 11540 114661 11543
rect 114060 11512 114661 11540
rect 114060 11500 114066 11512
rect 114649 11509 114661 11512
rect 114695 11509 114707 11543
rect 131850 11540 131856 11552
rect 131811 11512 131856 11540
rect 114649 11503 114707 11509
rect 131850 11500 131856 11512
rect 131908 11500 131914 11552
rect 147306 11500 147312 11552
rect 147364 11540 147370 11552
rect 150069 11543 150127 11549
rect 150069 11540 150081 11543
rect 147364 11512 150081 11540
rect 147364 11500 147370 11512
rect 150069 11509 150081 11512
rect 150115 11540 150127 11543
rect 151722 11540 151728 11552
rect 150115 11512 151728 11540
rect 150115 11509 150127 11512
rect 150069 11503 150127 11509
rect 151722 11500 151728 11512
rect 151780 11500 151786 11552
rect 178696 11540 178724 11648
rect 179325 11645 179337 11648
rect 179371 11645 179383 11679
rect 179984 11676 180012 11707
rect 180058 11704 180064 11756
rect 180116 11744 180122 11756
rect 180610 11744 180616 11756
rect 180116 11716 180616 11744
rect 180116 11704 180122 11716
rect 180610 11704 180616 11716
rect 180668 11704 180674 11756
rect 180794 11676 180800 11688
rect 179984 11648 180800 11676
rect 179325 11639 179383 11645
rect 180794 11636 180800 11648
rect 180852 11676 180858 11688
rect 181530 11676 181536 11688
rect 180852 11648 181536 11676
rect 180852 11636 180858 11648
rect 181530 11636 181536 11648
rect 181588 11636 181594 11688
rect 189552 11676 189580 11772
rect 189626 11704 189632 11756
rect 189684 11744 189690 11756
rect 190089 11747 190147 11753
rect 189684 11716 189729 11744
rect 189684 11704 189690 11716
rect 190089 11713 190101 11747
rect 190135 11744 190147 11747
rect 190733 11747 190791 11753
rect 190733 11744 190745 11747
rect 190135 11716 190745 11744
rect 190135 11713 190147 11716
rect 190089 11707 190147 11713
rect 190733 11713 190745 11716
rect 190779 11744 190791 11747
rect 190822 11744 190828 11756
rect 190779 11716 190828 11744
rect 190779 11713 190791 11716
rect 190733 11707 190791 11713
rect 190104 11676 190132 11707
rect 190822 11704 190828 11716
rect 190880 11704 190886 11756
rect 191834 11744 191840 11756
rect 191795 11716 191840 11744
rect 191834 11704 191840 11716
rect 191892 11704 191898 11756
rect 194060 11753 194088 11852
rect 194410 11840 194416 11852
rect 194468 11840 194474 11892
rect 194686 11840 194692 11892
rect 194744 11880 194750 11892
rect 196253 11883 196311 11889
rect 196253 11880 196265 11883
rect 194744 11852 196265 11880
rect 194744 11840 194750 11852
rect 196253 11849 196265 11852
rect 196299 11849 196311 11883
rect 202874 11880 202880 11892
rect 202835 11852 202880 11880
rect 196253 11843 196311 11849
rect 202874 11840 202880 11852
rect 202932 11840 202938 11892
rect 204073 11883 204131 11889
rect 204073 11849 204085 11883
rect 204119 11880 204131 11883
rect 204530 11880 204536 11892
rect 204119 11852 204536 11880
rect 204119 11849 204131 11852
rect 204073 11843 204131 11849
rect 204530 11840 204536 11852
rect 204588 11840 204594 11892
rect 205177 11883 205235 11889
rect 205177 11849 205189 11883
rect 205223 11880 205235 11883
rect 206554 11880 206560 11892
rect 205223 11852 206560 11880
rect 205223 11849 205235 11852
rect 205177 11843 205235 11849
rect 206554 11840 206560 11852
rect 206612 11840 206618 11892
rect 227806 11840 227812 11892
rect 227864 11880 227870 11892
rect 228269 11883 228327 11889
rect 228269 11880 228281 11883
rect 227864 11852 228281 11880
rect 227864 11840 227870 11852
rect 228269 11849 228281 11852
rect 228315 11880 228327 11883
rect 228818 11880 228824 11892
rect 228315 11852 228824 11880
rect 228315 11849 228327 11852
rect 228269 11843 228327 11849
rect 228818 11840 228824 11852
rect 228876 11880 228882 11892
rect 229465 11883 229523 11889
rect 228876 11852 229094 11880
rect 228876 11840 228882 11852
rect 196802 11812 196808 11824
rect 195546 11784 196808 11812
rect 196802 11772 196808 11784
rect 196860 11772 196866 11824
rect 202325 11815 202383 11821
rect 202325 11781 202337 11815
rect 202371 11812 202383 11815
rect 203150 11812 203156 11824
rect 202371 11784 203156 11812
rect 202371 11781 202383 11784
rect 202325 11775 202383 11781
rect 203150 11772 203156 11784
rect 203208 11772 203214 11824
rect 203981 11815 204039 11821
rect 203981 11781 203993 11815
rect 204027 11812 204039 11815
rect 205269 11815 205327 11821
rect 205269 11812 205281 11815
rect 204027 11784 205281 11812
rect 204027 11781 204039 11784
rect 203981 11775 204039 11781
rect 205269 11781 205281 11784
rect 205315 11812 205327 11815
rect 205542 11812 205548 11824
rect 205315 11784 205548 11812
rect 205315 11781 205327 11784
rect 205269 11775 205327 11781
rect 205542 11772 205548 11784
rect 205600 11772 205606 11824
rect 227714 11772 227720 11824
rect 227772 11812 227778 11824
rect 228361 11815 228419 11821
rect 228361 11812 228373 11815
rect 227772 11784 228373 11812
rect 227772 11772 227778 11784
rect 228361 11781 228373 11784
rect 228407 11781 228419 11815
rect 229066 11812 229094 11852
rect 229465 11849 229477 11883
rect 229511 11880 229523 11883
rect 229922 11880 229928 11892
rect 229511 11852 229928 11880
rect 229511 11849 229523 11852
rect 229465 11843 229523 11849
rect 229922 11840 229928 11852
rect 229980 11840 229986 11892
rect 230382 11880 230388 11892
rect 230343 11852 230388 11880
rect 230382 11840 230388 11852
rect 230440 11840 230446 11892
rect 231026 11840 231032 11892
rect 231084 11880 231090 11892
rect 231581 11883 231639 11889
rect 231581 11880 231593 11883
rect 231084 11852 231593 11880
rect 231084 11840 231090 11852
rect 231581 11849 231593 11852
rect 231627 11849 231639 11883
rect 231581 11843 231639 11849
rect 231670 11840 231676 11892
rect 231728 11880 231734 11892
rect 238757 11883 238815 11889
rect 238757 11880 238769 11883
rect 231728 11852 238769 11880
rect 231728 11840 231734 11852
rect 238757 11849 238769 11852
rect 238803 11849 238815 11883
rect 240318 11880 240324 11892
rect 240279 11852 240324 11880
rect 238757 11843 238815 11849
rect 240318 11840 240324 11852
rect 240376 11840 240382 11892
rect 241054 11880 241060 11892
rect 241015 11852 241060 11880
rect 241054 11840 241060 11852
rect 241112 11840 241118 11892
rect 241790 11880 241796 11892
rect 241751 11852 241796 11880
rect 241790 11840 241796 11852
rect 241848 11840 241854 11892
rect 251821 11883 251879 11889
rect 251821 11849 251833 11883
rect 251867 11880 251879 11883
rect 252922 11880 252928 11892
rect 251867 11852 252928 11880
rect 251867 11849 251879 11852
rect 251821 11843 251879 11849
rect 252922 11840 252928 11852
rect 252980 11840 252986 11892
rect 254121 11883 254179 11889
rect 254121 11849 254133 11883
rect 254167 11880 254179 11883
rect 254670 11880 254676 11892
rect 254167 11852 254676 11880
rect 254167 11849 254179 11852
rect 254121 11843 254179 11849
rect 254670 11840 254676 11852
rect 254728 11840 254734 11892
rect 254762 11840 254768 11892
rect 254820 11880 254826 11892
rect 254949 11883 255007 11889
rect 254949 11880 254961 11883
rect 254820 11852 254961 11880
rect 254820 11840 254826 11852
rect 254949 11849 254961 11852
rect 254995 11849 255007 11883
rect 254949 11843 255007 11849
rect 255038 11840 255044 11892
rect 255096 11880 255102 11892
rect 255593 11883 255651 11889
rect 255593 11880 255605 11883
rect 255096 11852 255605 11880
rect 255096 11840 255102 11852
rect 255593 11849 255605 11852
rect 255639 11849 255651 11883
rect 255593 11843 255651 11849
rect 264977 11883 265035 11889
rect 264977 11849 264989 11883
rect 265023 11880 265035 11883
rect 266814 11880 266820 11892
rect 265023 11852 266820 11880
rect 265023 11849 265035 11852
rect 264977 11843 265035 11849
rect 266814 11840 266820 11852
rect 266872 11840 266878 11892
rect 267369 11883 267427 11889
rect 267369 11849 267381 11883
rect 267415 11880 267427 11883
rect 268197 11883 268255 11889
rect 267415 11852 267734 11880
rect 267415 11849 267427 11852
rect 267369 11843 267427 11849
rect 229557 11815 229615 11821
rect 229557 11812 229569 11815
rect 229066 11784 229569 11812
rect 228361 11775 228419 11781
rect 229557 11781 229569 11784
rect 229603 11781 229615 11815
rect 229557 11775 229615 11781
rect 194045 11747 194103 11753
rect 194045 11713 194057 11747
rect 194091 11713 194103 11747
rect 194045 11707 194103 11713
rect 196437 11747 196495 11753
rect 196437 11713 196449 11747
rect 196483 11744 196495 11747
rect 197906 11744 197912 11756
rect 196483 11716 197912 11744
rect 196483 11713 196495 11716
rect 196437 11707 196495 11713
rect 197906 11704 197912 11716
rect 197964 11704 197970 11756
rect 201034 11704 201040 11756
rect 201092 11744 201098 11756
rect 202233 11747 202291 11753
rect 202233 11744 202245 11747
rect 201092 11716 202245 11744
rect 201092 11704 201098 11716
rect 202233 11713 202245 11716
rect 202279 11713 202291 11747
rect 203058 11744 203064 11756
rect 203019 11716 203064 11744
rect 202233 11707 202291 11713
rect 203058 11704 203064 11716
rect 203116 11704 203122 11756
rect 206370 11744 206376 11756
rect 203168 11716 206376 11744
rect 192110 11676 192116 11688
rect 189552 11648 190132 11676
rect 192071 11648 192116 11676
rect 192110 11636 192116 11648
rect 192168 11636 192174 11688
rect 194318 11676 194324 11688
rect 194279 11648 194324 11676
rect 194318 11636 194324 11648
rect 194376 11636 194382 11688
rect 194410 11636 194416 11688
rect 194468 11676 194474 11688
rect 195793 11679 195851 11685
rect 194468 11648 195376 11676
rect 194468 11636 194474 11648
rect 178773 11611 178831 11617
rect 178773 11577 178785 11611
rect 178819 11608 178831 11611
rect 180334 11608 180340 11620
rect 178819 11580 180340 11608
rect 178819 11577 178831 11580
rect 178773 11571 178831 11577
rect 180334 11568 180340 11580
rect 180392 11568 180398 11620
rect 190181 11611 190239 11617
rect 190181 11577 190193 11611
rect 190227 11608 190239 11611
rect 195348 11608 195376 11648
rect 195793 11645 195805 11679
rect 195839 11676 195851 11679
rect 197354 11676 197360 11688
rect 195839 11648 197360 11676
rect 195839 11645 195851 11648
rect 195793 11639 195851 11645
rect 197354 11636 197360 11648
rect 197412 11676 197418 11688
rect 201310 11676 201316 11688
rect 197412 11648 201316 11676
rect 197412 11636 197418 11648
rect 201310 11636 201316 11648
rect 201368 11636 201374 11688
rect 202874 11636 202880 11688
rect 202932 11676 202938 11688
rect 203168 11676 203196 11716
rect 206370 11704 206376 11716
rect 206428 11704 206434 11756
rect 228376 11744 228404 11775
rect 230842 11772 230848 11824
rect 230900 11812 230906 11824
rect 238665 11815 238723 11821
rect 230900 11784 231072 11812
rect 230900 11772 230906 11784
rect 229370 11744 229376 11756
rect 228376 11716 229376 11744
rect 229370 11704 229376 11716
rect 229428 11704 229434 11756
rect 231044 11753 231072 11784
rect 238665 11781 238677 11815
rect 238711 11812 238723 11815
rect 240134 11812 240140 11824
rect 238711 11784 240140 11812
rect 238711 11781 238723 11784
rect 238665 11775 238723 11781
rect 240134 11772 240140 11784
rect 240192 11772 240198 11824
rect 241514 11812 241520 11824
rect 240244 11784 241520 11812
rect 230293 11747 230351 11753
rect 230293 11713 230305 11747
rect 230339 11744 230351 11747
rect 230937 11747 230995 11753
rect 230937 11744 230949 11747
rect 230339 11716 230949 11744
rect 230339 11713 230351 11716
rect 230293 11707 230351 11713
rect 230937 11713 230949 11716
rect 230983 11713 230995 11747
rect 230937 11707 230995 11713
rect 231029 11747 231087 11753
rect 231029 11713 231041 11747
rect 231075 11713 231087 11747
rect 231029 11707 231087 11713
rect 202932 11648 203196 11676
rect 202932 11636 202938 11648
rect 203518 11636 203524 11688
rect 203576 11676 203582 11688
rect 204257 11679 204315 11685
rect 204257 11676 204269 11679
rect 203576 11648 204269 11676
rect 203576 11636 203582 11648
rect 204257 11645 204269 11648
rect 204303 11676 204315 11679
rect 205453 11679 205511 11685
rect 205453 11676 205465 11679
rect 204303 11648 205465 11676
rect 204303 11645 204315 11648
rect 204257 11639 204315 11645
rect 205453 11645 205465 11648
rect 205499 11676 205511 11679
rect 207842 11676 207848 11688
rect 205499 11648 207848 11676
rect 205499 11645 205511 11648
rect 205453 11639 205511 11645
rect 207842 11636 207848 11648
rect 207900 11636 207906 11688
rect 227254 11636 227260 11688
rect 227312 11676 227318 11688
rect 228453 11679 228511 11685
rect 228453 11676 228465 11679
rect 227312 11648 228465 11676
rect 227312 11636 227318 11648
rect 228453 11645 228465 11648
rect 228499 11676 228511 11679
rect 229741 11679 229799 11685
rect 229741 11676 229753 11679
rect 228499 11648 229753 11676
rect 228499 11645 228511 11648
rect 228453 11639 228511 11645
rect 229741 11645 229753 11648
rect 229787 11676 229799 11679
rect 229787 11648 230888 11676
rect 229787 11645 229799 11648
rect 229741 11639 229799 11645
rect 197446 11608 197452 11620
rect 190227 11580 191972 11608
rect 195348 11580 197452 11608
rect 190227 11577 190239 11580
rect 190181 11571 190239 11577
rect 180518 11540 180524 11552
rect 178696 11512 180524 11540
rect 180518 11500 180524 11512
rect 180576 11500 180582 11552
rect 189442 11540 189448 11552
rect 189403 11512 189448 11540
rect 189442 11500 189448 11512
rect 189500 11500 189506 11552
rect 191944 11540 191972 11580
rect 197446 11568 197452 11580
rect 197504 11568 197510 11620
rect 203426 11568 203432 11620
rect 203484 11608 203490 11620
rect 204898 11608 204904 11620
rect 203484 11580 204904 11608
rect 203484 11568 203490 11580
rect 204898 11568 204904 11580
rect 204956 11568 204962 11620
rect 227901 11611 227959 11617
rect 227901 11577 227913 11611
rect 227947 11608 227959 11611
rect 230290 11608 230296 11620
rect 227947 11580 230296 11608
rect 227947 11577 227959 11580
rect 227901 11571 227959 11577
rect 230290 11568 230296 11580
rect 230348 11568 230354 11620
rect 193306 11540 193312 11552
rect 191944 11512 193312 11540
rect 193306 11500 193312 11512
rect 193364 11500 193370 11552
rect 193490 11500 193496 11552
rect 193548 11540 193554 11552
rect 193585 11543 193643 11549
rect 193585 11540 193597 11543
rect 193548 11512 193597 11540
rect 193548 11500 193554 11512
rect 193585 11509 193597 11512
rect 193631 11540 193643 11543
rect 195790 11540 195796 11552
rect 193631 11512 195796 11540
rect 193631 11509 193643 11512
rect 193585 11503 193643 11509
rect 195790 11500 195796 11512
rect 195848 11500 195854 11552
rect 195882 11500 195888 11552
rect 195940 11540 195946 11552
rect 196986 11540 196992 11552
rect 195940 11512 196992 11540
rect 195940 11500 195946 11512
rect 196986 11500 196992 11512
rect 197044 11500 197050 11552
rect 201494 11500 201500 11552
rect 201552 11540 201558 11552
rect 203613 11543 203671 11549
rect 203613 11540 203625 11543
rect 201552 11512 203625 11540
rect 201552 11500 201558 11512
rect 203613 11509 203625 11512
rect 203659 11509 203671 11543
rect 204806 11540 204812 11552
rect 204767 11512 204812 11540
rect 203613 11503 203671 11509
rect 204806 11500 204812 11512
rect 204864 11500 204870 11552
rect 229097 11543 229155 11549
rect 229097 11509 229109 11543
rect 229143 11540 229155 11543
rect 229370 11540 229376 11552
rect 229143 11512 229376 11540
rect 229143 11509 229155 11512
rect 229097 11503 229155 11509
rect 229370 11500 229376 11512
rect 229428 11500 229434 11552
rect 230860 11540 230888 11648
rect 230952 11608 230980 11707
rect 231210 11704 231216 11756
rect 231268 11744 231274 11756
rect 240244 11753 240272 11784
rect 241514 11772 241520 11784
rect 241572 11772 241578 11824
rect 244826 11812 244832 11824
rect 242636 11784 244832 11812
rect 231765 11747 231823 11753
rect 231765 11744 231777 11747
rect 231268 11716 231777 11744
rect 231268 11704 231274 11716
rect 231765 11713 231777 11716
rect 231811 11713 231823 11747
rect 231765 11707 231823 11713
rect 240229 11747 240287 11753
rect 240229 11713 240241 11747
rect 240275 11713 240287 11747
rect 241241 11747 241299 11753
rect 241241 11744 241253 11747
rect 240229 11707 240287 11713
rect 240612 11716 241253 11744
rect 239306 11636 239312 11688
rect 239364 11676 239370 11688
rect 239950 11676 239956 11688
rect 239364 11648 239956 11676
rect 239364 11636 239370 11648
rect 239950 11636 239956 11648
rect 240008 11676 240014 11688
rect 240413 11679 240471 11685
rect 240413 11676 240425 11679
rect 240008 11648 240425 11676
rect 240008 11636 240014 11648
rect 240413 11645 240425 11648
rect 240459 11645 240471 11679
rect 240413 11639 240471 11645
rect 232130 11608 232136 11620
rect 230952 11580 232136 11608
rect 232130 11568 232136 11580
rect 232188 11568 232194 11620
rect 239861 11611 239919 11617
rect 239861 11577 239873 11611
rect 239907 11608 239919 11611
rect 240612 11608 240640 11716
rect 241241 11713 241253 11716
rect 241287 11713 241299 11747
rect 241241 11707 241299 11713
rect 241701 11747 241759 11753
rect 241701 11713 241713 11747
rect 241747 11713 241759 11747
rect 242526 11744 242532 11756
rect 242487 11716 242532 11744
rect 241701 11707 241759 11713
rect 241716 11676 241744 11707
rect 242526 11704 242532 11716
rect 242584 11704 242590 11756
rect 241974 11676 241980 11688
rect 241716 11648 241980 11676
rect 241974 11636 241980 11648
rect 242032 11676 242038 11688
rect 242636 11676 242664 11784
rect 244826 11772 244832 11784
rect 244884 11772 244890 11824
rect 254029 11815 254087 11821
rect 254029 11781 254041 11815
rect 254075 11812 254087 11815
rect 254302 11812 254308 11824
rect 254075 11784 254308 11812
rect 254075 11781 254087 11784
rect 254029 11775 254087 11781
rect 254302 11772 254308 11784
rect 254360 11772 254366 11824
rect 264425 11815 264483 11821
rect 264425 11781 264437 11815
rect 264471 11812 264483 11815
rect 267706 11812 267734 11852
rect 268197 11849 268209 11883
rect 268243 11880 268255 11883
rect 270678 11880 270684 11892
rect 268243 11852 270684 11880
rect 268243 11849 268255 11852
rect 268197 11843 268255 11849
rect 270678 11840 270684 11852
rect 270736 11840 270742 11892
rect 270770 11840 270776 11892
rect 270828 11880 270834 11892
rect 271417 11883 271475 11889
rect 271417 11880 271429 11883
rect 270828 11852 271429 11880
rect 270828 11840 270834 11852
rect 271417 11849 271429 11852
rect 271463 11849 271475 11883
rect 271417 11843 271475 11849
rect 268286 11812 268292 11824
rect 264471 11784 266386 11812
rect 267706 11784 268292 11812
rect 264471 11781 264483 11784
rect 264425 11775 264483 11781
rect 268286 11772 268292 11784
rect 268344 11772 268350 11824
rect 269850 11772 269856 11824
rect 269908 11772 269914 11824
rect 252002 11744 252008 11756
rect 251963 11716 252008 11744
rect 252002 11704 252008 11716
rect 252060 11704 252066 11756
rect 252373 11747 252431 11753
rect 252373 11713 252385 11747
rect 252419 11744 252431 11747
rect 252738 11744 252744 11756
rect 252419 11716 252744 11744
rect 252419 11713 252431 11716
rect 252373 11707 252431 11713
rect 252738 11704 252744 11716
rect 252796 11704 252802 11756
rect 253014 11704 253020 11756
rect 253072 11744 253078 11756
rect 254857 11747 254915 11753
rect 254857 11744 254869 11747
rect 253072 11716 254869 11744
rect 253072 11704 253078 11716
rect 254857 11713 254869 11716
rect 254903 11744 254915 11747
rect 255501 11747 255559 11753
rect 255501 11744 255513 11747
rect 254903 11716 255513 11744
rect 254903 11713 254915 11716
rect 254857 11707 254915 11713
rect 255501 11713 255513 11716
rect 255547 11744 255559 11747
rect 256234 11744 256240 11756
rect 255547 11716 256240 11744
rect 255547 11713 255559 11716
rect 255501 11707 255559 11713
rect 256234 11704 256240 11716
rect 256292 11744 256298 11756
rect 257246 11744 257252 11756
rect 256292 11716 257252 11744
rect 256292 11704 256298 11716
rect 257246 11704 257252 11716
rect 257304 11704 257310 11756
rect 264330 11744 264336 11756
rect 264291 11716 264336 11744
rect 264330 11704 264336 11716
rect 264388 11704 264394 11756
rect 265158 11744 265164 11756
rect 265119 11716 265164 11744
rect 265158 11704 265164 11716
rect 265216 11704 265222 11756
rect 265250 11704 265256 11756
rect 265308 11744 265314 11756
rect 265621 11747 265679 11753
rect 265621 11744 265633 11747
rect 265308 11716 265633 11744
rect 265308 11704 265314 11716
rect 265621 11713 265633 11716
rect 265667 11713 265679 11747
rect 268470 11744 268476 11756
rect 265621 11707 265679 11713
rect 268304 11716 268476 11744
rect 242032 11648 242664 11676
rect 242032 11636 242038 11648
rect 242710 11636 242716 11688
rect 242768 11676 242774 11688
rect 244550 11676 244556 11688
rect 242768 11648 244556 11676
rect 242768 11636 242774 11648
rect 244550 11636 244556 11648
rect 244608 11636 244614 11688
rect 252094 11636 252100 11688
rect 252152 11676 252158 11688
rect 254213 11679 254271 11685
rect 254213 11676 254225 11679
rect 252152 11648 254225 11676
rect 252152 11636 252158 11648
rect 254213 11645 254225 11648
rect 254259 11676 254271 11679
rect 255590 11676 255596 11688
rect 254259 11648 255596 11676
rect 254259 11645 254271 11648
rect 254213 11639 254271 11645
rect 255590 11636 255596 11648
rect 255648 11676 255654 11688
rect 256418 11676 256424 11688
rect 255648 11648 256424 11676
rect 255648 11636 255654 11648
rect 256418 11636 256424 11648
rect 256476 11636 256482 11688
rect 263962 11636 263968 11688
rect 264020 11676 264026 11688
rect 268304 11685 268332 11716
rect 268470 11704 268476 11716
rect 268528 11704 268534 11756
rect 269114 11744 269120 11756
rect 269075 11716 269120 11744
rect 269114 11704 269120 11716
rect 269172 11704 269178 11756
rect 271322 11744 271328 11756
rect 271283 11716 271328 11744
rect 271322 11704 271328 11716
rect 271380 11704 271386 11756
rect 265897 11679 265955 11685
rect 265897 11676 265909 11679
rect 264020 11648 265909 11676
rect 264020 11636 264026 11648
rect 265897 11645 265909 11648
rect 265943 11645 265955 11679
rect 265897 11639 265955 11645
rect 268289 11679 268347 11685
rect 268289 11645 268301 11679
rect 268335 11645 268347 11679
rect 268289 11639 268347 11645
rect 268381 11679 268439 11685
rect 268381 11645 268393 11679
rect 268427 11645 268439 11679
rect 268381 11639 268439 11645
rect 239907 11580 240640 11608
rect 240704 11580 248414 11608
rect 239907 11577 239919 11580
rect 239861 11571 239919 11577
rect 231670 11540 231676 11552
rect 230860 11512 231676 11540
rect 231670 11500 231676 11512
rect 231728 11500 231734 11552
rect 239398 11500 239404 11552
rect 239456 11540 239462 11552
rect 240704 11540 240732 11580
rect 239456 11512 240732 11540
rect 239456 11500 239462 11512
rect 241238 11500 241244 11552
rect 241296 11540 241302 11552
rect 242345 11543 242403 11549
rect 242345 11540 242357 11543
rect 241296 11512 242357 11540
rect 241296 11500 241302 11512
rect 242345 11509 242357 11512
rect 242391 11509 242403 11543
rect 248386 11540 248414 11580
rect 251634 11568 251640 11620
rect 251692 11608 251698 11620
rect 252925 11611 252983 11617
rect 252925 11608 252937 11611
rect 251692 11580 252937 11608
rect 251692 11568 251698 11580
rect 252925 11577 252937 11580
rect 252971 11608 252983 11611
rect 252971 11580 260834 11608
rect 252971 11577 252983 11580
rect 252925 11571 252983 11577
rect 249058 11540 249064 11552
rect 248386 11512 249064 11540
rect 242345 11503 242403 11509
rect 249058 11500 249064 11512
rect 249116 11500 249122 11552
rect 253290 11500 253296 11552
rect 253348 11540 253354 11552
rect 253661 11543 253719 11549
rect 253661 11540 253673 11543
rect 253348 11512 253673 11540
rect 253348 11500 253354 11512
rect 253661 11509 253673 11512
rect 253707 11509 253719 11543
rect 260806 11540 260834 11580
rect 268010 11568 268016 11620
rect 268068 11608 268074 11620
rect 268396 11608 268424 11639
rect 268068 11580 268424 11608
rect 268068 11568 268074 11580
rect 261754 11540 261760 11552
rect 260806 11512 261760 11540
rect 253661 11503 253719 11509
rect 261754 11500 261760 11512
rect 261812 11500 261818 11552
rect 262674 11500 262680 11552
rect 262732 11540 262738 11552
rect 266262 11540 266268 11552
rect 262732 11512 266268 11540
rect 262732 11500 262738 11512
rect 266262 11500 266268 11512
rect 266320 11500 266326 11552
rect 266354 11500 266360 11552
rect 266412 11540 266418 11552
rect 267829 11543 267887 11549
rect 267829 11540 267841 11543
rect 266412 11512 267841 11540
rect 266412 11500 266418 11512
rect 267829 11509 267841 11512
rect 267875 11509 267887 11543
rect 268488 11540 268516 11704
rect 269390 11676 269396 11688
rect 269351 11648 269396 11676
rect 269390 11636 269396 11648
rect 269448 11636 269454 11688
rect 269942 11636 269948 11688
rect 270000 11676 270006 11688
rect 270865 11679 270923 11685
rect 270865 11676 270877 11679
rect 270000 11648 270877 11676
rect 270000 11636 270006 11648
rect 270865 11645 270877 11648
rect 270911 11676 270923 11679
rect 273162 11676 273168 11688
rect 270911 11648 273168 11676
rect 270911 11645 270923 11648
rect 270865 11639 270923 11645
rect 273162 11636 273168 11648
rect 273220 11636 273226 11688
rect 275094 11540 275100 11552
rect 268488 11512 275100 11540
rect 267829 11503 267887 11509
rect 275094 11500 275100 11512
rect 275152 11500 275158 11552
rect 1104 11450 305808 11472
rect 1104 11398 39049 11450
rect 39101 11398 39113 11450
rect 39165 11398 39177 11450
rect 39229 11398 39241 11450
rect 39293 11398 39305 11450
rect 39357 11398 115247 11450
rect 115299 11398 115311 11450
rect 115363 11398 115375 11450
rect 115427 11398 115439 11450
rect 115491 11398 115503 11450
rect 115555 11398 191445 11450
rect 191497 11398 191509 11450
rect 191561 11398 191573 11450
rect 191625 11398 191637 11450
rect 191689 11398 191701 11450
rect 191753 11398 267643 11450
rect 267695 11398 267707 11450
rect 267759 11398 267771 11450
rect 267823 11398 267835 11450
rect 267887 11398 267899 11450
rect 267951 11398 305808 11450
rect 1104 11376 305808 11398
rect 28813 11339 28871 11345
rect 28813 11305 28825 11339
rect 28859 11336 28871 11339
rect 29914 11336 29920 11348
rect 28859 11308 29920 11336
rect 28859 11305 28871 11308
rect 28813 11299 28871 11305
rect 29914 11296 29920 11308
rect 29972 11296 29978 11348
rect 30006 11296 30012 11348
rect 30064 11336 30070 11348
rect 30064 11308 31754 11336
rect 30064 11296 30070 11308
rect 28902 11228 28908 11280
rect 28960 11268 28966 11280
rect 31726 11268 31754 11308
rect 32398 11296 32404 11348
rect 32456 11336 32462 11348
rect 33318 11336 33324 11348
rect 32456 11308 33324 11336
rect 32456 11296 32462 11308
rect 33318 11296 33324 11308
rect 33376 11296 33382 11348
rect 33594 11336 33600 11348
rect 33555 11308 33600 11336
rect 33594 11296 33600 11308
rect 33652 11296 33658 11348
rect 40313 11339 40371 11345
rect 40313 11305 40325 11339
rect 40359 11336 40371 11339
rect 40402 11336 40408 11348
rect 40359 11308 40408 11336
rect 40359 11305 40371 11308
rect 40313 11299 40371 11305
rect 40402 11296 40408 11308
rect 40460 11296 40466 11348
rect 41046 11336 41052 11348
rect 41007 11308 41052 11336
rect 41046 11296 41052 11308
rect 41104 11296 41110 11348
rect 41598 11336 41604 11348
rect 41559 11308 41604 11336
rect 41598 11296 41604 11308
rect 41656 11296 41662 11348
rect 55030 11296 55036 11348
rect 55088 11336 55094 11348
rect 55309 11339 55367 11345
rect 55309 11336 55321 11339
rect 55088 11308 55321 11336
rect 55088 11296 55094 11308
rect 55309 11305 55321 11308
rect 55355 11305 55367 11339
rect 55309 11299 55367 11305
rect 56229 11339 56287 11345
rect 56229 11305 56241 11339
rect 56275 11336 56287 11339
rect 57698 11336 57704 11348
rect 56275 11308 57704 11336
rect 56275 11305 56287 11308
rect 56229 11299 56287 11305
rect 57698 11296 57704 11308
rect 57756 11296 57762 11348
rect 76374 11296 76380 11348
rect 76432 11336 76438 11348
rect 76469 11339 76527 11345
rect 76469 11336 76481 11339
rect 76432 11308 76481 11336
rect 76432 11296 76438 11308
rect 76469 11305 76481 11308
rect 76515 11305 76527 11339
rect 76469 11299 76527 11305
rect 78217 11339 78275 11345
rect 78217 11305 78229 11339
rect 78263 11336 78275 11339
rect 78766 11336 78772 11348
rect 78263 11308 78772 11336
rect 78263 11305 78275 11308
rect 78217 11299 78275 11305
rect 78766 11296 78772 11308
rect 78824 11296 78830 11348
rect 84470 11296 84476 11348
rect 84528 11336 84534 11348
rect 86221 11339 86279 11345
rect 86221 11336 86233 11339
rect 84528 11308 86233 11336
rect 84528 11296 84534 11308
rect 86221 11305 86233 11308
rect 86267 11305 86279 11339
rect 86221 11299 86279 11305
rect 86957 11339 87015 11345
rect 86957 11305 86969 11339
rect 87003 11336 87015 11339
rect 87138 11336 87144 11348
rect 87003 11308 87144 11336
rect 87003 11305 87015 11308
rect 86957 11299 87015 11305
rect 87138 11296 87144 11308
rect 87196 11296 87202 11348
rect 88245 11339 88303 11345
rect 88245 11305 88257 11339
rect 88291 11336 88303 11339
rect 89070 11336 89076 11348
rect 88291 11308 89076 11336
rect 88291 11305 88303 11308
rect 88245 11299 88303 11305
rect 89070 11296 89076 11308
rect 89128 11296 89134 11348
rect 102870 11336 102876 11348
rect 102831 11308 102876 11336
rect 102870 11296 102876 11308
rect 102928 11296 102934 11348
rect 115106 11296 115112 11348
rect 115164 11336 115170 11348
rect 116029 11339 116087 11345
rect 116029 11336 116041 11339
rect 115164 11308 116041 11336
rect 115164 11296 115170 11308
rect 116029 11305 116041 11308
rect 116075 11305 116087 11339
rect 116029 11299 116087 11305
rect 117133 11339 117191 11345
rect 117133 11305 117145 11339
rect 117179 11336 117191 11339
rect 117682 11336 117688 11348
rect 117179 11308 117688 11336
rect 117179 11305 117191 11308
rect 117133 11299 117191 11305
rect 117682 11296 117688 11308
rect 117740 11296 117746 11348
rect 130378 11296 130384 11348
rect 130436 11336 130442 11348
rect 130473 11339 130531 11345
rect 130473 11336 130485 11339
rect 130436 11308 130485 11336
rect 130436 11296 130442 11308
rect 130473 11305 130485 11308
rect 130519 11305 130531 11339
rect 131206 11336 131212 11348
rect 131167 11308 131212 11336
rect 130473 11299 130531 11305
rect 131206 11296 131212 11308
rect 131264 11296 131270 11348
rect 131761 11339 131819 11345
rect 131761 11305 131773 11339
rect 131807 11336 131819 11339
rect 132862 11336 132868 11348
rect 131807 11308 132868 11336
rect 131807 11305 131819 11308
rect 131761 11299 131819 11305
rect 132862 11296 132868 11308
rect 132920 11296 132926 11348
rect 148042 11336 148048 11348
rect 148003 11308 148048 11336
rect 148042 11296 148048 11308
rect 148100 11296 148106 11348
rect 150802 11336 150808 11348
rect 150763 11308 150808 11336
rect 150802 11296 150808 11308
rect 150860 11296 150866 11348
rect 157242 11296 157248 11348
rect 157300 11336 157306 11348
rect 157337 11339 157395 11345
rect 157337 11336 157349 11339
rect 157300 11308 157349 11336
rect 157300 11296 157306 11308
rect 157337 11305 157349 11308
rect 157383 11305 157395 11339
rect 157337 11299 157395 11305
rect 162029 11339 162087 11345
rect 162029 11305 162041 11339
rect 162075 11336 162087 11339
rect 162118 11336 162124 11348
rect 162075 11308 162124 11336
rect 162075 11305 162087 11308
rect 162029 11299 162087 11305
rect 162118 11296 162124 11308
rect 162176 11296 162182 11348
rect 162670 11336 162676 11348
rect 162631 11308 162676 11336
rect 162670 11296 162676 11308
rect 162728 11296 162734 11348
rect 163406 11296 163412 11348
rect 163464 11336 163470 11348
rect 163593 11339 163651 11345
rect 163593 11336 163605 11339
rect 163464 11308 163605 11336
rect 163464 11296 163470 11308
rect 163593 11305 163605 11308
rect 163639 11305 163651 11339
rect 163593 11299 163651 11305
rect 165890 11296 165896 11348
rect 165948 11336 165954 11348
rect 239398 11336 239404 11348
rect 165948 11308 239404 11336
rect 165948 11296 165954 11308
rect 239398 11296 239404 11308
rect 239456 11296 239462 11348
rect 239766 11296 239772 11348
rect 239824 11336 239830 11348
rect 239953 11339 240011 11345
rect 239953 11336 239965 11339
rect 239824 11308 239965 11336
rect 239824 11296 239830 11308
rect 239953 11305 239965 11308
rect 239999 11305 240011 11339
rect 239953 11299 240011 11305
rect 240042 11296 240048 11348
rect 240100 11336 240106 11348
rect 240873 11339 240931 11345
rect 240873 11336 240885 11339
rect 240100 11308 240885 11336
rect 240100 11296 240106 11308
rect 240873 11305 240885 11308
rect 240919 11305 240931 11339
rect 240873 11299 240931 11305
rect 240962 11296 240968 11348
rect 241020 11336 241026 11348
rect 241425 11339 241483 11345
rect 241425 11336 241437 11339
rect 241020 11308 241437 11336
rect 241020 11296 241026 11308
rect 241425 11305 241437 11308
rect 241471 11305 241483 11339
rect 241425 11299 241483 11305
rect 242066 11296 242072 11348
rect 242124 11336 242130 11348
rect 242161 11339 242219 11345
rect 242161 11336 242173 11339
rect 242124 11308 242173 11336
rect 242124 11296 242130 11308
rect 242161 11305 242173 11308
rect 242207 11305 242219 11339
rect 242161 11299 242219 11305
rect 252462 11296 252468 11348
rect 252520 11336 252526 11348
rect 252557 11339 252615 11345
rect 252557 11336 252569 11339
rect 252520 11308 252569 11336
rect 252520 11296 252526 11308
rect 252557 11305 252569 11308
rect 252603 11305 252615 11339
rect 253106 11336 253112 11348
rect 253067 11308 253112 11336
rect 252557 11299 252615 11305
rect 253106 11296 253112 11308
rect 253164 11296 253170 11348
rect 253753 11339 253811 11345
rect 253753 11305 253765 11339
rect 253799 11336 253811 11339
rect 254026 11336 254032 11348
rect 253799 11308 254032 11336
rect 253799 11305 253811 11308
rect 253753 11299 253811 11305
rect 254026 11296 254032 11308
rect 254084 11296 254090 11348
rect 265434 11296 265440 11348
rect 265492 11336 265498 11348
rect 265529 11339 265587 11345
rect 265529 11336 265541 11339
rect 265492 11308 265541 11336
rect 265492 11296 265498 11308
rect 265529 11305 265541 11308
rect 265575 11305 265587 11339
rect 265529 11299 265587 11305
rect 266262 11296 266268 11348
rect 266320 11336 266326 11348
rect 268013 11339 268071 11345
rect 266320 11308 267964 11336
rect 266320 11296 266326 11308
rect 36446 11268 36452 11280
rect 28960 11240 29776 11268
rect 31726 11240 36452 11268
rect 28960 11228 28966 11240
rect 27062 11160 27068 11212
rect 27120 11200 27126 11212
rect 29454 11200 29460 11212
rect 27120 11172 29460 11200
rect 27120 11160 27126 11172
rect 29454 11160 29460 11172
rect 29512 11160 29518 11212
rect 29546 11160 29552 11212
rect 29604 11200 29610 11212
rect 29641 11203 29699 11209
rect 29641 11200 29653 11203
rect 29604 11172 29653 11200
rect 29604 11160 29610 11172
rect 29641 11169 29653 11172
rect 29687 11169 29699 11203
rect 29748 11200 29776 11240
rect 36446 11228 36452 11240
rect 36504 11228 36510 11280
rect 41322 11228 41328 11280
rect 41380 11268 41386 11280
rect 42245 11271 42303 11277
rect 42245 11268 42257 11271
rect 41380 11240 42257 11268
rect 41380 11228 41386 11240
rect 42245 11237 42257 11240
rect 42291 11237 42303 11271
rect 42245 11231 42303 11237
rect 86770 11228 86776 11280
rect 86828 11268 86834 11280
rect 87601 11271 87659 11277
rect 87601 11268 87613 11271
rect 86828 11240 87613 11268
rect 86828 11228 86834 11240
rect 87601 11237 87613 11240
rect 87647 11237 87659 11271
rect 87601 11231 87659 11237
rect 102226 11228 102232 11280
rect 102284 11268 102290 11280
rect 103517 11271 103575 11277
rect 103517 11268 103529 11271
rect 102284 11240 103529 11268
rect 102284 11228 102290 11240
rect 103517 11237 103529 11240
rect 103563 11237 103575 11271
rect 103517 11231 103575 11237
rect 114186 11228 114192 11280
rect 114244 11268 114250 11280
rect 115385 11271 115443 11277
rect 115385 11268 115397 11271
rect 114244 11240 115397 11268
rect 114244 11228 114250 11240
rect 115385 11237 115397 11240
rect 115431 11237 115443 11271
rect 115385 11231 115443 11237
rect 147398 11228 147404 11280
rect 147456 11268 147462 11280
rect 149885 11271 149943 11277
rect 147456 11240 148732 11268
rect 147456 11228 147462 11240
rect 31386 11200 31392 11212
rect 29748 11172 31392 11200
rect 29641 11163 29699 11169
rect 31386 11160 31392 11172
rect 31444 11160 31450 11212
rect 32306 11200 32312 11212
rect 32267 11172 32312 11200
rect 32306 11160 32312 11172
rect 32364 11160 32370 11212
rect 32493 11203 32551 11209
rect 32493 11169 32505 11203
rect 32539 11200 32551 11203
rect 32582 11200 32588 11212
rect 32539 11172 32588 11200
rect 32539 11169 32551 11172
rect 32493 11163 32551 11169
rect 27614 11092 27620 11144
rect 27672 11132 27678 11144
rect 28997 11135 29055 11141
rect 28997 11132 29009 11135
rect 27672 11104 29009 11132
rect 27672 11092 27678 11104
rect 28997 11101 29009 11104
rect 29043 11101 29055 11135
rect 32214 11132 32220 11144
rect 32175 11104 32220 11132
rect 28997 11095 29055 11101
rect 32214 11092 32220 11104
rect 32272 11092 32278 11144
rect 27982 11024 27988 11076
rect 28040 11064 28046 11076
rect 29914 11064 29920 11076
rect 28040 11036 29776 11064
rect 29875 11036 29920 11064
rect 28040 11024 28046 11036
rect 29748 10996 29776 11036
rect 29914 11024 29920 11036
rect 29972 11024 29978 11076
rect 31662 11064 31668 11076
rect 31142 11036 31668 11064
rect 31662 11024 31668 11036
rect 31720 11024 31726 11076
rect 31754 11024 31760 11076
rect 31812 11064 31818 11076
rect 32508 11064 32536 11163
rect 32582 11160 32588 11172
rect 32640 11160 32646 11212
rect 45002 11200 45008 11212
rect 41800 11172 45008 11200
rect 33505 11135 33563 11141
rect 33505 11101 33517 11135
rect 33551 11132 33563 11135
rect 34698 11132 34704 11144
rect 33551 11104 34704 11132
rect 33551 11101 33563 11104
rect 33505 11095 33563 11101
rect 34698 11092 34704 11104
rect 34756 11092 34762 11144
rect 40494 11132 40500 11144
rect 40455 11104 40500 11132
rect 40494 11092 40500 11104
rect 40552 11092 40558 11144
rect 40957 11135 41015 11141
rect 40957 11101 40969 11135
rect 41003 11132 41015 11135
rect 41414 11132 41420 11144
rect 41003 11104 41420 11132
rect 41003 11101 41015 11104
rect 40957 11095 41015 11101
rect 41414 11092 41420 11104
rect 41472 11092 41478 11144
rect 41800 11141 41828 11172
rect 45002 11160 45008 11172
rect 45060 11160 45066 11212
rect 85482 11160 85488 11212
rect 85540 11200 85546 11212
rect 89162 11200 89168 11212
rect 85540 11172 89168 11200
rect 85540 11160 85546 11172
rect 41785 11135 41843 11141
rect 41785 11101 41797 11135
rect 41831 11101 41843 11135
rect 42426 11132 42432 11144
rect 42387 11104 42432 11132
rect 41785 11095 41843 11101
rect 42426 11092 42432 11104
rect 42484 11092 42490 11144
rect 55490 11132 55496 11144
rect 55451 11104 55496 11132
rect 55490 11092 55496 11104
rect 55548 11092 55554 11144
rect 56413 11135 56471 11141
rect 56413 11101 56425 11135
rect 56459 11132 56471 11135
rect 57238 11132 57244 11144
rect 56459 11104 57244 11132
rect 56459 11101 56471 11104
rect 56413 11095 56471 11101
rect 57238 11092 57244 11104
rect 57296 11092 57302 11144
rect 74718 11092 74724 11144
rect 74776 11132 74782 11144
rect 76653 11135 76711 11141
rect 76653 11132 76665 11135
rect 74776 11104 76665 11132
rect 74776 11092 74782 11104
rect 76653 11101 76665 11104
rect 76699 11101 76711 11135
rect 78398 11132 78404 11144
rect 78359 11104 78404 11132
rect 76653 11095 76711 11101
rect 78398 11092 78404 11104
rect 78456 11092 78462 11144
rect 86402 11132 86408 11144
rect 86363 11104 86408 11132
rect 86402 11092 86408 11104
rect 86460 11092 86466 11144
rect 86880 11141 86908 11172
rect 89162 11160 89168 11172
rect 89220 11160 89226 11212
rect 102042 11160 102048 11212
rect 102100 11200 102106 11212
rect 102321 11203 102379 11209
rect 102321 11200 102333 11203
rect 102100 11172 102333 11200
rect 102100 11160 102106 11172
rect 102321 11169 102333 11172
rect 102367 11169 102379 11203
rect 102321 11163 102379 11169
rect 102594 11160 102600 11212
rect 102652 11200 102658 11212
rect 102652 11172 103514 11200
rect 102652 11160 102658 11172
rect 86865 11135 86923 11141
rect 86865 11101 86877 11135
rect 86911 11101 86923 11135
rect 87782 11132 87788 11144
rect 87743 11104 87788 11132
rect 86865 11095 86923 11101
rect 87782 11092 87788 11104
rect 87840 11092 87846 11144
rect 88426 11132 88432 11144
rect 88387 11104 88432 11132
rect 88426 11092 88432 11104
rect 88484 11092 88490 11144
rect 102137 11135 102195 11141
rect 102137 11101 102149 11135
rect 102183 11132 102195 11135
rect 102410 11132 102416 11144
rect 102183 11104 102416 11132
rect 102183 11101 102195 11104
rect 102137 11095 102195 11101
rect 102410 11092 102416 11104
rect 102468 11092 102474 11144
rect 103054 11132 103060 11144
rect 103015 11104 103060 11132
rect 103054 11092 103060 11104
rect 103112 11092 103118 11144
rect 103486 11132 103514 11172
rect 130286 11160 130292 11212
rect 130344 11200 130350 11212
rect 132586 11200 132592 11212
rect 130344 11172 132592 11200
rect 130344 11160 130350 11172
rect 103701 11135 103759 11141
rect 103701 11132 103713 11135
rect 103486 11104 103713 11132
rect 103701 11101 103713 11104
rect 103747 11101 103759 11135
rect 103701 11095 103759 11101
rect 114738 11092 114744 11144
rect 114796 11132 114802 11144
rect 115293 11135 115351 11141
rect 115293 11132 115305 11135
rect 114796 11104 115305 11132
rect 114796 11092 114802 11104
rect 115293 11101 115305 11104
rect 115339 11132 115351 11135
rect 115750 11132 115756 11144
rect 115339 11104 115756 11132
rect 115339 11101 115351 11104
rect 115293 11095 115351 11101
rect 115750 11092 115756 11104
rect 115808 11092 115814 11144
rect 115842 11092 115848 11144
rect 115900 11132 115906 11144
rect 116213 11135 116271 11141
rect 116213 11132 116225 11135
rect 115900 11104 116225 11132
rect 115900 11092 115906 11104
rect 116213 11101 116225 11104
rect 116259 11101 116271 11135
rect 116213 11095 116271 11101
rect 117317 11135 117375 11141
rect 117317 11101 117329 11135
rect 117363 11132 117375 11135
rect 119706 11132 119712 11144
rect 117363 11104 119712 11132
rect 117363 11101 117375 11104
rect 117317 11095 117375 11101
rect 119706 11092 119712 11104
rect 119764 11092 119770 11144
rect 130657 11135 130715 11141
rect 130657 11101 130669 11135
rect 130703 11132 130715 11135
rect 130930 11132 130936 11144
rect 130703 11104 130936 11132
rect 130703 11101 130715 11104
rect 130657 11095 130715 11101
rect 130930 11092 130936 11104
rect 130988 11092 130994 11144
rect 131132 11141 131160 11172
rect 132586 11160 132592 11172
rect 132644 11160 132650 11212
rect 143258 11160 143264 11212
rect 143316 11200 143322 11212
rect 143316 11172 145880 11200
rect 143316 11160 143322 11172
rect 131117 11135 131175 11141
rect 131117 11101 131129 11135
rect 131163 11101 131175 11135
rect 131117 11095 131175 11101
rect 131945 11135 132003 11141
rect 131945 11101 131957 11135
rect 131991 11132 132003 11135
rect 133138 11132 133144 11144
rect 131991 11104 133144 11132
rect 131991 11101 132003 11104
rect 131945 11095 132003 11101
rect 133138 11092 133144 11104
rect 133196 11092 133202 11144
rect 142062 11132 142068 11144
rect 141975 11104 142068 11132
rect 142062 11092 142068 11104
rect 142120 11132 142126 11144
rect 145742 11132 145748 11144
rect 142120 11104 145748 11132
rect 142120 11092 142126 11104
rect 145742 11092 145748 11104
rect 145800 11092 145806 11144
rect 145852 11132 145880 11172
rect 147490 11160 147496 11212
rect 147548 11200 147554 11212
rect 148704 11209 148732 11240
rect 149885 11237 149897 11271
rect 149931 11268 149943 11271
rect 156414 11268 156420 11280
rect 149931 11240 156420 11268
rect 149931 11237 149943 11240
rect 149885 11231 149943 11237
rect 156414 11228 156420 11240
rect 156472 11228 156478 11280
rect 165430 11228 165436 11280
rect 165488 11268 165494 11280
rect 252738 11268 252744 11280
rect 165488 11240 192156 11268
rect 165488 11228 165494 11240
rect 148505 11203 148563 11209
rect 148505 11200 148517 11203
rect 147548 11172 148517 11200
rect 147548 11160 147554 11172
rect 148505 11169 148517 11172
rect 148551 11169 148563 11203
rect 148505 11163 148563 11169
rect 148689 11203 148747 11209
rect 148689 11169 148701 11203
rect 148735 11200 148747 11203
rect 151354 11200 151360 11212
rect 148735 11172 151360 11200
rect 148735 11169 148747 11172
rect 148689 11163 148747 11169
rect 151354 11160 151360 11172
rect 151412 11160 151418 11212
rect 165338 11200 165344 11212
rect 162872 11172 165344 11200
rect 150989 11135 151047 11141
rect 145852 11104 149560 11132
rect 31812 11036 32536 11064
rect 31812 11024 31818 11036
rect 81618 11024 81624 11076
rect 81676 11064 81682 11076
rect 87874 11064 87880 11076
rect 81676 11036 87880 11064
rect 81676 11024 81682 11036
rect 87874 11024 87880 11036
rect 87932 11024 87938 11076
rect 102428 11064 102456 11092
rect 113726 11064 113732 11076
rect 102428 11036 113732 11064
rect 113726 11024 113732 11036
rect 113784 11024 113790 11076
rect 140409 11067 140467 11073
rect 140409 11033 140421 11067
rect 140455 11064 140467 11067
rect 140682 11064 140688 11076
rect 140455 11036 140688 11064
rect 140455 11033 140467 11036
rect 140409 11027 140467 11033
rect 140682 11024 140688 11036
rect 140740 11064 140746 11076
rect 149532 11064 149560 11104
rect 150989 11101 151001 11135
rect 151035 11132 151047 11135
rect 153102 11132 153108 11144
rect 151035 11104 153108 11132
rect 151035 11101 151047 11104
rect 150989 11095 151047 11101
rect 153102 11092 153108 11104
rect 153160 11092 153166 11144
rect 162210 11132 162216 11144
rect 162171 11104 162216 11132
rect 162210 11092 162216 11104
rect 162268 11092 162274 11144
rect 162872 11141 162900 11172
rect 165338 11160 165344 11172
rect 165396 11160 165402 11212
rect 177577 11203 177635 11209
rect 177577 11169 177589 11203
rect 177623 11200 177635 11203
rect 177666 11200 177672 11212
rect 177623 11172 177672 11200
rect 177623 11169 177635 11172
rect 177577 11163 177635 11169
rect 177666 11160 177672 11172
rect 177724 11160 177730 11212
rect 177942 11160 177948 11212
rect 178000 11200 178006 11212
rect 178221 11203 178279 11209
rect 178221 11200 178233 11203
rect 178000 11172 178233 11200
rect 178000 11160 178006 11172
rect 178221 11169 178233 11172
rect 178267 11169 178279 11203
rect 180794 11200 180800 11212
rect 178221 11163 178279 11169
rect 178604 11172 180800 11200
rect 162857 11135 162915 11141
rect 162857 11101 162869 11135
rect 162903 11101 162915 11135
rect 163498 11132 163504 11144
rect 163459 11104 163504 11132
rect 162857 11095 162915 11101
rect 163498 11092 163504 11104
rect 163556 11092 163562 11144
rect 177485 11135 177543 11141
rect 177485 11101 177497 11135
rect 177531 11132 177543 11135
rect 178034 11132 178040 11144
rect 177531 11104 178040 11132
rect 177531 11101 177543 11104
rect 177485 11095 177543 11101
rect 178034 11092 178040 11104
rect 178092 11132 178098 11144
rect 178129 11135 178187 11141
rect 178129 11132 178141 11135
rect 178092 11104 178141 11132
rect 178092 11092 178098 11104
rect 178129 11101 178141 11104
rect 178175 11132 178187 11135
rect 178604 11132 178632 11172
rect 180794 11160 180800 11172
rect 180852 11160 180858 11212
rect 190273 11203 190331 11209
rect 190273 11169 190285 11203
rect 190319 11200 190331 11203
rect 191190 11200 191196 11212
rect 190319 11172 191196 11200
rect 190319 11169 190331 11172
rect 190273 11163 190331 11169
rect 191190 11160 191196 11172
rect 191248 11160 191254 11212
rect 191834 11160 191840 11212
rect 191892 11200 191898 11212
rect 192021 11203 192079 11209
rect 192021 11200 192033 11203
rect 191892 11172 192033 11200
rect 191892 11160 191898 11172
rect 192021 11169 192033 11172
rect 192067 11169 192079 11203
rect 192128 11200 192156 11240
rect 193324 11240 252744 11268
rect 193324 11200 193352 11240
rect 252738 11228 252744 11240
rect 252796 11228 252802 11280
rect 253198 11228 253204 11280
rect 253256 11268 253262 11280
rect 254397 11271 254455 11277
rect 254397 11268 254409 11271
rect 253256 11240 254409 11268
rect 253256 11228 253262 11240
rect 254397 11237 254409 11240
rect 254443 11237 254455 11271
rect 254397 11231 254455 11237
rect 265158 11228 265164 11280
rect 265216 11268 265222 11280
rect 266817 11271 266875 11277
rect 266817 11268 266829 11271
rect 265216 11240 266829 11268
rect 265216 11228 265222 11240
rect 266817 11237 266829 11240
rect 266863 11237 266875 11271
rect 267936 11268 267964 11308
rect 268013 11305 268025 11339
rect 268059 11336 268071 11339
rect 269298 11336 269304 11348
rect 268059 11308 269304 11336
rect 268059 11305 268071 11308
rect 268013 11299 268071 11305
rect 269298 11296 269304 11308
rect 269356 11296 269362 11348
rect 267936 11240 269436 11268
rect 266817 11231 266875 11237
rect 192128 11172 193352 11200
rect 192021 11163 192079 11169
rect 193490 11160 193496 11212
rect 193548 11200 193554 11212
rect 193769 11203 193827 11209
rect 193769 11200 193781 11203
rect 193548 11172 193781 11200
rect 193548 11160 193554 11172
rect 193769 11169 193781 11172
rect 193815 11200 193827 11203
rect 194410 11200 194416 11212
rect 193815 11172 194416 11200
rect 193815 11169 193827 11172
rect 193769 11163 193827 11169
rect 194410 11160 194416 11172
rect 194468 11160 194474 11212
rect 194594 11160 194600 11212
rect 194652 11200 194658 11212
rect 194965 11203 195023 11209
rect 194965 11200 194977 11203
rect 194652 11172 194977 11200
rect 194652 11160 194658 11172
rect 194965 11169 194977 11172
rect 195011 11169 195023 11203
rect 196434 11200 196440 11212
rect 194965 11163 195023 11169
rect 195440 11172 196440 11200
rect 178175 11104 178632 11132
rect 179141 11135 179199 11141
rect 178175 11101 178187 11104
rect 178129 11095 178187 11101
rect 179141 11101 179153 11135
rect 179187 11132 179199 11135
rect 180426 11132 180432 11144
rect 179187 11104 180432 11132
rect 179187 11101 179199 11104
rect 179141 11095 179199 11101
rect 180426 11092 180432 11104
rect 180484 11092 180490 11144
rect 188982 11092 188988 11144
rect 189040 11132 189046 11144
rect 190181 11135 190239 11141
rect 190181 11132 190193 11135
rect 189040 11104 190193 11132
rect 189040 11092 189046 11104
rect 190181 11101 190193 11104
rect 190227 11132 190239 11135
rect 190638 11132 190644 11144
rect 190227 11104 190644 11132
rect 190227 11101 190239 11104
rect 190181 11095 190239 11101
rect 190638 11092 190644 11104
rect 190696 11092 190702 11144
rect 190822 11132 190828 11144
rect 190783 11104 190828 11132
rect 190822 11092 190828 11104
rect 190880 11092 190886 11144
rect 190917 11135 190975 11141
rect 190917 11101 190929 11135
rect 190963 11132 190975 11135
rect 191926 11132 191932 11144
rect 190963 11104 191932 11132
rect 190963 11101 190975 11104
rect 190917 11095 190975 11101
rect 191926 11092 191932 11104
rect 191984 11092 191990 11144
rect 194781 11135 194839 11141
rect 194781 11101 194793 11135
rect 194827 11132 194839 11135
rect 194870 11132 194876 11144
rect 194827 11104 194876 11132
rect 194827 11101 194839 11104
rect 194781 11095 194839 11101
rect 194870 11092 194876 11104
rect 194928 11092 194934 11144
rect 195440 11132 195468 11172
rect 196434 11160 196440 11172
rect 196492 11160 196498 11212
rect 201034 11160 201040 11212
rect 201092 11200 201098 11212
rect 202877 11203 202935 11209
rect 201092 11172 202828 11200
rect 201092 11160 201098 11172
rect 195790 11132 195796 11144
rect 195164 11104 195468 11132
rect 195751 11104 195796 11132
rect 149609 11067 149667 11073
rect 149609 11064 149621 11067
rect 140740 11036 149468 11064
rect 149532 11036 149621 11064
rect 140740 11024 140746 11036
rect 31389 10999 31447 11005
rect 31389 10996 31401 10999
rect 29748 10968 31401 10996
rect 31389 10965 31401 10968
rect 31435 10965 31447 10999
rect 31846 10996 31852 11008
rect 31807 10968 31852 10996
rect 31389 10959 31447 10965
rect 31846 10956 31852 10968
rect 31904 10956 31910 11008
rect 148413 10999 148471 11005
rect 148413 10965 148425 10999
rect 148459 10996 148471 10999
rect 149054 10996 149060 11008
rect 148459 10968 149060 10996
rect 148459 10965 148471 10968
rect 148413 10959 148471 10965
rect 149054 10956 149060 10968
rect 149112 10956 149118 11008
rect 149440 10996 149468 11036
rect 149609 11033 149621 11036
rect 149655 11033 149667 11067
rect 156049 11067 156107 11073
rect 156049 11064 156061 11067
rect 149609 11027 149667 11033
rect 149716 11036 156061 11064
rect 149514 10996 149520 11008
rect 149440 10968 149520 10996
rect 149514 10956 149520 10968
rect 149572 10996 149578 11008
rect 149716 10996 149744 11036
rect 156049 11033 156061 11036
rect 156095 11064 156107 11067
rect 156138 11064 156144 11076
rect 156095 11036 156144 11064
rect 156095 11033 156107 11036
rect 156049 11027 156107 11033
rect 156138 11024 156144 11036
rect 156196 11024 156202 11076
rect 179414 11064 179420 11076
rect 178972 11036 179420 11064
rect 178972 11005 179000 11036
rect 179414 11024 179420 11036
rect 179472 11024 179478 11076
rect 189442 11024 189448 11076
rect 189500 11064 189506 11076
rect 192297 11067 192355 11073
rect 192297 11064 192309 11067
rect 189500 11036 192309 11064
rect 189500 11024 189506 11036
rect 192297 11033 192309 11036
rect 192343 11033 192355 11067
rect 192297 11027 192355 11033
rect 193306 11024 193312 11076
rect 193364 11024 193370 11076
rect 195164 11064 195192 11104
rect 195790 11092 195796 11104
rect 195848 11092 195854 11144
rect 202325 11135 202383 11141
rect 202325 11101 202337 11135
rect 202371 11132 202383 11135
rect 202690 11132 202696 11144
rect 202371 11104 202696 11132
rect 202371 11101 202383 11104
rect 202325 11095 202383 11101
rect 202690 11092 202696 11104
rect 202748 11092 202754 11144
rect 202800 11141 202828 11172
rect 202877 11169 202889 11203
rect 202923 11200 202935 11203
rect 203334 11200 203340 11212
rect 202923 11172 203340 11200
rect 202923 11169 202935 11172
rect 202877 11163 202935 11169
rect 203334 11160 203340 11172
rect 203392 11160 203398 11212
rect 204990 11200 204996 11212
rect 203536 11172 204996 11200
rect 202785 11135 202843 11141
rect 202785 11101 202797 11135
rect 202831 11132 202843 11135
rect 203429 11135 203487 11141
rect 203429 11132 203441 11135
rect 202831 11104 203441 11132
rect 202831 11101 202843 11104
rect 202785 11095 202843 11101
rect 203429 11101 203441 11104
rect 203475 11101 203487 11135
rect 203429 11095 203487 11101
rect 194888 11036 195192 11064
rect 149572 10968 149744 10996
rect 178957 10999 179015 11005
rect 149572 10956 149578 10968
rect 178957 10965 178969 10999
rect 179003 10965 179015 10999
rect 194410 10996 194416 11008
rect 194371 10968 194416 10996
rect 178957 10959 179015 10965
rect 194410 10956 194416 10968
rect 194468 10956 194474 11008
rect 194888 11005 194916 11036
rect 195238 11024 195244 11076
rect 195296 11064 195302 11076
rect 203536 11064 203564 11172
rect 204990 11160 204996 11172
rect 205048 11160 205054 11212
rect 238018 11160 238024 11212
rect 238076 11200 238082 11212
rect 242710 11200 242716 11212
rect 238076 11172 242716 11200
rect 238076 11160 238082 11172
rect 242710 11160 242716 11172
rect 242768 11160 242774 11212
rect 264977 11203 265035 11209
rect 264977 11169 264989 11203
rect 265023 11200 265035 11203
rect 267274 11200 267280 11212
rect 265023 11172 267280 11200
rect 265023 11169 265035 11172
rect 264977 11163 265035 11169
rect 267274 11160 267280 11172
rect 267332 11160 267338 11212
rect 267461 11203 267519 11209
rect 267461 11169 267473 11203
rect 267507 11200 267519 11203
rect 268010 11200 268016 11212
rect 267507 11172 268016 11200
rect 267507 11169 267519 11172
rect 267461 11163 267519 11169
rect 268010 11160 268016 11172
rect 268068 11160 268074 11212
rect 268470 11200 268476 11212
rect 268120 11172 268476 11200
rect 195296 11036 195652 11064
rect 195296 11024 195302 11036
rect 195624 11005 195652 11036
rect 202156 11036 203564 11064
rect 203628 11104 204852 11132
rect 202156 11005 202184 11036
rect 194873 10999 194931 11005
rect 194873 10965 194885 10999
rect 194919 10965 194931 10999
rect 194873 10959 194931 10965
rect 195609 10999 195667 11005
rect 195609 10965 195621 10999
rect 195655 10965 195667 10999
rect 195609 10959 195667 10965
rect 202141 10999 202199 11005
rect 202141 10965 202153 10999
rect 202187 10965 202199 10999
rect 202141 10959 202199 10965
rect 203521 10999 203579 11005
rect 203521 10965 203533 10999
rect 203567 10996 203579 10999
rect 203628 10996 203656 11104
rect 204070 11024 204076 11076
rect 204128 11064 204134 11076
rect 204824 11064 204852 11104
rect 204898 11092 204904 11144
rect 204956 11132 204962 11144
rect 229370 11132 229376 11144
rect 204956 11104 205001 11132
rect 229331 11104 229376 11132
rect 204956 11092 204962 11104
rect 229370 11092 229376 11104
rect 229428 11092 229434 11144
rect 239861 11135 239919 11141
rect 239861 11101 239873 11135
rect 239907 11132 239919 11135
rect 240781 11135 240839 11141
rect 240781 11132 240793 11135
rect 239907 11104 240793 11132
rect 239907 11101 239919 11104
rect 239861 11095 239919 11101
rect 240781 11101 240793 11104
rect 240827 11101 240839 11135
rect 240781 11095 240839 11101
rect 205450 11064 205456 11076
rect 204128 11036 204760 11064
rect 204824 11036 205456 11064
rect 204128 11024 204134 11036
rect 204732 11005 204760 11036
rect 205450 11024 205456 11036
rect 205508 11024 205514 11076
rect 230750 11064 230756 11076
rect 229204 11036 230756 11064
rect 229204 11005 229232 11036
rect 230750 11024 230756 11036
rect 230808 11024 230814 11076
rect 240796 11064 240824 11095
rect 240870 11092 240876 11144
rect 240928 11132 240934 11144
rect 241609 11135 241667 11141
rect 241609 11132 241621 11135
rect 240928 11104 241621 11132
rect 240928 11092 240934 11104
rect 241609 11101 241621 11104
rect 241655 11101 241667 11135
rect 241609 11095 241667 11101
rect 241974 11092 241980 11144
rect 242032 11132 242038 11144
rect 242069 11135 242127 11141
rect 242069 11132 242081 11135
rect 242032 11104 242081 11132
rect 242032 11092 242038 11104
rect 242069 11101 242081 11104
rect 242115 11101 242127 11135
rect 242069 11095 242127 11101
rect 251542 11092 251548 11144
rect 251600 11132 251606 11144
rect 252465 11135 252523 11141
rect 252465 11132 252477 11135
rect 251600 11104 252477 11132
rect 251600 11092 251606 11104
rect 252465 11101 252477 11104
rect 252511 11132 252523 11135
rect 253014 11132 253020 11144
rect 252511 11104 253020 11132
rect 252511 11101 252523 11104
rect 252465 11095 252523 11101
rect 253014 11092 253020 11104
rect 253072 11092 253078 11144
rect 253290 11132 253296 11144
rect 253251 11104 253296 11132
rect 253290 11092 253296 11104
rect 253348 11092 253354 11144
rect 253937 11135 253995 11141
rect 253937 11101 253949 11135
rect 253983 11132 253995 11135
rect 254394 11132 254400 11144
rect 253983 11104 254400 11132
rect 253983 11101 253995 11104
rect 253937 11095 253995 11101
rect 254394 11092 254400 11104
rect 254452 11092 254458 11144
rect 254581 11135 254639 11141
rect 254581 11101 254593 11135
rect 254627 11132 254639 11135
rect 254670 11132 254676 11144
rect 254627 11104 254676 11132
rect 254627 11101 254639 11104
rect 254581 11095 254639 11101
rect 254670 11092 254676 11104
rect 254728 11092 254734 11144
rect 264330 11092 264336 11144
rect 264388 11132 264394 11144
rect 264882 11132 264888 11144
rect 264388 11104 264888 11132
rect 264388 11092 264394 11104
rect 264882 11092 264888 11104
rect 264940 11092 264946 11144
rect 265618 11092 265624 11144
rect 265676 11132 265682 11144
rect 265713 11135 265771 11141
rect 265713 11132 265725 11135
rect 265676 11104 265725 11132
rect 265676 11092 265682 11104
rect 265713 11101 265725 11104
rect 265759 11101 265771 11135
rect 265713 11095 265771 11101
rect 267185 11135 267243 11141
rect 267185 11101 267197 11135
rect 267231 11132 267243 11135
rect 268120 11132 268148 11172
rect 268470 11160 268476 11172
rect 268528 11160 268534 11212
rect 268565 11203 268623 11209
rect 268565 11169 268577 11203
rect 268611 11200 268623 11203
rect 268930 11200 268936 11212
rect 268611 11172 268936 11200
rect 268611 11169 268623 11172
rect 268565 11163 268623 11169
rect 268930 11160 268936 11172
rect 268988 11160 268994 11212
rect 269408 11209 269436 11240
rect 269393 11203 269451 11209
rect 269393 11169 269405 11203
rect 269439 11200 269451 11203
rect 270589 11203 270647 11209
rect 270589 11200 270601 11203
rect 269439 11172 270601 11200
rect 269439 11169 269451 11172
rect 269393 11163 269451 11169
rect 270589 11169 270601 11172
rect 270635 11200 270647 11203
rect 272242 11200 272248 11212
rect 270635 11172 272248 11200
rect 270635 11169 270647 11172
rect 270589 11163 270647 11169
rect 272242 11160 272248 11172
rect 272300 11160 272306 11212
rect 267231 11104 268148 11132
rect 268197 11135 268255 11141
rect 267231 11101 267243 11104
rect 267185 11095 267243 11101
rect 268197 11101 268209 11135
rect 268243 11132 268255 11135
rect 269666 11132 269672 11144
rect 268243 11104 269672 11132
rect 268243 11101 268255 11104
rect 268197 11095 268255 11101
rect 269666 11092 269672 11104
rect 269724 11092 269730 11144
rect 270402 11132 270408 11144
rect 270363 11104 270408 11132
rect 270402 11092 270408 11104
rect 270460 11092 270466 11144
rect 270497 11135 270555 11141
rect 270497 11101 270509 11135
rect 270543 11132 270555 11135
rect 270862 11132 270868 11144
rect 270543 11104 270868 11132
rect 270543 11101 270555 11104
rect 270497 11095 270555 11101
rect 270862 11092 270868 11104
rect 270920 11092 270926 11144
rect 241992 11064 242020 11092
rect 240796 11036 242020 11064
rect 267277 11067 267335 11073
rect 267277 11033 267289 11067
rect 267323 11064 267335 11067
rect 268286 11064 268292 11076
rect 267323 11036 268292 11064
rect 267323 11033 267335 11036
rect 267277 11027 267335 11033
rect 268286 11024 268292 11036
rect 268344 11024 268350 11076
rect 268930 11024 268936 11076
rect 268988 11064 268994 11076
rect 269209 11067 269267 11073
rect 269209 11064 269221 11067
rect 268988 11036 269221 11064
rect 268988 11024 268994 11036
rect 269209 11033 269221 11036
rect 269255 11033 269267 11067
rect 269209 11027 269267 11033
rect 269301 11067 269359 11073
rect 269301 11033 269313 11067
rect 269347 11064 269359 11067
rect 269942 11064 269948 11076
rect 269347 11036 269948 11064
rect 269347 11033 269359 11036
rect 269301 11027 269359 11033
rect 269942 11024 269948 11036
rect 270000 11024 270006 11076
rect 203567 10968 203656 10996
rect 204717 10999 204775 11005
rect 203567 10965 203579 10968
rect 203521 10959 203579 10965
rect 204717 10965 204729 10999
rect 204763 10965 204775 10999
rect 204717 10959 204775 10965
rect 229189 10999 229247 11005
rect 229189 10965 229201 10999
rect 229235 10965 229247 10999
rect 268838 10996 268844 11008
rect 268799 10968 268844 10996
rect 229189 10959 229247 10965
rect 268838 10956 268844 10968
rect 268896 10956 268902 11008
rect 270034 10996 270040 11008
rect 269995 10968 270040 10996
rect 270034 10956 270040 10968
rect 270092 10956 270098 11008
rect 1104 10906 305808 10928
rect 1104 10854 77148 10906
rect 77200 10854 77212 10906
rect 77264 10854 77276 10906
rect 77328 10854 77340 10906
rect 77392 10854 77404 10906
rect 77456 10854 153346 10906
rect 153398 10854 153410 10906
rect 153462 10854 153474 10906
rect 153526 10854 153538 10906
rect 153590 10854 153602 10906
rect 153654 10854 229544 10906
rect 229596 10854 229608 10906
rect 229660 10854 229672 10906
rect 229724 10854 229736 10906
rect 229788 10854 229800 10906
rect 229852 10854 305808 10906
rect 1104 10832 305808 10854
rect 29641 10795 29699 10801
rect 29641 10761 29653 10795
rect 29687 10792 29699 10795
rect 29822 10792 29828 10804
rect 29687 10764 29828 10792
rect 29687 10761 29699 10764
rect 29641 10755 29699 10761
rect 29822 10752 29828 10764
rect 29880 10752 29886 10804
rect 30466 10752 30472 10804
rect 30524 10792 30530 10804
rect 30653 10795 30711 10801
rect 30653 10792 30665 10795
rect 30524 10764 30665 10792
rect 30524 10752 30530 10764
rect 30653 10761 30665 10764
rect 30699 10761 30711 10795
rect 30653 10755 30711 10761
rect 30742 10752 30748 10804
rect 30800 10792 30806 10804
rect 32125 10795 32183 10801
rect 32125 10792 32137 10795
rect 30800 10764 30845 10792
rect 30944 10764 32137 10792
rect 30800 10752 30806 10764
rect 29730 10684 29736 10736
rect 29788 10724 29794 10736
rect 29788 10696 30144 10724
rect 29788 10684 29794 10696
rect 28442 10616 28448 10668
rect 28500 10656 28506 10668
rect 29825 10659 29883 10665
rect 29825 10656 29837 10659
rect 28500 10628 29837 10656
rect 28500 10616 28506 10628
rect 29825 10625 29837 10628
rect 29871 10625 29883 10659
rect 30116 10656 30144 10696
rect 30190 10684 30196 10736
rect 30248 10724 30254 10736
rect 30944 10724 30972 10764
rect 32125 10761 32137 10764
rect 32171 10761 32183 10795
rect 32125 10755 32183 10761
rect 32674 10752 32680 10804
rect 32732 10792 32738 10804
rect 32769 10795 32827 10801
rect 32769 10792 32781 10795
rect 32732 10764 32781 10792
rect 32732 10752 32738 10764
rect 32769 10761 32781 10764
rect 32815 10761 32827 10795
rect 32769 10755 32827 10761
rect 33042 10752 33048 10804
rect 33100 10792 33106 10804
rect 33413 10795 33471 10801
rect 33413 10792 33425 10795
rect 33100 10764 33425 10792
rect 33100 10752 33106 10764
rect 33413 10761 33425 10764
rect 33459 10761 33471 10795
rect 101674 10792 101680 10804
rect 101635 10764 101680 10792
rect 33413 10755 33471 10761
rect 101674 10752 101680 10764
rect 101732 10752 101738 10804
rect 130470 10792 130476 10804
rect 130431 10764 130476 10792
rect 130470 10752 130476 10764
rect 130528 10752 130534 10804
rect 141970 10792 141976 10804
rect 141931 10764 141976 10792
rect 141970 10752 141976 10764
rect 142028 10752 142034 10804
rect 148594 10752 148600 10804
rect 148652 10792 148658 10804
rect 148873 10795 148931 10801
rect 148873 10792 148885 10795
rect 148652 10764 148885 10792
rect 148652 10752 148658 10764
rect 148873 10761 148885 10764
rect 148919 10761 148931 10795
rect 148873 10755 148931 10761
rect 148962 10752 148968 10804
rect 149020 10792 149026 10804
rect 150713 10795 150771 10801
rect 150713 10792 150725 10795
rect 149020 10764 150725 10792
rect 149020 10752 149026 10764
rect 150713 10761 150725 10764
rect 150759 10761 150771 10795
rect 150713 10755 150771 10761
rect 191098 10752 191104 10804
rect 191156 10792 191162 10804
rect 191837 10795 191895 10801
rect 191837 10792 191849 10795
rect 191156 10764 191849 10792
rect 191156 10752 191162 10764
rect 191837 10761 191849 10764
rect 191883 10761 191895 10795
rect 191837 10755 191895 10761
rect 192128 10764 193812 10792
rect 31754 10724 31760 10736
rect 30248 10696 30972 10724
rect 31036 10696 31760 10724
rect 30248 10684 30254 10696
rect 31036 10656 31064 10696
rect 31754 10684 31760 10696
rect 31812 10684 31818 10736
rect 31846 10684 31852 10736
rect 31904 10724 31910 10736
rect 140682 10724 140688 10736
rect 31904 10696 33640 10724
rect 140643 10696 140688 10724
rect 31904 10684 31910 10696
rect 32309 10659 32367 10665
rect 32309 10656 32321 10659
rect 30116 10628 31064 10656
rect 31726 10628 32321 10656
rect 29825 10619 29883 10625
rect 30852 10597 30880 10628
rect 30837 10591 30895 10597
rect 30837 10557 30849 10591
rect 30883 10557 30895 10591
rect 30837 10551 30895 10557
rect 30285 10523 30343 10529
rect 30285 10489 30297 10523
rect 30331 10520 30343 10523
rect 31726 10520 31754 10628
rect 32309 10625 32321 10628
rect 32355 10625 32367 10659
rect 32950 10656 32956 10668
rect 32911 10628 32956 10656
rect 32309 10619 32367 10625
rect 32950 10616 32956 10628
rect 33008 10616 33014 10668
rect 33612 10665 33640 10696
rect 140682 10684 140688 10696
rect 140740 10684 140746 10736
rect 151630 10724 151636 10736
rect 149072 10696 151636 10724
rect 33597 10659 33655 10665
rect 33597 10625 33609 10659
rect 33643 10625 33655 10659
rect 101858 10656 101864 10668
rect 101819 10628 101864 10656
rect 33597 10619 33655 10625
rect 101858 10616 101864 10628
rect 101916 10616 101922 10668
rect 130286 10616 130292 10668
rect 130344 10656 130350 10668
rect 149072 10665 149100 10696
rect 151630 10684 151636 10696
rect 151688 10684 151694 10736
rect 156138 10724 156144 10736
rect 156099 10696 156144 10724
rect 156138 10684 156144 10696
rect 156196 10684 156202 10736
rect 192128 10724 192156 10764
rect 187252 10696 192156 10724
rect 130381 10659 130439 10665
rect 130381 10656 130393 10659
rect 130344 10628 130393 10656
rect 130344 10616 130350 10628
rect 130381 10625 130393 10628
rect 130427 10625 130439 10659
rect 130381 10619 130439 10625
rect 149057 10659 149115 10665
rect 149057 10625 149069 10659
rect 149103 10625 149115 10659
rect 149057 10619 149115 10625
rect 150342 10616 150348 10668
rect 150400 10656 150406 10668
rect 187252 10665 187280 10696
rect 192202 10684 192208 10736
rect 192260 10724 192266 10736
rect 192260 10696 192708 10724
rect 192260 10684 192266 10696
rect 150621 10659 150679 10665
rect 150621 10656 150633 10659
rect 150400 10628 150633 10656
rect 150400 10616 150406 10628
rect 150621 10625 150633 10628
rect 150667 10625 150679 10659
rect 150621 10619 150679 10625
rect 187237 10659 187295 10665
rect 187237 10625 187249 10659
rect 187283 10625 187295 10659
rect 187237 10619 187295 10625
rect 190546 10616 190552 10668
rect 190604 10656 190610 10668
rect 191285 10659 191343 10665
rect 191285 10656 191297 10659
rect 190604 10628 191297 10656
rect 190604 10616 190610 10628
rect 191285 10625 191297 10628
rect 191331 10625 191343 10659
rect 191285 10619 191343 10625
rect 192021 10659 192079 10665
rect 192021 10625 192033 10659
rect 192067 10656 192079 10659
rect 192294 10656 192300 10668
rect 192067 10628 192300 10656
rect 192067 10625 192079 10628
rect 192021 10619 192079 10625
rect 192294 10616 192300 10628
rect 192352 10616 192358 10668
rect 192680 10665 192708 10696
rect 193214 10684 193220 10736
rect 193272 10724 193278 10736
rect 193493 10727 193551 10733
rect 193493 10724 193505 10727
rect 193272 10696 193505 10724
rect 193272 10684 193278 10696
rect 193493 10693 193505 10696
rect 193539 10693 193551 10727
rect 193784 10724 193812 10764
rect 193858 10752 193864 10804
rect 193916 10792 193922 10804
rect 194229 10795 194287 10801
rect 194229 10792 194241 10795
rect 193916 10764 194241 10792
rect 193916 10752 193922 10764
rect 194229 10761 194241 10764
rect 194275 10761 194287 10795
rect 194229 10755 194287 10761
rect 202877 10795 202935 10801
rect 202877 10761 202889 10795
rect 202923 10792 202935 10795
rect 205082 10792 205088 10804
rect 202923 10764 205088 10792
rect 202923 10761 202935 10764
rect 202877 10755 202935 10761
rect 205082 10752 205088 10764
rect 205140 10752 205146 10804
rect 253661 10795 253719 10801
rect 253661 10761 253673 10795
rect 253707 10792 253719 10795
rect 255222 10792 255228 10804
rect 253707 10764 255228 10792
rect 253707 10761 253719 10764
rect 253661 10755 253719 10761
rect 255222 10752 255228 10764
rect 255280 10752 255286 10804
rect 266538 10792 266544 10804
rect 266499 10764 266544 10792
rect 266538 10752 266544 10764
rect 266596 10752 266602 10804
rect 267737 10795 267795 10801
rect 267737 10761 267749 10795
rect 267783 10792 267795 10795
rect 268194 10792 268200 10804
rect 267783 10764 268200 10792
rect 267783 10761 267795 10764
rect 267737 10755 267795 10761
rect 268194 10752 268200 10764
rect 268252 10752 268258 10804
rect 268381 10795 268439 10801
rect 268381 10761 268393 10795
rect 268427 10792 268439 10795
rect 269390 10792 269396 10804
rect 268427 10764 269396 10792
rect 268427 10761 268439 10764
rect 268381 10755 268439 10761
rect 269390 10752 269396 10764
rect 269448 10752 269454 10804
rect 195054 10724 195060 10736
rect 193784 10696 195060 10724
rect 193493 10687 193551 10693
rect 195054 10684 195060 10696
rect 195112 10684 195118 10736
rect 264882 10684 264888 10736
rect 264940 10724 264946 10736
rect 270034 10724 270040 10736
rect 264940 10696 266492 10724
rect 264940 10684 264946 10696
rect 192665 10659 192723 10665
rect 192665 10625 192677 10659
rect 192711 10625 192723 10659
rect 194134 10656 194140 10668
rect 194095 10628 194140 10656
rect 192665 10619 192723 10625
rect 194134 10616 194140 10628
rect 194192 10656 194198 10668
rect 194962 10656 194968 10668
rect 194192 10628 194968 10656
rect 194192 10616 194198 10628
rect 194962 10616 194968 10628
rect 195020 10616 195026 10668
rect 203061 10659 203119 10665
rect 203061 10625 203073 10659
rect 203107 10656 203119 10659
rect 204806 10656 204812 10668
rect 203107 10628 204812 10656
rect 203107 10625 203119 10628
rect 203061 10619 203119 10625
rect 204806 10616 204812 10628
rect 204864 10616 204870 10668
rect 253845 10659 253903 10665
rect 253845 10625 253857 10659
rect 253891 10656 253903 10659
rect 254946 10656 254952 10668
rect 253891 10628 254952 10656
rect 253891 10625 253903 10628
rect 253845 10619 253903 10625
rect 254946 10616 254952 10628
rect 255004 10616 255010 10668
rect 265989 10659 266047 10665
rect 265989 10625 266001 10659
rect 266035 10656 266047 10659
rect 266354 10656 266360 10668
rect 266035 10628 266360 10656
rect 266035 10625 266047 10628
rect 265989 10619 266047 10625
rect 266354 10616 266360 10628
rect 266412 10616 266418 10668
rect 266464 10665 266492 10696
rect 267936 10696 270040 10724
rect 267936 10665 267964 10696
rect 270034 10684 270040 10696
rect 270092 10684 270098 10736
rect 266449 10659 266507 10665
rect 266449 10625 266461 10659
rect 266495 10656 266507 10659
rect 267093 10659 267151 10665
rect 267093 10656 267105 10659
rect 266495 10628 267105 10656
rect 266495 10625 266507 10628
rect 266449 10619 266507 10625
rect 267093 10625 267105 10628
rect 267139 10625 267151 10659
rect 267093 10619 267151 10625
rect 267921 10659 267979 10665
rect 267921 10625 267933 10659
rect 267967 10625 267979 10659
rect 267921 10619 267979 10625
rect 268565 10659 268623 10665
rect 268565 10625 268577 10659
rect 268611 10625 268623 10659
rect 268565 10619 268623 10625
rect 187510 10588 187516 10600
rect 187471 10560 187516 10588
rect 187510 10548 187516 10560
rect 187568 10548 187574 10600
rect 201034 10588 201040 10600
rect 192864 10560 201040 10588
rect 30331 10492 31754 10520
rect 191101 10523 191159 10529
rect 30331 10489 30343 10492
rect 30285 10483 30343 10489
rect 191101 10489 191113 10523
rect 191147 10520 191159 10523
rect 192110 10520 192116 10532
rect 191147 10492 192116 10520
rect 191147 10489 191159 10492
rect 191101 10483 191159 10489
rect 192110 10480 192116 10492
rect 192168 10480 192174 10532
rect 192864 10529 192892 10560
rect 201034 10548 201040 10560
rect 201092 10548 201098 10600
rect 268580 10588 268608 10619
rect 269022 10616 269028 10668
rect 269080 10656 269086 10668
rect 269117 10659 269175 10665
rect 269117 10656 269129 10659
rect 269080 10628 269129 10656
rect 269080 10616 269086 10628
rect 269117 10625 269129 10628
rect 269163 10625 269175 10659
rect 269117 10619 269175 10625
rect 269209 10659 269267 10665
rect 269209 10625 269221 10659
rect 269255 10656 269267 10659
rect 270310 10656 270316 10668
rect 269255 10628 270316 10656
rect 269255 10625 269267 10628
rect 269209 10619 269267 10625
rect 270310 10616 270316 10628
rect 270368 10616 270374 10668
rect 272518 10588 272524 10600
rect 268580 10560 272524 10588
rect 272518 10548 272524 10560
rect 272576 10548 272582 10600
rect 192849 10523 192907 10529
rect 192849 10489 192861 10523
rect 192895 10489 192907 10523
rect 192849 10483 192907 10489
rect 193677 10523 193735 10529
rect 193677 10489 193689 10523
rect 193723 10520 193735 10523
rect 267185 10523 267243 10529
rect 193723 10492 196848 10520
rect 193723 10489 193735 10492
rect 193677 10483 193735 10489
rect 157613 10455 157671 10461
rect 157613 10421 157625 10455
rect 157659 10452 157671 10455
rect 179138 10452 179144 10464
rect 157659 10424 179144 10452
rect 157659 10421 157671 10424
rect 157613 10415 157671 10421
rect 179138 10412 179144 10424
rect 179196 10412 179202 10464
rect 196820 10452 196848 10492
rect 267185 10489 267197 10523
rect 267231 10520 267243 10523
rect 268746 10520 268752 10532
rect 267231 10492 268752 10520
rect 267231 10489 267243 10492
rect 267185 10483 267243 10489
rect 268746 10480 268752 10492
rect 268804 10480 268810 10532
rect 203518 10452 203524 10464
rect 196820 10424 203524 10452
rect 203518 10412 203524 10424
rect 203576 10412 203582 10464
rect 265805 10455 265863 10461
rect 265805 10421 265817 10455
rect 265851 10452 265863 10455
rect 269574 10452 269580 10464
rect 265851 10424 269580 10452
rect 265851 10421 265863 10424
rect 265805 10415 265863 10421
rect 269574 10412 269580 10424
rect 269632 10412 269638 10464
rect 1104 10362 305808 10384
rect 1104 10310 39049 10362
rect 39101 10310 39113 10362
rect 39165 10310 39177 10362
rect 39229 10310 39241 10362
rect 39293 10310 39305 10362
rect 39357 10310 115247 10362
rect 115299 10310 115311 10362
rect 115363 10310 115375 10362
rect 115427 10310 115439 10362
rect 115491 10310 115503 10362
rect 115555 10310 191445 10362
rect 191497 10310 191509 10362
rect 191561 10310 191573 10362
rect 191625 10310 191637 10362
rect 191689 10310 191701 10362
rect 191753 10310 267643 10362
rect 267695 10310 267707 10362
rect 267759 10310 267771 10362
rect 267823 10310 267835 10362
rect 267887 10310 267899 10362
rect 267951 10310 305808 10362
rect 1104 10288 305808 10310
rect 30098 10208 30104 10260
rect 30156 10248 30162 10260
rect 30929 10251 30987 10257
rect 30929 10248 30941 10251
rect 30156 10220 30941 10248
rect 30156 10208 30162 10220
rect 30929 10217 30941 10220
rect 30975 10217 30987 10251
rect 31662 10248 31668 10260
rect 31623 10220 31668 10248
rect 30929 10211 30987 10217
rect 31662 10208 31668 10220
rect 31720 10208 31726 10260
rect 32122 10208 32128 10260
rect 32180 10248 32186 10260
rect 32861 10251 32919 10257
rect 32861 10248 32873 10251
rect 32180 10220 32873 10248
rect 32180 10208 32186 10220
rect 32861 10217 32873 10220
rect 32907 10217 32919 10251
rect 32861 10211 32919 10217
rect 33318 10208 33324 10260
rect 33376 10248 33382 10260
rect 33597 10251 33655 10257
rect 33597 10248 33609 10251
rect 33376 10220 33609 10248
rect 33376 10208 33382 10220
rect 33597 10217 33609 10220
rect 33643 10217 33655 10251
rect 33597 10211 33655 10217
rect 191282 10208 191288 10260
rect 191340 10248 191346 10260
rect 191837 10251 191895 10257
rect 191837 10248 191849 10251
rect 191340 10220 191849 10248
rect 191340 10208 191346 10220
rect 191837 10217 191849 10220
rect 191883 10217 191895 10251
rect 191837 10211 191895 10217
rect 192478 10208 192484 10260
rect 192536 10248 192542 10260
rect 193125 10251 193183 10257
rect 193125 10248 193137 10251
rect 192536 10220 193137 10248
rect 192536 10208 192542 10220
rect 193125 10217 193137 10220
rect 193171 10217 193183 10251
rect 193125 10211 193183 10217
rect 266906 10208 266912 10260
rect 266964 10248 266970 10260
rect 267737 10251 267795 10257
rect 267737 10248 267749 10251
rect 266964 10220 267749 10248
rect 266964 10208 266970 10220
rect 267737 10217 267749 10220
rect 267783 10217 267795 10251
rect 267737 10211 267795 10217
rect 268562 10208 268568 10260
rect 268620 10248 268626 10260
rect 269025 10251 269083 10257
rect 269025 10248 269037 10251
rect 268620 10220 269037 10248
rect 268620 10208 268626 10220
rect 269025 10217 269037 10220
rect 269071 10217 269083 10251
rect 269025 10211 269083 10217
rect 27522 10140 27528 10192
rect 27580 10180 27586 10192
rect 30285 10183 30343 10189
rect 30285 10180 30297 10183
rect 27580 10152 30297 10180
rect 27580 10140 27586 10152
rect 30285 10149 30297 10152
rect 30331 10149 30343 10183
rect 30285 10143 30343 10149
rect 31570 10140 31576 10192
rect 31628 10180 31634 10192
rect 32309 10183 32367 10189
rect 32309 10180 32321 10183
rect 31628 10152 32321 10180
rect 31628 10140 31634 10152
rect 32309 10149 32321 10152
rect 32355 10149 32367 10183
rect 32309 10143 32367 10149
rect 267093 10183 267151 10189
rect 267093 10149 267105 10183
rect 267139 10180 267151 10183
rect 268378 10180 268384 10192
rect 267139 10152 267734 10180
rect 267139 10149 267151 10152
rect 267093 10143 267151 10149
rect 267706 10124 267734 10152
rect 267844 10152 268384 10180
rect 157797 10115 157855 10121
rect 157797 10081 157809 10115
rect 157843 10112 157855 10115
rect 163590 10112 163596 10124
rect 157843 10084 163596 10112
rect 157843 10081 157855 10084
rect 157797 10075 157855 10081
rect 163590 10072 163596 10084
rect 163648 10072 163654 10124
rect 195882 10112 195888 10124
rect 192680 10084 195888 10112
rect 29454 10004 29460 10056
rect 29512 10044 29518 10056
rect 30469 10047 30527 10053
rect 30469 10044 30481 10047
rect 29512 10016 30481 10044
rect 29512 10004 29518 10016
rect 30469 10013 30481 10016
rect 30515 10013 30527 10047
rect 30469 10007 30527 10013
rect 30926 10004 30932 10056
rect 30984 10044 30990 10056
rect 31113 10047 31171 10053
rect 31113 10044 31125 10047
rect 30984 10016 31125 10044
rect 30984 10004 30990 10016
rect 31113 10013 31125 10016
rect 31159 10013 31171 10047
rect 31113 10007 31171 10013
rect 31573 10047 31631 10053
rect 31573 10013 31585 10047
rect 31619 10044 31631 10047
rect 32217 10047 32275 10053
rect 32217 10044 32229 10047
rect 31619 10016 32229 10044
rect 31619 10013 31631 10016
rect 31573 10007 31631 10013
rect 32217 10013 32229 10016
rect 32263 10013 32275 10047
rect 32217 10007 32275 10013
rect 33045 10047 33103 10053
rect 33045 10013 33057 10047
rect 33091 10044 33103 10047
rect 33410 10044 33416 10056
rect 33091 10016 33416 10044
rect 33091 10013 33103 10016
rect 33045 10007 33103 10013
rect 32232 9976 32260 10007
rect 33410 10004 33416 10016
rect 33468 10004 33474 10056
rect 33505 10047 33563 10053
rect 33505 10013 33517 10047
rect 33551 10044 33563 10047
rect 33686 10044 33692 10056
rect 33551 10016 33692 10044
rect 33551 10013 33563 10016
rect 33505 10007 33563 10013
rect 33520 9976 33548 10007
rect 33686 10004 33692 10016
rect 33744 10004 33750 10056
rect 140409 10047 140467 10053
rect 140409 10013 140421 10047
rect 140455 10044 140467 10047
rect 140682 10044 140688 10056
rect 140455 10016 140688 10044
rect 140455 10013 140467 10016
rect 140409 10007 140467 10013
rect 140682 10004 140688 10016
rect 140740 10004 140746 10056
rect 156049 10047 156107 10053
rect 156049 10013 156061 10047
rect 156095 10044 156107 10047
rect 156138 10044 156144 10056
rect 156095 10016 156144 10044
rect 156095 10013 156107 10016
rect 156049 10007 156107 10013
rect 156138 10004 156144 10016
rect 156196 10004 156202 10056
rect 192021 10047 192079 10053
rect 192021 10013 192033 10047
rect 192067 10044 192079 10047
rect 192570 10044 192576 10056
rect 192067 10016 192576 10044
rect 192067 10013 192079 10016
rect 192021 10007 192079 10013
rect 192570 10004 192576 10016
rect 192628 10004 192634 10056
rect 192680 10053 192708 10084
rect 195882 10072 195888 10084
rect 195940 10072 195946 10124
rect 267706 10084 267740 10124
rect 267734 10072 267740 10084
rect 267792 10072 267798 10124
rect 192665 10047 192723 10053
rect 192665 10013 192677 10047
rect 192711 10013 192723 10047
rect 192665 10007 192723 10013
rect 193309 10047 193367 10053
rect 193309 10013 193321 10047
rect 193355 10044 193367 10047
rect 194410 10044 194416 10056
rect 193355 10016 194416 10044
rect 193355 10013 193367 10016
rect 193309 10007 193367 10013
rect 194410 10004 194416 10016
rect 194468 10004 194474 10056
rect 267277 10047 267335 10053
rect 267277 10013 267289 10047
rect 267323 10044 267335 10047
rect 267844 10044 267872 10152
rect 268378 10140 268384 10152
rect 268436 10140 268442 10192
rect 268473 10183 268531 10189
rect 268473 10149 268485 10183
rect 268519 10180 268531 10183
rect 269482 10180 269488 10192
rect 268519 10152 269488 10180
rect 268519 10149 268531 10152
rect 268473 10143 268531 10149
rect 269482 10140 269488 10152
rect 269540 10140 269546 10192
rect 268838 10112 268844 10124
rect 267936 10084 268844 10112
rect 267936 10053 267964 10084
rect 268838 10072 268844 10084
rect 268896 10072 268902 10124
rect 267323 10016 267872 10044
rect 267921 10047 267979 10053
rect 267323 10013 267335 10016
rect 267277 10007 267335 10013
rect 267921 10013 267933 10047
rect 267967 10013 267979 10047
rect 267921 10007 267979 10013
rect 268102 10004 268108 10056
rect 268160 10044 268166 10056
rect 268381 10047 268439 10053
rect 268381 10044 268393 10047
rect 268160 10016 268393 10044
rect 268160 10004 268166 10016
rect 268381 10013 268393 10016
rect 268427 10044 268439 10047
rect 269022 10044 269028 10056
rect 268427 10016 269028 10044
rect 268427 10013 268439 10016
rect 268381 10007 268439 10013
rect 269022 10004 269028 10016
rect 269080 10004 269086 10056
rect 269206 10044 269212 10056
rect 269167 10016 269212 10044
rect 269206 10004 269212 10016
rect 269264 10004 269270 10056
rect 304442 10044 304448 10056
rect 304403 10016 304448 10044
rect 304442 10004 304448 10016
rect 304500 10004 304506 10056
rect 32232 9948 33548 9976
rect 252738 9936 252744 9988
rect 252796 9976 252802 9988
rect 304813 9979 304871 9985
rect 304813 9976 304825 9979
rect 252796 9948 304825 9976
rect 252796 9936 252802 9948
rect 304813 9945 304825 9948
rect 304859 9945 304871 9979
rect 304813 9939 304871 9945
rect 117406 9868 117412 9920
rect 117464 9908 117470 9920
rect 141697 9911 141755 9917
rect 141697 9908 141709 9911
rect 117464 9880 141709 9908
rect 117464 9868 117470 9880
rect 141697 9877 141709 9880
rect 141743 9877 141755 9911
rect 141697 9871 141755 9877
rect 192481 9911 192539 9917
rect 192481 9877 192493 9911
rect 192527 9908 192539 9911
rect 194318 9908 194324 9920
rect 192527 9880 194324 9908
rect 192527 9877 192539 9880
rect 192481 9871 192539 9877
rect 194318 9868 194324 9880
rect 194376 9868 194382 9920
rect 267734 9868 267740 9920
rect 267792 9908 267798 9920
rect 270954 9908 270960 9920
rect 267792 9880 270960 9908
rect 267792 9868 267798 9880
rect 270954 9868 270960 9880
rect 271012 9868 271018 9920
rect 1104 9818 305808 9840
rect 1104 9766 77148 9818
rect 77200 9766 77212 9818
rect 77264 9766 77276 9818
rect 77328 9766 77340 9818
rect 77392 9766 77404 9818
rect 77456 9766 153346 9818
rect 153398 9766 153410 9818
rect 153462 9766 153474 9818
rect 153526 9766 153538 9818
rect 153590 9766 153602 9818
rect 153654 9766 229544 9818
rect 229596 9766 229608 9818
rect 229660 9766 229672 9818
rect 229724 9766 229736 9818
rect 229788 9766 229800 9818
rect 229852 9766 305808 9818
rect 1104 9744 305808 9766
rect 31202 9596 31208 9648
rect 31260 9636 31266 9648
rect 32861 9639 32919 9645
rect 32861 9636 32873 9639
rect 31260 9608 32873 9636
rect 31260 9596 31266 9608
rect 32861 9605 32873 9608
rect 32907 9605 32919 9639
rect 140682 9636 140688 9648
rect 140643 9608 140688 9636
rect 32861 9599 32919 9605
rect 140682 9596 140688 9608
rect 140740 9596 140746 9648
rect 156138 9636 156144 9648
rect 156099 9608 156144 9636
rect 156138 9596 156144 9608
rect 156196 9596 156202 9648
rect 157889 9639 157947 9645
rect 157889 9605 157901 9639
rect 157935 9636 157947 9639
rect 158622 9636 158628 9648
rect 157935 9608 158628 9636
rect 157935 9605 157947 9608
rect 157889 9599 157947 9605
rect 158622 9596 158628 9608
rect 158680 9596 158686 9648
rect 190638 9596 190644 9648
rect 190696 9636 190702 9648
rect 193033 9639 193091 9645
rect 190696 9608 192984 9636
rect 190696 9596 190702 9608
rect 27338 9528 27344 9580
rect 27396 9568 27402 9580
rect 31297 9571 31355 9577
rect 31297 9568 31309 9571
rect 27396 9540 31309 9568
rect 27396 9528 27402 9540
rect 31297 9537 31309 9540
rect 31343 9537 31355 9571
rect 31297 9531 31355 9537
rect 32125 9571 32183 9577
rect 32125 9537 32137 9571
rect 32171 9568 32183 9571
rect 32769 9571 32827 9577
rect 32769 9568 32781 9571
rect 32171 9540 32781 9568
rect 32171 9537 32183 9540
rect 32125 9531 32183 9537
rect 32769 9537 32781 9540
rect 32815 9568 32827 9571
rect 33686 9568 33692 9580
rect 32815 9540 33692 9568
rect 32815 9537 32827 9540
rect 32769 9531 32827 9537
rect 33686 9528 33692 9540
rect 33744 9528 33750 9580
rect 192956 9577 192984 9608
rect 193033 9605 193045 9639
rect 193079 9636 193091 9639
rect 193306 9636 193312 9648
rect 193079 9608 193312 9636
rect 193079 9605 193091 9608
rect 193033 9599 193091 9605
rect 193306 9596 193312 9608
rect 193364 9596 193370 9648
rect 267921 9639 267979 9645
rect 267921 9605 267933 9639
rect 267967 9636 267979 9639
rect 269850 9636 269856 9648
rect 267967 9608 269856 9636
rect 267967 9605 267979 9608
rect 267921 9599 267979 9605
rect 269850 9596 269856 9608
rect 269908 9596 269914 9648
rect 192481 9571 192539 9577
rect 192481 9537 192493 9571
rect 192527 9537 192539 9571
rect 192481 9531 192539 9537
rect 192941 9571 192999 9577
rect 192941 9537 192953 9571
rect 192987 9568 192999 9571
rect 194134 9568 194140 9580
rect 192987 9540 194140 9568
rect 192987 9537 192999 9540
rect 192941 9531 192999 9537
rect 30558 9460 30564 9512
rect 30616 9500 30622 9512
rect 32217 9503 32275 9509
rect 32217 9500 32229 9503
rect 30616 9472 32229 9500
rect 30616 9460 30622 9472
rect 32217 9469 32229 9472
rect 32263 9469 32275 9503
rect 192496 9500 192524 9531
rect 194134 9528 194140 9540
rect 194192 9528 194198 9580
rect 267829 9571 267887 9577
rect 267829 9537 267841 9571
rect 267875 9568 267887 9571
rect 268102 9568 268108 9580
rect 267875 9540 268108 9568
rect 267875 9537 267887 9540
rect 267829 9531 267887 9537
rect 268102 9528 268108 9540
rect 268160 9528 268166 9580
rect 195974 9500 195980 9512
rect 192496 9472 195980 9500
rect 32217 9463 32275 9469
rect 195974 9460 195980 9472
rect 196032 9460 196038 9512
rect 29914 9392 29920 9444
rect 29972 9432 29978 9444
rect 31113 9435 31171 9441
rect 31113 9432 31125 9435
rect 29972 9404 31125 9432
rect 29972 9392 29978 9404
rect 31113 9401 31125 9404
rect 31159 9401 31171 9435
rect 31113 9395 31171 9401
rect 192297 9435 192355 9441
rect 192297 9401 192309 9435
rect 192343 9432 192355 9435
rect 194502 9432 194508 9444
rect 192343 9404 194508 9432
rect 192343 9401 192355 9404
rect 192297 9395 192355 9401
rect 194502 9392 194508 9404
rect 194560 9392 194566 9444
rect 104250 9324 104256 9376
rect 104308 9364 104314 9376
rect 141973 9367 142031 9373
rect 141973 9364 141985 9367
rect 104308 9336 141985 9364
rect 104308 9324 104314 9336
rect 141973 9333 141985 9336
rect 142019 9364 142031 9367
rect 148318 9364 148324 9376
rect 142019 9336 148324 9364
rect 142019 9333 142031 9336
rect 141973 9327 142031 9333
rect 148318 9324 148324 9336
rect 148376 9324 148382 9376
rect 1104 9274 305808 9296
rect 1104 9222 39049 9274
rect 39101 9222 39113 9274
rect 39165 9222 39177 9274
rect 39229 9222 39241 9274
rect 39293 9222 39305 9274
rect 39357 9222 115247 9274
rect 115299 9222 115311 9274
rect 115363 9222 115375 9274
rect 115427 9222 115439 9274
rect 115491 9222 115503 9274
rect 115555 9222 191445 9274
rect 191497 9222 191509 9274
rect 191561 9222 191573 9274
rect 191625 9222 191637 9274
rect 191689 9222 191701 9274
rect 191753 9222 267643 9274
rect 267695 9222 267707 9274
rect 267759 9222 267771 9274
rect 267823 9222 267835 9274
rect 267887 9222 267899 9274
rect 267951 9222 305808 9274
rect 1104 9200 305808 9222
rect 1104 8730 305808 8752
rect 1104 8678 77148 8730
rect 77200 8678 77212 8730
rect 77264 8678 77276 8730
rect 77328 8678 77340 8730
rect 77392 8678 77404 8730
rect 77456 8678 153346 8730
rect 153398 8678 153410 8730
rect 153462 8678 153474 8730
rect 153526 8678 153538 8730
rect 153590 8678 153602 8730
rect 153654 8678 229544 8730
rect 229596 8678 229608 8730
rect 229660 8678 229672 8730
rect 229724 8678 229736 8730
rect 229788 8678 229800 8730
rect 229852 8678 305808 8730
rect 1104 8656 305808 8678
rect 1581 8483 1639 8489
rect 1581 8449 1593 8483
rect 1627 8480 1639 8483
rect 1627 8452 1992 8480
rect 1627 8449 1639 8452
rect 1581 8443 1639 8449
rect 1394 8344 1400 8356
rect 1355 8316 1400 8344
rect 1394 8304 1400 8316
rect 1452 8304 1458 8356
rect 1964 8353 1992 8452
rect 1949 8347 2007 8353
rect 1949 8313 1961 8347
rect 1995 8344 2007 8347
rect 2317 8347 2375 8353
rect 2317 8344 2329 8347
rect 1995 8316 2329 8344
rect 1995 8313 2007 8316
rect 1949 8307 2007 8313
rect 2317 8313 2329 8316
rect 2363 8344 2375 8347
rect 2685 8347 2743 8353
rect 2685 8344 2697 8347
rect 2363 8316 2697 8344
rect 2363 8313 2375 8316
rect 2317 8307 2375 8313
rect 2685 8313 2697 8316
rect 2731 8344 2743 8347
rect 3053 8347 3111 8353
rect 3053 8344 3065 8347
rect 2731 8316 3065 8344
rect 2731 8313 2743 8316
rect 2685 8307 2743 8313
rect 3053 8313 3065 8316
rect 3099 8344 3111 8347
rect 187510 8344 187516 8356
rect 3099 8316 187516 8344
rect 3099 8313 3111 8316
rect 3053 8307 3111 8313
rect 187510 8304 187516 8316
rect 187568 8304 187574 8356
rect 1104 8186 305808 8208
rect 1104 8134 39049 8186
rect 39101 8134 39113 8186
rect 39165 8134 39177 8186
rect 39229 8134 39241 8186
rect 39293 8134 39305 8186
rect 39357 8134 115247 8186
rect 115299 8134 115311 8186
rect 115363 8134 115375 8186
rect 115427 8134 115439 8186
rect 115491 8134 115503 8186
rect 115555 8134 191445 8186
rect 191497 8134 191509 8186
rect 191561 8134 191573 8186
rect 191625 8134 191637 8186
rect 191689 8134 191701 8186
rect 191753 8134 267643 8186
rect 267695 8134 267707 8186
rect 267759 8134 267771 8186
rect 267823 8134 267835 8186
rect 267887 8134 267899 8186
rect 267951 8134 305808 8186
rect 1104 8112 305808 8134
rect 1104 7642 305808 7664
rect 1104 7590 77148 7642
rect 77200 7590 77212 7642
rect 77264 7590 77276 7642
rect 77328 7590 77340 7642
rect 77392 7590 77404 7642
rect 77456 7590 153346 7642
rect 153398 7590 153410 7642
rect 153462 7590 153474 7642
rect 153526 7590 153538 7642
rect 153590 7590 153602 7642
rect 153654 7590 229544 7642
rect 229596 7590 229608 7642
rect 229660 7590 229672 7642
rect 229724 7590 229736 7642
rect 229788 7590 229800 7642
rect 229852 7590 305808 7642
rect 1104 7568 305808 7590
rect 1104 7098 305808 7120
rect 1104 7046 39049 7098
rect 39101 7046 39113 7098
rect 39165 7046 39177 7098
rect 39229 7046 39241 7098
rect 39293 7046 39305 7098
rect 39357 7046 115247 7098
rect 115299 7046 115311 7098
rect 115363 7046 115375 7098
rect 115427 7046 115439 7098
rect 115491 7046 115503 7098
rect 115555 7046 191445 7098
rect 191497 7046 191509 7098
rect 191561 7046 191573 7098
rect 191625 7046 191637 7098
rect 191689 7046 191701 7098
rect 191753 7046 267643 7098
rect 267695 7046 267707 7098
rect 267759 7046 267771 7098
rect 267823 7046 267835 7098
rect 267887 7046 267899 7098
rect 267951 7046 305808 7098
rect 1104 7024 305808 7046
rect 1104 6554 305808 6576
rect 1104 6502 77148 6554
rect 77200 6502 77212 6554
rect 77264 6502 77276 6554
rect 77328 6502 77340 6554
rect 77392 6502 77404 6554
rect 77456 6502 153346 6554
rect 153398 6502 153410 6554
rect 153462 6502 153474 6554
rect 153526 6502 153538 6554
rect 153590 6502 153602 6554
rect 153654 6502 229544 6554
rect 229596 6502 229608 6554
rect 229660 6502 229672 6554
rect 229724 6502 229736 6554
rect 229788 6502 229800 6554
rect 229852 6502 305808 6554
rect 1104 6480 305808 6502
rect 303982 6304 303988 6316
rect 303943 6276 303988 6304
rect 303982 6264 303988 6276
rect 304040 6264 304046 6316
rect 249058 6196 249064 6248
rect 249116 6236 249122 6248
rect 304261 6239 304319 6245
rect 304261 6236 304273 6239
rect 249116 6208 304273 6236
rect 249116 6196 249122 6208
rect 304261 6205 304273 6208
rect 304307 6205 304319 6239
rect 304261 6199 304319 6205
rect 1104 6010 305808 6032
rect 1104 5958 39049 6010
rect 39101 5958 39113 6010
rect 39165 5958 39177 6010
rect 39229 5958 39241 6010
rect 39293 5958 39305 6010
rect 39357 5958 115247 6010
rect 115299 5958 115311 6010
rect 115363 5958 115375 6010
rect 115427 5958 115439 6010
rect 115491 5958 115503 6010
rect 115555 5958 191445 6010
rect 191497 5958 191509 6010
rect 191561 5958 191573 6010
rect 191625 5958 191637 6010
rect 191689 5958 191701 6010
rect 191753 5958 267643 6010
rect 267695 5958 267707 6010
rect 267759 5958 267771 6010
rect 267823 5958 267835 6010
rect 267887 5958 267899 6010
rect 267951 5958 305808 6010
rect 1104 5936 305808 5958
rect 1104 5466 305808 5488
rect 1104 5414 77148 5466
rect 77200 5414 77212 5466
rect 77264 5414 77276 5466
rect 77328 5414 77340 5466
rect 77392 5414 77404 5466
rect 77456 5414 153346 5466
rect 153398 5414 153410 5466
rect 153462 5414 153474 5466
rect 153526 5414 153538 5466
rect 153590 5414 153602 5466
rect 153654 5414 229544 5466
rect 229596 5414 229608 5466
rect 229660 5414 229672 5466
rect 229724 5414 229736 5466
rect 229788 5414 229800 5466
rect 229852 5414 305808 5466
rect 1104 5392 305808 5414
rect 1104 4922 305808 4944
rect 1104 4870 39049 4922
rect 39101 4870 39113 4922
rect 39165 4870 39177 4922
rect 39229 4870 39241 4922
rect 39293 4870 39305 4922
rect 39357 4870 115247 4922
rect 115299 4870 115311 4922
rect 115363 4870 115375 4922
rect 115427 4870 115439 4922
rect 115491 4870 115503 4922
rect 115555 4870 191445 4922
rect 191497 4870 191509 4922
rect 191561 4870 191573 4922
rect 191625 4870 191637 4922
rect 191689 4870 191701 4922
rect 191753 4870 267643 4922
rect 267695 4870 267707 4922
rect 267759 4870 267771 4922
rect 267823 4870 267835 4922
rect 267887 4870 267899 4922
rect 267951 4870 305808 4922
rect 1104 4848 305808 4870
rect 1104 4378 305808 4400
rect 1104 4326 77148 4378
rect 77200 4326 77212 4378
rect 77264 4326 77276 4378
rect 77328 4326 77340 4378
rect 77392 4326 77404 4378
rect 77456 4326 153346 4378
rect 153398 4326 153410 4378
rect 153462 4326 153474 4378
rect 153526 4326 153538 4378
rect 153590 4326 153602 4378
rect 153654 4326 229544 4378
rect 229596 4326 229608 4378
rect 229660 4326 229672 4378
rect 229724 4326 229736 4378
rect 229788 4326 229800 4378
rect 229852 4326 305808 4378
rect 1104 4304 305808 4326
rect 1104 3834 305808 3856
rect 1104 3782 39049 3834
rect 39101 3782 39113 3834
rect 39165 3782 39177 3834
rect 39229 3782 39241 3834
rect 39293 3782 39305 3834
rect 39357 3782 115247 3834
rect 115299 3782 115311 3834
rect 115363 3782 115375 3834
rect 115427 3782 115439 3834
rect 115491 3782 115503 3834
rect 115555 3782 191445 3834
rect 191497 3782 191509 3834
rect 191561 3782 191573 3834
rect 191625 3782 191637 3834
rect 191689 3782 191701 3834
rect 191753 3782 267643 3834
rect 267695 3782 267707 3834
rect 267759 3782 267771 3834
rect 267823 3782 267835 3834
rect 267887 3782 267899 3834
rect 267951 3782 305808 3834
rect 1104 3760 305808 3782
rect 1104 3290 305808 3312
rect 1104 3238 77148 3290
rect 77200 3238 77212 3290
rect 77264 3238 77276 3290
rect 77328 3238 77340 3290
rect 77392 3238 77404 3290
rect 77456 3238 153346 3290
rect 153398 3238 153410 3290
rect 153462 3238 153474 3290
rect 153526 3238 153538 3290
rect 153590 3238 153602 3290
rect 153654 3238 229544 3290
rect 229596 3238 229608 3290
rect 229660 3238 229672 3290
rect 229724 3238 229736 3290
rect 229788 3238 229800 3290
rect 229852 3238 305808 3290
rect 1104 3216 305808 3238
rect 1104 2746 305808 2768
rect 1104 2694 39049 2746
rect 39101 2694 39113 2746
rect 39165 2694 39177 2746
rect 39229 2694 39241 2746
rect 39293 2694 39305 2746
rect 39357 2694 115247 2746
rect 115299 2694 115311 2746
rect 115363 2694 115375 2746
rect 115427 2694 115439 2746
rect 115491 2694 115503 2746
rect 115555 2694 191445 2746
rect 191497 2694 191509 2746
rect 191561 2694 191573 2746
rect 191625 2694 191637 2746
rect 191689 2694 191701 2746
rect 191753 2694 267643 2746
rect 267695 2694 267707 2746
rect 267759 2694 267771 2746
rect 267823 2694 267835 2746
rect 267887 2694 267899 2746
rect 267951 2694 305808 2746
rect 1104 2672 305808 2694
rect 149422 2592 149428 2644
rect 149480 2632 149486 2644
rect 302234 2632 302240 2644
rect 149480 2604 302240 2632
rect 149480 2592 149486 2604
rect 302234 2592 302240 2604
rect 302292 2592 302298 2644
rect 1104 2202 305808 2224
rect 1104 2150 77148 2202
rect 77200 2150 77212 2202
rect 77264 2150 77276 2202
rect 77328 2150 77340 2202
rect 77392 2150 77404 2202
rect 77456 2150 153346 2202
rect 153398 2150 153410 2202
rect 153462 2150 153474 2202
rect 153526 2150 153538 2202
rect 153590 2150 153602 2202
rect 153654 2150 229544 2202
rect 229596 2150 229608 2202
rect 229660 2150 229672 2202
rect 229724 2150 229736 2202
rect 229788 2150 229800 2202
rect 229852 2150 305808 2202
rect 1104 2128 305808 2150
<< via1 >>
rect 29000 13744 29052 13796
rect 32956 13744 33008 13796
rect 46204 13744 46256 13796
rect 63408 13744 63460 13796
rect 69296 13744 69348 13796
rect 75368 13744 75420 13796
rect 76012 13744 76064 13796
rect 90640 13744 90692 13796
rect 102416 13744 102468 13796
rect 113824 13744 113876 13796
rect 125508 13744 125560 13796
rect 131856 13744 131908 13796
rect 161664 13744 161716 13796
rect 166080 13744 166132 13796
rect 167368 13744 167420 13796
rect 174176 13744 174228 13796
rect 177764 13744 177816 13796
rect 181904 13744 181956 13796
rect 189908 13812 189960 13864
rect 189356 13744 189408 13796
rect 193220 13744 193272 13796
rect 195980 13744 196032 13796
rect 302792 13744 302844 13796
rect 27160 13676 27212 13728
rect 36544 13676 36596 13728
rect 42524 13676 42576 13728
rect 47860 13676 47912 13728
rect 51632 13676 51684 13728
rect 54116 13676 54168 13728
rect 66168 13676 66220 13728
rect 72424 13676 72476 13728
rect 73896 13676 73948 13728
rect 76380 13676 76432 13728
rect 83096 13676 83148 13728
rect 86408 13676 86460 13728
rect 91836 13676 91888 13728
rect 101956 13676 102008 13728
rect 114652 13676 114704 13728
rect 127440 13676 127492 13728
rect 127532 13676 127584 13728
rect 129740 13676 129792 13728
rect 133604 13676 133656 13728
rect 136824 13676 136876 13728
rect 148140 13676 148192 13728
rect 150440 13676 150492 13728
rect 157156 13676 157208 13728
rect 301412 13676 301464 13728
rect 39049 13574 39101 13626
rect 39113 13574 39165 13626
rect 39177 13574 39229 13626
rect 39241 13574 39293 13626
rect 39305 13574 39357 13626
rect 115247 13574 115299 13626
rect 115311 13574 115363 13626
rect 115375 13574 115427 13626
rect 115439 13574 115491 13626
rect 115503 13574 115555 13626
rect 191445 13574 191497 13626
rect 191509 13574 191561 13626
rect 191573 13574 191625 13626
rect 191637 13574 191689 13626
rect 191701 13574 191753 13626
rect 267643 13574 267695 13626
rect 267707 13574 267759 13626
rect 267771 13574 267823 13626
rect 267835 13574 267887 13626
rect 267899 13574 267951 13626
rect 1584 13515 1636 13524
rect 1584 13481 1593 13515
rect 1593 13481 1627 13515
rect 1627 13481 1636 13515
rect 1584 13472 1636 13481
rect 4620 13515 4672 13524
rect 4620 13481 4629 13515
rect 4629 13481 4663 13515
rect 4663 13481 4672 13515
rect 4620 13472 4672 13481
rect 7656 13515 7708 13524
rect 7656 13481 7665 13515
rect 7665 13481 7699 13515
rect 7699 13481 7708 13515
rect 7656 13472 7708 13481
rect 10784 13515 10836 13524
rect 10784 13481 10793 13515
rect 10793 13481 10827 13515
rect 10827 13481 10836 13515
rect 10784 13472 10836 13481
rect 13820 13472 13872 13524
rect 16856 13515 16908 13524
rect 16856 13481 16865 13515
rect 16865 13481 16899 13515
rect 16899 13481 16908 13515
rect 16856 13472 16908 13481
rect 19984 13515 20036 13524
rect 19984 13481 19993 13515
rect 19993 13481 20027 13515
rect 20027 13481 20036 13515
rect 19984 13472 20036 13481
rect 23020 13515 23072 13524
rect 23020 13481 23029 13515
rect 23029 13481 23063 13515
rect 23063 13481 23072 13515
rect 23020 13472 23072 13481
rect 27620 13472 27672 13524
rect 27712 13472 27764 13524
rect 30472 13472 30524 13524
rect 36544 13472 36596 13524
rect 46204 13472 46256 13524
rect 47584 13515 47636 13524
rect 47584 13481 47593 13515
rect 47593 13481 47627 13515
rect 47627 13481 47636 13515
rect 47584 13472 47636 13481
rect 50528 13472 50580 13524
rect 53012 13472 53064 13524
rect 55588 13472 55640 13524
rect 57888 13472 57940 13524
rect 61752 13472 61804 13524
rect 63408 13472 63460 13524
rect 142896 13515 142948 13524
rect 27160 13404 27212 13456
rect 44180 13404 44232 13456
rect 4804 13311 4856 13320
rect 4804 13277 4813 13311
rect 4813 13277 4847 13311
rect 4847 13277 4856 13311
rect 4804 13268 4856 13277
rect 14280 13311 14332 13320
rect 14280 13277 14289 13311
rect 14289 13277 14323 13311
rect 14323 13277 14332 13311
rect 14280 13268 14332 13277
rect 17040 13311 17092 13320
rect 17040 13277 17049 13311
rect 17049 13277 17083 13311
rect 17083 13277 17092 13311
rect 17040 13268 17092 13277
rect 20168 13311 20220 13320
rect 20168 13277 20177 13311
rect 20177 13277 20211 13311
rect 20211 13277 20220 13311
rect 20168 13268 20220 13277
rect 23204 13311 23256 13320
rect 23204 13277 23213 13311
rect 23213 13277 23247 13311
rect 23247 13277 23256 13311
rect 23204 13268 23256 13277
rect 26976 13336 27028 13388
rect 29828 13311 29880 13320
rect 29828 13277 29837 13311
rect 29837 13277 29871 13311
rect 29871 13277 29880 13311
rect 29828 13268 29880 13277
rect 32404 13311 32456 13320
rect 32404 13277 32413 13311
rect 32413 13277 32447 13311
rect 32447 13277 32456 13311
rect 32404 13268 32456 13277
rect 33784 13268 33836 13320
rect 44364 13404 44416 13456
rect 45560 13379 45612 13388
rect 45560 13345 45569 13379
rect 45569 13345 45603 13379
rect 45603 13345 45612 13379
rect 51632 13379 51684 13388
rect 45560 13336 45612 13345
rect 51632 13345 51641 13379
rect 51641 13345 51675 13379
rect 51675 13345 51684 13379
rect 51632 13336 51684 13345
rect 59820 13404 59872 13456
rect 63040 13447 63092 13456
rect 63040 13413 63049 13447
rect 63049 13413 63083 13447
rect 63083 13413 63092 13447
rect 63040 13404 63092 13413
rect 75368 13447 75420 13456
rect 72700 13379 72752 13388
rect 27528 13243 27580 13252
rect 27252 13132 27304 13184
rect 27528 13209 27537 13243
rect 27537 13209 27571 13243
rect 27571 13209 27580 13243
rect 27528 13200 27580 13209
rect 27712 13132 27764 13184
rect 30196 13200 30248 13252
rect 32680 13243 32732 13252
rect 30472 13132 30524 13184
rect 32680 13209 32689 13243
rect 32689 13209 32723 13243
rect 32723 13209 32732 13243
rect 32680 13200 32732 13209
rect 34520 13200 34572 13252
rect 35992 13200 36044 13252
rect 33600 13132 33652 13184
rect 34152 13175 34204 13184
rect 34152 13141 34161 13175
rect 34161 13141 34195 13175
rect 34195 13141 34204 13175
rect 34152 13132 34204 13141
rect 34336 13132 34388 13184
rect 37464 13132 37516 13184
rect 38936 13268 38988 13320
rect 37832 13243 37884 13252
rect 37832 13209 37841 13243
rect 37841 13209 37875 13243
rect 37875 13209 37884 13243
rect 37832 13200 37884 13209
rect 42524 13311 42576 13320
rect 39304 13175 39356 13184
rect 39304 13141 39313 13175
rect 39313 13141 39347 13175
rect 39347 13141 39356 13175
rect 39304 13132 39356 13141
rect 39948 13132 40000 13184
rect 42524 13277 42533 13311
rect 42533 13277 42567 13311
rect 42567 13277 42576 13311
rect 42524 13268 42576 13277
rect 44272 13268 44324 13320
rect 51356 13311 51408 13320
rect 40408 13243 40460 13252
rect 40408 13209 40417 13243
rect 40417 13209 40451 13243
rect 40451 13209 40460 13243
rect 40408 13200 40460 13209
rect 41420 13200 41472 13252
rect 42892 13200 42944 13252
rect 43260 13200 43312 13252
rect 42432 13132 42484 13184
rect 45008 13175 45060 13184
rect 45008 13141 45017 13175
rect 45017 13141 45051 13175
rect 45051 13141 45060 13175
rect 45008 13132 45060 13141
rect 45376 13175 45428 13184
rect 45376 13141 45385 13175
rect 45385 13141 45419 13175
rect 45419 13141 45428 13175
rect 45376 13132 45428 13141
rect 51356 13277 51365 13311
rect 51365 13277 51399 13311
rect 51399 13277 51408 13311
rect 51356 13268 51408 13277
rect 47860 13200 47912 13252
rect 54392 13268 54444 13320
rect 54760 13268 54812 13320
rect 55588 13311 55640 13320
rect 55588 13277 55597 13311
rect 55597 13277 55631 13311
rect 55631 13277 55640 13311
rect 55588 13268 55640 13277
rect 57888 13311 57940 13320
rect 57888 13277 57897 13311
rect 57897 13277 57931 13311
rect 57931 13277 57940 13311
rect 57888 13268 57940 13277
rect 60648 13311 60700 13320
rect 60648 13277 60657 13311
rect 60657 13277 60691 13311
rect 60691 13277 60700 13311
rect 60648 13268 60700 13277
rect 53288 13243 53340 13252
rect 53288 13209 53297 13243
rect 53297 13209 53331 13243
rect 53331 13209 53340 13243
rect 53288 13200 53340 13209
rect 55864 13243 55916 13252
rect 54668 13132 54720 13184
rect 55864 13209 55873 13243
rect 55873 13209 55907 13243
rect 55907 13209 55916 13243
rect 55864 13200 55916 13209
rect 56600 13200 56652 13252
rect 57336 13175 57388 13184
rect 57336 13141 57345 13175
rect 57345 13141 57379 13175
rect 57379 13141 57388 13175
rect 57336 13132 57388 13141
rect 57704 13200 57756 13252
rect 58624 13200 58676 13252
rect 61476 13200 61528 13252
rect 59636 13175 59688 13184
rect 59636 13141 59645 13175
rect 59645 13141 59679 13175
rect 59679 13141 59688 13175
rect 66168 13311 66220 13320
rect 66168 13277 66177 13311
rect 66177 13277 66211 13311
rect 66211 13277 66220 13311
rect 66168 13268 66220 13277
rect 69296 13311 69348 13320
rect 69296 13277 69305 13311
rect 69305 13277 69339 13311
rect 69339 13277 69348 13311
rect 69296 13268 69348 13277
rect 72700 13345 72709 13379
rect 72709 13345 72743 13379
rect 72743 13345 72752 13379
rect 72700 13336 72752 13345
rect 75368 13413 75377 13447
rect 75377 13413 75411 13447
rect 75411 13413 75420 13447
rect 75368 13404 75420 13413
rect 75644 13404 75696 13456
rect 80244 13379 80296 13388
rect 80244 13345 80253 13379
rect 80253 13345 80287 13379
rect 80287 13345 80296 13379
rect 80244 13336 80296 13345
rect 81624 13379 81676 13388
rect 81624 13345 81633 13379
rect 81633 13345 81667 13379
rect 81667 13345 81676 13379
rect 93860 13404 93912 13456
rect 81624 13336 81676 13345
rect 61752 13200 61804 13252
rect 59636 13132 59688 13141
rect 61660 13132 61712 13184
rect 65892 13132 65944 13184
rect 65984 13175 66036 13184
rect 65984 13141 65993 13175
rect 65993 13141 66027 13175
rect 66027 13141 66036 13175
rect 69112 13175 69164 13184
rect 65984 13132 66036 13141
rect 69112 13141 69121 13175
rect 69121 13141 69155 13175
rect 69155 13141 69164 13175
rect 69112 13132 69164 13141
rect 72332 13132 72384 13184
rect 72424 13175 72476 13184
rect 72424 13141 72433 13175
rect 72433 13141 72467 13175
rect 72467 13141 72476 13175
rect 73896 13243 73948 13252
rect 73896 13209 73905 13243
rect 73905 13209 73939 13243
rect 73939 13209 73948 13243
rect 73896 13200 73948 13209
rect 75184 13200 75236 13252
rect 78404 13268 78456 13320
rect 81440 13268 81492 13320
rect 83096 13311 83148 13320
rect 76472 13243 76524 13252
rect 76472 13209 76481 13243
rect 76481 13209 76515 13243
rect 76515 13209 76524 13243
rect 76472 13200 76524 13209
rect 78772 13243 78824 13252
rect 72424 13132 72476 13141
rect 77944 13175 77996 13184
rect 77944 13141 77953 13175
rect 77953 13141 77987 13175
rect 77987 13141 77996 13175
rect 78772 13209 78781 13243
rect 78781 13209 78815 13243
rect 78815 13209 78824 13243
rect 78772 13200 78824 13209
rect 79324 13200 79376 13252
rect 80060 13200 80112 13252
rect 83096 13277 83105 13311
rect 83105 13277 83139 13311
rect 83139 13277 83148 13311
rect 83096 13268 83148 13277
rect 83924 13311 83976 13320
rect 83924 13277 83933 13311
rect 83933 13277 83967 13311
rect 83967 13277 83976 13311
rect 83924 13268 83976 13277
rect 77944 13132 77996 13141
rect 80796 13132 80848 13184
rect 81440 13175 81492 13184
rect 81440 13141 81449 13175
rect 81449 13141 81483 13175
rect 81483 13141 81492 13175
rect 81440 13132 81492 13141
rect 83832 13200 83884 13252
rect 84476 13200 84528 13252
rect 85488 13200 85540 13252
rect 82912 13175 82964 13184
rect 82912 13141 82921 13175
rect 82921 13141 82955 13175
rect 82955 13141 82964 13175
rect 82912 13132 82964 13141
rect 83924 13132 83976 13184
rect 86040 13132 86092 13184
rect 87880 13268 87932 13320
rect 86776 13243 86828 13252
rect 86776 13209 86785 13243
rect 86785 13209 86819 13243
rect 86819 13209 86828 13243
rect 86776 13200 86828 13209
rect 88248 13175 88300 13184
rect 88248 13141 88257 13175
rect 88257 13141 88291 13175
rect 88291 13141 88300 13175
rect 88248 13132 88300 13141
rect 89076 13243 89128 13252
rect 89076 13209 89085 13243
rect 89085 13209 89119 13243
rect 89119 13209 89128 13243
rect 89076 13200 89128 13209
rect 89536 13200 89588 13252
rect 91652 13200 91704 13252
rect 91836 13243 91888 13252
rect 91836 13209 91845 13243
rect 91845 13209 91879 13243
rect 91879 13209 91888 13243
rect 91836 13200 91888 13209
rect 92020 13243 92072 13252
rect 92020 13209 92029 13243
rect 92029 13209 92063 13243
rect 92063 13209 92072 13243
rect 92020 13200 92072 13209
rect 90548 13175 90600 13184
rect 90548 13141 90557 13175
rect 90557 13141 90591 13175
rect 90591 13141 90600 13175
rect 99104 13336 99156 13388
rect 100760 13404 100812 13456
rect 109040 13404 109092 13456
rect 111708 13404 111760 13456
rect 118884 13404 118936 13456
rect 121276 13447 121328 13456
rect 118240 13336 118292 13388
rect 121276 13413 121285 13447
rect 121285 13413 121319 13447
rect 121319 13413 121328 13447
rect 121276 13404 121328 13413
rect 124128 13447 124180 13456
rect 124128 13413 124137 13447
rect 124137 13413 124171 13447
rect 124171 13413 124180 13447
rect 124128 13404 124180 13413
rect 127532 13404 127584 13456
rect 136640 13447 136692 13456
rect 136640 13413 136649 13447
rect 136649 13413 136683 13447
rect 136683 13413 136692 13447
rect 136640 13404 136692 13413
rect 139584 13404 139636 13456
rect 142896 13481 142905 13515
rect 142905 13481 142939 13515
rect 142939 13481 142948 13515
rect 142896 13472 142948 13481
rect 145748 13472 145800 13524
rect 148140 13472 148192 13524
rect 150808 13472 150860 13524
rect 96712 13175 96764 13184
rect 90548 13132 90600 13141
rect 96712 13141 96721 13175
rect 96721 13141 96755 13175
rect 96755 13141 96764 13175
rect 96712 13132 96764 13141
rect 97540 13175 97592 13184
rect 97540 13141 97549 13175
rect 97549 13141 97583 13175
rect 97583 13141 97592 13175
rect 97540 13132 97592 13141
rect 98000 13200 98052 13252
rect 99196 13200 99248 13252
rect 101404 13268 101456 13320
rect 99656 13243 99708 13252
rect 99656 13209 99665 13243
rect 99665 13209 99699 13243
rect 99699 13209 99708 13243
rect 99656 13200 99708 13209
rect 100944 13200 100996 13252
rect 101036 13132 101088 13184
rect 103336 13268 103388 13320
rect 104256 13311 104308 13320
rect 102232 13243 102284 13252
rect 102232 13209 102241 13243
rect 102241 13209 102275 13243
rect 102275 13209 102284 13243
rect 102232 13200 102284 13209
rect 104256 13277 104265 13311
rect 104265 13277 104299 13311
rect 104299 13277 104308 13311
rect 104256 13268 104308 13277
rect 109592 13311 109644 13320
rect 109592 13277 109601 13311
rect 109601 13277 109635 13311
rect 109635 13277 109644 13311
rect 109592 13268 109644 13277
rect 111432 13311 111484 13320
rect 111432 13277 111441 13311
rect 111441 13277 111475 13311
rect 111475 13277 111484 13311
rect 111432 13268 111484 13277
rect 114836 13311 114888 13320
rect 114836 13277 114845 13311
rect 114845 13277 114879 13311
rect 114879 13277 114888 13311
rect 114836 13268 114888 13277
rect 117412 13311 117464 13320
rect 117412 13277 117421 13311
rect 117421 13277 117455 13311
rect 117455 13277 117464 13311
rect 117412 13268 117464 13277
rect 118792 13268 118844 13320
rect 130292 13379 130344 13388
rect 130292 13345 130301 13379
rect 130301 13345 130335 13379
rect 130335 13345 130344 13379
rect 130292 13336 130344 13345
rect 142068 13336 142120 13388
rect 104072 13200 104124 13252
rect 104992 13200 105044 13252
rect 112536 13243 112588 13252
rect 112536 13209 112545 13243
rect 112545 13209 112579 13243
rect 112579 13209 112588 13243
rect 112536 13200 112588 13209
rect 114192 13200 114244 13252
rect 115112 13243 115164 13252
rect 115112 13209 115121 13243
rect 115121 13209 115155 13243
rect 115155 13209 115164 13243
rect 115112 13200 115164 13209
rect 116952 13200 117004 13252
rect 117688 13243 117740 13252
rect 117688 13209 117697 13243
rect 117697 13209 117731 13243
rect 117731 13209 117740 13243
rect 117688 13200 117740 13209
rect 103704 13175 103756 13184
rect 103704 13141 103713 13175
rect 103713 13141 103747 13175
rect 103747 13141 103756 13175
rect 103704 13132 103756 13141
rect 104440 13132 104492 13184
rect 104624 13132 104676 13184
rect 109592 13132 109644 13184
rect 114560 13132 114612 13184
rect 114928 13132 114980 13184
rect 115756 13132 115808 13184
rect 118056 13132 118108 13184
rect 127532 13311 127584 13320
rect 127532 13277 127541 13311
rect 127541 13277 127575 13311
rect 127575 13277 127584 13311
rect 127532 13268 127584 13277
rect 129372 13268 129424 13320
rect 136824 13311 136876 13320
rect 136824 13277 136833 13311
rect 136833 13277 136867 13311
rect 136867 13277 136876 13311
rect 136824 13268 136876 13277
rect 143080 13311 143132 13320
rect 125508 13243 125560 13252
rect 125508 13209 125517 13243
rect 125517 13209 125551 13243
rect 125551 13209 125560 13243
rect 125508 13200 125560 13209
rect 127808 13243 127860 13252
rect 127808 13209 127817 13243
rect 127817 13209 127851 13243
rect 127851 13209 127860 13243
rect 127808 13200 127860 13209
rect 119712 13175 119764 13184
rect 119712 13141 119721 13175
rect 119721 13141 119755 13175
rect 119755 13141 119764 13175
rect 119712 13132 119764 13141
rect 126152 13175 126204 13184
rect 126152 13141 126161 13175
rect 126161 13141 126195 13175
rect 126195 13141 126204 13175
rect 126152 13132 126204 13141
rect 126520 13175 126572 13184
rect 126520 13141 126529 13175
rect 126529 13141 126563 13175
rect 126563 13141 126572 13175
rect 126520 13132 126572 13141
rect 128084 13132 128136 13184
rect 131212 13200 131264 13252
rect 132868 13243 132920 13252
rect 132868 13209 132877 13243
rect 132877 13209 132911 13243
rect 132911 13209 132920 13243
rect 132868 13200 132920 13209
rect 133328 13200 133380 13252
rect 143080 13277 143089 13311
rect 143089 13277 143123 13311
rect 143123 13277 143132 13311
rect 143080 13268 143132 13277
rect 145748 13311 145800 13320
rect 145748 13277 145757 13311
rect 145757 13277 145791 13311
rect 145791 13277 145800 13311
rect 145748 13268 145800 13277
rect 157248 13472 157300 13524
rect 157984 13472 158036 13524
rect 159456 13472 159508 13524
rect 161572 13472 161624 13524
rect 162676 13472 162728 13524
rect 163504 13472 163556 13524
rect 176384 13472 176436 13524
rect 182732 13515 182784 13524
rect 154948 13404 155000 13456
rect 166448 13404 166500 13456
rect 170404 13447 170456 13456
rect 160928 13379 160980 13388
rect 160928 13345 160937 13379
rect 160937 13345 160971 13379
rect 160971 13345 160980 13379
rect 160928 13336 160980 13345
rect 165252 13336 165304 13388
rect 129188 13132 129240 13184
rect 131580 13132 131632 13184
rect 133696 13132 133748 13184
rect 134156 13132 134208 13184
rect 145932 13200 145984 13252
rect 146024 13243 146076 13252
rect 146024 13209 146033 13243
rect 146033 13209 146067 13243
rect 146067 13209 146076 13243
rect 146024 13200 146076 13209
rect 147588 13200 147640 13252
rect 145840 13132 145892 13184
rect 147496 13175 147548 13184
rect 147496 13141 147505 13175
rect 147505 13141 147539 13175
rect 147539 13141 147548 13175
rect 147496 13132 147548 13141
rect 155224 13268 155276 13320
rect 155868 13268 155920 13320
rect 156420 13311 156472 13320
rect 156420 13277 156429 13311
rect 156429 13277 156463 13311
rect 156463 13277 156472 13311
rect 156420 13268 156472 13277
rect 157800 13311 157852 13320
rect 157800 13277 157809 13311
rect 157809 13277 157843 13311
rect 157843 13277 157852 13311
rect 157800 13268 157852 13277
rect 158628 13311 158680 13320
rect 158628 13277 158637 13311
rect 158637 13277 158671 13311
rect 158671 13277 158680 13311
rect 158628 13268 158680 13277
rect 162676 13268 162728 13320
rect 163504 13311 163556 13320
rect 149244 13132 149296 13184
rect 150440 13200 150492 13252
rect 151084 13200 151136 13252
rect 152464 13200 152516 13252
rect 153752 13243 153804 13252
rect 152648 13175 152700 13184
rect 152648 13141 152657 13175
rect 152657 13141 152691 13175
rect 152691 13141 152700 13175
rect 153752 13209 153761 13243
rect 153761 13209 153795 13243
rect 153795 13209 153804 13243
rect 153752 13200 153804 13209
rect 154212 13200 154264 13252
rect 156604 13200 156656 13252
rect 158904 13243 158956 13252
rect 155224 13175 155276 13184
rect 152648 13132 152700 13141
rect 155224 13141 155233 13175
rect 155233 13141 155267 13175
rect 155267 13141 155276 13175
rect 155224 13132 155276 13141
rect 158904 13209 158913 13243
rect 158913 13209 158947 13243
rect 158947 13209 158956 13243
rect 158904 13200 158956 13209
rect 161204 13243 161256 13252
rect 159548 13132 159600 13184
rect 160376 13175 160428 13184
rect 160376 13141 160385 13175
rect 160385 13141 160419 13175
rect 160419 13141 160428 13175
rect 160376 13132 160428 13141
rect 161204 13209 161213 13243
rect 161213 13209 161247 13243
rect 161247 13209 161256 13243
rect 161204 13200 161256 13209
rect 162768 13200 162820 13252
rect 162032 13132 162084 13184
rect 162492 13132 162544 13184
rect 163504 13277 163513 13311
rect 163513 13277 163547 13311
rect 163547 13277 163556 13311
rect 163504 13268 163556 13277
rect 164884 13268 164936 13320
rect 170404 13413 170413 13447
rect 170413 13413 170447 13447
rect 170447 13413 170456 13447
rect 170404 13404 170456 13413
rect 173072 13447 173124 13456
rect 173072 13413 173081 13447
rect 173081 13413 173115 13447
rect 173115 13413 173124 13447
rect 173072 13404 173124 13413
rect 173808 13447 173860 13456
rect 173808 13413 173817 13447
rect 173817 13413 173851 13447
rect 173851 13413 173860 13447
rect 173808 13404 173860 13413
rect 175924 13404 175976 13456
rect 176016 13404 176068 13456
rect 177764 13404 177816 13456
rect 180432 13404 180484 13456
rect 163780 13243 163832 13252
rect 163780 13209 163789 13243
rect 163789 13209 163823 13243
rect 163823 13209 163832 13243
rect 163780 13200 163832 13209
rect 164608 13132 164660 13184
rect 165160 13200 165212 13252
rect 167368 13243 167420 13252
rect 167368 13209 167377 13243
rect 167377 13209 167411 13243
rect 167411 13209 167420 13243
rect 167368 13200 167420 13209
rect 174176 13311 174228 13320
rect 174176 13277 174185 13311
rect 174185 13277 174219 13311
rect 174219 13277 174228 13311
rect 174176 13268 174228 13277
rect 165252 13175 165304 13184
rect 165252 13141 165261 13175
rect 165261 13141 165295 13175
rect 165295 13141 165304 13175
rect 165252 13132 165304 13141
rect 165344 13132 165396 13184
rect 166448 13175 166500 13184
rect 166448 13141 166457 13175
rect 166457 13141 166491 13175
rect 166491 13141 166500 13175
rect 166448 13132 166500 13141
rect 175832 13268 175884 13320
rect 181904 13336 181956 13388
rect 182088 13379 182140 13388
rect 182088 13345 182097 13379
rect 182097 13345 182131 13379
rect 182131 13345 182140 13379
rect 182732 13481 182741 13515
rect 182741 13481 182775 13515
rect 182775 13481 182784 13515
rect 182732 13472 182784 13481
rect 185768 13515 185820 13524
rect 185768 13481 185777 13515
rect 185777 13481 185811 13515
rect 185811 13481 185820 13515
rect 185768 13472 185820 13481
rect 189356 13472 189408 13524
rect 188804 13404 188856 13456
rect 189540 13404 189592 13456
rect 190920 13472 190972 13524
rect 193496 13472 193548 13524
rect 188528 13379 188580 13388
rect 182088 13336 182140 13345
rect 176384 13311 176436 13320
rect 176384 13277 176393 13311
rect 176393 13277 176427 13311
rect 176427 13277 176436 13311
rect 176384 13268 176436 13277
rect 180616 13268 180668 13320
rect 188528 13345 188537 13379
rect 188537 13345 188571 13379
rect 188571 13345 188580 13379
rect 188528 13336 188580 13345
rect 191840 13404 191892 13456
rect 207112 13472 207164 13524
rect 210332 13515 210384 13524
rect 189908 13336 189960 13388
rect 201960 13404 202012 13456
rect 203432 13404 203484 13456
rect 206008 13404 206060 13456
rect 207756 13404 207808 13456
rect 197636 13336 197688 13388
rect 202052 13336 202104 13388
rect 189540 13311 189592 13320
rect 175740 13200 175792 13252
rect 177672 13200 177724 13252
rect 175004 13132 175056 13184
rect 179972 13200 180024 13252
rect 180892 13200 180944 13252
rect 180708 13175 180760 13184
rect 180708 13141 180717 13175
rect 180717 13141 180751 13175
rect 180751 13141 180760 13175
rect 180708 13132 180760 13141
rect 189540 13277 189549 13311
rect 189549 13277 189583 13311
rect 189583 13277 189592 13311
rect 189540 13268 189592 13277
rect 187792 13132 187844 13184
rect 187976 13175 188028 13184
rect 187976 13141 187985 13175
rect 187985 13141 188019 13175
rect 188019 13141 188028 13175
rect 187976 13132 188028 13141
rect 188344 13175 188396 13184
rect 188344 13141 188353 13175
rect 188353 13141 188387 13175
rect 188387 13141 188396 13175
rect 188344 13132 188396 13141
rect 189540 13132 189592 13184
rect 191380 13132 191432 13184
rect 192392 13200 192444 13252
rect 193404 13200 193456 13252
rect 193956 13200 194008 13252
rect 201500 13268 201552 13320
rect 202144 13311 202196 13320
rect 202144 13277 202153 13311
rect 202153 13277 202187 13311
rect 202187 13277 202196 13311
rect 202144 13268 202196 13277
rect 194600 13200 194652 13252
rect 194784 13200 194836 13252
rect 196440 13243 196492 13252
rect 196440 13209 196449 13243
rect 196449 13209 196483 13243
rect 196483 13209 196492 13243
rect 196440 13200 196492 13209
rect 197360 13200 197412 13252
rect 202420 13243 202472 13252
rect 197728 13132 197780 13184
rect 197912 13132 197964 13184
rect 198556 13175 198608 13184
rect 198556 13141 198565 13175
rect 198565 13141 198599 13175
rect 198599 13141 198608 13175
rect 198556 13132 198608 13141
rect 200488 13175 200540 13184
rect 200488 13141 200497 13175
rect 200497 13141 200531 13175
rect 200531 13141 200540 13175
rect 200488 13132 200540 13141
rect 200856 13175 200908 13184
rect 200856 13141 200865 13175
rect 200865 13141 200899 13175
rect 200899 13141 200908 13175
rect 200856 13132 200908 13141
rect 201316 13132 201368 13184
rect 202420 13209 202429 13243
rect 202429 13209 202463 13243
rect 202463 13209 202472 13243
rect 202420 13200 202472 13209
rect 203156 13200 203208 13252
rect 204260 13200 204312 13252
rect 205456 13200 205508 13252
rect 205640 13132 205692 13184
rect 205732 13132 205784 13184
rect 207204 13268 207256 13320
rect 206376 13200 206428 13252
rect 207572 13200 207624 13252
rect 210332 13481 210341 13515
rect 210341 13481 210375 13515
rect 210375 13481 210384 13515
rect 210332 13472 210384 13481
rect 213368 13515 213420 13524
rect 213368 13481 213377 13515
rect 213377 13481 213411 13515
rect 213411 13481 213420 13515
rect 213368 13472 213420 13481
rect 208032 13404 208084 13456
rect 213276 13404 213328 13456
rect 268936 13472 268988 13524
rect 269580 13472 269632 13524
rect 271788 13472 271840 13524
rect 274916 13515 274968 13524
rect 274916 13481 274925 13515
rect 274925 13481 274959 13515
rect 274959 13481 274968 13515
rect 274916 13472 274968 13481
rect 277860 13515 277912 13524
rect 277860 13481 277869 13515
rect 277869 13481 277903 13515
rect 277903 13481 277912 13515
rect 277860 13472 277912 13481
rect 280896 13515 280948 13524
rect 280896 13481 280905 13515
rect 280905 13481 280939 13515
rect 280939 13481 280948 13515
rect 280896 13472 280948 13481
rect 284300 13472 284352 13524
rect 287060 13472 287112 13524
rect 290096 13515 290148 13524
rect 290096 13481 290105 13515
rect 290105 13481 290139 13515
rect 290139 13481 290148 13515
rect 290096 13472 290148 13481
rect 293224 13515 293276 13524
rect 293224 13481 293233 13515
rect 293233 13481 293267 13515
rect 293267 13481 293276 13515
rect 293224 13472 293276 13481
rect 296260 13515 296312 13524
rect 296260 13481 296269 13515
rect 296269 13481 296303 13515
rect 296303 13481 296312 13515
rect 296260 13472 296312 13481
rect 299296 13515 299348 13524
rect 299296 13481 299305 13515
rect 299305 13481 299339 13515
rect 299339 13481 299348 13515
rect 299296 13472 299348 13481
rect 301412 13515 301464 13524
rect 301412 13481 301421 13515
rect 301421 13481 301455 13515
rect 301455 13481 301464 13515
rect 301412 13472 301464 13481
rect 216404 13447 216456 13456
rect 216404 13413 216413 13447
rect 216413 13413 216447 13447
rect 216447 13413 216456 13447
rect 216404 13404 216456 13413
rect 219440 13404 219492 13456
rect 207940 13268 207992 13320
rect 213552 13311 213604 13320
rect 213552 13277 213561 13311
rect 213561 13277 213595 13311
rect 213595 13277 213604 13311
rect 213552 13268 213604 13277
rect 216588 13311 216640 13320
rect 216588 13277 216597 13311
rect 216597 13277 216631 13311
rect 216631 13277 216640 13311
rect 224132 13404 224184 13456
rect 224040 13336 224092 13388
rect 226432 13404 226484 13456
rect 226616 13447 226668 13456
rect 226616 13413 226625 13447
rect 226625 13413 226659 13447
rect 226659 13413 226668 13447
rect 226616 13404 226668 13413
rect 226892 13404 226944 13456
rect 227904 13404 227956 13456
rect 229192 13404 229244 13456
rect 224408 13336 224460 13388
rect 227076 13379 227128 13388
rect 227076 13345 227085 13379
rect 227085 13345 227119 13379
rect 227119 13345 227128 13379
rect 227076 13336 227128 13345
rect 227168 13379 227220 13388
rect 227168 13345 227177 13379
rect 227177 13345 227211 13379
rect 227211 13345 227220 13379
rect 227168 13336 227220 13345
rect 216588 13268 216640 13277
rect 224224 13200 224276 13252
rect 207388 13132 207440 13184
rect 213552 13132 213604 13184
rect 222752 13175 222804 13184
rect 222752 13141 222761 13175
rect 222761 13141 222795 13175
rect 222795 13141 222804 13175
rect 222752 13132 222804 13141
rect 223672 13175 223724 13184
rect 223672 13141 223681 13175
rect 223681 13141 223715 13175
rect 223715 13141 223724 13175
rect 223672 13132 223724 13141
rect 224040 13175 224092 13184
rect 224040 13141 224049 13175
rect 224049 13141 224083 13175
rect 224083 13141 224092 13175
rect 224040 13132 224092 13141
rect 224132 13175 224184 13184
rect 224132 13141 224141 13175
rect 224141 13141 224175 13175
rect 224175 13141 224184 13175
rect 224408 13200 224460 13252
rect 227720 13268 227772 13320
rect 231952 13336 232004 13388
rect 230388 13268 230440 13320
rect 231860 13268 231912 13320
rect 232044 13268 232096 13320
rect 233148 13336 233200 13388
rect 233332 13336 233384 13388
rect 233056 13311 233108 13320
rect 233056 13277 233065 13311
rect 233065 13277 233099 13311
rect 233099 13277 233108 13311
rect 233056 13268 233108 13277
rect 228088 13200 228140 13252
rect 230756 13243 230808 13252
rect 230756 13209 230765 13243
rect 230765 13209 230799 13243
rect 230799 13209 230808 13243
rect 230756 13200 230808 13209
rect 237932 13336 237984 13388
rect 238116 13336 238168 13388
rect 239496 13404 239548 13456
rect 244648 13404 244700 13456
rect 245384 13404 245436 13456
rect 247132 13447 247184 13456
rect 247132 13413 247141 13447
rect 247141 13413 247175 13447
rect 247175 13413 247184 13447
rect 247132 13404 247184 13413
rect 251088 13404 251140 13456
rect 252468 13404 252520 13456
rect 254952 13404 255004 13456
rect 259460 13447 259512 13456
rect 259460 13413 259469 13447
rect 259469 13413 259503 13447
rect 259503 13413 259512 13447
rect 259460 13404 259512 13413
rect 263508 13404 263560 13456
rect 265532 13404 265584 13456
rect 270408 13404 270460 13456
rect 244096 13336 244148 13388
rect 238208 13311 238260 13320
rect 238208 13277 238217 13311
rect 238217 13277 238251 13311
rect 238251 13277 238260 13311
rect 238208 13268 238260 13277
rect 239772 13268 239824 13320
rect 250996 13336 251048 13388
rect 251088 13311 251140 13320
rect 251088 13277 251097 13311
rect 251097 13277 251131 13311
rect 251131 13277 251140 13311
rect 251088 13268 251140 13277
rect 224132 13132 224184 13141
rect 225420 13132 225472 13184
rect 225696 13175 225748 13184
rect 225696 13141 225705 13175
rect 225705 13141 225739 13175
rect 225739 13141 225748 13175
rect 225696 13132 225748 13141
rect 227076 13132 227128 13184
rect 227628 13132 227680 13184
rect 227904 13132 227956 13184
rect 232136 13132 232188 13184
rect 233240 13132 233292 13184
rect 234896 13175 234948 13184
rect 234896 13141 234905 13175
rect 234905 13141 234939 13175
rect 234939 13141 234948 13175
rect 234896 13132 234948 13141
rect 237012 13132 237064 13184
rect 238484 13243 238536 13252
rect 238484 13209 238493 13243
rect 238493 13209 238527 13243
rect 238527 13209 238536 13243
rect 241060 13243 241112 13252
rect 238484 13200 238536 13209
rect 241060 13209 241069 13243
rect 241069 13209 241103 13243
rect 241103 13209 241112 13243
rect 241060 13200 241112 13209
rect 241796 13200 241848 13252
rect 243636 13243 243688 13252
rect 242532 13175 242584 13184
rect 242532 13141 242541 13175
rect 242541 13141 242575 13175
rect 242575 13141 242584 13175
rect 242532 13132 242584 13141
rect 243636 13209 243645 13243
rect 243645 13209 243679 13243
rect 243679 13209 243688 13243
rect 243636 13200 243688 13209
rect 244924 13200 244976 13252
rect 251180 13132 251232 13184
rect 251364 13243 251416 13252
rect 251364 13209 251373 13243
rect 251373 13209 251407 13243
rect 251407 13209 251416 13243
rect 251364 13200 251416 13209
rect 252376 13200 252428 13252
rect 256240 13311 256292 13320
rect 253020 13200 253072 13252
rect 254952 13200 255004 13252
rect 253480 13132 253532 13184
rect 256240 13277 256249 13311
rect 256249 13277 256283 13311
rect 256283 13277 256292 13311
rect 256240 13268 256292 13277
rect 255320 13200 255372 13252
rect 256976 13200 257028 13252
rect 256332 13132 256384 13184
rect 264152 13336 264204 13388
rect 272984 13404 273036 13456
rect 268936 13268 268988 13320
rect 273168 13336 273220 13388
rect 273260 13268 273312 13320
rect 275100 13311 275152 13320
rect 275100 13277 275109 13311
rect 275109 13277 275143 13311
rect 275143 13277 275152 13311
rect 275100 13268 275152 13277
rect 261852 13243 261904 13252
rect 261852 13209 261861 13243
rect 261861 13209 261895 13243
rect 261895 13209 261904 13243
rect 261852 13200 261904 13209
rect 263416 13200 263468 13252
rect 263508 13200 263560 13252
rect 264428 13200 264480 13252
rect 264612 13200 264664 13252
rect 264980 13200 265032 13252
rect 257988 13175 258040 13184
rect 257988 13141 257997 13175
rect 257997 13141 258031 13175
rect 258031 13141 258040 13175
rect 257988 13132 258040 13141
rect 262956 13132 263008 13184
rect 263324 13132 263376 13184
rect 266912 13200 266964 13252
rect 267648 13132 267700 13184
rect 268752 13200 268804 13252
rect 270684 13200 270736 13252
rect 270776 13132 270828 13184
rect 270960 13200 271012 13252
rect 281080 13311 281132 13320
rect 281080 13277 281089 13311
rect 281089 13277 281123 13311
rect 281123 13277 281132 13311
rect 281080 13268 281132 13277
rect 284760 13311 284812 13320
rect 284760 13277 284769 13311
rect 284769 13277 284803 13311
rect 284803 13277 284812 13311
rect 284760 13268 284812 13277
rect 290280 13311 290332 13320
rect 290280 13277 290289 13311
rect 290289 13277 290323 13311
rect 290323 13277 290332 13311
rect 290280 13268 290332 13277
rect 305000 13336 305052 13388
rect 271788 13132 271840 13184
rect 272892 13132 272944 13184
rect 299480 13311 299532 13320
rect 299480 13277 299489 13311
rect 299489 13277 299523 13311
rect 299523 13277 299532 13311
rect 299480 13268 299532 13277
rect 303528 13268 303580 13320
rect 295892 13175 295944 13184
rect 295892 13141 295901 13175
rect 295901 13141 295935 13175
rect 295935 13141 295944 13175
rect 295892 13132 295944 13141
rect 77148 13030 77200 13082
rect 77212 13030 77264 13082
rect 77276 13030 77328 13082
rect 77340 13030 77392 13082
rect 77404 13030 77456 13082
rect 153346 13030 153398 13082
rect 153410 13030 153462 13082
rect 153474 13030 153526 13082
rect 153538 13030 153590 13082
rect 153602 13030 153654 13082
rect 229544 13030 229596 13082
rect 229608 13030 229660 13082
rect 229672 13030 229724 13082
rect 229736 13030 229788 13082
rect 229800 13030 229852 13082
rect 26056 12971 26108 12980
rect 26056 12937 26065 12971
rect 26065 12937 26099 12971
rect 26099 12937 26108 12971
rect 26056 12928 26108 12937
rect 20168 12860 20220 12912
rect 27344 12860 27396 12912
rect 32220 12928 32272 12980
rect 34152 12928 34204 12980
rect 35532 12971 35584 12980
rect 35532 12937 35541 12971
rect 35541 12937 35575 12971
rect 35575 12937 35584 12971
rect 35532 12928 35584 12937
rect 29000 12903 29052 12912
rect 23204 12724 23256 12776
rect 29000 12869 29009 12903
rect 29009 12869 29043 12903
rect 29043 12869 29052 12903
rect 29000 12860 29052 12869
rect 27988 12792 28040 12844
rect 28080 12767 28132 12776
rect 27160 12656 27212 12708
rect 28080 12733 28089 12767
rect 28089 12733 28123 12767
rect 28123 12733 28132 12767
rect 28080 12724 28132 12733
rect 30380 12860 30432 12912
rect 31576 12860 31628 12912
rect 34428 12860 34480 12912
rect 33692 12792 33744 12844
rect 37464 12860 37516 12912
rect 39672 12860 39724 12912
rect 41052 12860 41104 12912
rect 43260 12928 43312 12980
rect 44272 12928 44324 12980
rect 44548 12971 44600 12980
rect 44548 12937 44557 12971
rect 44557 12937 44591 12971
rect 44591 12937 44600 12971
rect 44548 12928 44600 12937
rect 53288 12928 53340 12980
rect 42984 12860 43036 12912
rect 54668 12928 54720 12980
rect 55864 12928 55916 12980
rect 57980 12928 58032 12980
rect 59636 12928 59688 12980
rect 72148 12971 72200 12980
rect 72148 12937 72157 12971
rect 72157 12937 72191 12971
rect 72191 12937 72200 12971
rect 72148 12928 72200 12937
rect 72332 12928 72384 12980
rect 74724 12928 74776 12980
rect 29644 12724 29696 12776
rect 29828 12767 29880 12776
rect 29828 12733 29837 12767
rect 29837 12733 29871 12767
rect 29871 12733 29880 12767
rect 29828 12724 29880 12733
rect 30104 12767 30156 12776
rect 30104 12733 30113 12767
rect 30113 12733 30147 12767
rect 30147 12733 30156 12767
rect 30104 12724 30156 12733
rect 28908 12588 28960 12640
rect 33048 12724 33100 12776
rect 33416 12724 33468 12776
rect 34336 12724 34388 12776
rect 39304 12792 39356 12844
rect 41512 12792 41564 12844
rect 34888 12767 34940 12776
rect 34888 12733 34897 12767
rect 34897 12733 34931 12767
rect 34931 12733 34940 12767
rect 34888 12724 34940 12733
rect 35348 12724 35400 12776
rect 39396 12724 39448 12776
rect 40960 12724 41012 12776
rect 43076 12724 43128 12776
rect 43168 12724 43220 12776
rect 45376 12792 45428 12844
rect 55496 12860 55548 12912
rect 57336 12860 57388 12912
rect 60648 12860 60700 12912
rect 65892 12860 65944 12912
rect 53748 12792 53800 12844
rect 54024 12835 54076 12844
rect 43812 12724 43864 12776
rect 45468 12724 45520 12776
rect 51356 12724 51408 12776
rect 54024 12801 54033 12835
rect 54033 12801 54067 12835
rect 54067 12801 54076 12835
rect 54024 12792 54076 12801
rect 54760 12835 54812 12844
rect 54116 12767 54168 12776
rect 54116 12733 54125 12767
rect 54125 12733 54159 12767
rect 54159 12733 54168 12767
rect 54116 12724 54168 12733
rect 54760 12801 54769 12835
rect 54769 12801 54803 12835
rect 54803 12801 54812 12835
rect 54760 12792 54812 12801
rect 57428 12792 57480 12844
rect 74816 12792 74868 12844
rect 75460 12792 75512 12844
rect 78404 12860 78456 12912
rect 79692 12792 79744 12844
rect 83924 12928 83976 12980
rect 80520 12860 80572 12912
rect 82912 12860 82964 12912
rect 86500 12928 86552 12980
rect 87144 12928 87196 12980
rect 90456 12928 90508 12980
rect 91652 12928 91704 12980
rect 98000 12928 98052 12980
rect 55036 12767 55088 12776
rect 55036 12733 55045 12767
rect 55045 12733 55079 12767
rect 55079 12733 55088 12767
rect 55036 12724 55088 12733
rect 78588 12724 78640 12776
rect 31392 12588 31444 12640
rect 32404 12588 32456 12640
rect 34152 12588 34204 12640
rect 38016 12631 38068 12640
rect 38016 12597 38025 12631
rect 38025 12597 38059 12631
rect 38059 12597 38068 12631
rect 38016 12588 38068 12597
rect 41236 12631 41288 12640
rect 41236 12597 41245 12631
rect 41245 12597 41279 12631
rect 41279 12597 41288 12631
rect 41236 12588 41288 12597
rect 41788 12631 41840 12640
rect 41788 12597 41797 12631
rect 41797 12597 41831 12631
rect 41831 12597 41840 12631
rect 41788 12588 41840 12597
rect 42800 12588 42852 12640
rect 43260 12588 43312 12640
rect 43812 12588 43864 12640
rect 53104 12588 53156 12640
rect 54116 12588 54168 12640
rect 55588 12588 55640 12640
rect 56324 12588 56376 12640
rect 56508 12631 56560 12640
rect 56508 12597 56517 12631
rect 56517 12597 56551 12631
rect 56551 12597 56560 12631
rect 56508 12588 56560 12597
rect 57244 12588 57296 12640
rect 72700 12588 72752 12640
rect 75000 12588 75052 12640
rect 75184 12588 75236 12640
rect 77852 12656 77904 12708
rect 78128 12656 78180 12708
rect 80796 12724 80848 12776
rect 77208 12588 77260 12640
rect 81440 12656 81492 12708
rect 81624 12588 81676 12640
rect 84844 12724 84896 12776
rect 85764 12631 85816 12640
rect 85764 12597 85773 12631
rect 85773 12597 85807 12631
rect 85807 12597 85816 12631
rect 85764 12588 85816 12597
rect 90548 12860 90600 12912
rect 90732 12860 90784 12912
rect 99472 12903 99524 12912
rect 99472 12869 99481 12903
rect 99481 12869 99515 12903
rect 99515 12869 99524 12903
rect 99472 12860 99524 12869
rect 99932 12860 99984 12912
rect 104624 12903 104676 12912
rect 104624 12869 104633 12903
rect 104633 12869 104667 12903
rect 104667 12869 104676 12903
rect 104624 12860 104676 12869
rect 104716 12903 104768 12912
rect 104716 12869 104725 12903
rect 104725 12869 104759 12903
rect 104759 12869 104768 12903
rect 104716 12860 104768 12869
rect 90180 12792 90232 12844
rect 90456 12835 90508 12844
rect 90456 12801 90465 12835
rect 90465 12801 90499 12835
rect 90499 12801 90508 12835
rect 90456 12792 90508 12801
rect 90640 12792 90692 12844
rect 86500 12767 86552 12776
rect 86500 12733 86509 12767
rect 86509 12733 86543 12767
rect 86543 12733 86552 12767
rect 86500 12724 86552 12733
rect 88248 12724 88300 12776
rect 89720 12724 89772 12776
rect 90088 12724 90140 12776
rect 105176 12792 105228 12844
rect 99196 12767 99248 12776
rect 99196 12733 99205 12767
rect 99205 12733 99239 12767
rect 99239 12733 99248 12767
rect 101404 12767 101456 12776
rect 99196 12724 99248 12733
rect 101404 12733 101413 12767
rect 101413 12733 101447 12767
rect 101447 12733 101456 12767
rect 101404 12724 101456 12733
rect 101680 12767 101732 12776
rect 101680 12733 101689 12767
rect 101689 12733 101723 12767
rect 101723 12733 101732 12767
rect 101680 12724 101732 12733
rect 87788 12588 87840 12640
rect 87972 12631 88024 12640
rect 87972 12597 87981 12631
rect 87981 12597 88015 12631
rect 88015 12597 88024 12631
rect 87972 12588 88024 12597
rect 88432 12588 88484 12640
rect 89904 12588 89956 12640
rect 99196 12588 99248 12640
rect 101036 12656 101088 12708
rect 103244 12656 103296 12708
rect 105912 12699 105964 12708
rect 105912 12665 105921 12699
rect 105921 12665 105955 12699
rect 105955 12665 105964 12699
rect 105912 12656 105964 12665
rect 111432 12928 111484 12980
rect 114560 12928 114612 12980
rect 114744 12928 114796 12980
rect 117412 12928 117464 12980
rect 118240 12971 118292 12980
rect 118240 12937 118249 12971
rect 118249 12937 118283 12971
rect 118283 12937 118292 12971
rect 118240 12928 118292 12937
rect 118700 12971 118752 12980
rect 118700 12937 118709 12971
rect 118709 12937 118743 12971
rect 118743 12937 118752 12971
rect 118700 12928 118752 12937
rect 126888 12928 126940 12980
rect 128084 12971 128136 12980
rect 128084 12937 128093 12971
rect 128093 12937 128127 12971
rect 128127 12937 128136 12971
rect 128084 12928 128136 12937
rect 128636 12928 128688 12980
rect 129188 12971 129240 12980
rect 129188 12937 129197 12971
rect 129197 12937 129231 12971
rect 129231 12937 129240 12971
rect 129188 12928 129240 12937
rect 133328 12928 133380 12980
rect 109592 12860 109644 12912
rect 113088 12835 113140 12844
rect 113088 12801 113097 12835
rect 113097 12801 113131 12835
rect 113131 12801 113140 12835
rect 113088 12792 113140 12801
rect 113824 12835 113876 12844
rect 113824 12801 113833 12835
rect 113833 12801 113867 12835
rect 113867 12801 113876 12835
rect 113824 12792 113876 12801
rect 114652 12835 114704 12844
rect 114652 12801 114661 12835
rect 114661 12801 114695 12835
rect 114695 12801 114704 12835
rect 115756 12860 115808 12912
rect 117320 12860 117372 12912
rect 126520 12860 126572 12912
rect 114652 12792 114704 12801
rect 118056 12792 118108 12844
rect 132408 12860 132460 12912
rect 133604 12903 133656 12912
rect 133604 12869 133613 12903
rect 133613 12869 133647 12903
rect 133647 12869 133656 12903
rect 133604 12860 133656 12869
rect 133880 12928 133932 12980
rect 147680 12928 147732 12980
rect 134156 12860 134208 12912
rect 143080 12860 143132 12912
rect 145932 12903 145984 12912
rect 127440 12835 127492 12844
rect 127440 12801 127449 12835
rect 127449 12801 127483 12835
rect 127483 12801 127492 12835
rect 127440 12792 127492 12801
rect 113916 12724 113968 12776
rect 114744 12724 114796 12776
rect 115664 12724 115716 12776
rect 115848 12767 115900 12776
rect 115848 12733 115857 12767
rect 115857 12733 115891 12767
rect 115891 12733 115900 12767
rect 115848 12724 115900 12733
rect 116768 12767 116820 12776
rect 114836 12656 114888 12708
rect 116768 12733 116777 12767
rect 116777 12733 116811 12767
rect 116811 12733 116820 12767
rect 116768 12724 116820 12733
rect 100760 12588 100812 12640
rect 103060 12588 103112 12640
rect 103612 12588 103664 12640
rect 111892 12631 111944 12640
rect 111892 12597 111901 12631
rect 111901 12597 111935 12631
rect 111935 12597 111944 12631
rect 111892 12588 111944 12597
rect 113088 12588 113140 12640
rect 114744 12631 114796 12640
rect 114744 12597 114753 12631
rect 114753 12597 114787 12631
rect 114787 12597 114796 12631
rect 114744 12588 114796 12597
rect 115848 12588 115900 12640
rect 127532 12724 127584 12776
rect 128084 12588 128136 12640
rect 129096 12835 129148 12844
rect 129096 12801 129105 12835
rect 129105 12801 129139 12835
rect 129139 12801 129148 12835
rect 129096 12792 129148 12801
rect 128360 12724 128412 12776
rect 130292 12792 130344 12844
rect 129740 12724 129792 12776
rect 131120 12767 131172 12776
rect 131120 12733 131129 12767
rect 131129 12733 131163 12767
rect 131163 12733 131172 12767
rect 131120 12724 131172 12733
rect 132592 12767 132644 12776
rect 132592 12733 132601 12767
rect 132601 12733 132635 12767
rect 132635 12733 132644 12767
rect 133696 12792 133748 12844
rect 145932 12869 145941 12903
rect 145941 12869 145975 12903
rect 145975 12869 145984 12903
rect 145932 12860 145984 12869
rect 152648 12928 152700 12980
rect 152832 12928 152884 12980
rect 157156 12971 157208 12980
rect 157156 12937 157165 12971
rect 157165 12937 157199 12971
rect 157199 12937 157208 12971
rect 157156 12928 157208 12937
rect 158628 12928 158680 12980
rect 145840 12835 145892 12844
rect 132592 12724 132644 12733
rect 143264 12767 143316 12776
rect 130292 12656 130344 12708
rect 133696 12656 133748 12708
rect 133144 12631 133196 12640
rect 133144 12597 133153 12631
rect 133153 12597 133187 12631
rect 133187 12597 133196 12631
rect 133144 12588 133196 12597
rect 133236 12588 133288 12640
rect 143264 12733 143273 12767
rect 143273 12733 143307 12767
rect 143307 12733 143316 12767
rect 143264 12724 143316 12733
rect 145840 12801 145849 12835
rect 145849 12801 145883 12835
rect 145883 12801 145892 12835
rect 145840 12792 145892 12801
rect 156604 12860 156656 12912
rect 147312 12792 147364 12844
rect 149336 12792 149388 12844
rect 147404 12724 147456 12776
rect 147772 12767 147824 12776
rect 133880 12656 133932 12708
rect 145748 12656 145800 12708
rect 147772 12733 147781 12767
rect 147781 12733 147815 12767
rect 147815 12733 147824 12767
rect 147772 12724 147824 12733
rect 148968 12724 149020 12776
rect 149244 12767 149296 12776
rect 149244 12733 149253 12767
rect 149253 12733 149287 12767
rect 149287 12733 149296 12767
rect 149244 12724 149296 12733
rect 150440 12792 150492 12844
rect 155868 12792 155920 12844
rect 157800 12792 157852 12844
rect 160376 12860 160428 12912
rect 161664 12792 161716 12844
rect 151544 12767 151596 12776
rect 151544 12733 151553 12767
rect 151553 12733 151587 12767
rect 151587 12733 151596 12767
rect 151544 12724 151596 12733
rect 150348 12656 150400 12708
rect 151636 12656 151688 12708
rect 148508 12588 148560 12640
rect 149980 12631 150032 12640
rect 149980 12597 149989 12631
rect 149989 12597 150023 12631
rect 150023 12597 150032 12631
rect 149980 12588 150032 12597
rect 151268 12588 151320 12640
rect 151360 12588 151412 12640
rect 152740 12724 152792 12776
rect 152832 12656 152884 12708
rect 153108 12656 153160 12708
rect 155040 12767 155092 12776
rect 155040 12733 155049 12767
rect 155049 12733 155083 12767
rect 155083 12733 155092 12767
rect 159456 12767 159508 12776
rect 155040 12724 155092 12733
rect 158812 12699 158864 12708
rect 158812 12665 158821 12699
rect 158821 12665 158855 12699
rect 158855 12665 158864 12699
rect 158812 12656 158864 12665
rect 159456 12733 159465 12767
rect 159465 12733 159499 12767
rect 159499 12733 159508 12767
rect 159456 12724 159508 12733
rect 159548 12724 159600 12776
rect 161572 12724 161624 12776
rect 154120 12588 154172 12640
rect 157892 12588 157944 12640
rect 160284 12588 160336 12640
rect 163504 12928 163556 12980
rect 163412 12860 163464 12912
rect 165252 12928 165304 12980
rect 162124 12767 162176 12776
rect 162124 12733 162133 12767
rect 162133 12733 162167 12767
rect 162167 12733 162176 12767
rect 162124 12724 162176 12733
rect 162860 12724 162912 12776
rect 167184 12928 167236 12980
rect 175004 12971 175056 12980
rect 175004 12937 175013 12971
rect 175013 12937 175047 12971
rect 175047 12937 175056 12971
rect 175004 12928 175056 12937
rect 175740 12928 175792 12980
rect 176384 12928 176436 12980
rect 165436 12792 165488 12844
rect 166172 12792 166224 12844
rect 166540 12835 166592 12844
rect 166540 12801 166549 12835
rect 166549 12801 166583 12835
rect 166583 12801 166592 12835
rect 166540 12792 166592 12801
rect 173808 12860 173860 12912
rect 175924 12860 175976 12912
rect 176936 12860 176988 12912
rect 177948 12860 178000 12912
rect 176384 12835 176436 12844
rect 164608 12767 164660 12776
rect 164608 12733 164617 12767
rect 164617 12733 164651 12767
rect 164651 12733 164660 12767
rect 164608 12724 164660 12733
rect 163688 12588 163740 12640
rect 164240 12656 164292 12708
rect 176384 12801 176393 12835
rect 176393 12801 176427 12835
rect 176427 12801 176436 12835
rect 176384 12792 176436 12801
rect 180156 12928 180208 12980
rect 180248 12928 180300 12980
rect 180340 12792 180392 12844
rect 181536 12835 181588 12844
rect 181536 12801 181545 12835
rect 181545 12801 181579 12835
rect 181579 12801 181588 12835
rect 188344 12928 188396 12980
rect 191380 12928 191432 12980
rect 192484 12928 192536 12980
rect 188528 12860 188580 12912
rect 190920 12903 190972 12912
rect 181536 12792 181588 12801
rect 188344 12792 188396 12844
rect 188804 12792 188856 12844
rect 189356 12835 189408 12844
rect 189356 12801 189365 12835
rect 189365 12801 189399 12835
rect 189399 12801 189408 12835
rect 189356 12792 189408 12801
rect 176752 12724 176804 12776
rect 180156 12724 180208 12776
rect 189540 12724 189592 12776
rect 190920 12869 190929 12903
rect 190929 12869 190963 12903
rect 190963 12869 190972 12903
rect 190920 12860 190972 12869
rect 191748 12860 191800 12912
rect 193956 12928 194008 12980
rect 194876 12928 194928 12980
rect 195980 12971 196032 12980
rect 195980 12937 195989 12971
rect 195989 12937 196023 12971
rect 196023 12937 196032 12971
rect 195980 12928 196032 12937
rect 197728 12928 197780 12980
rect 192576 12792 192628 12844
rect 195060 12835 195112 12844
rect 195060 12801 195069 12835
rect 195069 12801 195103 12835
rect 195103 12801 195112 12835
rect 195060 12792 195112 12801
rect 197360 12835 197412 12844
rect 197360 12801 197369 12835
rect 197369 12801 197403 12835
rect 197403 12801 197412 12835
rect 197360 12792 197412 12801
rect 197452 12835 197504 12844
rect 197452 12801 197461 12835
rect 197461 12801 197495 12835
rect 197495 12801 197504 12835
rect 198372 12835 198424 12844
rect 197452 12792 197504 12801
rect 192668 12724 192720 12776
rect 193036 12767 193088 12776
rect 193036 12733 193045 12767
rect 193045 12733 193079 12767
rect 193079 12733 193088 12767
rect 193036 12724 193088 12733
rect 166172 12588 166224 12640
rect 166632 12631 166684 12640
rect 166632 12597 166641 12631
rect 166641 12597 166675 12631
rect 166675 12597 166684 12631
rect 166632 12588 166684 12597
rect 180248 12656 180300 12708
rect 180524 12656 180576 12708
rect 182088 12656 182140 12708
rect 188620 12656 188672 12708
rect 189172 12656 189224 12708
rect 191748 12656 191800 12708
rect 191932 12656 191984 12708
rect 192484 12656 192536 12708
rect 194784 12724 194836 12776
rect 195796 12724 195848 12776
rect 197636 12767 197688 12776
rect 197636 12733 197645 12767
rect 197645 12733 197679 12767
rect 197679 12733 197688 12767
rect 197636 12724 197688 12733
rect 198372 12801 198381 12835
rect 198381 12801 198415 12835
rect 198415 12801 198424 12835
rect 198372 12792 198424 12801
rect 200672 12792 200724 12844
rect 201316 12835 201368 12844
rect 201316 12801 201325 12835
rect 201325 12801 201359 12835
rect 201359 12801 201368 12835
rect 201316 12792 201368 12801
rect 198556 12724 198608 12776
rect 200396 12724 200448 12776
rect 202972 12860 203024 12912
rect 203340 12860 203392 12912
rect 205640 12860 205692 12912
rect 206560 12971 206612 12980
rect 206560 12937 206569 12971
rect 206569 12937 206603 12971
rect 206603 12937 206612 12971
rect 206560 12928 206612 12937
rect 207388 12928 207440 12980
rect 207848 12928 207900 12980
rect 202880 12767 202932 12776
rect 177396 12588 177448 12640
rect 177856 12588 177908 12640
rect 179880 12588 179932 12640
rect 180616 12588 180668 12640
rect 181444 12588 181496 12640
rect 187792 12588 187844 12640
rect 188988 12588 189040 12640
rect 190552 12631 190604 12640
rect 190552 12597 190561 12631
rect 190561 12597 190595 12631
rect 190595 12597 190604 12631
rect 190552 12588 190604 12597
rect 192024 12588 192076 12640
rect 192116 12588 192168 12640
rect 193036 12588 193088 12640
rect 202144 12656 202196 12708
rect 202880 12733 202889 12767
rect 202889 12733 202923 12767
rect 202923 12733 202932 12767
rect 202880 12724 202932 12733
rect 202972 12724 203024 12776
rect 204168 12724 204220 12776
rect 205088 12767 205140 12776
rect 205088 12733 205097 12767
rect 205097 12733 205131 12767
rect 205131 12733 205140 12767
rect 205088 12724 205140 12733
rect 205180 12724 205232 12776
rect 210608 12860 210660 12912
rect 219808 12928 219860 12980
rect 207664 12792 207716 12844
rect 216588 12792 216640 12844
rect 228272 12860 228324 12912
rect 230388 12860 230440 12912
rect 219808 12792 219860 12844
rect 223672 12792 223724 12844
rect 226800 12792 226852 12844
rect 227904 12835 227956 12844
rect 227904 12801 227913 12835
rect 227913 12801 227947 12835
rect 227947 12801 227956 12835
rect 227904 12792 227956 12801
rect 230296 12835 230348 12844
rect 230296 12801 230305 12835
rect 230305 12801 230339 12835
rect 230339 12801 230348 12835
rect 230296 12792 230348 12801
rect 238208 12928 238260 12980
rect 231032 12903 231084 12912
rect 231032 12869 231041 12903
rect 231041 12869 231075 12903
rect 231075 12869 231084 12903
rect 231032 12860 231084 12869
rect 232320 12860 232372 12912
rect 238300 12860 238352 12912
rect 233056 12835 233108 12844
rect 207296 12699 207348 12708
rect 194416 12588 194468 12640
rect 195980 12588 196032 12640
rect 198188 12631 198240 12640
rect 198188 12597 198197 12631
rect 198197 12597 198231 12631
rect 198231 12597 198240 12631
rect 198188 12588 198240 12597
rect 201132 12631 201184 12640
rect 201132 12597 201141 12631
rect 201141 12597 201175 12631
rect 201175 12597 201184 12631
rect 201132 12588 201184 12597
rect 201960 12588 202012 12640
rect 204260 12588 204312 12640
rect 204536 12588 204588 12640
rect 205180 12588 205232 12640
rect 205272 12588 205324 12640
rect 207296 12665 207305 12699
rect 207305 12665 207339 12699
rect 207339 12665 207348 12699
rect 207296 12656 207348 12665
rect 210608 12588 210660 12640
rect 219808 12656 219860 12708
rect 226892 12588 226944 12640
rect 228272 12724 228324 12776
rect 230204 12724 230256 12776
rect 233056 12801 233065 12835
rect 233065 12801 233099 12835
rect 233099 12801 233108 12835
rect 233056 12792 233108 12801
rect 237012 12835 237064 12844
rect 237012 12801 237021 12835
rect 237021 12801 237055 12835
rect 237055 12801 237064 12835
rect 237012 12792 237064 12801
rect 238392 12792 238444 12844
rect 239036 12860 239088 12912
rect 240048 12860 240100 12912
rect 251088 12928 251140 12980
rect 254676 12928 254728 12980
rect 256240 12928 256292 12980
rect 264612 12971 264664 12980
rect 240968 12903 241020 12912
rect 240968 12869 240977 12903
rect 240977 12869 241011 12903
rect 241011 12869 241020 12903
rect 240968 12860 241020 12869
rect 242072 12792 242124 12844
rect 242256 12792 242308 12844
rect 244648 12860 244700 12912
rect 244924 12860 244976 12912
rect 245384 12860 245436 12912
rect 251640 12860 251692 12912
rect 252468 12903 252520 12912
rect 252468 12869 252477 12903
rect 252477 12869 252511 12903
rect 252511 12869 252520 12903
rect 252468 12860 252520 12869
rect 244556 12835 244608 12844
rect 244556 12801 244565 12835
rect 244565 12801 244599 12835
rect 244599 12801 244608 12835
rect 244556 12792 244608 12801
rect 244832 12792 244884 12844
rect 251180 12792 251232 12844
rect 251548 12835 251600 12844
rect 251548 12801 251557 12835
rect 251557 12801 251591 12835
rect 251591 12801 251600 12835
rect 251548 12792 251600 12801
rect 256608 12792 256660 12844
rect 237840 12656 237892 12708
rect 237932 12656 237984 12708
rect 229560 12588 229612 12640
rect 230112 12631 230164 12640
rect 230112 12597 230121 12631
rect 230121 12597 230155 12631
rect 230155 12597 230164 12631
rect 230112 12588 230164 12597
rect 230204 12588 230256 12640
rect 232320 12588 232372 12640
rect 232504 12631 232556 12640
rect 232504 12597 232513 12631
rect 232513 12597 232547 12631
rect 232547 12597 232556 12631
rect 232504 12588 232556 12597
rect 233148 12588 233200 12640
rect 238484 12588 238536 12640
rect 238852 12588 238904 12640
rect 239128 12588 239180 12640
rect 240324 12588 240376 12640
rect 242164 12656 242216 12708
rect 242440 12631 242492 12640
rect 242440 12597 242449 12631
rect 242449 12597 242483 12631
rect 242483 12597 242492 12631
rect 242440 12588 242492 12597
rect 242900 12588 242952 12640
rect 244648 12656 244700 12708
rect 248328 12656 248380 12708
rect 250168 12699 250220 12708
rect 250168 12665 250177 12699
rect 250177 12665 250211 12699
rect 250211 12665 250220 12699
rect 250168 12656 250220 12665
rect 252100 12724 252152 12776
rect 253664 12767 253716 12776
rect 253664 12733 253673 12767
rect 253673 12733 253707 12767
rect 253707 12733 253716 12767
rect 253664 12724 253716 12733
rect 253940 12767 253992 12776
rect 253940 12733 253949 12767
rect 253949 12733 253983 12767
rect 253983 12733 253992 12767
rect 253940 12724 253992 12733
rect 255136 12724 255188 12776
rect 256332 12767 256384 12776
rect 256332 12733 256341 12767
rect 256341 12733 256375 12767
rect 256375 12733 256384 12767
rect 256332 12724 256384 12733
rect 256424 12767 256476 12776
rect 256424 12733 256433 12767
rect 256433 12733 256467 12767
rect 256467 12733 256476 12767
rect 256424 12724 256476 12733
rect 251824 12656 251876 12708
rect 255044 12656 255096 12708
rect 251916 12588 251968 12640
rect 252008 12631 252060 12640
rect 252008 12597 252017 12631
rect 252017 12597 252051 12631
rect 252051 12597 252060 12631
rect 257252 12860 257304 12912
rect 261760 12903 261812 12912
rect 261760 12869 261769 12903
rect 261769 12869 261803 12903
rect 261803 12869 261812 12903
rect 261760 12860 261812 12869
rect 263324 12860 263376 12912
rect 264612 12937 264621 12971
rect 264621 12937 264655 12971
rect 264655 12937 264664 12971
rect 264612 12928 264664 12937
rect 268384 12928 268436 12980
rect 302608 12971 302660 12980
rect 265532 12903 265584 12912
rect 261852 12792 261904 12844
rect 264336 12792 264388 12844
rect 264428 12792 264480 12844
rect 265532 12869 265541 12903
rect 265541 12869 265575 12903
rect 265575 12869 265584 12903
rect 265532 12860 265584 12869
rect 266544 12860 266596 12912
rect 257160 12724 257212 12776
rect 262312 12724 262364 12776
rect 271052 12860 271104 12912
rect 271788 12903 271840 12912
rect 271788 12869 271797 12903
rect 271797 12869 271831 12903
rect 271831 12869 271840 12903
rect 271788 12860 271840 12869
rect 272800 12860 272852 12912
rect 273168 12860 273220 12912
rect 268292 12792 268344 12844
rect 269028 12792 269080 12844
rect 257068 12656 257120 12708
rect 262680 12699 262732 12708
rect 252008 12588 252060 12597
rect 262220 12588 262272 12640
rect 262680 12665 262689 12699
rect 262689 12665 262723 12699
rect 262723 12665 262732 12699
rect 262680 12656 262732 12665
rect 267004 12724 267056 12776
rect 267556 12724 267608 12776
rect 268016 12767 268068 12776
rect 268016 12733 268025 12767
rect 268025 12733 268059 12767
rect 268059 12733 268068 12767
rect 268016 12724 268068 12733
rect 268384 12724 268436 12776
rect 270868 12792 270920 12844
rect 272616 12792 272668 12844
rect 295892 12860 295944 12912
rect 302608 12937 302617 12971
rect 302617 12937 302651 12971
rect 302651 12937 302660 12971
rect 302608 12928 302660 12937
rect 305368 12928 305420 12980
rect 305000 12903 305052 12912
rect 269396 12767 269448 12776
rect 269396 12733 269405 12767
rect 269405 12733 269439 12767
rect 269439 12733 269448 12767
rect 269396 12724 269448 12733
rect 263508 12656 263560 12708
rect 263968 12631 264020 12640
rect 263968 12597 263977 12631
rect 263977 12597 264011 12631
rect 264011 12597 264020 12631
rect 263968 12588 264020 12597
rect 267004 12631 267056 12640
rect 267004 12597 267013 12631
rect 267013 12597 267047 12631
rect 267047 12597 267056 12631
rect 267004 12588 267056 12597
rect 267096 12588 267148 12640
rect 267556 12588 267608 12640
rect 269120 12588 269172 12640
rect 272248 12724 272300 12776
rect 272892 12724 272944 12776
rect 272800 12656 272852 12708
rect 273168 12724 273220 12776
rect 290280 12792 290332 12844
rect 302792 12835 302844 12844
rect 302792 12801 302801 12835
rect 302801 12801 302835 12835
rect 302835 12801 302844 12835
rect 302792 12792 302844 12801
rect 305000 12869 305009 12903
rect 305009 12869 305043 12903
rect 305043 12869 305052 12903
rect 305460 12903 305512 12912
rect 305000 12860 305052 12869
rect 305460 12869 305469 12903
rect 305469 12869 305503 12903
rect 305503 12869 305512 12903
rect 305460 12860 305512 12869
rect 270868 12631 270920 12640
rect 270868 12597 270877 12631
rect 270877 12597 270911 12631
rect 270911 12597 270920 12631
rect 270868 12588 270920 12597
rect 271144 12588 271196 12640
rect 272524 12631 272576 12640
rect 272524 12597 272533 12631
rect 272533 12597 272567 12631
rect 272567 12597 272576 12631
rect 272524 12588 272576 12597
rect 272616 12588 272668 12640
rect 281080 12588 281132 12640
rect 39049 12486 39101 12538
rect 39113 12486 39165 12538
rect 39177 12486 39229 12538
rect 39241 12486 39293 12538
rect 39305 12486 39357 12538
rect 115247 12486 115299 12538
rect 115311 12486 115363 12538
rect 115375 12486 115427 12538
rect 115439 12486 115491 12538
rect 115503 12486 115555 12538
rect 191445 12486 191497 12538
rect 191509 12486 191561 12538
rect 191573 12486 191625 12538
rect 191637 12486 191689 12538
rect 191701 12486 191753 12538
rect 267643 12486 267695 12538
rect 267707 12486 267759 12538
rect 267771 12486 267823 12538
rect 267835 12486 267887 12538
rect 267899 12486 267951 12538
rect 26976 12384 27028 12436
rect 28080 12384 28132 12436
rect 14280 12316 14332 12368
rect 28816 12384 28868 12436
rect 32588 12384 32640 12436
rect 34520 12384 34572 12436
rect 35992 12384 36044 12436
rect 4804 12044 4856 12096
rect 26884 12248 26936 12300
rect 28080 12248 28132 12300
rect 28724 12291 28776 12300
rect 28724 12257 28733 12291
rect 28733 12257 28767 12291
rect 28767 12257 28776 12291
rect 28724 12248 28776 12257
rect 34888 12316 34940 12368
rect 37832 12384 37884 12436
rect 38936 12384 38988 12436
rect 39396 12384 39448 12436
rect 40960 12384 41012 12436
rect 43168 12427 43220 12436
rect 43168 12393 43177 12427
rect 43177 12393 43211 12427
rect 43211 12393 43220 12427
rect 43168 12384 43220 12393
rect 43812 12427 43864 12436
rect 43812 12393 43821 12427
rect 43821 12393 43855 12427
rect 43855 12393 43864 12427
rect 43812 12384 43864 12393
rect 54024 12384 54076 12436
rect 55496 12384 55548 12436
rect 56692 12384 56744 12436
rect 57980 12427 58032 12436
rect 57980 12393 57989 12427
rect 57989 12393 58023 12427
rect 58023 12393 58032 12427
rect 57980 12384 58032 12393
rect 75092 12384 75144 12436
rect 79324 12427 79376 12436
rect 29000 12248 29052 12300
rect 29552 12291 29604 12300
rect 29552 12257 29561 12291
rect 29561 12257 29595 12291
rect 29595 12257 29604 12291
rect 29552 12248 29604 12257
rect 17040 12180 17092 12232
rect 27436 12223 27488 12232
rect 27436 12189 27445 12223
rect 27445 12189 27479 12223
rect 27479 12189 27488 12223
rect 27436 12180 27488 12189
rect 29368 12180 29420 12232
rect 34152 12223 34204 12232
rect 34152 12189 34161 12223
rect 34161 12189 34195 12223
rect 34195 12189 34204 12223
rect 34152 12180 34204 12189
rect 34704 12223 34756 12232
rect 34704 12189 34713 12223
rect 34713 12189 34747 12223
rect 34747 12189 34756 12223
rect 35348 12223 35400 12232
rect 34704 12180 34756 12189
rect 35348 12189 35357 12223
rect 35357 12189 35391 12223
rect 35391 12189 35400 12223
rect 35348 12180 35400 12189
rect 27068 12087 27120 12096
rect 27068 12053 27077 12087
rect 27077 12053 27111 12087
rect 27111 12053 27120 12087
rect 27068 12044 27120 12053
rect 27160 12044 27212 12096
rect 27988 12044 28040 12096
rect 29460 12112 29512 12164
rect 29828 12155 29880 12164
rect 29828 12121 29837 12155
rect 29837 12121 29871 12155
rect 29871 12121 29880 12155
rect 29828 12112 29880 12121
rect 31208 12112 31260 12164
rect 32036 12155 32088 12164
rect 32036 12121 32045 12155
rect 32045 12121 32079 12155
rect 32079 12121 32088 12155
rect 32036 12112 32088 12121
rect 43720 12316 43772 12368
rect 40960 12248 41012 12300
rect 38016 12180 38068 12232
rect 40316 12180 40368 12232
rect 40592 12223 40644 12232
rect 40592 12189 40601 12223
rect 40601 12189 40635 12223
rect 40635 12189 40644 12223
rect 40592 12180 40644 12189
rect 76012 12316 76064 12368
rect 53840 12248 53892 12300
rect 43720 12223 43772 12232
rect 43720 12189 43729 12223
rect 43729 12189 43763 12223
rect 43763 12189 43772 12223
rect 43720 12180 43772 12189
rect 41604 12112 41656 12164
rect 41788 12112 41840 12164
rect 28908 12044 28960 12096
rect 31116 12044 31168 12096
rect 32312 12044 32364 12096
rect 32956 12044 33008 12096
rect 36452 12087 36504 12096
rect 36452 12053 36461 12087
rect 36461 12053 36495 12087
rect 36495 12053 36504 12087
rect 36452 12044 36504 12053
rect 40500 12044 40552 12096
rect 40684 12087 40736 12096
rect 40684 12053 40693 12087
rect 40693 12053 40727 12087
rect 40727 12053 40736 12087
rect 40684 12044 40736 12053
rect 56416 12248 56468 12300
rect 74816 12248 74868 12300
rect 77208 12316 77260 12368
rect 78404 12316 78456 12368
rect 55312 12180 55364 12232
rect 56508 12180 56560 12232
rect 76932 12291 76984 12300
rect 76932 12257 76941 12291
rect 76941 12257 76975 12291
rect 76975 12257 76984 12291
rect 78128 12291 78180 12300
rect 76932 12248 76984 12257
rect 78128 12257 78137 12291
rect 78137 12257 78171 12291
rect 78171 12257 78180 12291
rect 78128 12248 78180 12257
rect 52644 12155 52696 12164
rect 52644 12121 52653 12155
rect 52653 12121 52687 12155
rect 52687 12121 52696 12155
rect 52644 12112 52696 12121
rect 53104 12112 53156 12164
rect 77944 12223 77996 12232
rect 77944 12189 77953 12223
rect 77953 12189 77987 12223
rect 77987 12189 77996 12223
rect 77944 12180 77996 12189
rect 79324 12393 79333 12427
rect 79333 12393 79367 12427
rect 79367 12393 79376 12427
rect 79324 12384 79376 12393
rect 80520 12384 80572 12436
rect 85488 12384 85540 12436
rect 86408 12427 86460 12436
rect 86408 12393 86417 12427
rect 86417 12393 86451 12427
rect 86451 12393 86460 12427
rect 86408 12384 86460 12393
rect 87880 12384 87932 12436
rect 90180 12427 90232 12436
rect 90180 12393 90189 12427
rect 90189 12393 90223 12427
rect 90223 12393 90232 12427
rect 90180 12384 90232 12393
rect 99472 12384 99524 12436
rect 99932 12384 99984 12436
rect 104992 12384 105044 12436
rect 105176 12427 105228 12436
rect 105176 12393 105185 12427
rect 105185 12393 105219 12427
rect 105219 12393 105228 12427
rect 105176 12384 105228 12393
rect 112536 12384 112588 12436
rect 115020 12384 115072 12436
rect 116952 12384 117004 12436
rect 127808 12384 127860 12436
rect 129096 12384 129148 12436
rect 130936 12384 130988 12436
rect 132408 12384 132460 12436
rect 147772 12384 147824 12436
rect 152464 12384 152516 12436
rect 78588 12180 78640 12232
rect 86132 12316 86184 12368
rect 87420 12316 87472 12368
rect 81440 12248 81492 12300
rect 84660 12291 84712 12300
rect 84660 12257 84669 12291
rect 84669 12257 84703 12291
rect 84703 12257 84712 12291
rect 84660 12248 84712 12257
rect 83832 12180 83884 12232
rect 85764 12248 85816 12300
rect 86316 12248 86368 12300
rect 88156 12291 88208 12300
rect 88156 12257 88165 12291
rect 88165 12257 88199 12291
rect 88199 12257 88208 12291
rect 88156 12248 88208 12257
rect 85488 12223 85540 12232
rect 85488 12189 85497 12223
rect 85497 12189 85531 12223
rect 85531 12189 85540 12223
rect 85488 12180 85540 12189
rect 86040 12180 86092 12232
rect 88248 12180 88300 12232
rect 89168 12248 89220 12300
rect 88984 12180 89036 12232
rect 92020 12180 92072 12232
rect 99104 12248 99156 12300
rect 102048 12248 102100 12300
rect 103244 12248 103296 12300
rect 103336 12248 103388 12300
rect 115756 12316 115808 12368
rect 97540 12180 97592 12232
rect 103704 12180 103756 12232
rect 100760 12155 100812 12164
rect 55864 12044 55916 12096
rect 56048 12087 56100 12096
rect 56048 12053 56057 12087
rect 56057 12053 56091 12087
rect 56091 12053 56100 12087
rect 56048 12044 56100 12053
rect 57336 12044 57388 12096
rect 76288 12087 76340 12096
rect 76288 12053 76297 12087
rect 76297 12053 76331 12087
rect 76331 12053 76340 12087
rect 76288 12044 76340 12053
rect 80244 12044 80296 12096
rect 84016 12087 84068 12096
rect 84016 12053 84025 12087
rect 84025 12053 84059 12087
rect 84059 12053 84068 12087
rect 84016 12044 84068 12053
rect 84660 12044 84712 12096
rect 86316 12044 86368 12096
rect 87512 12044 87564 12096
rect 87788 12044 87840 12096
rect 87972 12044 88024 12096
rect 88708 12044 88760 12096
rect 100760 12121 100769 12155
rect 100769 12121 100803 12155
rect 100803 12121 100812 12155
rect 100760 12112 100812 12121
rect 101036 12112 101088 12164
rect 101956 12155 102008 12164
rect 101956 12121 101965 12155
rect 101965 12121 101999 12155
rect 101999 12121 102008 12155
rect 101956 12112 102008 12121
rect 102140 12155 102192 12164
rect 102140 12121 102149 12155
rect 102149 12121 102183 12155
rect 102183 12121 102192 12155
rect 111892 12180 111944 12232
rect 114284 12180 114336 12232
rect 118884 12248 118936 12300
rect 141976 12316 142028 12368
rect 147588 12316 147640 12368
rect 151636 12316 151688 12368
rect 102140 12112 102192 12121
rect 113824 12112 113876 12164
rect 100392 12087 100444 12096
rect 100392 12053 100401 12087
rect 100401 12053 100435 12087
rect 100435 12053 100444 12087
rect 100392 12044 100444 12053
rect 102324 12044 102376 12096
rect 102600 12087 102652 12096
rect 102600 12053 102609 12087
rect 102609 12053 102643 12087
rect 102643 12053 102652 12087
rect 102600 12044 102652 12053
rect 103060 12087 103112 12096
rect 103060 12053 103069 12087
rect 103069 12053 103103 12087
rect 103103 12053 103112 12087
rect 103060 12044 103112 12053
rect 113916 12044 113968 12096
rect 115664 12044 115716 12096
rect 116400 12044 116452 12096
rect 118056 12180 118108 12232
rect 118332 12223 118384 12232
rect 118332 12189 118341 12223
rect 118341 12189 118375 12223
rect 118375 12189 118384 12223
rect 118332 12180 118384 12189
rect 126152 12180 126204 12232
rect 128636 12223 128688 12232
rect 128636 12189 128645 12223
rect 128645 12189 128679 12223
rect 128679 12189 128688 12223
rect 128636 12180 128688 12189
rect 131028 12248 131080 12300
rect 133236 12248 133288 12300
rect 149060 12248 149112 12300
rect 118240 12112 118292 12164
rect 130476 12180 130528 12232
rect 132408 12180 132460 12232
rect 132592 12223 132644 12232
rect 132592 12189 132601 12223
rect 132601 12189 132635 12223
rect 132635 12189 132644 12223
rect 132592 12180 132644 12189
rect 137744 12223 137796 12232
rect 137744 12189 137753 12223
rect 137753 12189 137787 12223
rect 137787 12189 137796 12223
rect 137744 12180 137796 12189
rect 148048 12180 148100 12232
rect 149336 12180 149388 12232
rect 149428 12223 149480 12232
rect 149428 12189 149437 12223
rect 149437 12189 149471 12223
rect 149471 12189 149480 12223
rect 149428 12180 149480 12189
rect 151360 12180 151412 12232
rect 152740 12316 152792 12368
rect 132500 12112 132552 12164
rect 138020 12155 138072 12164
rect 138020 12121 138029 12155
rect 138029 12121 138063 12155
rect 138063 12121 138072 12155
rect 138020 12112 138072 12121
rect 153752 12384 153804 12436
rect 157248 12384 157300 12436
rect 160928 12384 160980 12436
rect 161572 12384 161624 12436
rect 155040 12316 155092 12368
rect 158904 12316 158956 12368
rect 166448 12384 166500 12436
rect 176476 12384 176528 12436
rect 179512 12384 179564 12436
rect 189172 12384 189224 12436
rect 189632 12384 189684 12436
rect 190828 12384 190880 12436
rect 194048 12384 194100 12436
rect 165436 12316 165488 12368
rect 166080 12359 166132 12368
rect 166080 12325 166089 12359
rect 166089 12325 166123 12359
rect 166123 12325 166132 12359
rect 166080 12316 166132 12325
rect 154120 12248 154172 12300
rect 160376 12248 160428 12300
rect 161480 12291 161532 12300
rect 161480 12257 161489 12291
rect 161489 12257 161523 12291
rect 161523 12257 161532 12291
rect 162492 12291 162544 12300
rect 161480 12248 161532 12257
rect 162492 12257 162501 12291
rect 162501 12257 162535 12291
rect 162535 12257 162544 12291
rect 162492 12248 162544 12257
rect 162676 12291 162728 12300
rect 162676 12257 162685 12291
rect 162685 12257 162719 12291
rect 162719 12257 162728 12291
rect 162676 12248 162728 12257
rect 163596 12291 163648 12300
rect 163596 12257 163605 12291
rect 163605 12257 163639 12291
rect 163639 12257 163648 12291
rect 163596 12248 163648 12257
rect 177764 12316 177816 12368
rect 180892 12359 180944 12368
rect 180892 12325 180901 12359
rect 180901 12325 180935 12359
rect 180935 12325 180944 12359
rect 180892 12316 180944 12325
rect 192576 12359 192628 12368
rect 177120 12291 177172 12300
rect 177120 12257 177129 12291
rect 177129 12257 177163 12291
rect 177163 12257 177172 12291
rect 177120 12248 177172 12257
rect 158812 12180 158864 12232
rect 161756 12180 161808 12232
rect 187976 12248 188028 12300
rect 177856 12180 177908 12232
rect 179144 12223 179196 12232
rect 179144 12189 179153 12223
rect 179153 12189 179187 12223
rect 179187 12189 179196 12223
rect 179144 12180 179196 12189
rect 180708 12180 180760 12232
rect 189540 12223 189592 12232
rect 131580 12044 131632 12096
rect 155868 12112 155920 12164
rect 156420 12112 156472 12164
rect 162584 12112 162636 12164
rect 162676 12112 162728 12164
rect 164332 12112 164384 12164
rect 165896 12155 165948 12164
rect 165896 12121 165905 12155
rect 165905 12121 165939 12155
rect 165939 12121 165948 12155
rect 165896 12112 165948 12121
rect 166540 12112 166592 12164
rect 179420 12155 179472 12164
rect 149520 12044 149572 12096
rect 151636 12087 151688 12096
rect 151636 12053 151645 12087
rect 151645 12053 151679 12087
rect 151679 12053 151688 12087
rect 151636 12044 151688 12053
rect 151728 12044 151780 12096
rect 152188 12044 152240 12096
rect 152556 12044 152608 12096
rect 161112 12044 161164 12096
rect 162216 12044 162268 12096
rect 162860 12044 162912 12096
rect 176660 12044 176712 12096
rect 178040 12087 178092 12096
rect 178040 12053 178049 12087
rect 178049 12053 178083 12087
rect 178083 12053 178092 12087
rect 178040 12044 178092 12053
rect 179420 12121 179429 12155
rect 179429 12121 179463 12155
rect 179463 12121 179472 12155
rect 179420 12112 179472 12121
rect 181444 12112 181496 12164
rect 189540 12189 189549 12223
rect 189549 12189 189583 12223
rect 189583 12189 189592 12223
rect 189540 12180 189592 12189
rect 192576 12325 192585 12359
rect 192585 12325 192619 12359
rect 192619 12325 192628 12359
rect 192576 12316 192628 12325
rect 191840 12248 191892 12300
rect 192668 12248 192720 12300
rect 194416 12223 194468 12232
rect 190828 12112 190880 12164
rect 191104 12155 191156 12164
rect 191104 12121 191113 12155
rect 191113 12121 191147 12155
rect 191147 12121 191156 12155
rect 191104 12112 191156 12121
rect 191196 12112 191248 12164
rect 180156 12044 180208 12096
rect 193404 12155 193456 12164
rect 193404 12121 193413 12155
rect 193413 12121 193447 12155
rect 193447 12121 193456 12155
rect 193404 12112 193456 12121
rect 193036 12087 193088 12096
rect 193036 12053 193045 12087
rect 193045 12053 193079 12087
rect 193079 12053 193088 12087
rect 193036 12044 193088 12053
rect 193680 12044 193732 12096
rect 194416 12189 194425 12223
rect 194425 12189 194459 12223
rect 194459 12189 194468 12223
rect 194416 12180 194468 12189
rect 194692 12155 194744 12164
rect 194692 12121 194701 12155
rect 194701 12121 194735 12155
rect 194735 12121 194744 12155
rect 194692 12112 194744 12121
rect 197452 12316 197504 12368
rect 202420 12384 202472 12436
rect 205640 12384 205692 12436
rect 207664 12384 207716 12436
rect 230112 12384 230164 12436
rect 231860 12384 231912 12436
rect 239036 12384 239088 12436
rect 240140 12384 240192 12436
rect 228824 12316 228876 12368
rect 231124 12316 231176 12368
rect 232504 12316 232556 12368
rect 194968 12044 195020 12096
rect 200488 12248 200540 12300
rect 197452 12223 197504 12232
rect 197452 12189 197461 12223
rect 197461 12189 197495 12223
rect 197495 12189 197504 12223
rect 197452 12180 197504 12189
rect 198372 12180 198424 12232
rect 200580 12180 200632 12232
rect 201040 12223 201092 12232
rect 201040 12189 201049 12223
rect 201049 12189 201083 12223
rect 201083 12189 201092 12223
rect 201040 12180 201092 12189
rect 202052 12248 202104 12300
rect 203524 12291 203576 12300
rect 203524 12257 203533 12291
rect 203533 12257 203567 12291
rect 203567 12257 203576 12291
rect 203524 12248 203576 12257
rect 204536 12180 204588 12232
rect 229928 12223 229980 12232
rect 229928 12189 229937 12223
rect 229937 12189 229971 12223
rect 229971 12189 229980 12223
rect 229928 12180 229980 12189
rect 231308 12180 231360 12232
rect 204996 12155 205048 12164
rect 204996 12121 205005 12155
rect 205005 12121 205039 12155
rect 205039 12121 205048 12155
rect 204996 12112 205048 12121
rect 196808 12087 196860 12096
rect 196808 12053 196817 12087
rect 196817 12053 196851 12087
rect 196851 12053 196860 12087
rect 196808 12044 196860 12053
rect 196992 12087 197044 12096
rect 196992 12053 197001 12087
rect 197001 12053 197035 12087
rect 197035 12053 197044 12087
rect 196992 12044 197044 12053
rect 197360 12087 197412 12096
rect 197360 12053 197369 12087
rect 197369 12053 197403 12087
rect 197403 12053 197412 12087
rect 197360 12044 197412 12053
rect 203064 12044 203116 12096
rect 203432 12044 203484 12096
rect 204260 12044 204312 12096
rect 230848 12112 230900 12164
rect 231124 12112 231176 12164
rect 231676 12248 231728 12300
rect 238852 12248 238904 12300
rect 239312 12291 239364 12300
rect 239312 12257 239321 12291
rect 239321 12257 239355 12291
rect 239355 12257 239364 12291
rect 239312 12248 239364 12257
rect 232136 12223 232188 12232
rect 232136 12189 232145 12223
rect 232145 12189 232179 12223
rect 232179 12189 232188 12223
rect 232136 12180 232188 12189
rect 233056 12180 233108 12232
rect 238024 12223 238076 12232
rect 238024 12189 238033 12223
rect 238033 12189 238067 12223
rect 238067 12189 238076 12223
rect 238024 12180 238076 12189
rect 238392 12180 238444 12232
rect 239128 12223 239180 12232
rect 239128 12189 239137 12223
rect 239137 12189 239171 12223
rect 239171 12189 239180 12223
rect 239128 12180 239180 12189
rect 239496 12180 239548 12232
rect 239956 12248 240008 12300
rect 242256 12316 242308 12368
rect 242440 12248 242492 12300
rect 242992 12316 243044 12368
rect 242900 12291 242952 12300
rect 242900 12257 242909 12291
rect 242909 12257 242943 12291
rect 242943 12257 242952 12291
rect 242900 12248 242952 12257
rect 242164 12180 242216 12232
rect 243636 12384 243688 12436
rect 244188 12427 244240 12436
rect 244188 12393 244197 12427
rect 244197 12393 244231 12427
rect 244231 12393 244240 12427
rect 244188 12384 244240 12393
rect 251364 12384 251416 12436
rect 251916 12384 251968 12436
rect 251456 12316 251508 12368
rect 252100 12359 252152 12368
rect 252100 12325 252109 12359
rect 252109 12325 252143 12359
rect 252143 12325 252152 12359
rect 252100 12316 252152 12325
rect 254308 12359 254360 12368
rect 254308 12325 254317 12359
rect 254317 12325 254351 12359
rect 254351 12325 254360 12359
rect 254308 12316 254360 12325
rect 255228 12316 255280 12368
rect 243176 12248 243228 12300
rect 248328 12248 248380 12300
rect 249248 12248 249300 12300
rect 251272 12223 251324 12232
rect 251272 12189 251281 12223
rect 251281 12189 251315 12223
rect 251315 12189 251324 12223
rect 251916 12223 251968 12232
rect 251272 12180 251324 12189
rect 251916 12189 251925 12223
rect 251925 12189 251959 12223
rect 251959 12189 251968 12223
rect 251916 12180 251968 12189
rect 255136 12223 255188 12232
rect 255136 12189 255145 12223
rect 255145 12189 255179 12223
rect 255179 12189 255188 12223
rect 255136 12180 255188 12189
rect 249064 12155 249116 12164
rect 228824 12044 228876 12096
rect 231216 12044 231268 12096
rect 249064 12121 249073 12155
rect 249073 12121 249107 12155
rect 249107 12121 249116 12155
rect 249064 12112 249116 12121
rect 249248 12155 249300 12164
rect 249248 12121 249257 12155
rect 249257 12121 249291 12155
rect 249291 12121 249300 12155
rect 249248 12112 249300 12121
rect 253112 12112 253164 12164
rect 255596 12248 255648 12300
rect 256516 12384 256568 12436
rect 262496 12427 262548 12436
rect 262496 12393 262505 12427
rect 262505 12393 262539 12427
rect 262539 12393 262548 12427
rect 262496 12384 262548 12393
rect 265532 12384 265584 12436
rect 256976 12316 257028 12368
rect 264980 12316 265032 12368
rect 268016 12384 268068 12436
rect 268384 12384 268436 12436
rect 271052 12427 271104 12436
rect 271052 12393 271061 12427
rect 271061 12393 271095 12427
rect 271095 12393 271104 12427
rect 271052 12384 271104 12393
rect 305460 12427 305512 12436
rect 305460 12393 305469 12427
rect 305469 12393 305503 12427
rect 305503 12393 305512 12427
rect 305460 12384 305512 12393
rect 261852 12248 261904 12300
rect 262404 12248 262456 12300
rect 256240 12223 256292 12232
rect 256240 12189 256249 12223
rect 256249 12189 256283 12223
rect 256283 12189 256292 12223
rect 256240 12180 256292 12189
rect 256332 12180 256384 12232
rect 263048 12180 263100 12232
rect 264152 12248 264204 12300
rect 265164 12248 265216 12300
rect 264336 12180 264388 12232
rect 265624 12248 265676 12300
rect 269120 12248 269172 12300
rect 269672 12248 269724 12300
rect 271144 12248 271196 12300
rect 272248 12291 272300 12300
rect 272248 12257 272257 12291
rect 272257 12257 272291 12291
rect 272291 12257 272300 12291
rect 272248 12248 272300 12257
rect 272800 12248 272852 12300
rect 231400 12087 231452 12096
rect 231400 12053 231409 12087
rect 231409 12053 231443 12087
rect 231443 12053 231452 12087
rect 231400 12044 231452 12053
rect 231768 12044 231820 12096
rect 233056 12044 233108 12096
rect 240876 12087 240928 12096
rect 240876 12053 240885 12087
rect 240885 12053 240919 12087
rect 240919 12053 240928 12087
rect 240876 12044 240928 12053
rect 241520 12044 241572 12096
rect 242532 12044 242584 12096
rect 244096 12044 244148 12096
rect 254400 12044 254452 12096
rect 255044 12044 255096 12096
rect 255228 12087 255280 12096
rect 255228 12053 255237 12087
rect 255237 12053 255271 12087
rect 255271 12053 255280 12087
rect 255228 12044 255280 12053
rect 256332 12044 256384 12096
rect 265164 12112 265216 12164
rect 268108 12180 268160 12232
rect 268660 12180 268712 12232
rect 266820 12155 266872 12164
rect 266820 12121 266829 12155
rect 266829 12121 266863 12155
rect 266863 12121 266872 12155
rect 266820 12112 266872 12121
rect 267280 12112 267332 12164
rect 268200 12112 268252 12164
rect 269488 12112 269540 12164
rect 267004 12044 267056 12096
rect 268476 12044 268528 12096
rect 268660 12044 268712 12096
rect 271328 12180 271380 12232
rect 272892 12180 272944 12232
rect 270408 12044 270460 12096
rect 284760 12044 284812 12096
rect 77148 11942 77200 11994
rect 77212 11942 77264 11994
rect 77276 11942 77328 11994
rect 77340 11942 77392 11994
rect 77404 11942 77456 11994
rect 153346 11942 153398 11994
rect 153410 11942 153462 11994
rect 153474 11942 153526 11994
rect 153538 11942 153590 11994
rect 153602 11942 153654 11994
rect 229544 11942 229596 11994
rect 229608 11942 229660 11994
rect 229672 11942 229724 11994
rect 229736 11942 229788 11994
rect 229800 11942 229852 11994
rect 29092 11840 29144 11892
rect 29460 11840 29512 11892
rect 30932 11840 30984 11892
rect 32220 11840 32272 11892
rect 33784 11883 33836 11892
rect 33784 11849 33793 11883
rect 33793 11849 33827 11883
rect 33827 11849 33836 11883
rect 33784 11840 33836 11849
rect 34428 11883 34480 11892
rect 34428 11849 34437 11883
rect 34437 11849 34471 11883
rect 34471 11849 34480 11883
rect 34428 11840 34480 11849
rect 38384 11883 38436 11892
rect 27712 11772 27764 11824
rect 28724 11772 28776 11824
rect 29000 11772 29052 11824
rect 28908 11679 28960 11688
rect 28908 11645 28917 11679
rect 28917 11645 28951 11679
rect 28951 11645 28960 11679
rect 28908 11636 28960 11645
rect 30012 11772 30064 11824
rect 32036 11772 32088 11824
rect 38384 11849 38393 11883
rect 38393 11849 38427 11883
rect 38427 11849 38436 11883
rect 38384 11840 38436 11849
rect 39580 11840 39632 11892
rect 29552 11704 29604 11756
rect 32404 11704 32456 11756
rect 29920 11679 29972 11688
rect 29920 11645 29929 11679
rect 29929 11645 29963 11679
rect 29963 11645 29972 11679
rect 29920 11636 29972 11645
rect 28448 11543 28500 11552
rect 28448 11509 28457 11543
rect 28457 11509 28491 11543
rect 28491 11509 28500 11543
rect 28448 11500 28500 11509
rect 32588 11636 32640 11688
rect 34704 11704 34756 11756
rect 39948 11840 40000 11892
rect 41420 11840 41472 11892
rect 42892 11840 42944 11892
rect 52644 11840 52696 11892
rect 53656 11883 53708 11892
rect 53656 11849 53665 11883
rect 53665 11849 53699 11883
rect 53699 11849 53708 11883
rect 53656 11840 53708 11849
rect 54392 11883 54444 11892
rect 54392 11849 54401 11883
rect 54401 11849 54435 11883
rect 54435 11849 54444 11883
rect 54392 11840 54444 11849
rect 55312 11883 55364 11892
rect 55312 11849 55321 11883
rect 55321 11849 55355 11883
rect 55355 11849 55364 11883
rect 55312 11840 55364 11849
rect 56600 11840 56652 11892
rect 58624 11840 58676 11892
rect 75460 11840 75512 11892
rect 75644 11840 75696 11892
rect 76472 11840 76524 11892
rect 77852 11883 77904 11892
rect 77852 11849 77861 11883
rect 77861 11849 77895 11883
rect 77895 11849 77904 11883
rect 77852 11840 77904 11849
rect 78496 11883 78548 11892
rect 78496 11849 78505 11883
rect 78505 11849 78539 11883
rect 78539 11849 78548 11883
rect 78496 11840 78548 11849
rect 84292 11840 84344 11892
rect 86040 11883 86092 11892
rect 34060 11636 34112 11688
rect 31116 11568 31168 11620
rect 40684 11772 40736 11824
rect 41236 11772 41288 11824
rect 53748 11772 53800 11824
rect 40316 11704 40368 11756
rect 42800 11704 42852 11756
rect 42984 11704 43036 11756
rect 53012 11747 53064 11756
rect 40960 11636 41012 11688
rect 41420 11636 41472 11688
rect 53012 11713 53021 11747
rect 53021 11713 53055 11747
rect 53055 11713 53064 11747
rect 53012 11704 53064 11713
rect 57428 11772 57480 11824
rect 84936 11772 84988 11824
rect 54668 11636 54720 11688
rect 55588 11679 55640 11688
rect 55588 11645 55597 11679
rect 55597 11645 55631 11679
rect 55631 11645 55640 11679
rect 55588 11636 55640 11645
rect 55864 11636 55916 11688
rect 76012 11704 76064 11756
rect 76288 11704 76340 11756
rect 78588 11704 78640 11756
rect 81440 11704 81492 11756
rect 86040 11849 86049 11883
rect 86049 11849 86083 11883
rect 86083 11849 86092 11883
rect 86040 11840 86092 11849
rect 86132 11840 86184 11892
rect 87880 11883 87932 11892
rect 87880 11849 87889 11883
rect 87889 11849 87923 11883
rect 87923 11849 87932 11883
rect 87880 11840 87932 11849
rect 89536 11840 89588 11892
rect 99656 11840 99708 11892
rect 100944 11883 100996 11892
rect 100944 11849 100953 11883
rect 100953 11849 100987 11883
rect 100987 11849 100996 11883
rect 100944 11840 100996 11849
rect 103060 11840 103112 11892
rect 103520 11840 103572 11892
rect 113824 11883 113876 11892
rect 85304 11772 85356 11824
rect 113824 11849 113833 11883
rect 113833 11849 113867 11883
rect 113867 11849 113876 11883
rect 113824 11840 113876 11849
rect 114284 11840 114336 11892
rect 115664 11840 115716 11892
rect 116768 11840 116820 11892
rect 117320 11840 117372 11892
rect 118792 11840 118844 11892
rect 129372 11883 129424 11892
rect 129372 11849 129381 11883
rect 129381 11849 129415 11883
rect 129415 11849 129424 11883
rect 129372 11840 129424 11849
rect 130292 11840 130344 11892
rect 130936 11883 130988 11892
rect 130936 11849 130945 11883
rect 130945 11849 130979 11883
rect 130979 11849 130988 11883
rect 130936 11840 130988 11849
rect 131120 11840 131172 11892
rect 137744 11840 137796 11892
rect 151084 11883 151136 11892
rect 75000 11636 75052 11688
rect 76932 11636 76984 11688
rect 84016 11636 84068 11688
rect 85764 11704 85816 11756
rect 86960 11747 87012 11756
rect 86960 11713 86969 11747
rect 86969 11713 87003 11747
rect 87003 11713 87012 11747
rect 86960 11704 87012 11713
rect 86316 11679 86368 11688
rect 86316 11645 86325 11679
rect 86325 11645 86359 11679
rect 86359 11645 86368 11679
rect 86316 11636 86368 11645
rect 89168 11704 89220 11756
rect 100392 11747 100444 11756
rect 100392 11713 100401 11747
rect 100401 11713 100435 11747
rect 100435 11713 100444 11747
rect 100392 11704 100444 11713
rect 102140 11704 102192 11756
rect 103612 11704 103664 11756
rect 56048 11568 56100 11620
rect 90456 11636 90508 11688
rect 100760 11636 100812 11688
rect 102048 11679 102100 11688
rect 102048 11645 102057 11679
rect 102057 11645 102091 11679
rect 102091 11645 102100 11679
rect 102048 11636 102100 11645
rect 102324 11636 102376 11688
rect 103520 11636 103572 11688
rect 114560 11772 114612 11824
rect 114008 11747 114060 11756
rect 114008 11713 114017 11747
rect 114017 11713 114051 11747
rect 114051 11713 114060 11747
rect 114008 11704 114060 11713
rect 138020 11772 138072 11824
rect 149980 11772 150032 11824
rect 151084 11849 151093 11883
rect 151093 11849 151127 11883
rect 151127 11849 151136 11883
rect 151084 11840 151136 11849
rect 152004 11883 152056 11892
rect 152004 11849 152013 11883
rect 152013 11849 152047 11883
rect 152047 11849 152056 11883
rect 152004 11840 152056 11849
rect 154212 11840 154264 11892
rect 115020 11704 115072 11756
rect 116400 11747 116452 11756
rect 116400 11713 116409 11747
rect 116409 11713 116443 11747
rect 116443 11713 116452 11747
rect 116400 11704 116452 11713
rect 115664 11636 115716 11688
rect 115756 11636 115808 11688
rect 118332 11704 118384 11756
rect 128360 11704 128412 11756
rect 130292 11704 130344 11756
rect 131580 11704 131632 11756
rect 129740 11636 129792 11688
rect 131028 11679 131080 11688
rect 131028 11645 131037 11679
rect 131037 11645 131071 11679
rect 131071 11645 131080 11679
rect 131028 11636 131080 11645
rect 132500 11704 132552 11756
rect 147680 11704 147732 11756
rect 151268 11747 151320 11756
rect 151268 11713 151277 11747
rect 151277 11713 151311 11747
rect 151311 11713 151320 11747
rect 151268 11704 151320 11713
rect 152188 11747 152240 11756
rect 152188 11713 152197 11747
rect 152197 11713 152231 11747
rect 152231 11713 152240 11747
rect 152188 11704 152240 11713
rect 152740 11704 152792 11756
rect 161112 11747 161164 11756
rect 161112 11713 161121 11747
rect 161121 11713 161155 11747
rect 161155 11713 161164 11747
rect 161112 11704 161164 11713
rect 161756 11747 161808 11756
rect 161756 11713 161765 11747
rect 161765 11713 161799 11747
rect 161799 11713 161808 11747
rect 161756 11704 161808 11713
rect 137744 11636 137796 11688
rect 148324 11679 148376 11688
rect 148324 11645 148333 11679
rect 148333 11645 148367 11679
rect 148367 11645 148376 11679
rect 148324 11636 148376 11645
rect 148600 11679 148652 11688
rect 148600 11645 148609 11679
rect 148609 11645 148643 11679
rect 148643 11645 148652 11679
rect 148600 11636 148652 11645
rect 143264 11568 143316 11620
rect 146024 11568 146076 11620
rect 161204 11568 161256 11620
rect 161296 11568 161348 11620
rect 162032 11840 162084 11892
rect 162768 11840 162820 11892
rect 163780 11840 163832 11892
rect 164332 11840 164384 11892
rect 164884 11883 164936 11892
rect 164884 11849 164893 11883
rect 164893 11849 164927 11883
rect 164927 11849 164936 11883
rect 164884 11840 164936 11849
rect 176752 11840 176804 11892
rect 177396 11840 177448 11892
rect 177856 11840 177908 11892
rect 179880 11840 179932 11892
rect 179972 11840 180024 11892
rect 180156 11840 180208 11892
rect 188344 11840 188396 11892
rect 191748 11840 191800 11892
rect 191840 11840 191892 11892
rect 162584 11772 162636 11824
rect 189540 11772 189592 11824
rect 193864 11772 193916 11824
rect 163688 11747 163740 11756
rect 163688 11713 163697 11747
rect 163697 11713 163731 11747
rect 163731 11713 163740 11747
rect 163688 11704 163740 11713
rect 163504 11636 163556 11688
rect 166632 11704 166684 11756
rect 176660 11747 176712 11756
rect 176660 11713 176669 11747
rect 176669 11713 176703 11747
rect 176703 11713 176712 11747
rect 176660 11704 176712 11713
rect 179880 11704 179932 11756
rect 177120 11636 177172 11688
rect 165896 11568 165948 11620
rect 31392 11543 31444 11552
rect 31392 11509 31401 11543
rect 31401 11509 31435 11543
rect 31435 11509 31444 11543
rect 31392 11500 31444 11509
rect 32956 11500 33008 11552
rect 55496 11500 55548 11552
rect 84844 11500 84896 11552
rect 86408 11500 86460 11552
rect 101864 11500 101916 11552
rect 104072 11500 104124 11552
rect 114008 11500 114060 11552
rect 131856 11543 131908 11552
rect 131856 11509 131865 11543
rect 131865 11509 131899 11543
rect 131899 11509 131908 11543
rect 131856 11500 131908 11509
rect 147312 11500 147364 11552
rect 151728 11500 151780 11552
rect 180064 11704 180116 11756
rect 180616 11704 180668 11756
rect 180800 11636 180852 11688
rect 181536 11636 181588 11688
rect 189632 11747 189684 11756
rect 189632 11713 189641 11747
rect 189641 11713 189675 11747
rect 189675 11713 189684 11747
rect 189632 11704 189684 11713
rect 190828 11704 190880 11756
rect 191840 11747 191892 11756
rect 191840 11713 191849 11747
rect 191849 11713 191883 11747
rect 191883 11713 191892 11747
rect 191840 11704 191892 11713
rect 194416 11840 194468 11892
rect 194692 11840 194744 11892
rect 202880 11883 202932 11892
rect 202880 11849 202889 11883
rect 202889 11849 202923 11883
rect 202923 11849 202932 11883
rect 202880 11840 202932 11849
rect 204536 11840 204588 11892
rect 206560 11840 206612 11892
rect 227812 11840 227864 11892
rect 228824 11840 228876 11892
rect 196808 11772 196860 11824
rect 203156 11772 203208 11824
rect 205548 11772 205600 11824
rect 227720 11772 227772 11824
rect 229928 11840 229980 11892
rect 230388 11883 230440 11892
rect 230388 11849 230397 11883
rect 230397 11849 230431 11883
rect 230431 11849 230440 11883
rect 230388 11840 230440 11849
rect 231032 11840 231084 11892
rect 231676 11840 231728 11892
rect 240324 11883 240376 11892
rect 240324 11849 240333 11883
rect 240333 11849 240367 11883
rect 240367 11849 240376 11883
rect 240324 11840 240376 11849
rect 241060 11883 241112 11892
rect 241060 11849 241069 11883
rect 241069 11849 241103 11883
rect 241103 11849 241112 11883
rect 241060 11840 241112 11849
rect 241796 11883 241848 11892
rect 241796 11849 241805 11883
rect 241805 11849 241839 11883
rect 241839 11849 241848 11883
rect 241796 11840 241848 11849
rect 252928 11840 252980 11892
rect 254676 11840 254728 11892
rect 254768 11840 254820 11892
rect 255044 11840 255096 11892
rect 266820 11840 266872 11892
rect 197912 11704 197964 11756
rect 201040 11704 201092 11756
rect 203064 11747 203116 11756
rect 203064 11713 203073 11747
rect 203073 11713 203107 11747
rect 203107 11713 203116 11747
rect 203064 11704 203116 11713
rect 192116 11679 192168 11688
rect 192116 11645 192125 11679
rect 192125 11645 192159 11679
rect 192159 11645 192168 11679
rect 192116 11636 192168 11645
rect 194324 11679 194376 11688
rect 194324 11645 194333 11679
rect 194333 11645 194367 11679
rect 194367 11645 194376 11679
rect 194324 11636 194376 11645
rect 194416 11636 194468 11688
rect 180340 11568 180392 11620
rect 197360 11636 197412 11688
rect 201316 11636 201368 11688
rect 202880 11636 202932 11688
rect 206376 11704 206428 11756
rect 230848 11772 230900 11824
rect 229376 11704 229428 11756
rect 240140 11772 240192 11824
rect 203524 11636 203576 11688
rect 207848 11636 207900 11688
rect 227260 11636 227312 11688
rect 180524 11500 180576 11552
rect 189448 11543 189500 11552
rect 189448 11509 189457 11543
rect 189457 11509 189491 11543
rect 189491 11509 189500 11543
rect 189448 11500 189500 11509
rect 197452 11568 197504 11620
rect 203432 11568 203484 11620
rect 204904 11568 204956 11620
rect 230296 11568 230348 11620
rect 193312 11500 193364 11552
rect 193496 11500 193548 11552
rect 195796 11500 195848 11552
rect 195888 11500 195940 11552
rect 196992 11500 197044 11552
rect 201500 11500 201552 11552
rect 204812 11543 204864 11552
rect 204812 11509 204821 11543
rect 204821 11509 204855 11543
rect 204855 11509 204864 11543
rect 204812 11500 204864 11509
rect 229376 11500 229428 11552
rect 231216 11704 231268 11756
rect 241520 11772 241572 11824
rect 239312 11636 239364 11688
rect 239956 11636 240008 11688
rect 232136 11568 232188 11620
rect 242532 11747 242584 11756
rect 242532 11713 242541 11747
rect 242541 11713 242575 11747
rect 242575 11713 242584 11747
rect 242532 11704 242584 11713
rect 241980 11636 242032 11688
rect 244832 11772 244884 11824
rect 254308 11772 254360 11824
rect 270684 11840 270736 11892
rect 270776 11840 270828 11892
rect 268292 11772 268344 11824
rect 269856 11772 269908 11824
rect 252008 11747 252060 11756
rect 252008 11713 252017 11747
rect 252017 11713 252051 11747
rect 252051 11713 252060 11747
rect 252008 11704 252060 11713
rect 252744 11747 252796 11756
rect 252744 11713 252753 11747
rect 252753 11713 252787 11747
rect 252787 11713 252796 11747
rect 252744 11704 252796 11713
rect 253020 11704 253072 11756
rect 256240 11704 256292 11756
rect 257252 11704 257304 11756
rect 264336 11747 264388 11756
rect 264336 11713 264345 11747
rect 264345 11713 264379 11747
rect 264379 11713 264388 11747
rect 264336 11704 264388 11713
rect 265164 11747 265216 11756
rect 265164 11713 265173 11747
rect 265173 11713 265207 11747
rect 265207 11713 265216 11747
rect 265164 11704 265216 11713
rect 265256 11704 265308 11756
rect 242716 11636 242768 11688
rect 244556 11636 244608 11688
rect 252100 11636 252152 11688
rect 255596 11636 255648 11688
rect 256424 11636 256476 11688
rect 263968 11636 264020 11688
rect 268476 11704 268528 11756
rect 269120 11747 269172 11756
rect 269120 11713 269129 11747
rect 269129 11713 269163 11747
rect 269163 11713 269172 11747
rect 269120 11704 269172 11713
rect 271328 11747 271380 11756
rect 271328 11713 271337 11747
rect 271337 11713 271371 11747
rect 271371 11713 271380 11747
rect 271328 11704 271380 11713
rect 231676 11500 231728 11552
rect 239404 11500 239456 11552
rect 241244 11500 241296 11552
rect 251640 11568 251692 11620
rect 249064 11500 249116 11552
rect 253296 11500 253348 11552
rect 268016 11568 268068 11620
rect 261760 11500 261812 11552
rect 262680 11500 262732 11552
rect 266268 11500 266320 11552
rect 266360 11500 266412 11552
rect 269396 11679 269448 11688
rect 269396 11645 269405 11679
rect 269405 11645 269439 11679
rect 269439 11645 269448 11679
rect 269396 11636 269448 11645
rect 269948 11636 270000 11688
rect 273168 11636 273220 11688
rect 275100 11500 275152 11552
rect 39049 11398 39101 11450
rect 39113 11398 39165 11450
rect 39177 11398 39229 11450
rect 39241 11398 39293 11450
rect 39305 11398 39357 11450
rect 115247 11398 115299 11450
rect 115311 11398 115363 11450
rect 115375 11398 115427 11450
rect 115439 11398 115491 11450
rect 115503 11398 115555 11450
rect 191445 11398 191497 11450
rect 191509 11398 191561 11450
rect 191573 11398 191625 11450
rect 191637 11398 191689 11450
rect 191701 11398 191753 11450
rect 267643 11398 267695 11450
rect 267707 11398 267759 11450
rect 267771 11398 267823 11450
rect 267835 11398 267887 11450
rect 267899 11398 267951 11450
rect 29920 11296 29972 11348
rect 30012 11296 30064 11348
rect 28908 11228 28960 11280
rect 32404 11296 32456 11348
rect 33324 11296 33376 11348
rect 33600 11339 33652 11348
rect 33600 11305 33609 11339
rect 33609 11305 33643 11339
rect 33643 11305 33652 11339
rect 33600 11296 33652 11305
rect 40408 11296 40460 11348
rect 41052 11339 41104 11348
rect 41052 11305 41061 11339
rect 41061 11305 41095 11339
rect 41095 11305 41104 11339
rect 41052 11296 41104 11305
rect 41604 11339 41656 11348
rect 41604 11305 41613 11339
rect 41613 11305 41647 11339
rect 41647 11305 41656 11339
rect 41604 11296 41656 11305
rect 55036 11296 55088 11348
rect 57704 11296 57756 11348
rect 76380 11296 76432 11348
rect 78772 11296 78824 11348
rect 84476 11296 84528 11348
rect 87144 11296 87196 11348
rect 89076 11296 89128 11348
rect 102876 11339 102928 11348
rect 102876 11305 102885 11339
rect 102885 11305 102919 11339
rect 102919 11305 102928 11339
rect 102876 11296 102928 11305
rect 115112 11296 115164 11348
rect 117688 11296 117740 11348
rect 130384 11296 130436 11348
rect 131212 11339 131264 11348
rect 131212 11305 131221 11339
rect 131221 11305 131255 11339
rect 131255 11305 131264 11339
rect 131212 11296 131264 11305
rect 132868 11296 132920 11348
rect 148048 11339 148100 11348
rect 148048 11305 148057 11339
rect 148057 11305 148091 11339
rect 148091 11305 148100 11339
rect 148048 11296 148100 11305
rect 150808 11339 150860 11348
rect 150808 11305 150817 11339
rect 150817 11305 150851 11339
rect 150851 11305 150860 11339
rect 150808 11296 150860 11305
rect 157248 11296 157300 11348
rect 162124 11296 162176 11348
rect 162676 11339 162728 11348
rect 162676 11305 162685 11339
rect 162685 11305 162719 11339
rect 162719 11305 162728 11339
rect 162676 11296 162728 11305
rect 163412 11296 163464 11348
rect 165896 11296 165948 11348
rect 239404 11296 239456 11348
rect 239772 11296 239824 11348
rect 240048 11296 240100 11348
rect 240968 11296 241020 11348
rect 242072 11296 242124 11348
rect 252468 11296 252520 11348
rect 253112 11339 253164 11348
rect 253112 11305 253121 11339
rect 253121 11305 253155 11339
rect 253155 11305 253164 11339
rect 253112 11296 253164 11305
rect 254032 11296 254084 11348
rect 265440 11296 265492 11348
rect 266268 11296 266320 11348
rect 27068 11160 27120 11212
rect 29460 11160 29512 11212
rect 29552 11160 29604 11212
rect 36452 11228 36504 11280
rect 41328 11228 41380 11280
rect 86776 11228 86828 11280
rect 102232 11228 102284 11280
rect 114192 11228 114244 11280
rect 147404 11228 147456 11280
rect 31392 11160 31444 11212
rect 32312 11203 32364 11212
rect 32312 11169 32321 11203
rect 32321 11169 32355 11203
rect 32355 11169 32364 11203
rect 32312 11160 32364 11169
rect 27620 11092 27672 11144
rect 32220 11135 32272 11144
rect 32220 11101 32229 11135
rect 32229 11101 32263 11135
rect 32263 11101 32272 11135
rect 32220 11092 32272 11101
rect 27988 11024 28040 11076
rect 29920 11067 29972 11076
rect 29920 11033 29929 11067
rect 29929 11033 29963 11067
rect 29963 11033 29972 11067
rect 29920 11024 29972 11033
rect 31668 11024 31720 11076
rect 31760 11024 31812 11076
rect 32588 11160 32640 11212
rect 34704 11092 34756 11144
rect 40500 11135 40552 11144
rect 40500 11101 40509 11135
rect 40509 11101 40543 11135
rect 40543 11101 40552 11135
rect 40500 11092 40552 11101
rect 41420 11092 41472 11144
rect 45008 11160 45060 11212
rect 85488 11160 85540 11212
rect 42432 11135 42484 11144
rect 42432 11101 42441 11135
rect 42441 11101 42475 11135
rect 42475 11101 42484 11135
rect 42432 11092 42484 11101
rect 55496 11135 55548 11144
rect 55496 11101 55505 11135
rect 55505 11101 55539 11135
rect 55539 11101 55548 11135
rect 55496 11092 55548 11101
rect 57244 11092 57296 11144
rect 74724 11092 74776 11144
rect 78404 11135 78456 11144
rect 78404 11101 78413 11135
rect 78413 11101 78447 11135
rect 78447 11101 78456 11135
rect 78404 11092 78456 11101
rect 86408 11135 86460 11144
rect 86408 11101 86417 11135
rect 86417 11101 86451 11135
rect 86451 11101 86460 11135
rect 86408 11092 86460 11101
rect 89168 11160 89220 11212
rect 102048 11160 102100 11212
rect 102600 11160 102652 11212
rect 87788 11135 87840 11144
rect 87788 11101 87797 11135
rect 87797 11101 87831 11135
rect 87831 11101 87840 11135
rect 87788 11092 87840 11101
rect 88432 11135 88484 11144
rect 88432 11101 88441 11135
rect 88441 11101 88475 11135
rect 88475 11101 88484 11135
rect 88432 11092 88484 11101
rect 102416 11092 102468 11144
rect 103060 11135 103112 11144
rect 103060 11101 103069 11135
rect 103069 11101 103103 11135
rect 103103 11101 103112 11135
rect 103060 11092 103112 11101
rect 130292 11160 130344 11212
rect 114744 11092 114796 11144
rect 115756 11092 115808 11144
rect 115848 11092 115900 11144
rect 119712 11092 119764 11144
rect 130936 11092 130988 11144
rect 132592 11160 132644 11212
rect 143264 11160 143316 11212
rect 133144 11092 133196 11144
rect 142068 11135 142120 11144
rect 142068 11101 142077 11135
rect 142077 11101 142111 11135
rect 142111 11101 142120 11135
rect 142068 11092 142120 11101
rect 145748 11092 145800 11144
rect 147496 11160 147548 11212
rect 156420 11228 156472 11280
rect 165436 11228 165488 11280
rect 151360 11160 151412 11212
rect 81624 11024 81676 11076
rect 87880 11024 87932 11076
rect 113732 11024 113784 11076
rect 140688 11024 140740 11076
rect 153108 11092 153160 11144
rect 162216 11135 162268 11144
rect 162216 11101 162225 11135
rect 162225 11101 162259 11135
rect 162259 11101 162268 11135
rect 162216 11092 162268 11101
rect 165344 11160 165396 11212
rect 177672 11160 177724 11212
rect 177948 11160 178000 11212
rect 163504 11135 163556 11144
rect 163504 11101 163513 11135
rect 163513 11101 163547 11135
rect 163547 11101 163556 11135
rect 163504 11092 163556 11101
rect 178040 11092 178092 11144
rect 180800 11160 180852 11212
rect 191196 11160 191248 11212
rect 191840 11160 191892 11212
rect 252744 11228 252796 11280
rect 253204 11228 253256 11280
rect 265164 11228 265216 11280
rect 269304 11296 269356 11348
rect 193496 11160 193548 11212
rect 194416 11160 194468 11212
rect 194600 11160 194652 11212
rect 180432 11092 180484 11144
rect 188988 11092 189040 11144
rect 190644 11092 190696 11144
rect 190828 11135 190880 11144
rect 190828 11101 190837 11135
rect 190837 11101 190871 11135
rect 190871 11101 190880 11135
rect 190828 11092 190880 11101
rect 191932 11092 191984 11144
rect 194876 11092 194928 11144
rect 196440 11160 196492 11212
rect 201040 11160 201092 11212
rect 195796 11135 195848 11144
rect 31852 10999 31904 11008
rect 31852 10965 31861 10999
rect 31861 10965 31895 10999
rect 31895 10965 31904 10999
rect 31852 10956 31904 10965
rect 149060 10956 149112 11008
rect 149520 10956 149572 11008
rect 156144 11024 156196 11076
rect 179420 11024 179472 11076
rect 189448 11024 189500 11076
rect 193312 11024 193364 11076
rect 195796 11101 195805 11135
rect 195805 11101 195839 11135
rect 195839 11101 195848 11135
rect 195796 11092 195848 11101
rect 202696 11092 202748 11144
rect 203340 11160 203392 11212
rect 194416 10999 194468 11008
rect 194416 10965 194425 10999
rect 194425 10965 194459 10999
rect 194459 10965 194468 10999
rect 194416 10956 194468 10965
rect 195244 11024 195296 11076
rect 204996 11160 205048 11212
rect 238024 11160 238076 11212
rect 242716 11160 242768 11212
rect 267280 11160 267332 11212
rect 268016 11160 268068 11212
rect 204076 11024 204128 11076
rect 204904 11135 204956 11144
rect 204904 11101 204913 11135
rect 204913 11101 204947 11135
rect 204947 11101 204956 11135
rect 229376 11135 229428 11144
rect 204904 11092 204956 11101
rect 229376 11101 229385 11135
rect 229385 11101 229419 11135
rect 229419 11101 229428 11135
rect 229376 11092 229428 11101
rect 205456 11024 205508 11076
rect 230756 11024 230808 11076
rect 240876 11092 240928 11144
rect 241980 11092 242032 11144
rect 251548 11092 251600 11144
rect 253020 11092 253072 11144
rect 253296 11135 253348 11144
rect 253296 11101 253305 11135
rect 253305 11101 253339 11135
rect 253339 11101 253348 11135
rect 253296 11092 253348 11101
rect 254400 11092 254452 11144
rect 254676 11092 254728 11144
rect 264336 11092 264388 11144
rect 264888 11135 264940 11144
rect 264888 11101 264897 11135
rect 264897 11101 264931 11135
rect 264931 11101 264940 11135
rect 264888 11092 264940 11101
rect 265624 11092 265676 11144
rect 268476 11160 268528 11212
rect 268936 11160 268988 11212
rect 272248 11160 272300 11212
rect 269672 11092 269724 11144
rect 270408 11135 270460 11144
rect 270408 11101 270417 11135
rect 270417 11101 270451 11135
rect 270451 11101 270460 11135
rect 270408 11092 270460 11101
rect 270868 11092 270920 11144
rect 268292 11024 268344 11076
rect 268936 11024 268988 11076
rect 269948 11024 270000 11076
rect 268844 10999 268896 11008
rect 268844 10965 268853 10999
rect 268853 10965 268887 10999
rect 268887 10965 268896 10999
rect 268844 10956 268896 10965
rect 270040 10999 270092 11008
rect 270040 10965 270049 10999
rect 270049 10965 270083 10999
rect 270083 10965 270092 10999
rect 270040 10956 270092 10965
rect 77148 10854 77200 10906
rect 77212 10854 77264 10906
rect 77276 10854 77328 10906
rect 77340 10854 77392 10906
rect 77404 10854 77456 10906
rect 153346 10854 153398 10906
rect 153410 10854 153462 10906
rect 153474 10854 153526 10906
rect 153538 10854 153590 10906
rect 153602 10854 153654 10906
rect 229544 10854 229596 10906
rect 229608 10854 229660 10906
rect 229672 10854 229724 10906
rect 229736 10854 229788 10906
rect 229800 10854 229852 10906
rect 29828 10752 29880 10804
rect 30472 10752 30524 10804
rect 30748 10795 30800 10804
rect 30748 10761 30757 10795
rect 30757 10761 30791 10795
rect 30791 10761 30800 10795
rect 30748 10752 30800 10761
rect 29736 10684 29788 10736
rect 28448 10616 28500 10668
rect 30196 10684 30248 10736
rect 32680 10752 32732 10804
rect 33048 10752 33100 10804
rect 101680 10795 101732 10804
rect 101680 10761 101689 10795
rect 101689 10761 101723 10795
rect 101723 10761 101732 10795
rect 101680 10752 101732 10761
rect 130476 10795 130528 10804
rect 130476 10761 130485 10795
rect 130485 10761 130519 10795
rect 130519 10761 130528 10795
rect 130476 10752 130528 10761
rect 141976 10795 142028 10804
rect 141976 10761 141985 10795
rect 141985 10761 142019 10795
rect 142019 10761 142028 10795
rect 141976 10752 142028 10761
rect 148600 10752 148652 10804
rect 148968 10752 149020 10804
rect 191104 10752 191156 10804
rect 31760 10684 31812 10736
rect 31852 10684 31904 10736
rect 140688 10727 140740 10736
rect 32956 10659 33008 10668
rect 32956 10625 32965 10659
rect 32965 10625 32999 10659
rect 32999 10625 33008 10659
rect 32956 10616 33008 10625
rect 140688 10693 140697 10727
rect 140697 10693 140731 10727
rect 140731 10693 140740 10727
rect 140688 10684 140740 10693
rect 101864 10659 101916 10668
rect 101864 10625 101873 10659
rect 101873 10625 101907 10659
rect 101907 10625 101916 10659
rect 101864 10616 101916 10625
rect 130292 10616 130344 10668
rect 151636 10684 151688 10736
rect 156144 10727 156196 10736
rect 156144 10693 156153 10727
rect 156153 10693 156187 10727
rect 156187 10693 156196 10727
rect 156144 10684 156196 10693
rect 150348 10616 150400 10668
rect 192208 10684 192260 10736
rect 190552 10616 190604 10668
rect 192300 10616 192352 10668
rect 193220 10684 193272 10736
rect 193864 10752 193916 10804
rect 205088 10752 205140 10804
rect 255228 10752 255280 10804
rect 266544 10795 266596 10804
rect 266544 10761 266553 10795
rect 266553 10761 266587 10795
rect 266587 10761 266596 10795
rect 266544 10752 266596 10761
rect 268200 10752 268252 10804
rect 269396 10752 269448 10804
rect 195060 10684 195112 10736
rect 264888 10684 264940 10736
rect 194140 10659 194192 10668
rect 194140 10625 194149 10659
rect 194149 10625 194183 10659
rect 194183 10625 194192 10659
rect 194140 10616 194192 10625
rect 194968 10616 195020 10668
rect 204812 10616 204864 10668
rect 254952 10616 255004 10668
rect 266360 10616 266412 10668
rect 270040 10684 270092 10736
rect 187516 10591 187568 10600
rect 187516 10557 187525 10591
rect 187525 10557 187559 10591
rect 187559 10557 187568 10591
rect 187516 10548 187568 10557
rect 192116 10480 192168 10532
rect 201040 10548 201092 10600
rect 269028 10616 269080 10668
rect 270316 10616 270368 10668
rect 272524 10548 272576 10600
rect 179144 10412 179196 10464
rect 268752 10480 268804 10532
rect 203524 10412 203576 10464
rect 269580 10412 269632 10464
rect 39049 10310 39101 10362
rect 39113 10310 39165 10362
rect 39177 10310 39229 10362
rect 39241 10310 39293 10362
rect 39305 10310 39357 10362
rect 115247 10310 115299 10362
rect 115311 10310 115363 10362
rect 115375 10310 115427 10362
rect 115439 10310 115491 10362
rect 115503 10310 115555 10362
rect 191445 10310 191497 10362
rect 191509 10310 191561 10362
rect 191573 10310 191625 10362
rect 191637 10310 191689 10362
rect 191701 10310 191753 10362
rect 267643 10310 267695 10362
rect 267707 10310 267759 10362
rect 267771 10310 267823 10362
rect 267835 10310 267887 10362
rect 267899 10310 267951 10362
rect 30104 10208 30156 10260
rect 31668 10251 31720 10260
rect 31668 10217 31677 10251
rect 31677 10217 31711 10251
rect 31711 10217 31720 10251
rect 31668 10208 31720 10217
rect 32128 10208 32180 10260
rect 33324 10208 33376 10260
rect 191288 10208 191340 10260
rect 192484 10208 192536 10260
rect 266912 10208 266964 10260
rect 268568 10208 268620 10260
rect 27528 10140 27580 10192
rect 31576 10140 31628 10192
rect 163596 10072 163648 10124
rect 29460 10004 29512 10056
rect 30932 10004 30984 10056
rect 33416 10004 33468 10056
rect 33692 10004 33744 10056
rect 140688 10004 140740 10056
rect 156144 10004 156196 10056
rect 192576 10004 192628 10056
rect 195888 10072 195940 10124
rect 267740 10072 267792 10124
rect 194416 10004 194468 10056
rect 268384 10140 268436 10192
rect 269488 10140 269540 10192
rect 268844 10072 268896 10124
rect 268108 10004 268160 10056
rect 269028 10004 269080 10056
rect 269212 10047 269264 10056
rect 269212 10013 269221 10047
rect 269221 10013 269255 10047
rect 269255 10013 269264 10047
rect 269212 10004 269264 10013
rect 304448 10047 304500 10056
rect 304448 10013 304457 10047
rect 304457 10013 304491 10047
rect 304491 10013 304500 10047
rect 304448 10004 304500 10013
rect 252744 9936 252796 9988
rect 117412 9868 117464 9920
rect 194324 9868 194376 9920
rect 267740 9868 267792 9920
rect 270960 9868 271012 9920
rect 77148 9766 77200 9818
rect 77212 9766 77264 9818
rect 77276 9766 77328 9818
rect 77340 9766 77392 9818
rect 77404 9766 77456 9818
rect 153346 9766 153398 9818
rect 153410 9766 153462 9818
rect 153474 9766 153526 9818
rect 153538 9766 153590 9818
rect 153602 9766 153654 9818
rect 229544 9766 229596 9818
rect 229608 9766 229660 9818
rect 229672 9766 229724 9818
rect 229736 9766 229788 9818
rect 229800 9766 229852 9818
rect 31208 9596 31260 9648
rect 140688 9639 140740 9648
rect 140688 9605 140697 9639
rect 140697 9605 140731 9639
rect 140731 9605 140740 9639
rect 140688 9596 140740 9605
rect 156144 9639 156196 9648
rect 156144 9605 156153 9639
rect 156153 9605 156187 9639
rect 156187 9605 156196 9639
rect 156144 9596 156196 9605
rect 158628 9596 158680 9648
rect 190644 9596 190696 9648
rect 27344 9528 27396 9580
rect 33692 9528 33744 9580
rect 193312 9596 193364 9648
rect 269856 9596 269908 9648
rect 30564 9460 30616 9512
rect 194140 9528 194192 9580
rect 268108 9528 268160 9580
rect 195980 9460 196032 9512
rect 29920 9392 29972 9444
rect 194508 9392 194560 9444
rect 104256 9324 104308 9376
rect 148324 9324 148376 9376
rect 39049 9222 39101 9274
rect 39113 9222 39165 9274
rect 39177 9222 39229 9274
rect 39241 9222 39293 9274
rect 39305 9222 39357 9274
rect 115247 9222 115299 9274
rect 115311 9222 115363 9274
rect 115375 9222 115427 9274
rect 115439 9222 115491 9274
rect 115503 9222 115555 9274
rect 191445 9222 191497 9274
rect 191509 9222 191561 9274
rect 191573 9222 191625 9274
rect 191637 9222 191689 9274
rect 191701 9222 191753 9274
rect 267643 9222 267695 9274
rect 267707 9222 267759 9274
rect 267771 9222 267823 9274
rect 267835 9222 267887 9274
rect 267899 9222 267951 9274
rect 77148 8678 77200 8730
rect 77212 8678 77264 8730
rect 77276 8678 77328 8730
rect 77340 8678 77392 8730
rect 77404 8678 77456 8730
rect 153346 8678 153398 8730
rect 153410 8678 153462 8730
rect 153474 8678 153526 8730
rect 153538 8678 153590 8730
rect 153602 8678 153654 8730
rect 229544 8678 229596 8730
rect 229608 8678 229660 8730
rect 229672 8678 229724 8730
rect 229736 8678 229788 8730
rect 229800 8678 229852 8730
rect 1400 8347 1452 8356
rect 1400 8313 1409 8347
rect 1409 8313 1443 8347
rect 1443 8313 1452 8347
rect 1400 8304 1452 8313
rect 187516 8304 187568 8356
rect 39049 8134 39101 8186
rect 39113 8134 39165 8186
rect 39177 8134 39229 8186
rect 39241 8134 39293 8186
rect 39305 8134 39357 8186
rect 115247 8134 115299 8186
rect 115311 8134 115363 8186
rect 115375 8134 115427 8186
rect 115439 8134 115491 8186
rect 115503 8134 115555 8186
rect 191445 8134 191497 8186
rect 191509 8134 191561 8186
rect 191573 8134 191625 8186
rect 191637 8134 191689 8186
rect 191701 8134 191753 8186
rect 267643 8134 267695 8186
rect 267707 8134 267759 8186
rect 267771 8134 267823 8186
rect 267835 8134 267887 8186
rect 267899 8134 267951 8186
rect 77148 7590 77200 7642
rect 77212 7590 77264 7642
rect 77276 7590 77328 7642
rect 77340 7590 77392 7642
rect 77404 7590 77456 7642
rect 153346 7590 153398 7642
rect 153410 7590 153462 7642
rect 153474 7590 153526 7642
rect 153538 7590 153590 7642
rect 153602 7590 153654 7642
rect 229544 7590 229596 7642
rect 229608 7590 229660 7642
rect 229672 7590 229724 7642
rect 229736 7590 229788 7642
rect 229800 7590 229852 7642
rect 39049 7046 39101 7098
rect 39113 7046 39165 7098
rect 39177 7046 39229 7098
rect 39241 7046 39293 7098
rect 39305 7046 39357 7098
rect 115247 7046 115299 7098
rect 115311 7046 115363 7098
rect 115375 7046 115427 7098
rect 115439 7046 115491 7098
rect 115503 7046 115555 7098
rect 191445 7046 191497 7098
rect 191509 7046 191561 7098
rect 191573 7046 191625 7098
rect 191637 7046 191689 7098
rect 191701 7046 191753 7098
rect 267643 7046 267695 7098
rect 267707 7046 267759 7098
rect 267771 7046 267823 7098
rect 267835 7046 267887 7098
rect 267899 7046 267951 7098
rect 77148 6502 77200 6554
rect 77212 6502 77264 6554
rect 77276 6502 77328 6554
rect 77340 6502 77392 6554
rect 77404 6502 77456 6554
rect 153346 6502 153398 6554
rect 153410 6502 153462 6554
rect 153474 6502 153526 6554
rect 153538 6502 153590 6554
rect 153602 6502 153654 6554
rect 229544 6502 229596 6554
rect 229608 6502 229660 6554
rect 229672 6502 229724 6554
rect 229736 6502 229788 6554
rect 229800 6502 229852 6554
rect 303988 6307 304040 6316
rect 303988 6273 303997 6307
rect 303997 6273 304031 6307
rect 304031 6273 304040 6307
rect 303988 6264 304040 6273
rect 249064 6196 249116 6248
rect 39049 5958 39101 6010
rect 39113 5958 39165 6010
rect 39177 5958 39229 6010
rect 39241 5958 39293 6010
rect 39305 5958 39357 6010
rect 115247 5958 115299 6010
rect 115311 5958 115363 6010
rect 115375 5958 115427 6010
rect 115439 5958 115491 6010
rect 115503 5958 115555 6010
rect 191445 5958 191497 6010
rect 191509 5958 191561 6010
rect 191573 5958 191625 6010
rect 191637 5958 191689 6010
rect 191701 5958 191753 6010
rect 267643 5958 267695 6010
rect 267707 5958 267759 6010
rect 267771 5958 267823 6010
rect 267835 5958 267887 6010
rect 267899 5958 267951 6010
rect 77148 5414 77200 5466
rect 77212 5414 77264 5466
rect 77276 5414 77328 5466
rect 77340 5414 77392 5466
rect 77404 5414 77456 5466
rect 153346 5414 153398 5466
rect 153410 5414 153462 5466
rect 153474 5414 153526 5466
rect 153538 5414 153590 5466
rect 153602 5414 153654 5466
rect 229544 5414 229596 5466
rect 229608 5414 229660 5466
rect 229672 5414 229724 5466
rect 229736 5414 229788 5466
rect 229800 5414 229852 5466
rect 39049 4870 39101 4922
rect 39113 4870 39165 4922
rect 39177 4870 39229 4922
rect 39241 4870 39293 4922
rect 39305 4870 39357 4922
rect 115247 4870 115299 4922
rect 115311 4870 115363 4922
rect 115375 4870 115427 4922
rect 115439 4870 115491 4922
rect 115503 4870 115555 4922
rect 191445 4870 191497 4922
rect 191509 4870 191561 4922
rect 191573 4870 191625 4922
rect 191637 4870 191689 4922
rect 191701 4870 191753 4922
rect 267643 4870 267695 4922
rect 267707 4870 267759 4922
rect 267771 4870 267823 4922
rect 267835 4870 267887 4922
rect 267899 4870 267951 4922
rect 77148 4326 77200 4378
rect 77212 4326 77264 4378
rect 77276 4326 77328 4378
rect 77340 4326 77392 4378
rect 77404 4326 77456 4378
rect 153346 4326 153398 4378
rect 153410 4326 153462 4378
rect 153474 4326 153526 4378
rect 153538 4326 153590 4378
rect 153602 4326 153654 4378
rect 229544 4326 229596 4378
rect 229608 4326 229660 4378
rect 229672 4326 229724 4378
rect 229736 4326 229788 4378
rect 229800 4326 229852 4378
rect 39049 3782 39101 3834
rect 39113 3782 39165 3834
rect 39177 3782 39229 3834
rect 39241 3782 39293 3834
rect 39305 3782 39357 3834
rect 115247 3782 115299 3834
rect 115311 3782 115363 3834
rect 115375 3782 115427 3834
rect 115439 3782 115491 3834
rect 115503 3782 115555 3834
rect 191445 3782 191497 3834
rect 191509 3782 191561 3834
rect 191573 3782 191625 3834
rect 191637 3782 191689 3834
rect 191701 3782 191753 3834
rect 267643 3782 267695 3834
rect 267707 3782 267759 3834
rect 267771 3782 267823 3834
rect 267835 3782 267887 3834
rect 267899 3782 267951 3834
rect 77148 3238 77200 3290
rect 77212 3238 77264 3290
rect 77276 3238 77328 3290
rect 77340 3238 77392 3290
rect 77404 3238 77456 3290
rect 153346 3238 153398 3290
rect 153410 3238 153462 3290
rect 153474 3238 153526 3290
rect 153538 3238 153590 3290
rect 153602 3238 153654 3290
rect 229544 3238 229596 3290
rect 229608 3238 229660 3290
rect 229672 3238 229724 3290
rect 229736 3238 229788 3290
rect 229800 3238 229852 3290
rect 39049 2694 39101 2746
rect 39113 2694 39165 2746
rect 39177 2694 39229 2746
rect 39241 2694 39293 2746
rect 39305 2694 39357 2746
rect 115247 2694 115299 2746
rect 115311 2694 115363 2746
rect 115375 2694 115427 2746
rect 115439 2694 115491 2746
rect 115503 2694 115555 2746
rect 191445 2694 191497 2746
rect 191509 2694 191561 2746
rect 191573 2694 191625 2746
rect 191637 2694 191689 2746
rect 191701 2694 191753 2746
rect 267643 2694 267695 2746
rect 267707 2694 267759 2746
rect 267771 2694 267823 2746
rect 267835 2694 267887 2746
rect 267899 2694 267951 2746
rect 149428 2592 149480 2644
rect 302240 2592 302292 2644
rect 77148 2150 77200 2202
rect 77212 2150 77264 2202
rect 77276 2150 77328 2202
rect 77340 2150 77392 2202
rect 77404 2150 77456 2202
rect 153346 2150 153398 2202
rect 153410 2150 153462 2202
rect 153474 2150 153526 2202
rect 153538 2150 153590 2202
rect 153602 2150 153654 2202
rect 229544 2150 229596 2202
rect 229608 2150 229660 2202
rect 229672 2150 229724 2202
rect 229736 2150 229788 2202
rect 229800 2150 229852 2202
<< metal2 >>
rect 1490 15314 1546 16000
rect 4526 15314 4582 16000
rect 7562 15314 7618 16000
rect 10690 15314 10746 16000
rect 1490 15286 1624 15314
rect 1490 15200 1546 15286
rect 1596 13530 1624 15286
rect 4526 15286 4660 15314
rect 4526 15200 4582 15286
rect 4632 13530 4660 15286
rect 7562 15286 7696 15314
rect 7562 15200 7618 15286
rect 7668 13530 7696 15286
rect 10690 15286 10824 15314
rect 10690 15200 10746 15286
rect 10796 13530 10824 15286
rect 13726 15200 13782 16000
rect 16762 15314 16818 16000
rect 19890 15314 19946 16000
rect 22926 15314 22982 16000
rect 25962 15314 26018 16000
rect 16762 15286 16896 15314
rect 16762 15200 16818 15286
rect 1584 13524 1636 13530
rect 1584 13466 1636 13472
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 7656 13524 7708 13530
rect 7656 13466 7708 13472
rect 10784 13524 10836 13530
rect 13740 13512 13768 15200
rect 16868 13530 16896 15286
rect 19890 15286 20024 15314
rect 19890 15200 19946 15286
rect 19996 13530 20024 15286
rect 22926 15286 23060 15314
rect 22926 15200 22982 15286
rect 23032 13530 23060 15286
rect 25962 15286 26096 15314
rect 25962 15200 26018 15286
rect 13820 13524 13872 13530
rect 13740 13484 13820 13512
rect 10784 13466 10836 13472
rect 13820 13466 13872 13472
rect 16856 13524 16908 13530
rect 16856 13466 16908 13472
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 23020 13524 23072 13530
rect 23020 13466 23072 13472
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 20168 13320 20220 13326
rect 20168 13262 20220 13268
rect 23204 13320 23256 13326
rect 23204 13262 23256 13268
rect 4816 12102 4844 13262
rect 14292 12374 14320 13262
rect 14280 12368 14332 12374
rect 14280 12310 14332 12316
rect 17052 12238 17080 13262
rect 20180 12918 20208 13262
rect 20168 12912 20220 12918
rect 20168 12854 20220 12860
rect 23216 12782 23244 13262
rect 26068 12986 26096 15286
rect 29090 15200 29146 16000
rect 32126 15200 32182 16000
rect 35254 15314 35310 16000
rect 38290 15314 38346 16000
rect 35254 15286 35572 15314
rect 35254 15200 35310 15286
rect 29000 13796 29052 13802
rect 29000 13738 29052 13744
rect 27160 13728 27212 13734
rect 27160 13670 27212 13676
rect 27172 13462 27200 13670
rect 27448 13654 27752 13682
rect 27160 13456 27212 13462
rect 27160 13398 27212 13404
rect 26976 13388 27028 13394
rect 26976 13330 27028 13336
rect 26056 12980 26108 12986
rect 26056 12922 26108 12928
rect 23204 12776 23256 12782
rect 23204 12718 23256 12724
rect 26988 12442 27016 13330
rect 27172 12714 27200 13398
rect 27252 13184 27304 13190
rect 27252 13126 27304 13132
rect 27264 13002 27292 13126
rect 27448 13002 27476 13654
rect 27724 13530 27752 13654
rect 27620 13524 27672 13530
rect 27620 13466 27672 13472
rect 27712 13524 27764 13530
rect 27712 13466 27764 13472
rect 27528 13252 27580 13258
rect 27528 13194 27580 13200
rect 27264 12974 27476 13002
rect 27344 12912 27396 12918
rect 27344 12854 27396 12860
rect 27160 12708 27212 12714
rect 27160 12650 27212 12656
rect 26976 12436 27028 12442
rect 26976 12378 27028 12384
rect 26884 12300 26936 12306
rect 26884 12242 26936 12248
rect 17040 12232 17092 12238
rect 17040 12174 17092 12180
rect 26896 12186 26924 12242
rect 26896 12158 27200 12186
rect 27172 12102 27200 12158
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 27068 12096 27120 12102
rect 27068 12038 27120 12044
rect 27160 12096 27212 12102
rect 27160 12038 27212 12044
rect 27080 11218 27108 12038
rect 27068 11212 27120 11218
rect 27068 11154 27120 11160
rect 27356 9586 27384 12854
rect 27448 12238 27476 12974
rect 27436 12232 27488 12238
rect 27436 12174 27488 12180
rect 27540 10198 27568 13194
rect 27632 11150 27660 13466
rect 27712 13184 27764 13190
rect 27712 13126 27764 13132
rect 27724 11830 27752 13126
rect 29012 12918 29040 13738
rect 29000 12912 29052 12918
rect 29000 12854 29052 12860
rect 27988 12844 28040 12850
rect 27988 12786 28040 12792
rect 28000 12102 28028 12786
rect 28080 12776 28132 12782
rect 28080 12718 28132 12724
rect 28092 12442 28120 12718
rect 28908 12640 28960 12646
rect 28908 12582 28960 12588
rect 28080 12436 28132 12442
rect 28080 12378 28132 12384
rect 28816 12436 28868 12442
rect 28816 12378 28868 12384
rect 28092 12306 28120 12378
rect 28828 12322 28856 12378
rect 28736 12306 28856 12322
rect 28080 12300 28132 12306
rect 28080 12242 28132 12248
rect 28724 12300 28856 12306
rect 28776 12294 28856 12300
rect 28724 12242 28776 12248
rect 27988 12096 28040 12102
rect 27988 12038 28040 12044
rect 27712 11824 27764 11830
rect 27712 11766 27764 11772
rect 27620 11144 27672 11150
rect 27620 11086 27672 11092
rect 28000 11082 28028 12038
rect 28736 11830 28764 12242
rect 28920 12102 28948 12582
rect 29000 12300 29052 12306
rect 29000 12242 29052 12248
rect 28908 12096 28960 12102
rect 28908 12038 28960 12044
rect 29012 11830 29040 12242
rect 29104 11898 29132 15200
rect 30472 13524 30524 13530
rect 30472 13466 30524 13472
rect 30484 13410 30512 13466
rect 30392 13382 30512 13410
rect 29828 13320 29880 13326
rect 29828 13262 29880 13268
rect 29840 12782 29868 13262
rect 30196 13252 30248 13258
rect 30196 13194 30248 13200
rect 29644 12776 29696 12782
rect 29644 12718 29696 12724
rect 29828 12776 29880 12782
rect 29828 12718 29880 12724
rect 30104 12776 30156 12782
rect 30104 12718 30156 12724
rect 29656 12434 29684 12718
rect 29656 12406 29776 12434
rect 29552 12300 29604 12306
rect 29552 12242 29604 12248
rect 29368 12232 29420 12238
rect 29366 12200 29368 12209
rect 29420 12200 29422 12209
rect 29366 12135 29422 12144
rect 29460 12164 29512 12170
rect 29460 12106 29512 12112
rect 29472 11898 29500 12106
rect 29092 11892 29144 11898
rect 29092 11834 29144 11840
rect 29460 11892 29512 11898
rect 29460 11834 29512 11840
rect 28724 11824 28776 11830
rect 28724 11766 28776 11772
rect 29000 11824 29052 11830
rect 29000 11766 29052 11772
rect 29564 11762 29592 12242
rect 29552 11756 29604 11762
rect 29552 11698 29604 11704
rect 28908 11688 28960 11694
rect 28908 11630 28960 11636
rect 28448 11552 28500 11558
rect 28448 11494 28500 11500
rect 27988 11076 28040 11082
rect 27988 11018 28040 11024
rect 28460 10674 28488 11494
rect 28920 11286 28948 11630
rect 28908 11280 28960 11286
rect 28908 11222 28960 11228
rect 29564 11218 29592 11698
rect 29460 11212 29512 11218
rect 29460 11154 29512 11160
rect 29552 11212 29604 11218
rect 29552 11154 29604 11160
rect 28448 10668 28500 10674
rect 28448 10610 28500 10616
rect 27528 10192 27580 10198
rect 27528 10134 27580 10140
rect 29472 10062 29500 11154
rect 29748 10742 29776 12406
rect 29828 12164 29880 12170
rect 29828 12106 29880 12112
rect 29840 10810 29868 12106
rect 30012 11824 30064 11830
rect 30012 11766 30064 11772
rect 29920 11688 29972 11694
rect 29920 11630 29972 11636
rect 29932 11354 29960 11630
rect 30024 11354 30052 11766
rect 29920 11348 29972 11354
rect 29920 11290 29972 11296
rect 30012 11348 30064 11354
rect 30012 11290 30064 11296
rect 29920 11076 29972 11082
rect 29920 11018 29972 11024
rect 29828 10804 29880 10810
rect 29828 10746 29880 10752
rect 29736 10736 29788 10742
rect 29736 10678 29788 10684
rect 29460 10056 29512 10062
rect 29460 9998 29512 10004
rect 27344 9580 27396 9586
rect 27344 9522 27396 9528
rect 29932 9450 29960 11018
rect 30116 10266 30144 12718
rect 30208 10742 30236 13194
rect 30392 12918 30420 13382
rect 30472 13184 30524 13190
rect 30472 13126 30524 13132
rect 30380 12912 30432 12918
rect 30380 12854 30432 12860
rect 30392 11370 30420 12854
rect 30484 12434 30512 13126
rect 31576 12912 31628 12918
rect 31576 12854 31628 12860
rect 31392 12640 31444 12646
rect 31392 12582 31444 12588
rect 30484 12406 30604 12434
rect 30392 11342 30512 11370
rect 30484 10810 30512 11342
rect 30472 10804 30524 10810
rect 30472 10746 30524 10752
rect 30196 10736 30248 10742
rect 30196 10678 30248 10684
rect 30104 10260 30156 10266
rect 30104 10202 30156 10208
rect 30576 9518 30604 12406
rect 31404 12209 31432 12582
rect 30746 12200 30802 12209
rect 31390 12200 31446 12209
rect 30746 12135 30802 12144
rect 31208 12164 31260 12170
rect 30760 10810 30788 12135
rect 31390 12135 31446 12144
rect 31208 12106 31260 12112
rect 31116 12096 31168 12102
rect 31116 12038 31168 12044
rect 30932 11892 30984 11898
rect 30932 11834 30984 11840
rect 30748 10804 30800 10810
rect 30748 10746 30800 10752
rect 30944 10062 30972 11834
rect 31128 11626 31156 12038
rect 31116 11620 31168 11626
rect 31116 11562 31168 11568
rect 30932 10056 30984 10062
rect 30932 9998 30984 10004
rect 31220 9654 31248 12106
rect 31392 11552 31444 11558
rect 31392 11494 31444 11500
rect 31404 11218 31432 11494
rect 31392 11212 31444 11218
rect 31392 11154 31444 11160
rect 31588 10198 31616 12854
rect 32036 12164 32088 12170
rect 32036 12106 32088 12112
rect 32048 11830 32076 12106
rect 32036 11824 32088 11830
rect 32036 11766 32088 11772
rect 31668 11076 31720 11082
rect 31668 11018 31720 11024
rect 31760 11076 31812 11082
rect 31760 11018 31812 11024
rect 31680 10266 31708 11018
rect 31772 10742 31800 11018
rect 31852 11008 31904 11014
rect 31852 10950 31904 10956
rect 31864 10742 31892 10950
rect 31760 10736 31812 10742
rect 31760 10678 31812 10684
rect 31852 10736 31904 10742
rect 31852 10678 31904 10684
rect 32140 10266 32168 15200
rect 32956 13796 33008 13802
rect 32956 13738 33008 13744
rect 32404 13320 32456 13326
rect 32404 13262 32456 13268
rect 32220 12980 32272 12986
rect 32220 12922 32272 12928
rect 32232 11898 32260 12922
rect 32416 12646 32444 13262
rect 32680 13252 32732 13258
rect 32680 13194 32732 13200
rect 32404 12640 32456 12646
rect 32404 12582 32456 12588
rect 32588 12436 32640 12442
rect 32588 12378 32640 12384
rect 32312 12096 32364 12102
rect 32312 12038 32364 12044
rect 32220 11892 32272 11898
rect 32220 11834 32272 11840
rect 32232 11150 32260 11834
rect 32324 11218 32352 12038
rect 32404 11756 32456 11762
rect 32404 11698 32456 11704
rect 32416 11354 32444 11698
rect 32600 11694 32628 12378
rect 32588 11688 32640 11694
rect 32588 11630 32640 11636
rect 32404 11348 32456 11354
rect 32404 11290 32456 11296
rect 32600 11218 32628 11630
rect 32312 11212 32364 11218
rect 32312 11154 32364 11160
rect 32588 11212 32640 11218
rect 32588 11154 32640 11160
rect 32220 11144 32272 11150
rect 32220 11086 32272 11092
rect 32692 10810 32720 13194
rect 32968 12102 32996 13738
rect 33784 13320 33836 13326
rect 33784 13262 33836 13268
rect 33600 13184 33652 13190
rect 33600 13126 33652 13132
rect 33048 12776 33100 12782
rect 33048 12718 33100 12724
rect 33416 12776 33468 12782
rect 33416 12718 33468 12724
rect 32956 12096 33008 12102
rect 32956 12038 33008 12044
rect 32956 11552 33008 11558
rect 32956 11494 33008 11500
rect 32680 10804 32732 10810
rect 32680 10746 32732 10752
rect 32968 10674 32996 11494
rect 33060 10810 33088 12718
rect 33324 11348 33376 11354
rect 33324 11290 33376 11296
rect 33048 10804 33100 10810
rect 33048 10746 33100 10752
rect 32956 10668 33008 10674
rect 32956 10610 33008 10616
rect 33336 10266 33364 11290
rect 31668 10260 31720 10266
rect 31668 10202 31720 10208
rect 32128 10260 32180 10266
rect 32128 10202 32180 10208
rect 33324 10260 33376 10266
rect 33324 10202 33376 10208
rect 31576 10192 31628 10198
rect 31576 10134 31628 10140
rect 33428 10062 33456 12718
rect 33612 11354 33640 13126
rect 33692 12844 33744 12850
rect 33692 12786 33744 12792
rect 33600 11348 33652 11354
rect 33600 11290 33652 11296
rect 33704 10062 33732 12786
rect 33796 11898 33824 13262
rect 34520 13252 34572 13258
rect 34520 13194 34572 13200
rect 34152 13184 34204 13190
rect 34152 13126 34204 13132
rect 34336 13184 34388 13190
rect 34336 13126 34388 13132
rect 34164 12986 34192 13126
rect 34152 12980 34204 12986
rect 34152 12922 34204 12928
rect 34164 12832 34192 12922
rect 34072 12804 34192 12832
rect 33784 11892 33836 11898
rect 33784 11834 33836 11840
rect 34072 11694 34100 12804
rect 34348 12782 34376 13126
rect 34428 12912 34480 12918
rect 34428 12854 34480 12860
rect 34336 12776 34388 12782
rect 34336 12718 34388 12724
rect 34152 12640 34204 12646
rect 34152 12582 34204 12588
rect 34164 12238 34192 12582
rect 34152 12232 34204 12238
rect 34152 12174 34204 12180
rect 34440 11898 34468 12854
rect 34532 12442 34560 13194
rect 35544 12986 35572 15286
rect 38290 15286 38424 15314
rect 38290 15200 38346 15286
rect 36544 13728 36596 13734
rect 36544 13670 36596 13676
rect 36556 13530 36584 13670
rect 36544 13524 36596 13530
rect 36544 13466 36596 13472
rect 35992 13252 36044 13258
rect 35992 13194 36044 13200
rect 37832 13252 37884 13258
rect 37832 13194 37884 13200
rect 35532 12980 35584 12986
rect 35532 12922 35584 12928
rect 34888 12776 34940 12782
rect 34888 12718 34940 12724
rect 35348 12776 35400 12782
rect 35348 12718 35400 12724
rect 34520 12436 34572 12442
rect 34520 12378 34572 12384
rect 34900 12374 34928 12718
rect 34888 12368 34940 12374
rect 34888 12310 34940 12316
rect 35360 12238 35388 12718
rect 36004 12442 36032 13194
rect 37464 13184 37516 13190
rect 37464 13126 37516 13132
rect 37476 12918 37504 13126
rect 37464 12912 37516 12918
rect 37464 12854 37516 12860
rect 37844 12442 37872 13194
rect 38016 12640 38068 12646
rect 38016 12582 38068 12588
rect 35992 12436 36044 12442
rect 35992 12378 36044 12384
rect 37832 12436 37884 12442
rect 37832 12378 37884 12384
rect 38028 12238 38056 12582
rect 34704 12232 34756 12238
rect 34704 12174 34756 12180
rect 35348 12232 35400 12238
rect 35348 12174 35400 12180
rect 38016 12232 38068 12238
rect 38016 12174 38068 12180
rect 34428 11892 34480 11898
rect 34428 11834 34480 11840
rect 34716 11762 34744 12174
rect 36452 12096 36504 12102
rect 36452 12038 36504 12044
rect 34704 11756 34756 11762
rect 34704 11698 34756 11704
rect 34060 11688 34112 11694
rect 34060 11630 34112 11636
rect 34716 11150 34744 11698
rect 36464 11286 36492 12038
rect 38396 11898 38424 15286
rect 41326 15200 41382 16000
rect 44454 15314 44510 16000
rect 47490 15314 47546 16000
rect 44454 15286 44588 15314
rect 44454 15200 44510 15286
rect 39049 13628 39357 13637
rect 39049 13626 39055 13628
rect 39111 13626 39135 13628
rect 39191 13626 39215 13628
rect 39271 13626 39295 13628
rect 39351 13626 39357 13628
rect 39111 13574 39113 13626
rect 39293 13574 39295 13626
rect 39049 13572 39055 13574
rect 39111 13572 39135 13574
rect 39191 13572 39215 13574
rect 39271 13572 39295 13574
rect 39351 13572 39357 13574
rect 39049 13563 39357 13572
rect 38936 13320 38988 13326
rect 38936 13262 38988 13268
rect 38948 12442 38976 13262
rect 40408 13252 40460 13258
rect 40408 13194 40460 13200
rect 39304 13184 39356 13190
rect 39304 13126 39356 13132
rect 39948 13184 40000 13190
rect 39948 13126 40000 13132
rect 39316 12850 39344 13126
rect 39672 12912 39724 12918
rect 39672 12854 39724 12860
rect 39304 12844 39356 12850
rect 39304 12786 39356 12792
rect 39396 12776 39448 12782
rect 39396 12718 39448 12724
rect 39049 12540 39357 12549
rect 39049 12538 39055 12540
rect 39111 12538 39135 12540
rect 39191 12538 39215 12540
rect 39271 12538 39295 12540
rect 39351 12538 39357 12540
rect 39111 12486 39113 12538
rect 39293 12486 39295 12538
rect 39049 12484 39055 12486
rect 39111 12484 39135 12486
rect 39191 12484 39215 12486
rect 39271 12484 39295 12486
rect 39351 12484 39357 12486
rect 39049 12475 39357 12484
rect 39408 12442 39436 12718
rect 38936 12436 38988 12442
rect 38936 12378 38988 12384
rect 39396 12436 39448 12442
rect 39396 12378 39448 12384
rect 38384 11892 38436 11898
rect 38384 11834 38436 11840
rect 39580 11892 39632 11898
rect 39684 11880 39712 12854
rect 39960 11898 39988 13126
rect 40316 12232 40368 12238
rect 40316 12174 40368 12180
rect 39632 11852 39712 11880
rect 39948 11892 40000 11898
rect 39580 11834 39632 11840
rect 39948 11834 40000 11840
rect 40328 11762 40356 12174
rect 40316 11756 40368 11762
rect 40316 11698 40368 11704
rect 39049 11452 39357 11461
rect 39049 11450 39055 11452
rect 39111 11450 39135 11452
rect 39191 11450 39215 11452
rect 39271 11450 39295 11452
rect 39351 11450 39357 11452
rect 39111 11398 39113 11450
rect 39293 11398 39295 11450
rect 39049 11396 39055 11398
rect 39111 11396 39135 11398
rect 39191 11396 39215 11398
rect 39271 11396 39295 11398
rect 39351 11396 39357 11398
rect 39049 11387 39357 11396
rect 40420 11354 40448 13194
rect 41052 12912 41104 12918
rect 41052 12854 41104 12860
rect 40960 12776 41012 12782
rect 40960 12718 41012 12724
rect 40972 12442 41000 12718
rect 40960 12436 41012 12442
rect 40960 12378 41012 12384
rect 40972 12306 41000 12378
rect 40960 12300 41012 12306
rect 40960 12242 41012 12248
rect 40592 12232 40644 12238
rect 40590 12200 40592 12209
rect 40644 12200 40646 12209
rect 40590 12135 40646 12144
rect 40500 12096 40552 12102
rect 40500 12038 40552 12044
rect 40684 12096 40736 12102
rect 40684 12038 40736 12044
rect 40408 11348 40460 11354
rect 40408 11290 40460 11296
rect 36452 11280 36504 11286
rect 36452 11222 36504 11228
rect 40512 11150 40540 12038
rect 40696 11830 40724 12038
rect 40684 11824 40736 11830
rect 40684 11766 40736 11772
rect 40972 11694 41000 12242
rect 40960 11688 41012 11694
rect 40960 11630 41012 11636
rect 41064 11354 41092 12854
rect 41236 12640 41288 12646
rect 41236 12582 41288 12588
rect 41248 11830 41276 12582
rect 41236 11824 41288 11830
rect 41236 11766 41288 11772
rect 41052 11348 41104 11354
rect 41052 11290 41104 11296
rect 41340 11286 41368 15200
rect 42524 13728 42576 13734
rect 42524 13670 42576 13676
rect 42536 13326 42564 13670
rect 44180 13456 44232 13462
rect 44364 13456 44416 13462
rect 44232 13416 44364 13444
rect 44180 13398 44232 13404
rect 44364 13398 44416 13404
rect 42524 13320 42576 13326
rect 42524 13262 42576 13268
rect 44272 13320 44324 13326
rect 44272 13262 44324 13268
rect 41420 13252 41472 13258
rect 41420 13194 41472 13200
rect 42892 13252 42944 13258
rect 42892 13194 42944 13200
rect 43260 13252 43312 13258
rect 43260 13194 43312 13200
rect 41432 11898 41460 13194
rect 42432 13184 42484 13190
rect 42432 13126 42484 13132
rect 41512 12844 41564 12850
rect 41512 12786 41564 12792
rect 41420 11892 41472 11898
rect 41420 11834 41472 11840
rect 41420 11688 41472 11694
rect 41524 11676 41552 12786
rect 41788 12640 41840 12646
rect 41788 12582 41840 12588
rect 41800 12170 41828 12582
rect 42444 12209 42472 13126
rect 42800 12640 42852 12646
rect 42800 12582 42852 12588
rect 42430 12200 42486 12209
rect 41604 12164 41656 12170
rect 41604 12106 41656 12112
rect 41788 12164 41840 12170
rect 42430 12135 42486 12144
rect 41788 12106 41840 12112
rect 41472 11648 41552 11676
rect 41420 11630 41472 11636
rect 41328 11280 41380 11286
rect 41328 11222 41380 11228
rect 41432 11150 41460 11630
rect 41616 11354 41644 12106
rect 41604 11348 41656 11354
rect 41604 11290 41656 11296
rect 42444 11150 42472 12135
rect 42812 11762 42840 12582
rect 42904 11898 42932 13194
rect 43272 12986 43300 13194
rect 44284 12986 44312 13262
rect 44560 12986 44588 15286
rect 47490 15286 47624 15314
rect 47490 15200 47546 15286
rect 46204 13796 46256 13802
rect 46204 13738 46256 13744
rect 46216 13530 46244 13738
rect 47596 13530 47624 15286
rect 50526 15200 50582 16000
rect 53654 15200 53710 16000
rect 56690 15200 56746 16000
rect 59818 15200 59874 16000
rect 62854 15314 62910 16000
rect 65890 15314 65946 16000
rect 69018 15314 69074 16000
rect 72054 15314 72110 16000
rect 62854 15286 63080 15314
rect 62854 15200 62910 15286
rect 47860 13728 47912 13734
rect 47860 13670 47912 13676
rect 46204 13524 46256 13530
rect 46204 13466 46256 13472
rect 47584 13524 47636 13530
rect 47584 13466 47636 13472
rect 45560 13388 45612 13394
rect 45560 13330 45612 13336
rect 45008 13184 45060 13190
rect 45008 13126 45060 13132
rect 45376 13184 45428 13190
rect 45376 13126 45428 13132
rect 43260 12980 43312 12986
rect 43260 12922 43312 12928
rect 44272 12980 44324 12986
rect 44272 12922 44324 12928
rect 44548 12980 44600 12986
rect 44548 12922 44600 12928
rect 42984 12912 43036 12918
rect 42984 12854 43036 12860
rect 42892 11892 42944 11898
rect 42892 11834 42944 11840
rect 42996 11762 43024 12854
rect 43088 12838 43300 12866
rect 43088 12782 43116 12838
rect 43076 12776 43128 12782
rect 43076 12718 43128 12724
rect 43168 12776 43220 12782
rect 43168 12718 43220 12724
rect 43180 12442 43208 12718
rect 43272 12646 43300 12838
rect 43812 12776 43864 12782
rect 43812 12718 43864 12724
rect 43824 12646 43852 12718
rect 43260 12640 43312 12646
rect 43260 12582 43312 12588
rect 43812 12640 43864 12646
rect 43812 12582 43864 12588
rect 43824 12442 43852 12582
rect 43168 12436 43220 12442
rect 43168 12378 43220 12384
rect 43812 12436 43864 12442
rect 43812 12378 43864 12384
rect 43720 12368 43772 12374
rect 43720 12310 43772 12316
rect 43732 12238 43760 12310
rect 43720 12232 43772 12238
rect 43720 12174 43772 12180
rect 42800 11756 42852 11762
rect 42800 11698 42852 11704
rect 42984 11756 43036 11762
rect 42984 11698 43036 11704
rect 45020 11218 45048 13126
rect 45388 12850 45416 13126
rect 45376 12844 45428 12850
rect 45376 12786 45428 12792
rect 45468 12776 45520 12782
rect 45572 12764 45600 13330
rect 47872 13258 47900 13670
rect 50540 13530 50568 15200
rect 51632 13728 51684 13734
rect 51632 13670 51684 13676
rect 50528 13524 50580 13530
rect 50528 13466 50580 13472
rect 51644 13394 51672 13670
rect 53012 13524 53064 13530
rect 53012 13466 53064 13472
rect 51632 13388 51684 13394
rect 51632 13330 51684 13336
rect 51356 13320 51408 13326
rect 51356 13262 51408 13268
rect 47860 13252 47912 13258
rect 47860 13194 47912 13200
rect 51368 12782 51396 13262
rect 45520 12736 45600 12764
rect 51356 12776 51408 12782
rect 45468 12718 45520 12724
rect 51356 12718 51408 12724
rect 52644 12164 52696 12170
rect 52644 12106 52696 12112
rect 52656 11898 52684 12106
rect 52644 11892 52696 11898
rect 52644 11834 52696 11840
rect 53024 11762 53052 13466
rect 53288 13252 53340 13258
rect 53288 13194 53340 13200
rect 53300 12986 53328 13194
rect 53288 12980 53340 12986
rect 53288 12922 53340 12928
rect 53104 12640 53156 12646
rect 53104 12582 53156 12588
rect 53116 12170 53144 12582
rect 53104 12164 53156 12170
rect 53104 12106 53156 12112
rect 53668 11898 53696 15200
rect 54116 13728 54168 13734
rect 54116 13670 54168 13676
rect 53748 12844 53800 12850
rect 53748 12786 53800 12792
rect 54024 12844 54076 12850
rect 54024 12786 54076 12792
rect 53760 12322 53788 12786
rect 54036 12442 54064 12786
rect 54128 12782 54156 13670
rect 55588 13524 55640 13530
rect 55588 13466 55640 13472
rect 55600 13326 55628 13466
rect 54392 13320 54444 13326
rect 54392 13262 54444 13268
rect 54760 13320 54812 13326
rect 54760 13262 54812 13268
rect 55588 13320 55640 13326
rect 55588 13262 55640 13268
rect 54116 12776 54168 12782
rect 54116 12718 54168 12724
rect 54128 12646 54156 12718
rect 54116 12640 54168 12646
rect 54116 12582 54168 12588
rect 54024 12436 54076 12442
rect 54024 12378 54076 12384
rect 53760 12306 53880 12322
rect 53760 12300 53892 12306
rect 53760 12294 53840 12300
rect 53656 11892 53708 11898
rect 53656 11834 53708 11840
rect 53760 11830 53788 12294
rect 53840 12242 53892 12248
rect 54404 11898 54432 13262
rect 54668 13184 54720 13190
rect 54668 13126 54720 13132
rect 54680 12986 54708 13126
rect 54668 12980 54720 12986
rect 54668 12922 54720 12928
rect 54392 11892 54444 11898
rect 54392 11834 54444 11840
rect 53748 11824 53800 11830
rect 53748 11766 53800 11772
rect 53012 11756 53064 11762
rect 53012 11698 53064 11704
rect 54680 11694 54708 12922
rect 54772 12850 54800 13262
rect 55864 13252 55916 13258
rect 55864 13194 55916 13200
rect 56600 13252 56652 13258
rect 56600 13194 56652 13200
rect 55876 12986 55904 13194
rect 55864 12980 55916 12986
rect 55864 12922 55916 12928
rect 55496 12912 55548 12918
rect 55496 12854 55548 12860
rect 54760 12844 54812 12850
rect 54760 12786 54812 12792
rect 55036 12776 55088 12782
rect 55036 12718 55088 12724
rect 54668 11688 54720 11694
rect 54668 11630 54720 11636
rect 55048 11354 55076 12718
rect 55508 12442 55536 12854
rect 55588 12640 55640 12646
rect 55588 12582 55640 12588
rect 56324 12640 56376 12646
rect 56324 12582 56376 12588
rect 56508 12640 56560 12646
rect 56508 12582 56560 12588
rect 55496 12436 55548 12442
rect 55496 12378 55548 12384
rect 55312 12232 55364 12238
rect 55312 12174 55364 12180
rect 55324 11898 55352 12174
rect 55312 11892 55364 11898
rect 55312 11834 55364 11840
rect 55600 11694 55628 12582
rect 56336 12434 56364 12582
rect 56336 12406 56456 12434
rect 56428 12306 56456 12406
rect 56416 12300 56468 12306
rect 56416 12242 56468 12248
rect 56520 12238 56548 12582
rect 56508 12232 56560 12238
rect 56508 12174 56560 12180
rect 55864 12096 55916 12102
rect 55864 12038 55916 12044
rect 56048 12096 56100 12102
rect 56048 12038 56100 12044
rect 55876 11694 55904 12038
rect 55588 11688 55640 11694
rect 55588 11630 55640 11636
rect 55864 11688 55916 11694
rect 55864 11630 55916 11636
rect 56060 11626 56088 12038
rect 56612 11898 56640 13194
rect 56704 12442 56732 15200
rect 57888 13524 57940 13530
rect 57888 13466 57940 13472
rect 57900 13326 57928 13466
rect 59832 13462 59860 15200
rect 61752 13524 61804 13530
rect 61752 13466 61804 13472
rect 59820 13456 59872 13462
rect 59820 13398 59872 13404
rect 57888 13320 57940 13326
rect 57888 13262 57940 13268
rect 60648 13320 60700 13326
rect 60648 13262 60700 13268
rect 57704 13252 57756 13258
rect 57704 13194 57756 13200
rect 58624 13252 58676 13258
rect 58624 13194 58676 13200
rect 57336 13184 57388 13190
rect 57336 13126 57388 13132
rect 57348 12918 57376 13126
rect 57336 12912 57388 12918
rect 57336 12854 57388 12860
rect 57244 12640 57296 12646
rect 57244 12582 57296 12588
rect 56692 12436 56744 12442
rect 56692 12378 56744 12384
rect 56600 11892 56652 11898
rect 56600 11834 56652 11840
rect 56048 11620 56100 11626
rect 56048 11562 56100 11568
rect 55496 11552 55548 11558
rect 55496 11494 55548 11500
rect 55036 11348 55088 11354
rect 55036 11290 55088 11296
rect 45008 11212 45060 11218
rect 45008 11154 45060 11160
rect 55508 11150 55536 11494
rect 57256 11150 57284 12582
rect 57348 12102 57376 12854
rect 57428 12844 57480 12850
rect 57428 12786 57480 12792
rect 57336 12096 57388 12102
rect 57336 12038 57388 12044
rect 57440 11830 57468 12786
rect 57428 11824 57480 11830
rect 57428 11766 57480 11772
rect 57716 11354 57744 13194
rect 57980 12980 58032 12986
rect 57980 12922 58032 12928
rect 57992 12442 58020 12922
rect 57980 12436 58032 12442
rect 57980 12378 58032 12384
rect 58636 11898 58664 13194
rect 59636 13184 59688 13190
rect 59636 13126 59688 13132
rect 59648 12986 59676 13126
rect 59636 12980 59688 12986
rect 59636 12922 59688 12928
rect 60660 12918 60688 13262
rect 61488 13258 61700 13274
rect 61764 13258 61792 13466
rect 63052 13462 63080 15286
rect 65890 15286 66024 15314
rect 65890 15200 65946 15286
rect 63408 13796 63460 13802
rect 63408 13738 63460 13744
rect 63420 13530 63448 13738
rect 63408 13524 63460 13530
rect 63408 13466 63460 13472
rect 63040 13456 63092 13462
rect 63040 13398 63092 13404
rect 61476 13252 61700 13258
rect 61528 13246 61700 13252
rect 61476 13194 61528 13200
rect 61672 13190 61700 13246
rect 61752 13252 61804 13258
rect 61752 13194 61804 13200
rect 65996 13190 66024 15286
rect 69018 15286 69152 15314
rect 69018 15200 69074 15286
rect 66168 13728 66220 13734
rect 66168 13670 66220 13676
rect 66180 13326 66208 13670
rect 66168 13320 66220 13326
rect 66168 13262 66220 13268
rect 69124 13190 69152 15286
rect 72054 15286 72188 15314
rect 72054 15200 72110 15286
rect 69296 13796 69348 13802
rect 69296 13738 69348 13744
rect 69308 13326 69336 13738
rect 69296 13320 69348 13326
rect 69296 13262 69348 13268
rect 61660 13184 61712 13190
rect 61660 13126 61712 13132
rect 65892 13184 65944 13190
rect 65892 13126 65944 13132
rect 65984 13184 66036 13190
rect 65984 13126 66036 13132
rect 69112 13184 69164 13190
rect 69112 13126 69164 13132
rect 65904 12918 65932 13126
rect 72160 12986 72188 15286
rect 75090 15200 75146 16000
rect 78218 15314 78274 16000
rect 81254 15314 81310 16000
rect 78218 15286 78536 15314
rect 78218 15200 78274 15286
rect 72424 13728 72476 13734
rect 72424 13670 72476 13676
rect 73896 13728 73948 13734
rect 73896 13670 73948 13676
rect 72436 13190 72464 13670
rect 72700 13388 72752 13394
rect 72700 13330 72752 13336
rect 72332 13184 72384 13190
rect 72332 13126 72384 13132
rect 72424 13184 72476 13190
rect 72424 13126 72476 13132
rect 72344 12986 72372 13126
rect 72148 12980 72200 12986
rect 72148 12922 72200 12928
rect 72332 12980 72384 12986
rect 72332 12922 72384 12928
rect 60648 12912 60700 12918
rect 60648 12854 60700 12860
rect 65892 12912 65944 12918
rect 65892 12854 65944 12860
rect 72712 12646 72740 13330
rect 73908 13258 73936 13670
rect 73896 13252 73948 13258
rect 73896 13194 73948 13200
rect 74724 12980 74776 12986
rect 74724 12922 74776 12928
rect 72700 12640 72752 12646
rect 72700 12582 72752 12588
rect 58624 11892 58676 11898
rect 58624 11834 58676 11840
rect 57704 11348 57756 11354
rect 57704 11290 57756 11296
rect 74736 11150 74764 12922
rect 74816 12844 74868 12850
rect 74816 12786 74868 12792
rect 74828 12306 74856 12786
rect 75000 12640 75052 12646
rect 75000 12582 75052 12588
rect 74816 12300 74868 12306
rect 74816 12242 74868 12248
rect 75012 11694 75040 12582
rect 75104 12442 75132 15200
rect 75368 13796 75420 13802
rect 75368 13738 75420 13744
rect 76012 13796 76064 13802
rect 76012 13738 76064 13744
rect 75380 13462 75408 13738
rect 75368 13456 75420 13462
rect 75368 13398 75420 13404
rect 75644 13456 75696 13462
rect 75644 13398 75696 13404
rect 75184 13252 75236 13258
rect 75184 13194 75236 13200
rect 75196 12646 75224 13194
rect 75460 12844 75512 12850
rect 75460 12786 75512 12792
rect 75184 12640 75236 12646
rect 75184 12582 75236 12588
rect 75092 12436 75144 12442
rect 75092 12378 75144 12384
rect 75472 11898 75500 12786
rect 75656 11898 75684 13398
rect 76024 12374 76052 13738
rect 76380 13728 76432 13734
rect 76380 13670 76432 13676
rect 76012 12368 76064 12374
rect 76012 12310 76064 12316
rect 75460 11892 75512 11898
rect 75460 11834 75512 11840
rect 75644 11892 75696 11898
rect 75644 11834 75696 11840
rect 76024 11762 76052 12310
rect 76288 12096 76340 12102
rect 76288 12038 76340 12044
rect 76300 11762 76328 12038
rect 76012 11756 76064 11762
rect 76012 11698 76064 11704
rect 76288 11756 76340 11762
rect 76288 11698 76340 11704
rect 75000 11688 75052 11694
rect 75000 11630 75052 11636
rect 76392 11354 76420 13670
rect 78404 13320 78456 13326
rect 78404 13262 78456 13268
rect 76472 13252 76524 13258
rect 76472 13194 76524 13200
rect 76484 11898 76512 13194
rect 77944 13184 77996 13190
rect 77944 13126 77996 13132
rect 77148 13084 77456 13093
rect 77148 13082 77154 13084
rect 77210 13082 77234 13084
rect 77290 13082 77314 13084
rect 77370 13082 77394 13084
rect 77450 13082 77456 13084
rect 77210 13030 77212 13082
rect 77392 13030 77394 13082
rect 77148 13028 77154 13030
rect 77210 13028 77234 13030
rect 77290 13028 77314 13030
rect 77370 13028 77394 13030
rect 77450 13028 77456 13030
rect 77148 13019 77456 13028
rect 77852 12708 77904 12714
rect 77852 12650 77904 12656
rect 77208 12640 77260 12646
rect 77208 12582 77260 12588
rect 77220 12374 77248 12582
rect 77208 12368 77260 12374
rect 77208 12310 77260 12316
rect 76932 12300 76984 12306
rect 76932 12242 76984 12248
rect 76472 11892 76524 11898
rect 76472 11834 76524 11840
rect 76944 11694 76972 12242
rect 77148 11996 77456 12005
rect 77148 11994 77154 11996
rect 77210 11994 77234 11996
rect 77290 11994 77314 11996
rect 77370 11994 77394 11996
rect 77450 11994 77456 11996
rect 77210 11942 77212 11994
rect 77392 11942 77394 11994
rect 77148 11940 77154 11942
rect 77210 11940 77234 11942
rect 77290 11940 77314 11942
rect 77370 11940 77394 11942
rect 77450 11940 77456 11942
rect 77148 11931 77456 11940
rect 77864 11898 77892 12650
rect 77956 12238 77984 13126
rect 78416 12918 78444 13262
rect 78404 12912 78456 12918
rect 78404 12854 78456 12860
rect 78128 12708 78180 12714
rect 78128 12650 78180 12656
rect 78140 12306 78168 12650
rect 78404 12368 78456 12374
rect 78404 12310 78456 12316
rect 78128 12300 78180 12306
rect 78128 12242 78180 12248
rect 77944 12232 77996 12238
rect 77944 12174 77996 12180
rect 77852 11892 77904 11898
rect 77852 11834 77904 11840
rect 76932 11688 76984 11694
rect 76932 11630 76984 11636
rect 76380 11348 76432 11354
rect 76380 11290 76432 11296
rect 78416 11150 78444 12310
rect 78508 11898 78536 15286
rect 81254 15286 81388 15314
rect 81254 15200 81310 15286
rect 81360 13410 81388 15286
rect 84290 15200 84346 16000
rect 87418 15200 87474 16000
rect 90454 15200 90510 16000
rect 93582 15314 93638 16000
rect 96618 15314 96674 16000
rect 93582 15286 93808 15314
rect 93582 15200 93638 15286
rect 83096 13728 83148 13734
rect 83096 13670 83148 13676
rect 80244 13388 80296 13394
rect 81360 13382 81480 13410
rect 80244 13330 80296 13336
rect 79980 13258 80100 13274
rect 78772 13252 78824 13258
rect 78772 13194 78824 13200
rect 79324 13252 79376 13258
rect 79324 13194 79376 13200
rect 79980 13252 80112 13258
rect 79980 13246 80060 13252
rect 78588 12776 78640 12782
rect 78588 12718 78640 12724
rect 78600 12238 78628 12718
rect 78588 12232 78640 12238
rect 78588 12174 78640 12180
rect 78496 11892 78548 11898
rect 78496 11834 78548 11840
rect 78600 11762 78628 12174
rect 78588 11756 78640 11762
rect 78588 11698 78640 11704
rect 78784 11354 78812 13194
rect 79336 12442 79364 13194
rect 79980 12866 80008 13246
rect 80060 13194 80112 13200
rect 79704 12850 80008 12866
rect 79692 12844 80008 12850
rect 79744 12838 80008 12844
rect 79692 12786 79744 12792
rect 79324 12436 79376 12442
rect 79324 12378 79376 12384
rect 80256 12102 80284 13330
rect 81452 13326 81480 13382
rect 81624 13388 81676 13394
rect 81624 13330 81676 13336
rect 81440 13320 81492 13326
rect 81440 13262 81492 13268
rect 80796 13184 80848 13190
rect 80796 13126 80848 13132
rect 81440 13184 81492 13190
rect 81440 13126 81492 13132
rect 80520 12912 80572 12918
rect 80520 12854 80572 12860
rect 80532 12442 80560 12854
rect 80808 12782 80836 13126
rect 80796 12776 80848 12782
rect 80796 12718 80848 12724
rect 81452 12714 81480 13126
rect 81440 12708 81492 12714
rect 81440 12650 81492 12656
rect 80520 12436 80572 12442
rect 80520 12378 80572 12384
rect 81452 12306 81480 12650
rect 81636 12646 81664 13330
rect 83108 13326 83136 13670
rect 83096 13320 83148 13326
rect 83096 13262 83148 13268
rect 83924 13320 83976 13326
rect 83924 13262 83976 13268
rect 83832 13252 83884 13258
rect 83832 13194 83884 13200
rect 82912 13184 82964 13190
rect 82912 13126 82964 13132
rect 82924 12918 82952 13126
rect 82912 12912 82964 12918
rect 82912 12854 82964 12860
rect 81624 12640 81676 12646
rect 81624 12582 81676 12588
rect 81440 12300 81492 12306
rect 81440 12242 81492 12248
rect 80244 12096 80296 12102
rect 80244 12038 80296 12044
rect 81452 11762 81480 12242
rect 81440 11756 81492 11762
rect 81440 11698 81492 11704
rect 78772 11348 78824 11354
rect 78772 11290 78824 11296
rect 34704 11144 34756 11150
rect 34704 11086 34756 11092
rect 40500 11144 40552 11150
rect 40500 11086 40552 11092
rect 41420 11144 41472 11150
rect 41420 11086 41472 11092
rect 42432 11144 42484 11150
rect 42432 11086 42484 11092
rect 55496 11144 55548 11150
rect 55496 11086 55548 11092
rect 57244 11144 57296 11150
rect 57244 11086 57296 11092
rect 74724 11144 74776 11150
rect 74724 11086 74776 11092
rect 78404 11144 78456 11150
rect 78404 11086 78456 11092
rect 81636 11082 81664 12582
rect 83844 12238 83872 13194
rect 83936 13190 83964 13262
rect 83924 13184 83976 13190
rect 83924 13126 83976 13132
rect 83936 12986 83964 13126
rect 83924 12980 83976 12986
rect 83924 12922 83976 12928
rect 83832 12232 83884 12238
rect 83832 12174 83884 12180
rect 84016 12096 84068 12102
rect 84016 12038 84068 12044
rect 84028 11694 84056 12038
rect 84304 11898 84332 15200
rect 86408 13728 86460 13734
rect 86408 13670 86460 13676
rect 84476 13252 84528 13258
rect 84476 13194 84528 13200
rect 85488 13252 85540 13258
rect 85488 13194 85540 13200
rect 84292 11892 84344 11898
rect 84292 11834 84344 11840
rect 84016 11688 84068 11694
rect 84016 11630 84068 11636
rect 84488 11354 84516 13194
rect 84844 12776 84896 12782
rect 84844 12718 84896 12724
rect 84660 12300 84712 12306
rect 84660 12242 84712 12248
rect 84672 12102 84700 12242
rect 84660 12096 84712 12102
rect 84660 12038 84712 12044
rect 84856 11558 84884 12718
rect 85500 12442 85528 13194
rect 86040 13184 86092 13190
rect 86040 13126 86092 13132
rect 85764 12640 85816 12646
rect 85764 12582 85816 12588
rect 85488 12436 85540 12442
rect 85488 12378 85540 12384
rect 85776 12306 85804 12582
rect 85764 12300 85816 12306
rect 85764 12242 85816 12248
rect 85488 12232 85540 12238
rect 85488 12174 85540 12180
rect 84936 11824 84988 11830
rect 85304 11824 85356 11830
rect 84988 11772 85304 11778
rect 84936 11766 85356 11772
rect 84948 11750 85344 11766
rect 84844 11552 84896 11558
rect 84844 11494 84896 11500
rect 84476 11348 84528 11354
rect 84476 11290 84528 11296
rect 85500 11218 85528 12174
rect 85776 11762 85804 12242
rect 86052 12238 86080 13126
rect 86420 12442 86448 13670
rect 86776 13252 86828 13258
rect 86776 13194 86828 13200
rect 86500 12980 86552 12986
rect 86500 12922 86552 12928
rect 86512 12782 86540 12922
rect 86500 12776 86552 12782
rect 86500 12718 86552 12724
rect 86408 12436 86460 12442
rect 86408 12378 86460 12384
rect 86132 12368 86184 12374
rect 86132 12310 86184 12316
rect 86040 12232 86092 12238
rect 86040 12174 86092 12180
rect 86052 11898 86080 12174
rect 86144 11898 86172 12310
rect 86316 12300 86368 12306
rect 86316 12242 86368 12248
rect 86328 12102 86356 12242
rect 86316 12096 86368 12102
rect 86316 12038 86368 12044
rect 86040 11892 86092 11898
rect 86040 11834 86092 11840
rect 86132 11892 86184 11898
rect 86132 11834 86184 11840
rect 85764 11756 85816 11762
rect 85764 11698 85816 11704
rect 86328 11694 86356 12038
rect 86316 11688 86368 11694
rect 86316 11630 86368 11636
rect 86408 11552 86460 11558
rect 86408 11494 86460 11500
rect 85488 11212 85540 11218
rect 85488 11154 85540 11160
rect 86420 11150 86448 11494
rect 86788 11286 86816 13194
rect 86958 13152 87014 13161
rect 86958 13087 87014 13096
rect 86972 11762 87000 13087
rect 87144 12980 87196 12986
rect 87144 12922 87196 12928
rect 86960 11756 87012 11762
rect 86960 11698 87012 11704
rect 87156 11354 87184 12922
rect 87432 12374 87460 15200
rect 87880 13320 87932 13326
rect 87880 13262 87932 13268
rect 87786 12744 87842 12753
rect 87786 12679 87842 12688
rect 87800 12646 87828 12679
rect 87788 12640 87840 12646
rect 87788 12582 87840 12588
rect 87892 12442 87920 13262
rect 89076 13252 89128 13258
rect 89076 13194 89128 13200
rect 89536 13252 89588 13258
rect 89536 13194 89588 13200
rect 88248 13184 88300 13190
rect 88248 13126 88300 13132
rect 88260 12782 88288 13126
rect 88248 12776 88300 12782
rect 88248 12718 88300 12724
rect 87972 12640 88024 12646
rect 87972 12582 88024 12588
rect 87880 12436 87932 12442
rect 87880 12378 87932 12384
rect 87420 12368 87472 12374
rect 87420 12310 87472 12316
rect 87984 12186 88012 12582
rect 88154 12336 88210 12345
rect 88154 12271 88156 12280
rect 88208 12271 88210 12280
rect 88156 12242 88208 12248
rect 88260 12238 88288 12718
rect 88432 12640 88484 12646
rect 88432 12582 88484 12588
rect 87524 12158 88012 12186
rect 88248 12232 88300 12238
rect 88248 12174 88300 12180
rect 87524 12102 87552 12158
rect 87984 12102 88012 12158
rect 87512 12096 87564 12102
rect 87512 12038 87564 12044
rect 87788 12096 87840 12102
rect 87788 12038 87840 12044
rect 87972 12096 88024 12102
rect 87972 12038 88024 12044
rect 87144 11348 87196 11354
rect 87144 11290 87196 11296
rect 86776 11280 86828 11286
rect 86776 11222 86828 11228
rect 87800 11150 87828 12038
rect 87880 11892 87932 11898
rect 87880 11834 87932 11840
rect 86408 11144 86460 11150
rect 86408 11086 86460 11092
rect 87788 11144 87840 11150
rect 87788 11086 87840 11092
rect 87892 11082 87920 11834
rect 88444 11150 88472 12582
rect 88984 12232 89036 12238
rect 88720 12180 88984 12186
rect 88720 12174 89036 12180
rect 88720 12158 89024 12174
rect 88720 12102 88748 12158
rect 88708 12096 88760 12102
rect 88708 12038 88760 12044
rect 89088 11354 89116 13194
rect 89168 12300 89220 12306
rect 89168 12242 89220 12248
rect 89180 11762 89208 12242
rect 89548 11898 89576 13194
rect 90468 12986 90496 15200
rect 90640 13796 90692 13802
rect 90640 13738 90692 13744
rect 90548 13184 90600 13190
rect 90548 13126 90600 13132
rect 90456 12980 90508 12986
rect 90456 12922 90508 12928
rect 90560 12918 90588 13126
rect 90548 12912 90600 12918
rect 90548 12854 90600 12860
rect 90652 12850 90680 13738
rect 91836 13728 91888 13734
rect 91836 13670 91888 13676
rect 91848 13258 91876 13670
rect 93780 13546 93808 15286
rect 96618 15286 96752 15314
rect 96618 15200 96674 15286
rect 93780 13518 93900 13546
rect 93872 13462 93900 13518
rect 93860 13456 93912 13462
rect 93860 13398 93912 13404
rect 91652 13252 91704 13258
rect 91652 13194 91704 13200
rect 91836 13252 91888 13258
rect 91836 13194 91888 13200
rect 92020 13252 92072 13258
rect 92020 13194 92072 13200
rect 91664 12986 91692 13194
rect 91848 13161 91876 13194
rect 91834 13152 91890 13161
rect 91834 13087 91890 13096
rect 91652 12980 91704 12986
rect 91652 12922 91704 12928
rect 90732 12912 90784 12918
rect 90732 12854 90784 12860
rect 90180 12844 90232 12850
rect 90180 12786 90232 12792
rect 90456 12844 90508 12850
rect 90456 12786 90508 12792
rect 90640 12844 90692 12850
rect 90640 12786 90692 12792
rect 89720 12776 89772 12782
rect 90088 12776 90140 12782
rect 89772 12736 90088 12764
rect 89720 12718 89772 12724
rect 90088 12718 90140 12724
rect 89904 12640 89956 12646
rect 89904 12582 89956 12588
rect 89916 12345 89944 12582
rect 90192 12442 90220 12786
rect 90180 12436 90232 12442
rect 90180 12378 90232 12384
rect 89902 12336 89958 12345
rect 89902 12271 89958 12280
rect 89536 11892 89588 11898
rect 89536 11834 89588 11840
rect 89168 11756 89220 11762
rect 89168 11698 89220 11704
rect 89076 11348 89128 11354
rect 89076 11290 89128 11296
rect 89180 11218 89208 11698
rect 90468 11694 90496 12786
rect 90744 12753 90772 12854
rect 90730 12744 90786 12753
rect 90730 12679 90786 12688
rect 92032 12238 92060 13194
rect 96724 13190 96752 15286
rect 99654 15200 99710 16000
rect 102782 15314 102838 16000
rect 105818 15314 105874 16000
rect 108854 15314 108910 16000
rect 111982 15314 112038 16000
rect 102782 15286 102916 15314
rect 102782 15200 102838 15286
rect 99668 13410 99696 15200
rect 102416 13796 102468 13802
rect 102416 13738 102468 13744
rect 101956 13728 102008 13734
rect 101956 13670 102008 13676
rect 99104 13388 99156 13394
rect 99104 13330 99156 13336
rect 99392 13382 99696 13410
rect 100760 13456 100812 13462
rect 100760 13398 100812 13404
rect 98000 13252 98052 13258
rect 98000 13194 98052 13200
rect 96712 13184 96764 13190
rect 96712 13126 96764 13132
rect 97540 13184 97592 13190
rect 97540 13126 97592 13132
rect 97552 12238 97580 13126
rect 98012 12986 98040 13194
rect 98000 12980 98052 12986
rect 98000 12922 98052 12928
rect 99116 12306 99144 13330
rect 99196 13252 99248 13258
rect 99196 13194 99248 13200
rect 99208 12782 99236 13194
rect 99196 12776 99248 12782
rect 99196 12718 99248 12724
rect 99196 12640 99248 12646
rect 99392 12628 99420 13382
rect 99656 13252 99708 13258
rect 99656 13194 99708 13200
rect 99472 12912 99524 12918
rect 99472 12854 99524 12860
rect 99248 12600 99420 12628
rect 99196 12582 99248 12588
rect 99484 12442 99512 12854
rect 99472 12436 99524 12442
rect 99472 12378 99524 12384
rect 99104 12300 99156 12306
rect 99104 12242 99156 12248
rect 92020 12232 92072 12238
rect 92020 12174 92072 12180
rect 97540 12232 97592 12238
rect 97540 12174 97592 12180
rect 99668 11898 99696 13194
rect 99932 12912 99984 12918
rect 99932 12854 99984 12860
rect 99944 12442 99972 12854
rect 100772 12646 100800 13398
rect 101404 13320 101456 13326
rect 101404 13262 101456 13268
rect 100944 13252 100996 13258
rect 100944 13194 100996 13200
rect 100760 12640 100812 12646
rect 100760 12582 100812 12588
rect 99932 12436 99984 12442
rect 99932 12378 99984 12384
rect 100772 12170 100800 12582
rect 100760 12164 100812 12170
rect 100760 12106 100812 12112
rect 100392 12096 100444 12102
rect 100392 12038 100444 12044
rect 99656 11892 99708 11898
rect 99656 11834 99708 11840
rect 100404 11762 100432 12038
rect 100392 11756 100444 11762
rect 100392 11698 100444 11704
rect 100772 11694 100800 12106
rect 100956 11898 100984 13194
rect 101036 13184 101088 13190
rect 101036 13126 101088 13132
rect 101048 12714 101076 13126
rect 101416 12782 101444 13262
rect 101404 12776 101456 12782
rect 101404 12718 101456 12724
rect 101680 12776 101732 12782
rect 101680 12718 101732 12724
rect 101036 12708 101088 12714
rect 101036 12650 101088 12656
rect 101048 12170 101076 12650
rect 101036 12164 101088 12170
rect 101036 12106 101088 12112
rect 100944 11892 100996 11898
rect 100944 11834 100996 11840
rect 90456 11688 90508 11694
rect 90456 11630 90508 11636
rect 100760 11688 100812 11694
rect 100760 11630 100812 11636
rect 89168 11212 89220 11218
rect 89168 11154 89220 11160
rect 88432 11144 88484 11150
rect 88432 11086 88484 11092
rect 81624 11076 81676 11082
rect 81624 11018 81676 11024
rect 87880 11076 87932 11082
rect 87880 11018 87932 11024
rect 77148 10908 77456 10917
rect 77148 10906 77154 10908
rect 77210 10906 77234 10908
rect 77290 10906 77314 10908
rect 77370 10906 77394 10908
rect 77450 10906 77456 10908
rect 77210 10854 77212 10906
rect 77392 10854 77394 10906
rect 77148 10852 77154 10854
rect 77210 10852 77234 10854
rect 77290 10852 77314 10854
rect 77370 10852 77394 10854
rect 77450 10852 77456 10854
rect 77148 10843 77456 10852
rect 101692 10810 101720 12718
rect 101968 12170 101996 13670
rect 102232 13252 102284 13258
rect 102232 13194 102284 13200
rect 102048 12300 102100 12306
rect 102048 12242 102100 12248
rect 101956 12164 102008 12170
rect 101956 12106 102008 12112
rect 102060 11694 102088 12242
rect 102140 12164 102192 12170
rect 102140 12106 102192 12112
rect 102152 11762 102180 12106
rect 102140 11756 102192 11762
rect 102140 11698 102192 11704
rect 102048 11688 102100 11694
rect 102048 11630 102100 11636
rect 101864 11552 101916 11558
rect 101864 11494 101916 11500
rect 101680 10804 101732 10810
rect 101680 10746 101732 10752
rect 101876 10674 101904 11494
rect 102060 11218 102088 11630
rect 102244 11286 102272 13194
rect 102324 12096 102376 12102
rect 102324 12038 102376 12044
rect 102336 11694 102364 12038
rect 102324 11688 102376 11694
rect 102324 11630 102376 11636
rect 102232 11280 102284 11286
rect 102232 11222 102284 11228
rect 102048 11212 102100 11218
rect 102048 11154 102100 11160
rect 102428 11150 102456 13738
rect 102600 12096 102652 12102
rect 102600 12038 102652 12044
rect 102612 11218 102640 12038
rect 102888 11354 102916 15286
rect 105818 15286 105952 15314
rect 105818 15200 105874 15286
rect 103336 13320 103388 13326
rect 103336 13262 103388 13268
rect 104256 13320 104308 13326
rect 104256 13262 104308 13268
rect 103244 12708 103296 12714
rect 103244 12650 103296 12656
rect 103060 12640 103112 12646
rect 103060 12582 103112 12588
rect 103072 12102 103100 12582
rect 103256 12306 103284 12650
rect 103348 12306 103376 13262
rect 104072 13252 104124 13258
rect 104072 13194 104124 13200
rect 103704 13184 103756 13190
rect 103704 13126 103756 13132
rect 103612 12640 103664 12646
rect 103612 12582 103664 12588
rect 103244 12300 103296 12306
rect 103244 12242 103296 12248
rect 103336 12300 103388 12306
rect 103336 12242 103388 12248
rect 103060 12096 103112 12102
rect 103060 12038 103112 12044
rect 103072 11898 103100 12038
rect 103060 11892 103112 11898
rect 103060 11834 103112 11840
rect 103520 11892 103572 11898
rect 103520 11834 103572 11840
rect 102876 11348 102928 11354
rect 102876 11290 102928 11296
rect 102600 11212 102652 11218
rect 102600 11154 102652 11160
rect 103072 11150 103100 11834
rect 103532 11694 103560 11834
rect 103624 11762 103652 12582
rect 103716 12238 103744 13126
rect 103704 12232 103756 12238
rect 103704 12174 103756 12180
rect 103612 11756 103664 11762
rect 103612 11698 103664 11704
rect 103520 11688 103572 11694
rect 103520 11630 103572 11636
rect 104084 11558 104112 13194
rect 104072 11552 104124 11558
rect 104072 11494 104124 11500
rect 102416 11144 102468 11150
rect 102416 11086 102468 11092
rect 103060 11144 103112 11150
rect 103060 11086 103112 11092
rect 101864 10668 101916 10674
rect 101864 10610 101916 10616
rect 39049 10364 39357 10373
rect 39049 10362 39055 10364
rect 39111 10362 39135 10364
rect 39191 10362 39215 10364
rect 39271 10362 39295 10364
rect 39351 10362 39357 10364
rect 39111 10310 39113 10362
rect 39293 10310 39295 10362
rect 39049 10308 39055 10310
rect 39111 10308 39135 10310
rect 39191 10308 39215 10310
rect 39271 10308 39295 10310
rect 39351 10308 39357 10310
rect 39049 10299 39357 10308
rect 33416 10056 33468 10062
rect 33416 9998 33468 10004
rect 33692 10056 33744 10062
rect 33692 9998 33744 10004
rect 31208 9648 31260 9654
rect 31208 9590 31260 9596
rect 33704 9586 33732 9998
rect 77148 9820 77456 9829
rect 77148 9818 77154 9820
rect 77210 9818 77234 9820
rect 77290 9818 77314 9820
rect 77370 9818 77394 9820
rect 77450 9818 77456 9820
rect 77210 9766 77212 9818
rect 77392 9766 77394 9818
rect 77148 9764 77154 9766
rect 77210 9764 77234 9766
rect 77290 9764 77314 9766
rect 77370 9764 77394 9766
rect 77450 9764 77456 9766
rect 77148 9755 77456 9764
rect 33692 9580 33744 9586
rect 33692 9522 33744 9528
rect 30564 9512 30616 9518
rect 30564 9454 30616 9460
rect 29920 9444 29972 9450
rect 29920 9386 29972 9392
rect 104268 9382 104296 13262
rect 104452 13246 104756 13274
rect 104452 13190 104480 13246
rect 104440 13184 104492 13190
rect 104440 13126 104492 13132
rect 104624 13184 104676 13190
rect 104624 13126 104676 13132
rect 104636 12918 104664 13126
rect 104728 12918 104756 13246
rect 104992 13252 105044 13258
rect 104992 13194 105044 13200
rect 104624 12912 104676 12918
rect 104624 12854 104676 12860
rect 104716 12912 104768 12918
rect 104716 12854 104768 12860
rect 105004 12442 105032 13194
rect 105176 12844 105228 12850
rect 105176 12786 105228 12792
rect 105188 12442 105216 12786
rect 105924 12714 105952 15286
rect 108854 15286 108988 15314
rect 108854 15200 108910 15286
rect 108960 13546 108988 15286
rect 111812 15286 112038 15314
rect 111812 13546 111840 15286
rect 111982 15200 112038 15286
rect 115018 15200 115074 16000
rect 118146 15314 118202 16000
rect 121182 15314 121238 16000
rect 118146 15286 118648 15314
rect 118146 15200 118202 15286
rect 113824 13796 113876 13802
rect 113824 13738 113876 13744
rect 108960 13518 109080 13546
rect 109052 13462 109080 13518
rect 111720 13518 111840 13546
rect 111720 13462 111748 13518
rect 109040 13456 109092 13462
rect 109040 13398 109092 13404
rect 111708 13456 111760 13462
rect 111708 13398 111760 13404
rect 109592 13320 109644 13326
rect 109592 13262 109644 13268
rect 111432 13320 111484 13326
rect 111432 13262 111484 13268
rect 109604 13190 109632 13262
rect 109592 13184 109644 13190
rect 109592 13126 109644 13132
rect 109604 12918 109632 13126
rect 111444 12986 111472 13262
rect 112536 13252 112588 13258
rect 112536 13194 112588 13200
rect 111432 12980 111484 12986
rect 111432 12922 111484 12928
rect 109592 12912 109644 12918
rect 109592 12854 109644 12860
rect 105912 12708 105964 12714
rect 105912 12650 105964 12656
rect 111892 12640 111944 12646
rect 111892 12582 111944 12588
rect 104992 12436 105044 12442
rect 104992 12378 105044 12384
rect 105176 12436 105228 12442
rect 105176 12378 105228 12384
rect 111904 12238 111932 12582
rect 112548 12442 112576 13194
rect 113836 12850 113864 13738
rect 114652 13728 114704 13734
rect 114652 13670 114704 13676
rect 114192 13252 114244 13258
rect 114192 13194 114244 13200
rect 113088 12844 113140 12850
rect 113088 12786 113140 12792
rect 113824 12844 113876 12850
rect 113824 12786 113876 12792
rect 113100 12646 113128 12786
rect 113088 12640 113140 12646
rect 113088 12582 113140 12588
rect 112536 12436 112588 12442
rect 112536 12378 112588 12384
rect 113836 12322 113864 12786
rect 113916 12776 113968 12782
rect 113916 12718 113968 12724
rect 113744 12294 113864 12322
rect 111892 12232 111944 12238
rect 111892 12174 111944 12180
rect 113744 11082 113772 12294
rect 113824 12164 113876 12170
rect 113824 12106 113876 12112
rect 113836 11898 113864 12106
rect 113928 12102 113956 12718
rect 113916 12096 113968 12102
rect 113916 12038 113968 12044
rect 113824 11892 113876 11898
rect 113824 11834 113876 11840
rect 114008 11756 114060 11762
rect 114008 11698 114060 11704
rect 114020 11558 114048 11698
rect 114008 11552 114060 11558
rect 114008 11494 114060 11500
rect 114204 11286 114232 13194
rect 114560 13184 114612 13190
rect 114560 13126 114612 13132
rect 114572 12986 114600 13126
rect 114560 12980 114612 12986
rect 114560 12922 114612 12928
rect 114664 12850 114692 13670
rect 114836 13320 114888 13326
rect 114836 13262 114888 13268
rect 114744 12980 114796 12986
rect 114744 12922 114796 12928
rect 114652 12844 114704 12850
rect 114652 12786 114704 12792
rect 114664 12322 114692 12786
rect 114756 12782 114784 12922
rect 114744 12776 114796 12782
rect 114744 12718 114796 12724
rect 114848 12714 114876 13262
rect 114928 13184 114980 13190
rect 114928 13126 114980 13132
rect 114836 12708 114888 12714
rect 114836 12650 114888 12656
rect 114744 12640 114796 12646
rect 114744 12582 114796 12588
rect 114572 12294 114692 12322
rect 114284 12232 114336 12238
rect 114284 12174 114336 12180
rect 114296 11898 114324 12174
rect 114284 11892 114336 11898
rect 114284 11834 114336 11840
rect 114572 11830 114600 12294
rect 114560 11824 114612 11830
rect 114560 11766 114612 11772
rect 114192 11280 114244 11286
rect 114192 11222 114244 11228
rect 114756 11150 114784 12582
rect 114940 12322 114968 13126
rect 115032 12442 115060 15200
rect 118620 13682 118648 15286
rect 121182 15286 121316 15314
rect 121182 15200 121238 15286
rect 118620 13654 118740 13682
rect 115247 13628 115555 13637
rect 115247 13626 115253 13628
rect 115309 13626 115333 13628
rect 115389 13626 115413 13628
rect 115469 13626 115493 13628
rect 115549 13626 115555 13628
rect 115309 13574 115311 13626
rect 115491 13574 115493 13626
rect 115247 13572 115253 13574
rect 115309 13572 115333 13574
rect 115389 13572 115413 13574
rect 115469 13572 115493 13574
rect 115549 13572 115555 13574
rect 115247 13563 115555 13572
rect 118240 13388 118292 13394
rect 118240 13330 118292 13336
rect 117412 13320 117464 13326
rect 117412 13262 117464 13268
rect 115112 13252 115164 13258
rect 115112 13194 115164 13200
rect 116952 13252 117004 13258
rect 116952 13194 117004 13200
rect 115020 12436 115072 12442
rect 115020 12378 115072 12384
rect 114940 12294 115060 12322
rect 115032 11762 115060 12294
rect 115020 11756 115072 11762
rect 115020 11698 115072 11704
rect 115124 11354 115152 13194
rect 115756 13184 115808 13190
rect 115756 13126 115808 13132
rect 115768 12918 115796 13126
rect 115756 12912 115808 12918
rect 115756 12854 115808 12860
rect 115664 12776 115716 12782
rect 115848 12776 115900 12782
rect 115664 12718 115716 12724
rect 115768 12724 115848 12730
rect 115768 12718 115900 12724
rect 116768 12776 116820 12782
rect 116768 12718 116820 12724
rect 115247 12540 115555 12549
rect 115247 12538 115253 12540
rect 115309 12538 115333 12540
rect 115389 12538 115413 12540
rect 115469 12538 115493 12540
rect 115549 12538 115555 12540
rect 115309 12486 115311 12538
rect 115491 12486 115493 12538
rect 115247 12484 115253 12486
rect 115309 12484 115333 12486
rect 115389 12484 115413 12486
rect 115469 12484 115493 12486
rect 115549 12484 115555 12486
rect 115247 12475 115555 12484
rect 115676 12102 115704 12718
rect 115768 12702 115888 12718
rect 115768 12374 115796 12702
rect 115848 12640 115900 12646
rect 115848 12582 115900 12588
rect 115756 12368 115808 12374
rect 115756 12310 115808 12316
rect 115664 12096 115716 12102
rect 115664 12038 115716 12044
rect 115676 11898 115704 12038
rect 115664 11892 115716 11898
rect 115664 11834 115716 11840
rect 115768 11778 115796 12310
rect 115676 11750 115796 11778
rect 115676 11694 115704 11750
rect 115664 11688 115716 11694
rect 115664 11630 115716 11636
rect 115756 11688 115808 11694
rect 115756 11630 115808 11636
rect 115247 11452 115555 11461
rect 115247 11450 115253 11452
rect 115309 11450 115333 11452
rect 115389 11450 115413 11452
rect 115469 11450 115493 11452
rect 115549 11450 115555 11452
rect 115309 11398 115311 11450
rect 115491 11398 115493 11450
rect 115247 11396 115253 11398
rect 115309 11396 115333 11398
rect 115389 11396 115413 11398
rect 115469 11396 115493 11398
rect 115549 11396 115555 11398
rect 115247 11387 115555 11396
rect 115112 11348 115164 11354
rect 115112 11290 115164 11296
rect 115768 11150 115796 11630
rect 115860 11150 115888 12582
rect 116400 12096 116452 12102
rect 116400 12038 116452 12044
rect 116412 11762 116440 12038
rect 116780 11898 116808 12718
rect 116964 12442 116992 13194
rect 117424 12986 117452 13262
rect 117688 13252 117740 13258
rect 117688 13194 117740 13200
rect 117412 12980 117464 12986
rect 117412 12922 117464 12928
rect 117320 12912 117372 12918
rect 117320 12854 117372 12860
rect 116952 12436 117004 12442
rect 116952 12378 117004 12384
rect 117332 11898 117360 12854
rect 116768 11892 116820 11898
rect 116768 11834 116820 11840
rect 117320 11892 117372 11898
rect 117320 11834 117372 11840
rect 116400 11756 116452 11762
rect 116400 11698 116452 11704
rect 114744 11144 114796 11150
rect 114744 11086 114796 11092
rect 115756 11144 115808 11150
rect 115756 11086 115808 11092
rect 115848 11144 115900 11150
rect 115848 11086 115900 11092
rect 113732 11076 113784 11082
rect 113732 11018 113784 11024
rect 115247 10364 115555 10373
rect 115247 10362 115253 10364
rect 115309 10362 115333 10364
rect 115389 10362 115413 10364
rect 115469 10362 115493 10364
rect 115549 10362 115555 10364
rect 115309 10310 115311 10362
rect 115491 10310 115493 10362
rect 115247 10308 115253 10310
rect 115309 10308 115333 10310
rect 115389 10308 115413 10310
rect 115469 10308 115493 10310
rect 115549 10308 115555 10310
rect 115247 10299 115555 10308
rect 117424 9926 117452 12922
rect 117700 11354 117728 13194
rect 118056 13184 118108 13190
rect 118056 13126 118108 13132
rect 118068 12850 118096 13126
rect 118252 12986 118280 13330
rect 118712 12986 118740 13654
rect 121288 13462 121316 15286
rect 124218 15200 124274 16000
rect 127346 15314 127402 16000
rect 126992 15286 127402 15314
rect 124232 13682 124260 15200
rect 125508 13796 125560 13802
rect 125508 13738 125560 13744
rect 124140 13654 124260 13682
rect 124140 13462 124168 13654
rect 118884 13456 118936 13462
rect 118884 13398 118936 13404
rect 121276 13456 121328 13462
rect 121276 13398 121328 13404
rect 124128 13456 124180 13462
rect 124128 13398 124180 13404
rect 118792 13320 118844 13326
rect 118792 13262 118844 13268
rect 118240 12980 118292 12986
rect 118240 12922 118292 12928
rect 118700 12980 118752 12986
rect 118700 12922 118752 12928
rect 118056 12844 118108 12850
rect 118056 12786 118108 12792
rect 118068 12238 118096 12786
rect 118056 12232 118108 12238
rect 118056 12174 118108 12180
rect 118252 12170 118280 12922
rect 118332 12232 118384 12238
rect 118332 12174 118384 12180
rect 118240 12164 118292 12170
rect 118240 12106 118292 12112
rect 118344 11762 118372 12174
rect 118804 11898 118832 13262
rect 118896 12306 118924 13398
rect 125520 13258 125548 13738
rect 125508 13252 125560 13258
rect 125508 13194 125560 13200
rect 119712 13184 119764 13190
rect 119712 13126 119764 13132
rect 126152 13184 126204 13190
rect 126152 13126 126204 13132
rect 126520 13184 126572 13190
rect 126520 13126 126572 13132
rect 118884 12300 118936 12306
rect 118884 12242 118936 12248
rect 118792 11892 118844 11898
rect 118792 11834 118844 11840
rect 118332 11756 118384 11762
rect 118332 11698 118384 11704
rect 117688 11348 117740 11354
rect 117688 11290 117740 11296
rect 119724 11150 119752 13126
rect 126164 12238 126192 13126
rect 126532 12918 126560 13126
rect 126992 13002 127020 15286
rect 127346 15200 127402 15286
rect 130382 15200 130438 16000
rect 133418 15314 133474 16000
rect 133418 15286 133828 15314
rect 133418 15200 133474 15286
rect 127440 13728 127492 13734
rect 127440 13670 127492 13676
rect 127532 13728 127584 13734
rect 127532 13670 127584 13676
rect 129740 13728 129792 13734
rect 129740 13670 129792 13676
rect 126900 12986 127020 13002
rect 126888 12980 127020 12986
rect 126940 12974 127020 12980
rect 126888 12922 126940 12928
rect 126520 12912 126572 12918
rect 126520 12854 126572 12860
rect 127452 12850 127480 13670
rect 127544 13462 127572 13670
rect 127532 13456 127584 13462
rect 127532 13398 127584 13404
rect 127532 13320 127584 13326
rect 127532 13262 127584 13268
rect 129372 13320 129424 13326
rect 129372 13262 129424 13268
rect 127440 12844 127492 12850
rect 127440 12786 127492 12792
rect 127544 12782 127572 13262
rect 127808 13252 127860 13258
rect 127808 13194 127860 13200
rect 127532 12776 127584 12782
rect 127532 12718 127584 12724
rect 127820 12442 127848 13194
rect 128084 13184 128136 13190
rect 128084 13126 128136 13132
rect 129188 13184 129240 13190
rect 129188 13126 129240 13132
rect 128096 12986 128124 13126
rect 129200 12986 129228 13126
rect 128084 12980 128136 12986
rect 128084 12922 128136 12928
rect 128636 12980 128688 12986
rect 128636 12922 128688 12928
rect 129188 12980 129240 12986
rect 129188 12922 129240 12928
rect 128360 12776 128412 12782
rect 128360 12718 128412 12724
rect 128084 12640 128136 12646
rect 128372 12594 128400 12718
rect 128136 12588 128400 12594
rect 128084 12582 128400 12588
rect 128096 12566 128400 12582
rect 127808 12436 127860 12442
rect 127808 12378 127860 12384
rect 126152 12232 126204 12238
rect 126152 12174 126204 12180
rect 128372 11762 128400 12566
rect 128648 12238 128676 12922
rect 129096 12844 129148 12850
rect 129096 12786 129148 12792
rect 129108 12442 129136 12786
rect 129096 12436 129148 12442
rect 129096 12378 129148 12384
rect 128636 12232 128688 12238
rect 128636 12174 128688 12180
rect 129384 11898 129412 13262
rect 129752 12782 129780 13670
rect 130292 13388 130344 13394
rect 130292 13330 130344 13336
rect 130304 12850 130332 13330
rect 130292 12844 130344 12850
rect 130292 12786 130344 12792
rect 129740 12776 129792 12782
rect 129740 12718 129792 12724
rect 129372 11892 129424 11898
rect 129372 11834 129424 11840
rect 128360 11756 128412 11762
rect 128360 11698 128412 11704
rect 129752 11694 129780 12718
rect 130292 12708 130344 12714
rect 130292 12650 130344 12656
rect 130304 11898 130332 12650
rect 130292 11892 130344 11898
rect 130292 11834 130344 11840
rect 130292 11756 130344 11762
rect 130292 11698 130344 11704
rect 129740 11688 129792 11694
rect 129740 11630 129792 11636
rect 130304 11218 130332 11698
rect 130396 11354 130424 15200
rect 131856 13796 131908 13802
rect 131856 13738 131908 13744
rect 131212 13252 131264 13258
rect 131212 13194 131264 13200
rect 131120 12776 131172 12782
rect 131120 12718 131172 12724
rect 130936 12436 130988 12442
rect 130936 12378 130988 12384
rect 130476 12232 130528 12238
rect 130476 12174 130528 12180
rect 130384 11348 130436 11354
rect 130384 11290 130436 11296
rect 130292 11212 130344 11218
rect 130292 11154 130344 11160
rect 119712 11144 119764 11150
rect 119712 11086 119764 11092
rect 130304 10674 130332 11154
rect 130488 10810 130516 12174
rect 130948 11898 130976 12378
rect 131028 12300 131080 12306
rect 131028 12242 131080 12248
rect 130936 11892 130988 11898
rect 130936 11834 130988 11840
rect 130948 11150 130976 11834
rect 131040 11694 131068 12242
rect 131132 11898 131160 12718
rect 131120 11892 131172 11898
rect 131120 11834 131172 11840
rect 131028 11688 131080 11694
rect 131028 11630 131080 11636
rect 131224 11354 131252 13194
rect 131580 13184 131632 13190
rect 131580 13126 131632 13132
rect 131592 12102 131620 13126
rect 131580 12096 131632 12102
rect 131580 12038 131632 12044
rect 131592 11762 131620 12038
rect 131580 11756 131632 11762
rect 131580 11698 131632 11704
rect 131868 11558 131896 13738
rect 133604 13728 133656 13734
rect 133604 13670 133656 13676
rect 132868 13252 132920 13258
rect 132868 13194 132920 13200
rect 133328 13252 133380 13258
rect 133328 13194 133380 13200
rect 132408 12912 132460 12918
rect 132408 12854 132460 12860
rect 132420 12442 132448 12854
rect 132592 12776 132644 12782
rect 132592 12718 132644 12724
rect 132408 12436 132460 12442
rect 132408 12378 132460 12384
rect 132604 12322 132632 12718
rect 132420 12294 132632 12322
rect 132420 12238 132448 12294
rect 132408 12232 132460 12238
rect 132408 12174 132460 12180
rect 132592 12232 132644 12238
rect 132592 12174 132644 12180
rect 132500 12164 132552 12170
rect 132500 12106 132552 12112
rect 132512 11762 132540 12106
rect 132500 11756 132552 11762
rect 132500 11698 132552 11704
rect 131856 11552 131908 11558
rect 131856 11494 131908 11500
rect 131212 11348 131264 11354
rect 131212 11290 131264 11296
rect 132604 11218 132632 12174
rect 132880 11354 132908 13194
rect 133340 12986 133368 13194
rect 133328 12980 133380 12986
rect 133328 12922 133380 12928
rect 133616 12918 133644 13670
rect 133800 13274 133828 15286
rect 136546 15200 136602 16000
rect 139582 15200 139638 16000
rect 142710 15314 142766 16000
rect 142710 15286 142936 15314
rect 142710 15200 142766 15286
rect 136560 13682 136588 15200
rect 136824 13728 136876 13734
rect 136560 13654 136680 13682
rect 136824 13670 136876 13676
rect 136652 13462 136680 13654
rect 136640 13456 136692 13462
rect 136640 13398 136692 13404
rect 136836 13326 136864 13670
rect 139596 13462 139624 15200
rect 142908 13530 142936 15286
rect 145746 15200 145802 16000
rect 148782 15314 148838 16000
rect 148520 15286 148838 15314
rect 145760 13530 145788 15200
rect 148140 13728 148192 13734
rect 148140 13670 148192 13676
rect 148152 13530 148180 13670
rect 142896 13524 142948 13530
rect 142896 13466 142948 13472
rect 145748 13524 145800 13530
rect 145748 13466 145800 13472
rect 148140 13524 148192 13530
rect 148140 13466 148192 13472
rect 139584 13456 139636 13462
rect 139584 13398 139636 13404
rect 142068 13388 142120 13394
rect 142068 13330 142120 13336
rect 136824 13320 136876 13326
rect 133800 13246 133920 13274
rect 136824 13262 136876 13268
rect 133696 13184 133748 13190
rect 133696 13126 133748 13132
rect 133604 12912 133656 12918
rect 133604 12854 133656 12860
rect 133708 12850 133736 13126
rect 133892 12986 133920 13246
rect 134156 13184 134208 13190
rect 134156 13126 134208 13132
rect 133880 12980 133932 12986
rect 133880 12922 133932 12928
rect 134168 12918 134196 13126
rect 134156 12912 134208 12918
rect 134156 12854 134208 12860
rect 133696 12844 133748 12850
rect 133696 12786 133748 12792
rect 133708 12714 133920 12730
rect 133696 12708 133932 12714
rect 133748 12702 133880 12708
rect 133696 12650 133748 12656
rect 133880 12650 133932 12656
rect 133144 12640 133196 12646
rect 133144 12582 133196 12588
rect 133236 12640 133288 12646
rect 133236 12582 133288 12588
rect 132868 11348 132920 11354
rect 132868 11290 132920 11296
rect 132592 11212 132644 11218
rect 132592 11154 132644 11160
rect 133156 11150 133184 12582
rect 133248 12306 133276 12582
rect 141976 12368 142028 12374
rect 141976 12310 142028 12316
rect 133236 12300 133288 12306
rect 133236 12242 133288 12248
rect 137744 12232 137796 12238
rect 137744 12174 137796 12180
rect 137756 11898 137784 12174
rect 138020 12164 138072 12170
rect 138020 12106 138072 12112
rect 137744 11892 137796 11898
rect 137744 11834 137796 11840
rect 137756 11694 137784 11834
rect 138032 11830 138060 12106
rect 138020 11824 138072 11830
rect 138020 11766 138072 11772
rect 137744 11688 137796 11694
rect 137744 11630 137796 11636
rect 130936 11144 130988 11150
rect 130936 11086 130988 11092
rect 133144 11144 133196 11150
rect 133144 11086 133196 11092
rect 140688 11076 140740 11082
rect 140688 11018 140740 11024
rect 130476 10804 130528 10810
rect 130476 10746 130528 10752
rect 140700 10742 140728 11018
rect 141988 10810 142016 12310
rect 142080 11150 142108 13330
rect 143080 13320 143132 13326
rect 143080 13262 143132 13268
rect 145748 13320 145800 13326
rect 145748 13262 145800 13268
rect 143092 12918 143120 13262
rect 143080 12912 143132 12918
rect 143080 12854 143132 12860
rect 143264 12776 143316 12782
rect 143264 12718 143316 12724
rect 143276 11626 143304 12718
rect 145760 12714 145788 13262
rect 145932 13252 145984 13258
rect 145932 13194 145984 13200
rect 146024 13252 146076 13258
rect 146024 13194 146076 13200
rect 147588 13252 147640 13258
rect 147588 13194 147640 13200
rect 145840 13184 145892 13190
rect 145840 13126 145892 13132
rect 145852 12850 145880 13126
rect 145944 12918 145972 13194
rect 145932 12912 145984 12918
rect 145932 12854 145984 12860
rect 145840 12844 145892 12850
rect 145840 12786 145892 12792
rect 145748 12708 145800 12714
rect 145748 12650 145800 12656
rect 143264 11620 143316 11626
rect 143264 11562 143316 11568
rect 143276 11218 143304 11562
rect 143264 11212 143316 11218
rect 143264 11154 143316 11160
rect 145760 11150 145788 12650
rect 146036 11626 146064 13194
rect 147496 13184 147548 13190
rect 147496 13126 147548 13132
rect 147312 12844 147364 12850
rect 147312 12786 147364 12792
rect 146024 11620 146076 11626
rect 146024 11562 146076 11568
rect 147324 11558 147352 12786
rect 147404 12776 147456 12782
rect 147404 12718 147456 12724
rect 147312 11552 147364 11558
rect 147312 11494 147364 11500
rect 147416 11286 147444 12718
rect 147404 11280 147456 11286
rect 147404 11222 147456 11228
rect 147508 11218 147536 13126
rect 147600 12374 147628 13194
rect 147680 12980 147732 12986
rect 147680 12922 147732 12928
rect 147588 12368 147640 12374
rect 147588 12310 147640 12316
rect 147692 11762 147720 12922
rect 147772 12776 147824 12782
rect 147772 12718 147824 12724
rect 147784 12442 147812 12718
rect 148520 12646 148548 15286
rect 148782 15200 148838 15286
rect 151910 15314 151966 16000
rect 151910 15286 152044 15314
rect 151910 15200 151966 15286
rect 150440 13728 150492 13734
rect 150440 13670 150492 13676
rect 150452 13258 150480 13670
rect 150808 13524 150860 13530
rect 150808 13466 150860 13472
rect 150440 13252 150492 13258
rect 150440 13194 150492 13200
rect 149244 13184 149296 13190
rect 149244 13126 149296 13132
rect 149256 12782 149284 13126
rect 150452 12850 150480 13194
rect 149336 12844 149388 12850
rect 149336 12786 149388 12792
rect 150440 12844 150492 12850
rect 150440 12786 150492 12792
rect 148968 12776 149020 12782
rect 149244 12776 149296 12782
rect 148968 12718 149020 12724
rect 149072 12736 149244 12764
rect 148508 12640 148560 12646
rect 148508 12582 148560 12588
rect 147772 12436 147824 12442
rect 147772 12378 147824 12384
rect 148048 12232 148100 12238
rect 148048 12174 148100 12180
rect 147680 11756 147732 11762
rect 147680 11698 147732 11704
rect 148060 11354 148088 12174
rect 148324 11688 148376 11694
rect 148324 11630 148376 11636
rect 148600 11688 148652 11694
rect 148600 11630 148652 11636
rect 148048 11348 148100 11354
rect 148048 11290 148100 11296
rect 147496 11212 147548 11218
rect 147496 11154 147548 11160
rect 142068 11144 142120 11150
rect 142068 11086 142120 11092
rect 145748 11144 145800 11150
rect 145748 11086 145800 11092
rect 141976 10804 142028 10810
rect 141976 10746 142028 10752
rect 140688 10736 140740 10742
rect 140688 10678 140740 10684
rect 130292 10668 130344 10674
rect 130292 10610 130344 10616
rect 140700 10062 140728 10678
rect 140688 10056 140740 10062
rect 140688 9998 140740 10004
rect 117412 9920 117464 9926
rect 117412 9862 117464 9868
rect 140700 9654 140728 9998
rect 140688 9648 140740 9654
rect 140688 9590 140740 9596
rect 148336 9382 148364 11630
rect 148612 10810 148640 11630
rect 148980 10810 149008 12718
rect 149072 12306 149100 12736
rect 149244 12718 149296 12724
rect 149060 12300 149112 12306
rect 149060 12242 149112 12248
rect 149072 11014 149100 12242
rect 149348 12238 149376 12786
rect 150348 12708 150400 12714
rect 150348 12650 150400 12656
rect 149980 12640 150032 12646
rect 149980 12582 150032 12588
rect 149336 12232 149388 12238
rect 149336 12174 149388 12180
rect 149428 12232 149480 12238
rect 149428 12174 149480 12180
rect 149060 11008 149112 11014
rect 149060 10950 149112 10956
rect 148600 10804 148652 10810
rect 148600 10746 148652 10752
rect 148968 10804 149020 10810
rect 148968 10746 149020 10752
rect 104256 9376 104308 9382
rect 104256 9318 104308 9324
rect 148324 9376 148376 9382
rect 148324 9318 148376 9324
rect 39049 9276 39357 9285
rect 39049 9274 39055 9276
rect 39111 9274 39135 9276
rect 39191 9274 39215 9276
rect 39271 9274 39295 9276
rect 39351 9274 39357 9276
rect 39111 9222 39113 9274
rect 39293 9222 39295 9274
rect 39049 9220 39055 9222
rect 39111 9220 39135 9222
rect 39191 9220 39215 9222
rect 39271 9220 39295 9222
rect 39351 9220 39357 9222
rect 39049 9211 39357 9220
rect 115247 9276 115555 9285
rect 115247 9274 115253 9276
rect 115309 9274 115333 9276
rect 115389 9274 115413 9276
rect 115469 9274 115493 9276
rect 115549 9274 115555 9276
rect 115309 9222 115311 9274
rect 115491 9222 115493 9274
rect 115247 9220 115253 9222
rect 115309 9220 115333 9222
rect 115389 9220 115413 9222
rect 115469 9220 115493 9222
rect 115549 9220 115555 9222
rect 115247 9211 115555 9220
rect 77148 8732 77456 8741
rect 77148 8730 77154 8732
rect 77210 8730 77234 8732
rect 77290 8730 77314 8732
rect 77370 8730 77394 8732
rect 77450 8730 77456 8732
rect 77210 8678 77212 8730
rect 77392 8678 77394 8730
rect 77148 8676 77154 8678
rect 77210 8676 77234 8678
rect 77290 8676 77314 8678
rect 77370 8676 77394 8678
rect 77450 8676 77456 8678
rect 77148 8667 77456 8676
rect 1400 8356 1452 8362
rect 1400 8298 1452 8304
rect 1412 8129 1440 8298
rect 39049 8188 39357 8197
rect 39049 8186 39055 8188
rect 39111 8186 39135 8188
rect 39191 8186 39215 8188
rect 39271 8186 39295 8188
rect 39351 8186 39357 8188
rect 39111 8134 39113 8186
rect 39293 8134 39295 8186
rect 39049 8132 39055 8134
rect 39111 8132 39135 8134
rect 39191 8132 39215 8134
rect 39271 8132 39295 8134
rect 39351 8132 39357 8134
rect 1398 8120 1454 8129
rect 39049 8123 39357 8132
rect 115247 8188 115555 8197
rect 115247 8186 115253 8188
rect 115309 8186 115333 8188
rect 115389 8186 115413 8188
rect 115469 8186 115493 8188
rect 115549 8186 115555 8188
rect 115309 8134 115311 8186
rect 115491 8134 115493 8186
rect 115247 8132 115253 8134
rect 115309 8132 115333 8134
rect 115389 8132 115413 8134
rect 115469 8132 115493 8134
rect 115549 8132 115555 8134
rect 115247 8123 115555 8132
rect 1398 8055 1454 8064
rect 77148 7644 77456 7653
rect 77148 7642 77154 7644
rect 77210 7642 77234 7644
rect 77290 7642 77314 7644
rect 77370 7642 77394 7644
rect 77450 7642 77456 7644
rect 77210 7590 77212 7642
rect 77392 7590 77394 7642
rect 77148 7588 77154 7590
rect 77210 7588 77234 7590
rect 77290 7588 77314 7590
rect 77370 7588 77394 7590
rect 77450 7588 77456 7590
rect 77148 7579 77456 7588
rect 39049 7100 39357 7109
rect 39049 7098 39055 7100
rect 39111 7098 39135 7100
rect 39191 7098 39215 7100
rect 39271 7098 39295 7100
rect 39351 7098 39357 7100
rect 39111 7046 39113 7098
rect 39293 7046 39295 7098
rect 39049 7044 39055 7046
rect 39111 7044 39135 7046
rect 39191 7044 39215 7046
rect 39271 7044 39295 7046
rect 39351 7044 39357 7046
rect 39049 7035 39357 7044
rect 115247 7100 115555 7109
rect 115247 7098 115253 7100
rect 115309 7098 115333 7100
rect 115389 7098 115413 7100
rect 115469 7098 115493 7100
rect 115549 7098 115555 7100
rect 115309 7046 115311 7098
rect 115491 7046 115493 7098
rect 115247 7044 115253 7046
rect 115309 7044 115333 7046
rect 115389 7044 115413 7046
rect 115469 7044 115493 7046
rect 115549 7044 115555 7046
rect 115247 7035 115555 7044
rect 77148 6556 77456 6565
rect 77148 6554 77154 6556
rect 77210 6554 77234 6556
rect 77290 6554 77314 6556
rect 77370 6554 77394 6556
rect 77450 6554 77456 6556
rect 77210 6502 77212 6554
rect 77392 6502 77394 6554
rect 77148 6500 77154 6502
rect 77210 6500 77234 6502
rect 77290 6500 77314 6502
rect 77370 6500 77394 6502
rect 77450 6500 77456 6502
rect 77148 6491 77456 6500
rect 39049 6012 39357 6021
rect 39049 6010 39055 6012
rect 39111 6010 39135 6012
rect 39191 6010 39215 6012
rect 39271 6010 39295 6012
rect 39351 6010 39357 6012
rect 39111 5958 39113 6010
rect 39293 5958 39295 6010
rect 39049 5956 39055 5958
rect 39111 5956 39135 5958
rect 39191 5956 39215 5958
rect 39271 5956 39295 5958
rect 39351 5956 39357 5958
rect 39049 5947 39357 5956
rect 115247 6012 115555 6021
rect 115247 6010 115253 6012
rect 115309 6010 115333 6012
rect 115389 6010 115413 6012
rect 115469 6010 115493 6012
rect 115549 6010 115555 6012
rect 115309 5958 115311 6010
rect 115491 5958 115493 6010
rect 115247 5956 115253 5958
rect 115309 5956 115333 5958
rect 115389 5956 115413 5958
rect 115469 5956 115493 5958
rect 115549 5956 115555 5958
rect 115247 5947 115555 5956
rect 77148 5468 77456 5477
rect 77148 5466 77154 5468
rect 77210 5466 77234 5468
rect 77290 5466 77314 5468
rect 77370 5466 77394 5468
rect 77450 5466 77456 5468
rect 77210 5414 77212 5466
rect 77392 5414 77394 5466
rect 77148 5412 77154 5414
rect 77210 5412 77234 5414
rect 77290 5412 77314 5414
rect 77370 5412 77394 5414
rect 77450 5412 77456 5414
rect 77148 5403 77456 5412
rect 39049 4924 39357 4933
rect 39049 4922 39055 4924
rect 39111 4922 39135 4924
rect 39191 4922 39215 4924
rect 39271 4922 39295 4924
rect 39351 4922 39357 4924
rect 39111 4870 39113 4922
rect 39293 4870 39295 4922
rect 39049 4868 39055 4870
rect 39111 4868 39135 4870
rect 39191 4868 39215 4870
rect 39271 4868 39295 4870
rect 39351 4868 39357 4870
rect 39049 4859 39357 4868
rect 115247 4924 115555 4933
rect 115247 4922 115253 4924
rect 115309 4922 115333 4924
rect 115389 4922 115413 4924
rect 115469 4922 115493 4924
rect 115549 4922 115555 4924
rect 115309 4870 115311 4922
rect 115491 4870 115493 4922
rect 115247 4868 115253 4870
rect 115309 4868 115333 4870
rect 115389 4868 115413 4870
rect 115469 4868 115493 4870
rect 115549 4868 115555 4870
rect 115247 4859 115555 4868
rect 77148 4380 77456 4389
rect 77148 4378 77154 4380
rect 77210 4378 77234 4380
rect 77290 4378 77314 4380
rect 77370 4378 77394 4380
rect 77450 4378 77456 4380
rect 77210 4326 77212 4378
rect 77392 4326 77394 4378
rect 77148 4324 77154 4326
rect 77210 4324 77234 4326
rect 77290 4324 77314 4326
rect 77370 4324 77394 4326
rect 77450 4324 77456 4326
rect 77148 4315 77456 4324
rect 39049 3836 39357 3845
rect 39049 3834 39055 3836
rect 39111 3834 39135 3836
rect 39191 3834 39215 3836
rect 39271 3834 39295 3836
rect 39351 3834 39357 3836
rect 39111 3782 39113 3834
rect 39293 3782 39295 3834
rect 39049 3780 39055 3782
rect 39111 3780 39135 3782
rect 39191 3780 39215 3782
rect 39271 3780 39295 3782
rect 39351 3780 39357 3782
rect 39049 3771 39357 3780
rect 115247 3836 115555 3845
rect 115247 3834 115253 3836
rect 115309 3834 115333 3836
rect 115389 3834 115413 3836
rect 115469 3834 115493 3836
rect 115549 3834 115555 3836
rect 115309 3782 115311 3834
rect 115491 3782 115493 3834
rect 115247 3780 115253 3782
rect 115309 3780 115333 3782
rect 115389 3780 115413 3782
rect 115469 3780 115493 3782
rect 115549 3780 115555 3782
rect 115247 3771 115555 3780
rect 77148 3292 77456 3301
rect 77148 3290 77154 3292
rect 77210 3290 77234 3292
rect 77290 3290 77314 3292
rect 77370 3290 77394 3292
rect 77450 3290 77456 3292
rect 77210 3238 77212 3290
rect 77392 3238 77394 3290
rect 77148 3236 77154 3238
rect 77210 3236 77234 3238
rect 77290 3236 77314 3238
rect 77370 3236 77394 3238
rect 77450 3236 77456 3238
rect 77148 3227 77456 3236
rect 39049 2748 39357 2757
rect 39049 2746 39055 2748
rect 39111 2746 39135 2748
rect 39191 2746 39215 2748
rect 39271 2746 39295 2748
rect 39351 2746 39357 2748
rect 39111 2694 39113 2746
rect 39293 2694 39295 2746
rect 39049 2692 39055 2694
rect 39111 2692 39135 2694
rect 39191 2692 39215 2694
rect 39271 2692 39295 2694
rect 39351 2692 39357 2694
rect 39049 2683 39357 2692
rect 115247 2748 115555 2757
rect 115247 2746 115253 2748
rect 115309 2746 115333 2748
rect 115389 2746 115413 2748
rect 115469 2746 115493 2748
rect 115549 2746 115555 2748
rect 115309 2694 115311 2746
rect 115491 2694 115493 2746
rect 115247 2692 115253 2694
rect 115309 2692 115333 2694
rect 115389 2692 115413 2694
rect 115469 2692 115493 2694
rect 115549 2692 115555 2694
rect 115247 2683 115555 2692
rect 149440 2650 149468 12174
rect 149520 12096 149572 12102
rect 149520 12038 149572 12044
rect 149532 11014 149560 12038
rect 149992 11830 150020 12582
rect 149980 11824 150032 11830
rect 149980 11766 150032 11772
rect 149520 11008 149572 11014
rect 149520 10950 149572 10956
rect 150360 10674 150388 12650
rect 150820 11354 150848 13466
rect 151084 13252 151136 13258
rect 151084 13194 151136 13200
rect 151096 11898 151124 13194
rect 151544 12776 151596 12782
rect 151544 12718 151596 12724
rect 151268 12640 151320 12646
rect 151268 12582 151320 12588
rect 151360 12640 151412 12646
rect 151360 12582 151412 12588
rect 151084 11892 151136 11898
rect 151084 11834 151136 11840
rect 151280 11762 151308 12582
rect 151372 12238 151400 12582
rect 151360 12232 151412 12238
rect 151360 12174 151412 12180
rect 151556 12186 151584 12718
rect 151636 12708 151688 12714
rect 151636 12650 151688 12656
rect 151648 12374 151676 12650
rect 151636 12368 151688 12374
rect 151636 12310 151688 12316
rect 151268 11756 151320 11762
rect 151268 11698 151320 11704
rect 150808 11348 150860 11354
rect 150808 11290 150860 11296
rect 151372 11218 151400 12174
rect 151556 12158 151768 12186
rect 151740 12102 151768 12158
rect 151636 12096 151688 12102
rect 151636 12038 151688 12044
rect 151728 12096 151780 12102
rect 151728 12038 151780 12044
rect 151360 11212 151412 11218
rect 151360 11154 151412 11160
rect 151648 10742 151676 12038
rect 151740 11558 151768 12038
rect 152016 11898 152044 15286
rect 154946 15200 155002 16000
rect 157982 15200 158038 16000
rect 161110 15314 161166 16000
rect 161110 15286 161336 15314
rect 161110 15200 161166 15286
rect 154960 13462 154988 15200
rect 157156 13728 157208 13734
rect 157156 13670 157208 13676
rect 154948 13456 155000 13462
rect 154948 13398 155000 13404
rect 155224 13320 155276 13326
rect 155224 13262 155276 13268
rect 155868 13320 155920 13326
rect 155868 13262 155920 13268
rect 156420 13320 156472 13326
rect 156420 13262 156472 13268
rect 152464 13252 152516 13258
rect 152464 13194 152516 13200
rect 153752 13252 153804 13258
rect 153752 13194 153804 13200
rect 154212 13252 154264 13258
rect 154212 13194 154264 13200
rect 152476 12442 152504 13194
rect 152648 13184 152700 13190
rect 152648 13126 152700 13132
rect 152660 12986 152688 13126
rect 153346 13084 153654 13093
rect 153346 13082 153352 13084
rect 153408 13082 153432 13084
rect 153488 13082 153512 13084
rect 153568 13082 153592 13084
rect 153648 13082 153654 13084
rect 153408 13030 153410 13082
rect 153590 13030 153592 13082
rect 153346 13028 153352 13030
rect 153408 13028 153432 13030
rect 153488 13028 153512 13030
rect 153568 13028 153592 13030
rect 153648 13028 153654 13030
rect 153346 13019 153654 13028
rect 152648 12980 152700 12986
rect 152648 12922 152700 12928
rect 152832 12980 152884 12986
rect 152832 12922 152884 12928
rect 152660 12832 152688 12922
rect 152568 12804 152688 12832
rect 152464 12436 152516 12442
rect 152464 12378 152516 12384
rect 152568 12102 152596 12804
rect 152740 12776 152792 12782
rect 152740 12718 152792 12724
rect 152752 12374 152780 12718
rect 152844 12714 152872 12922
rect 152832 12708 152884 12714
rect 152832 12650 152884 12656
rect 153108 12708 153160 12714
rect 153108 12650 153160 12656
rect 152740 12368 152792 12374
rect 152740 12310 152792 12316
rect 152188 12096 152240 12102
rect 152188 12038 152240 12044
rect 152556 12096 152608 12102
rect 152556 12038 152608 12044
rect 152004 11892 152056 11898
rect 152004 11834 152056 11840
rect 152200 11762 152228 12038
rect 152752 11762 152780 12310
rect 152188 11756 152240 11762
rect 152188 11698 152240 11704
rect 152740 11756 152792 11762
rect 152740 11698 152792 11704
rect 151728 11552 151780 11558
rect 151728 11494 151780 11500
rect 153120 11150 153148 12650
rect 153764 12442 153792 13194
rect 154120 12640 154172 12646
rect 154120 12582 154172 12588
rect 153752 12436 153804 12442
rect 153752 12378 153804 12384
rect 154132 12306 154160 12582
rect 154120 12300 154172 12306
rect 154120 12242 154172 12248
rect 153346 11996 153654 12005
rect 153346 11994 153352 11996
rect 153408 11994 153432 11996
rect 153488 11994 153512 11996
rect 153568 11994 153592 11996
rect 153648 11994 153654 11996
rect 153408 11942 153410 11994
rect 153590 11942 153592 11994
rect 153346 11940 153352 11942
rect 153408 11940 153432 11942
rect 153488 11940 153512 11942
rect 153568 11940 153592 11942
rect 153648 11940 153654 11942
rect 153346 11931 153654 11940
rect 154224 11898 154252 13194
rect 155236 13190 155264 13262
rect 155224 13184 155276 13190
rect 155224 13126 155276 13132
rect 155038 12880 155094 12889
rect 155880 12850 155908 13262
rect 155038 12815 155094 12824
rect 155868 12844 155920 12850
rect 155052 12782 155080 12815
rect 155868 12786 155920 12792
rect 155040 12776 155092 12782
rect 155040 12718 155092 12724
rect 155052 12374 155080 12718
rect 155040 12368 155092 12374
rect 155040 12310 155092 12316
rect 155880 12170 155908 12786
rect 156432 12170 156460 13262
rect 156604 13252 156656 13258
rect 156604 13194 156656 13200
rect 156616 12918 156644 13194
rect 157168 12986 157196 13670
rect 157996 13530 158024 15200
rect 157248 13524 157300 13530
rect 157248 13466 157300 13472
rect 157984 13524 158036 13530
rect 157984 13466 158036 13472
rect 159456 13524 159508 13530
rect 159456 13466 159508 13472
rect 157156 12980 157208 12986
rect 157156 12922 157208 12928
rect 156604 12912 156656 12918
rect 156604 12854 156656 12860
rect 157260 12442 157288 13466
rect 157800 13320 157852 13326
rect 157800 13262 157852 13268
rect 158628 13320 158680 13326
rect 158628 13262 158680 13268
rect 157812 12850 157840 13262
rect 158640 12986 158668 13262
rect 158904 13252 158956 13258
rect 158904 13194 158956 13200
rect 158628 12980 158680 12986
rect 158628 12922 158680 12928
rect 157800 12844 157852 12850
rect 157800 12786 157852 12792
rect 157892 12640 157944 12646
rect 157890 12608 157892 12617
rect 157944 12608 157946 12617
rect 157890 12543 157946 12552
rect 157248 12436 157300 12442
rect 157248 12378 157300 12384
rect 155868 12164 155920 12170
rect 155868 12106 155920 12112
rect 156420 12164 156472 12170
rect 156420 12106 156472 12112
rect 154212 11892 154264 11898
rect 154212 11834 154264 11840
rect 156432 11286 156460 12106
rect 157260 11354 157288 12378
rect 157248 11348 157300 11354
rect 157248 11290 157300 11296
rect 156420 11280 156472 11286
rect 156420 11222 156472 11228
rect 153108 11144 153160 11150
rect 153108 11086 153160 11092
rect 156144 11076 156196 11082
rect 156144 11018 156196 11024
rect 153346 10908 153654 10917
rect 153346 10906 153352 10908
rect 153408 10906 153432 10908
rect 153488 10906 153512 10908
rect 153568 10906 153592 10908
rect 153648 10906 153654 10908
rect 153408 10854 153410 10906
rect 153590 10854 153592 10906
rect 153346 10852 153352 10854
rect 153408 10852 153432 10854
rect 153488 10852 153512 10854
rect 153568 10852 153592 10854
rect 153648 10852 153654 10854
rect 153346 10843 153654 10852
rect 156156 10742 156184 11018
rect 151636 10736 151688 10742
rect 151636 10678 151688 10684
rect 156144 10736 156196 10742
rect 156144 10678 156196 10684
rect 150348 10668 150400 10674
rect 150348 10610 150400 10616
rect 156156 10062 156184 10678
rect 156144 10056 156196 10062
rect 156144 9998 156196 10004
rect 153346 9820 153654 9829
rect 153346 9818 153352 9820
rect 153408 9818 153432 9820
rect 153488 9818 153512 9820
rect 153568 9818 153592 9820
rect 153648 9818 153654 9820
rect 153408 9766 153410 9818
rect 153590 9766 153592 9818
rect 153346 9764 153352 9766
rect 153408 9764 153432 9766
rect 153488 9764 153512 9766
rect 153568 9764 153592 9766
rect 153648 9764 153654 9766
rect 153346 9755 153654 9764
rect 156156 9654 156184 9998
rect 158640 9654 158668 12922
rect 158812 12708 158864 12714
rect 158812 12650 158864 12656
rect 158824 12238 158852 12650
rect 158916 12374 158944 13194
rect 159468 12782 159496 13466
rect 160928 13388 160980 13394
rect 160928 13330 160980 13336
rect 159548 13184 159600 13190
rect 159548 13126 159600 13132
rect 160376 13184 160428 13190
rect 160376 13126 160428 13132
rect 159560 12782 159588 13126
rect 160388 12918 160416 13126
rect 160376 12912 160428 12918
rect 160376 12854 160428 12860
rect 159456 12776 159508 12782
rect 159456 12718 159508 12724
rect 159548 12776 159600 12782
rect 159548 12718 159600 12724
rect 160284 12640 160336 12646
rect 160282 12608 160284 12617
rect 160336 12608 160338 12617
rect 160282 12543 160338 12552
rect 158904 12368 158956 12374
rect 158904 12310 158956 12316
rect 160388 12306 160416 12854
rect 160940 12442 160968 13330
rect 161204 13252 161256 13258
rect 161204 13194 161256 13200
rect 160928 12436 160980 12442
rect 160928 12378 160980 12384
rect 160376 12300 160428 12306
rect 160376 12242 160428 12248
rect 158812 12232 158864 12238
rect 158812 12174 158864 12180
rect 161112 12096 161164 12102
rect 161112 12038 161164 12044
rect 161124 11762 161152 12038
rect 161112 11756 161164 11762
rect 161112 11698 161164 11704
rect 161216 11626 161244 13194
rect 161308 11626 161336 15286
rect 164146 15200 164202 16000
rect 167182 15200 167238 16000
rect 170310 15314 170366 16000
rect 173346 15314 173402 16000
rect 170310 15286 170444 15314
rect 170310 15200 170366 15286
rect 161664 13796 161716 13802
rect 161664 13738 161716 13744
rect 161572 13524 161624 13530
rect 161492 13484 161572 13512
rect 161492 12306 161520 13484
rect 161572 13466 161624 13472
rect 161676 12850 161704 13738
rect 162676 13524 162728 13530
rect 162676 13466 162728 13472
rect 163504 13524 163556 13530
rect 163504 13466 163556 13472
rect 162688 13326 162716 13466
rect 163516 13326 163544 13466
rect 162676 13320 162728 13326
rect 162676 13262 162728 13268
rect 163504 13320 163556 13326
rect 163504 13262 163556 13268
rect 162032 13184 162084 13190
rect 162032 13126 162084 13132
rect 162492 13184 162544 13190
rect 162492 13126 162544 13132
rect 161664 12844 161716 12850
rect 161664 12786 161716 12792
rect 161572 12776 161624 12782
rect 161572 12718 161624 12724
rect 161584 12442 161612 12718
rect 161572 12436 161624 12442
rect 161572 12378 161624 12384
rect 161480 12300 161532 12306
rect 161480 12242 161532 12248
rect 161756 12232 161808 12238
rect 161756 12174 161808 12180
rect 161768 11762 161796 12174
rect 162044 11898 162072 13126
rect 162124 12776 162176 12782
rect 162124 12718 162176 12724
rect 162032 11892 162084 11898
rect 162032 11834 162084 11840
rect 161756 11756 161808 11762
rect 161756 11698 161808 11704
rect 161204 11620 161256 11626
rect 161204 11562 161256 11568
rect 161296 11620 161348 11626
rect 161296 11562 161348 11568
rect 162136 11354 162164 12718
rect 162504 12306 162532 13126
rect 162688 12306 162716 13262
rect 162768 13252 162820 13258
rect 162768 13194 162820 13200
rect 162492 12300 162544 12306
rect 162492 12242 162544 12248
rect 162676 12300 162728 12306
rect 162676 12242 162728 12248
rect 162584 12164 162636 12170
rect 162584 12106 162636 12112
rect 162676 12164 162728 12170
rect 162676 12106 162728 12112
rect 162216 12096 162268 12102
rect 162216 12038 162268 12044
rect 162124 11348 162176 11354
rect 162124 11290 162176 11296
rect 162228 11150 162256 12038
rect 162596 11830 162624 12106
rect 162584 11824 162636 11830
rect 162584 11766 162636 11772
rect 162688 11354 162716 12106
rect 162780 11898 162808 13194
rect 163516 12986 163544 13262
rect 163780 13252 163832 13258
rect 163780 13194 163832 13200
rect 163504 12980 163556 12986
rect 163504 12922 163556 12928
rect 163412 12912 163464 12918
rect 163412 12854 163464 12860
rect 162860 12776 162912 12782
rect 162860 12718 162912 12724
rect 162872 12102 162900 12718
rect 162860 12096 162912 12102
rect 162860 12038 162912 12044
rect 162768 11892 162820 11898
rect 162768 11834 162820 11840
rect 163424 11354 163452 12854
rect 163688 12640 163740 12646
rect 163688 12582 163740 12588
rect 163594 12336 163650 12345
rect 163594 12271 163596 12280
rect 163648 12271 163650 12280
rect 163596 12242 163648 12248
rect 163504 11688 163556 11694
rect 163504 11630 163556 11636
rect 162676 11348 162728 11354
rect 162676 11290 162728 11296
rect 163412 11348 163464 11354
rect 163412 11290 163464 11296
rect 163516 11150 163544 11630
rect 162216 11144 162268 11150
rect 162216 11086 162268 11092
rect 163504 11144 163556 11150
rect 163504 11086 163556 11092
rect 163608 10130 163636 12242
rect 163700 11762 163728 12582
rect 163792 11898 163820 13194
rect 164160 12730 164188 15200
rect 166080 13796 166132 13802
rect 166080 13738 166132 13744
rect 165252 13388 165304 13394
rect 165252 13330 165304 13336
rect 164884 13320 164936 13326
rect 165264 13274 165292 13330
rect 164884 13262 164936 13268
rect 164608 13184 164660 13190
rect 164608 13126 164660 13132
rect 164620 12782 164648 13126
rect 164608 12776 164660 12782
rect 164160 12714 164280 12730
rect 164608 12718 164660 12724
rect 164160 12708 164292 12714
rect 164160 12702 164240 12708
rect 164240 12650 164292 12656
rect 164332 12164 164384 12170
rect 164332 12106 164384 12112
rect 164344 11898 164372 12106
rect 164896 11898 164924 13262
rect 165172 13258 165292 13274
rect 165160 13252 165292 13258
rect 165212 13246 165292 13252
rect 165160 13194 165212 13200
rect 165252 13184 165304 13190
rect 165252 13126 165304 13132
rect 165344 13184 165396 13190
rect 165344 13126 165396 13132
rect 165264 12986 165292 13126
rect 165252 12980 165304 12986
rect 165252 12922 165304 12928
rect 163780 11892 163832 11898
rect 163780 11834 163832 11840
rect 164332 11892 164384 11898
rect 164332 11834 164384 11840
rect 164884 11892 164936 11898
rect 164884 11834 164936 11840
rect 163688 11756 163740 11762
rect 163688 11698 163740 11704
rect 165356 11218 165384 13126
rect 165436 12844 165488 12850
rect 165436 12786 165488 12792
rect 165448 12374 165476 12786
rect 166092 12374 166120 13738
rect 166448 13456 166500 13462
rect 166448 13398 166500 13404
rect 166460 13190 166488 13398
rect 166448 13184 166500 13190
rect 166448 13126 166500 13132
rect 166172 12844 166224 12850
rect 166172 12786 166224 12792
rect 166184 12646 166212 12786
rect 166172 12640 166224 12646
rect 166172 12582 166224 12588
rect 166460 12442 166488 13126
rect 167196 12986 167224 15200
rect 167368 13796 167420 13802
rect 167368 13738 167420 13744
rect 167380 13258 167408 13738
rect 170416 13462 170444 15286
rect 173084 15286 173402 15314
rect 173084 13462 173112 15286
rect 173346 15200 173402 15286
rect 176474 15200 176530 16000
rect 179510 15200 179566 16000
rect 182546 15314 182602 16000
rect 185674 15314 185730 16000
rect 182546 15286 182772 15314
rect 182546 15200 182602 15286
rect 174176 13796 174228 13802
rect 174176 13738 174228 13744
rect 170404 13456 170456 13462
rect 170404 13398 170456 13404
rect 173072 13456 173124 13462
rect 173072 13398 173124 13404
rect 173808 13456 173860 13462
rect 173808 13398 173860 13404
rect 167368 13252 167420 13258
rect 167368 13194 167420 13200
rect 167184 12980 167236 12986
rect 167184 12922 167236 12928
rect 173820 12918 173848 13398
rect 174188 13326 174216 13738
rect 175844 13518 176056 13546
rect 175844 13326 175872 13518
rect 176028 13462 176056 13518
rect 176384 13524 176436 13530
rect 176384 13466 176436 13472
rect 175924 13456 175976 13462
rect 175924 13398 175976 13404
rect 176016 13456 176068 13462
rect 176016 13398 176068 13404
rect 174176 13320 174228 13326
rect 174176 13262 174228 13268
rect 175832 13320 175884 13326
rect 175832 13262 175884 13268
rect 175740 13252 175792 13258
rect 175740 13194 175792 13200
rect 175004 13184 175056 13190
rect 175004 13126 175056 13132
rect 175016 12986 175044 13126
rect 175752 12986 175780 13194
rect 175004 12980 175056 12986
rect 175004 12922 175056 12928
rect 175740 12980 175792 12986
rect 175740 12922 175792 12928
rect 175936 12918 175964 13398
rect 176396 13326 176424 13466
rect 176384 13320 176436 13326
rect 176384 13262 176436 13268
rect 176396 12986 176424 13262
rect 176384 12980 176436 12986
rect 176384 12922 176436 12928
rect 173808 12912 173860 12918
rect 173808 12854 173860 12860
rect 175924 12912 175976 12918
rect 175924 12854 175976 12860
rect 176396 12850 176424 12922
rect 166540 12844 166592 12850
rect 166540 12786 166592 12792
rect 176384 12844 176436 12850
rect 176384 12786 176436 12792
rect 166448 12436 166500 12442
rect 166448 12378 166500 12384
rect 165436 12368 165488 12374
rect 165436 12310 165488 12316
rect 166080 12368 166132 12374
rect 166080 12310 166132 12316
rect 165448 11286 165476 12310
rect 166552 12170 166580 12786
rect 166632 12640 166684 12646
rect 166632 12582 166684 12588
rect 165896 12164 165948 12170
rect 165896 12106 165948 12112
rect 166540 12164 166592 12170
rect 166540 12106 166592 12112
rect 165908 11626 165936 12106
rect 166644 11762 166672 12582
rect 176488 12442 176516 15200
rect 177764 13796 177816 13802
rect 177764 13738 177816 13744
rect 177776 13462 177804 13738
rect 177764 13456 177816 13462
rect 177764 13398 177816 13404
rect 177672 13252 177724 13258
rect 177672 13194 177724 13200
rect 176936 12912 176988 12918
rect 176936 12854 176988 12860
rect 176752 12776 176804 12782
rect 176752 12718 176804 12724
rect 176476 12436 176528 12442
rect 176476 12378 176528 12384
rect 176660 12096 176712 12102
rect 176660 12038 176712 12044
rect 176672 11762 176700 12038
rect 176764 11898 176792 12718
rect 176948 12458 176976 12854
rect 177396 12640 177448 12646
rect 177396 12582 177448 12588
rect 176948 12430 177160 12458
rect 177132 12306 177160 12430
rect 177120 12300 177172 12306
rect 177120 12242 177172 12248
rect 176752 11892 176804 11898
rect 176752 11834 176804 11840
rect 166632 11756 166684 11762
rect 166632 11698 166684 11704
rect 176660 11756 176712 11762
rect 176660 11698 176712 11704
rect 177132 11694 177160 12242
rect 177408 11898 177436 12582
rect 177396 11892 177448 11898
rect 177396 11834 177448 11840
rect 177120 11688 177172 11694
rect 177120 11630 177172 11636
rect 165896 11620 165948 11626
rect 165896 11562 165948 11568
rect 165908 11354 165936 11562
rect 165896 11348 165948 11354
rect 165896 11290 165948 11296
rect 165436 11280 165488 11286
rect 165436 11222 165488 11228
rect 177684 11218 177712 13194
rect 177776 12374 177804 13398
rect 177948 12912 178000 12918
rect 177948 12854 178000 12860
rect 177856 12640 177908 12646
rect 177856 12582 177908 12588
rect 177764 12368 177816 12374
rect 177764 12310 177816 12316
rect 177868 12238 177896 12582
rect 177856 12232 177908 12238
rect 177856 12174 177908 12180
rect 177868 11898 177896 12174
rect 177856 11892 177908 11898
rect 177856 11834 177908 11840
rect 177960 11218 177988 12854
rect 179524 12442 179552 15200
rect 181904 13796 181956 13802
rect 181904 13738 181956 13744
rect 180432 13456 180484 13462
rect 180432 13398 180484 13404
rect 179972 13252 180024 13258
rect 179972 13194 180024 13200
rect 179880 12640 179932 12646
rect 179880 12582 179932 12588
rect 179512 12436 179564 12442
rect 179512 12378 179564 12384
rect 179144 12232 179196 12238
rect 179144 12174 179196 12180
rect 178040 12096 178092 12102
rect 178040 12038 178092 12044
rect 165344 11212 165396 11218
rect 165344 11154 165396 11160
rect 177672 11212 177724 11218
rect 177672 11154 177724 11160
rect 177948 11212 178000 11218
rect 177948 11154 178000 11160
rect 178052 11150 178080 12038
rect 178040 11144 178092 11150
rect 178040 11086 178092 11092
rect 179156 10470 179184 12174
rect 179420 12164 179472 12170
rect 179420 12106 179472 12112
rect 179432 11082 179460 12106
rect 179892 11898 179920 12582
rect 179984 11898 180012 13194
rect 180156 12980 180208 12986
rect 180156 12922 180208 12928
rect 180248 12980 180300 12986
rect 180248 12922 180300 12928
rect 180168 12782 180196 12922
rect 180156 12776 180208 12782
rect 180156 12718 180208 12724
rect 180260 12714 180288 12922
rect 180340 12844 180392 12850
rect 180340 12786 180392 12792
rect 180248 12708 180300 12714
rect 180248 12650 180300 12656
rect 180156 12096 180208 12102
rect 180156 12038 180208 12044
rect 180168 11898 180196 12038
rect 179880 11892 179932 11898
rect 179880 11834 179932 11840
rect 179972 11892 180024 11898
rect 179972 11834 180024 11840
rect 180156 11892 180208 11898
rect 180156 11834 180208 11840
rect 179880 11756 179932 11762
rect 180064 11756 180116 11762
rect 179932 11716 180064 11744
rect 179880 11698 179932 11704
rect 180064 11698 180116 11704
rect 180352 11626 180380 12786
rect 180340 11620 180392 11626
rect 180340 11562 180392 11568
rect 180444 11150 180472 13398
rect 181916 13394 181944 13738
rect 182744 13530 182772 15286
rect 185674 15286 185808 15314
rect 185674 15200 185730 15286
rect 185780 13530 185808 15286
rect 188710 15200 188766 16000
rect 191746 15314 191802 16000
rect 191300 15286 191802 15314
rect 182732 13524 182784 13530
rect 182732 13466 182784 13472
rect 185768 13524 185820 13530
rect 185768 13466 185820 13472
rect 181904 13388 181956 13394
rect 181904 13330 181956 13336
rect 182088 13388 182140 13394
rect 182088 13330 182140 13336
rect 188528 13388 188580 13394
rect 188528 13330 188580 13336
rect 180616 13320 180668 13326
rect 180616 13262 180668 13268
rect 180524 12708 180576 12714
rect 180524 12650 180576 12656
rect 180536 11558 180564 12650
rect 180628 12646 180656 13262
rect 180892 13252 180944 13258
rect 180892 13194 180944 13200
rect 180708 13184 180760 13190
rect 180708 13126 180760 13132
rect 180616 12640 180668 12646
rect 180616 12582 180668 12588
rect 180720 12238 180748 13126
rect 180904 12374 180932 13194
rect 181536 12844 181588 12850
rect 181536 12786 181588 12792
rect 181444 12640 181496 12646
rect 181444 12582 181496 12588
rect 180892 12368 180944 12374
rect 180892 12310 180944 12316
rect 180708 12232 180760 12238
rect 180708 12174 180760 12180
rect 180616 11756 180668 11762
rect 180720 11744 180748 12174
rect 181456 12170 181484 12582
rect 181444 12164 181496 12170
rect 181444 12106 181496 12112
rect 180668 11716 180748 11744
rect 180616 11698 180668 11704
rect 181548 11694 181576 12786
rect 182100 12714 182128 13330
rect 187792 13184 187844 13190
rect 187792 13126 187844 13132
rect 187976 13184 188028 13190
rect 187976 13126 188028 13132
rect 188344 13184 188396 13190
rect 188344 13126 188396 13132
rect 182088 12708 182140 12714
rect 182088 12650 182140 12656
rect 187804 12646 187832 13126
rect 187792 12640 187844 12646
rect 187792 12582 187844 12588
rect 187988 12306 188016 13126
rect 188356 12986 188384 13126
rect 188344 12980 188396 12986
rect 188344 12922 188396 12928
rect 188540 12918 188568 13330
rect 188528 12912 188580 12918
rect 188528 12854 188580 12860
rect 188344 12844 188396 12850
rect 188344 12786 188396 12792
rect 187976 12300 188028 12306
rect 187976 12242 188028 12248
rect 188356 11898 188384 12786
rect 188620 12708 188672 12714
rect 188724 12696 188752 15200
rect 189908 13864 189960 13870
rect 189908 13806 189960 13812
rect 189356 13796 189408 13802
rect 189356 13738 189408 13744
rect 189368 13530 189396 13738
rect 189356 13524 189408 13530
rect 189356 13466 189408 13472
rect 188804 13456 188856 13462
rect 188804 13398 188856 13404
rect 188816 12850 188844 13398
rect 189368 12850 189396 13466
rect 189540 13456 189592 13462
rect 189592 13416 189672 13444
rect 189540 13398 189592 13404
rect 189540 13320 189592 13326
rect 189540 13262 189592 13268
rect 189552 13190 189580 13262
rect 189540 13184 189592 13190
rect 189540 13126 189592 13132
rect 188804 12844 188856 12850
rect 188804 12786 188856 12792
rect 189356 12844 189408 12850
rect 189356 12786 189408 12792
rect 189552 12782 189580 13126
rect 189540 12776 189592 12782
rect 189540 12718 189592 12724
rect 188672 12668 188752 12696
rect 189172 12708 189224 12714
rect 188620 12650 188672 12656
rect 189172 12650 189224 12656
rect 188988 12640 189040 12646
rect 188988 12582 189040 12588
rect 188344 11892 188396 11898
rect 188344 11834 188396 11840
rect 180800 11688 180852 11694
rect 180800 11630 180852 11636
rect 181536 11688 181588 11694
rect 181536 11630 181588 11636
rect 180524 11552 180576 11558
rect 180524 11494 180576 11500
rect 180812 11218 180840 11630
rect 180800 11212 180852 11218
rect 180800 11154 180852 11160
rect 189000 11150 189028 12582
rect 189184 12442 189212 12650
rect 189644 12442 189672 13416
rect 189920 13394 189948 13806
rect 190920 13524 190972 13530
rect 190920 13466 190972 13472
rect 189908 13388 189960 13394
rect 189908 13330 189960 13336
rect 190932 12918 190960 13466
rect 190920 12912 190972 12918
rect 190920 12854 190972 12860
rect 190552 12640 190604 12646
rect 190552 12582 190604 12588
rect 189172 12436 189224 12442
rect 189172 12378 189224 12384
rect 189632 12436 189684 12442
rect 189632 12378 189684 12384
rect 189540 12232 189592 12238
rect 189540 12174 189592 12180
rect 189552 11830 189580 12174
rect 189540 11824 189592 11830
rect 189540 11766 189592 11772
rect 189630 11792 189686 11801
rect 189630 11727 189632 11736
rect 189684 11727 189686 11736
rect 189632 11698 189684 11704
rect 189448 11552 189500 11558
rect 189448 11494 189500 11500
rect 180432 11144 180484 11150
rect 180432 11086 180484 11092
rect 188988 11144 189040 11150
rect 188988 11086 189040 11092
rect 189460 11082 189488 11494
rect 179420 11076 179472 11082
rect 179420 11018 179472 11024
rect 189448 11076 189500 11082
rect 189448 11018 189500 11024
rect 190564 10674 190592 12582
rect 190828 12436 190880 12442
rect 190828 12378 190880 12384
rect 190840 12170 190868 12378
rect 190828 12164 190880 12170
rect 190828 12106 190880 12112
rect 191104 12164 191156 12170
rect 191104 12106 191156 12112
rect 191196 12164 191248 12170
rect 191196 12106 191248 12112
rect 190828 11756 190880 11762
rect 190828 11698 190880 11704
rect 190840 11150 190868 11698
rect 190644 11144 190696 11150
rect 190644 11086 190696 11092
rect 190828 11144 190880 11150
rect 190828 11086 190880 11092
rect 190552 10668 190604 10674
rect 190552 10610 190604 10616
rect 187516 10600 187568 10606
rect 187516 10542 187568 10548
rect 179144 10464 179196 10470
rect 179144 10406 179196 10412
rect 163596 10124 163648 10130
rect 163596 10066 163648 10072
rect 156144 9648 156196 9654
rect 156144 9590 156196 9596
rect 158628 9648 158680 9654
rect 158628 9590 158680 9596
rect 153346 8732 153654 8741
rect 153346 8730 153352 8732
rect 153408 8730 153432 8732
rect 153488 8730 153512 8732
rect 153568 8730 153592 8732
rect 153648 8730 153654 8732
rect 153408 8678 153410 8730
rect 153590 8678 153592 8730
rect 153346 8676 153352 8678
rect 153408 8676 153432 8678
rect 153488 8676 153512 8678
rect 153568 8676 153592 8678
rect 153648 8676 153654 8678
rect 153346 8667 153654 8676
rect 187528 8362 187556 10542
rect 190656 9654 190684 11086
rect 191116 10810 191144 12106
rect 191208 11218 191236 12106
rect 191196 11212 191248 11218
rect 191196 11154 191248 11160
rect 191104 10804 191156 10810
rect 191104 10746 191156 10752
rect 191300 10266 191328 15286
rect 191746 15200 191802 15286
rect 194874 15314 194930 16000
rect 197910 15314 197966 16000
rect 201038 15314 201094 16000
rect 194874 15286 195284 15314
rect 194874 15200 194930 15286
rect 193220 13796 193272 13802
rect 193220 13738 193272 13744
rect 191445 13628 191753 13637
rect 191445 13626 191451 13628
rect 191507 13626 191531 13628
rect 191587 13626 191611 13628
rect 191667 13626 191691 13628
rect 191747 13626 191753 13628
rect 191507 13574 191509 13626
rect 191689 13574 191691 13626
rect 191445 13572 191451 13574
rect 191507 13572 191531 13574
rect 191587 13572 191611 13574
rect 191667 13572 191691 13574
rect 191747 13572 191753 13574
rect 191445 13563 191753 13572
rect 191840 13456 191892 13462
rect 191840 13398 191892 13404
rect 191380 13184 191432 13190
rect 191380 13126 191432 13132
rect 191392 12986 191420 13126
rect 191380 12980 191432 12986
rect 191380 12922 191432 12928
rect 191748 12912 191800 12918
rect 191748 12854 191800 12860
rect 191760 12714 191788 12854
rect 191748 12708 191800 12714
rect 191748 12650 191800 12656
rect 191852 12617 191880 13398
rect 192392 13252 192444 13258
rect 192392 13194 192444 13200
rect 191932 12708 191984 12714
rect 191932 12650 191984 12656
rect 192036 12702 192340 12730
rect 191838 12608 191894 12617
rect 191445 12540 191753 12549
rect 191838 12543 191894 12552
rect 191445 12538 191451 12540
rect 191507 12538 191531 12540
rect 191587 12538 191611 12540
rect 191667 12538 191691 12540
rect 191747 12538 191753 12540
rect 191507 12486 191509 12538
rect 191689 12486 191691 12538
rect 191445 12484 191451 12486
rect 191507 12484 191531 12486
rect 191587 12484 191611 12486
rect 191667 12484 191691 12486
rect 191747 12484 191753 12486
rect 191445 12475 191753 12484
rect 191944 12434 191972 12650
rect 192036 12646 192064 12702
rect 192024 12640 192076 12646
rect 192024 12582 192076 12588
rect 192116 12640 192168 12646
rect 192116 12582 192168 12588
rect 192206 12608 192262 12617
rect 192128 12434 192156 12582
rect 192206 12543 192262 12552
rect 191760 12406 191972 12434
rect 192036 12406 192156 12434
rect 191760 11898 191788 12406
rect 191840 12300 191892 12306
rect 191840 12242 191892 12248
rect 191852 11898 191880 12242
rect 191748 11892 191800 11898
rect 191748 11834 191800 11840
rect 191840 11892 191892 11898
rect 191840 11834 191892 11840
rect 191852 11762 191880 11834
rect 191840 11756 191892 11762
rect 191840 11698 191892 11704
rect 191445 11452 191753 11461
rect 191445 11450 191451 11452
rect 191507 11450 191531 11452
rect 191587 11450 191611 11452
rect 191667 11450 191691 11452
rect 191747 11450 191753 11452
rect 191507 11398 191509 11450
rect 191689 11398 191691 11450
rect 191445 11396 191451 11398
rect 191507 11396 191531 11398
rect 191587 11396 191611 11398
rect 191667 11396 191691 11398
rect 191747 11396 191753 11398
rect 191445 11387 191753 11396
rect 191852 11218 191880 11698
rect 192036 11234 192064 12406
rect 192116 11688 192168 11694
rect 192116 11630 192168 11636
rect 191840 11212 191892 11218
rect 191840 11154 191892 11160
rect 191944 11206 192064 11234
rect 191944 11150 191972 11206
rect 191932 11144 191984 11150
rect 191932 11086 191984 11092
rect 192128 10538 192156 11630
rect 192220 10742 192248 12543
rect 192208 10736 192260 10742
rect 192208 10678 192260 10684
rect 192312 10674 192340 12702
rect 192404 12434 192432 13194
rect 192484 12980 192536 12986
rect 192484 12922 192536 12928
rect 192496 12714 192524 12922
rect 192576 12844 192628 12850
rect 192576 12786 192628 12792
rect 192484 12708 192536 12714
rect 192484 12650 192536 12656
rect 192404 12406 192524 12434
rect 192300 10668 192352 10674
rect 192300 10610 192352 10616
rect 192116 10532 192168 10538
rect 192116 10474 192168 10480
rect 191445 10364 191753 10373
rect 191445 10362 191451 10364
rect 191507 10362 191531 10364
rect 191587 10362 191611 10364
rect 191667 10362 191691 10364
rect 191747 10362 191753 10364
rect 191507 10310 191509 10362
rect 191689 10310 191691 10362
rect 191445 10308 191451 10310
rect 191507 10308 191531 10310
rect 191587 10308 191611 10310
rect 191667 10308 191691 10310
rect 191747 10308 191753 10310
rect 191445 10299 191753 10308
rect 192496 10266 192524 12406
rect 192588 12374 192616 12786
rect 192668 12776 192720 12782
rect 192668 12718 192720 12724
rect 193036 12776 193088 12782
rect 193036 12718 193088 12724
rect 192576 12368 192628 12374
rect 192576 12310 192628 12316
rect 191288 10260 191340 10266
rect 191288 10202 191340 10208
rect 192484 10260 192536 10266
rect 192484 10202 192536 10208
rect 192588 10062 192616 12310
rect 192680 12306 192708 12718
rect 193048 12646 193076 12718
rect 193036 12640 193088 12646
rect 193036 12582 193088 12588
rect 193048 12345 193076 12582
rect 193034 12336 193090 12345
rect 192668 12300 192720 12306
rect 193034 12271 193090 12280
rect 192668 12242 192720 12248
rect 193036 12096 193088 12102
rect 193036 12038 193088 12044
rect 193048 11801 193076 12038
rect 193034 11792 193090 11801
rect 193034 11727 193090 11736
rect 193232 10742 193260 13738
rect 193496 13524 193548 13530
rect 193496 13466 193548 13472
rect 193404 13252 193456 13258
rect 193404 13194 193456 13200
rect 193416 12434 193444 13194
rect 193324 12406 193444 12434
rect 193324 11558 193352 12406
rect 193404 12164 193456 12170
rect 193404 12106 193456 12112
rect 193312 11552 193364 11558
rect 193312 11494 193364 11500
rect 193416 11370 193444 12106
rect 193508 12050 193536 13466
rect 193956 13252 194008 13258
rect 193956 13194 194008 13200
rect 194600 13252 194652 13258
rect 194600 13194 194652 13200
rect 194784 13252 194836 13258
rect 194784 13194 194836 13200
rect 193968 12986 193996 13194
rect 194612 13138 194640 13194
rect 194520 13110 194640 13138
rect 193956 12980 194008 12986
rect 193956 12922 194008 12928
rect 194416 12640 194468 12646
rect 194416 12582 194468 12588
rect 194048 12436 194100 12442
rect 194428 12434 194456 12582
rect 194100 12406 194456 12434
rect 194048 12378 194100 12384
rect 194416 12232 194468 12238
rect 194416 12174 194468 12180
rect 193680 12096 193732 12102
rect 193508 12044 193680 12050
rect 193508 12038 193732 12044
rect 193508 12022 193720 12038
rect 193508 11558 193536 12022
rect 194428 11898 194456 12174
rect 194416 11892 194468 11898
rect 194416 11834 194468 11840
rect 193864 11824 193916 11830
rect 193864 11766 193916 11772
rect 193496 11552 193548 11558
rect 193496 11494 193548 11500
rect 193416 11342 193536 11370
rect 193508 11218 193536 11342
rect 193496 11212 193548 11218
rect 193496 11154 193548 11160
rect 193312 11076 193364 11082
rect 193312 11018 193364 11024
rect 193220 10736 193272 10742
rect 193220 10678 193272 10684
rect 192576 10056 192628 10062
rect 192576 9998 192628 10004
rect 193324 9654 193352 11018
rect 193876 10810 193904 11766
rect 194324 11688 194376 11694
rect 194324 11630 194376 11636
rect 194416 11688 194468 11694
rect 194416 11630 194468 11636
rect 193864 10804 193916 10810
rect 193864 10746 193916 10752
rect 194140 10668 194192 10674
rect 194140 10610 194192 10616
rect 190644 9648 190696 9654
rect 190644 9590 190696 9596
rect 193312 9648 193364 9654
rect 193312 9590 193364 9596
rect 194152 9586 194180 10610
rect 194336 9926 194364 11630
rect 194428 11218 194456 11630
rect 194416 11212 194468 11218
rect 194416 11154 194468 11160
rect 194416 11008 194468 11014
rect 194416 10950 194468 10956
rect 194428 10062 194456 10950
rect 194416 10056 194468 10062
rect 194416 9998 194468 10004
rect 194324 9920 194376 9926
rect 194324 9862 194376 9868
rect 194140 9580 194192 9586
rect 194140 9522 194192 9528
rect 194520 9450 194548 13110
rect 194598 12880 194654 12889
rect 194598 12815 194654 12824
rect 194612 11218 194640 12815
rect 194796 12782 194824 13194
rect 194876 12980 194928 12986
rect 194876 12922 194928 12928
rect 194784 12776 194836 12782
rect 194784 12718 194836 12724
rect 194692 12164 194744 12170
rect 194692 12106 194744 12112
rect 194704 11898 194732 12106
rect 194692 11892 194744 11898
rect 194692 11834 194744 11840
rect 194600 11212 194652 11218
rect 194600 11154 194652 11160
rect 194888 11150 194916 12922
rect 195060 12844 195112 12850
rect 195060 12786 195112 12792
rect 195072 12753 195100 12786
rect 195058 12744 195114 12753
rect 195058 12679 195114 12688
rect 194968 12096 195020 12102
rect 194968 12038 195020 12044
rect 194876 11144 194928 11150
rect 194876 11086 194928 11092
rect 194980 10674 195008 12038
rect 195072 10742 195100 12679
rect 195256 11082 195284 15286
rect 197910 15286 198228 15314
rect 197910 15200 197966 15286
rect 195980 13796 196032 13802
rect 195980 13738 196032 13744
rect 195992 12986 196020 13738
rect 197636 13388 197688 13394
rect 197636 13330 197688 13336
rect 196440 13252 196492 13258
rect 196440 13194 196492 13200
rect 197360 13252 197412 13258
rect 197360 13194 197412 13200
rect 195980 12980 196032 12986
rect 195980 12922 196032 12928
rect 195794 12880 195850 12889
rect 195794 12815 195850 12824
rect 195808 12782 195836 12815
rect 195796 12776 195848 12782
rect 195796 12718 195848 12724
rect 195980 12640 196032 12646
rect 195980 12582 196032 12588
rect 195796 11552 195848 11558
rect 195796 11494 195848 11500
rect 195888 11552 195940 11558
rect 195888 11494 195940 11500
rect 195808 11150 195836 11494
rect 195796 11144 195848 11150
rect 195796 11086 195848 11092
rect 195244 11076 195296 11082
rect 195244 11018 195296 11024
rect 195060 10736 195112 10742
rect 195060 10678 195112 10684
rect 194968 10668 195020 10674
rect 194968 10610 195020 10616
rect 195900 10130 195928 11494
rect 195888 10124 195940 10130
rect 195888 10066 195940 10072
rect 195992 9518 196020 12582
rect 196452 11218 196480 13194
rect 197372 12889 197400 13194
rect 197358 12880 197414 12889
rect 197358 12815 197360 12824
rect 197412 12815 197414 12824
rect 197452 12844 197504 12850
rect 197360 12786 197412 12792
rect 197452 12786 197504 12792
rect 197464 12374 197492 12786
rect 197648 12782 197676 13330
rect 197728 13184 197780 13190
rect 197728 13126 197780 13132
rect 197912 13184 197964 13190
rect 197912 13126 197964 13132
rect 197740 12986 197768 13126
rect 197728 12980 197780 12986
rect 197728 12922 197780 12928
rect 197636 12776 197688 12782
rect 197636 12718 197688 12724
rect 197452 12368 197504 12374
rect 197452 12310 197504 12316
rect 197452 12232 197504 12238
rect 197452 12174 197504 12180
rect 196808 12096 196860 12102
rect 196808 12038 196860 12044
rect 196992 12096 197044 12102
rect 196992 12038 197044 12044
rect 197360 12096 197412 12102
rect 197360 12038 197412 12044
rect 196820 11830 196848 12038
rect 196808 11824 196860 11830
rect 196808 11766 196860 11772
rect 197004 11558 197032 12038
rect 197372 11694 197400 12038
rect 197360 11688 197412 11694
rect 197360 11630 197412 11636
rect 197464 11626 197492 12174
rect 197924 11762 197952 13126
rect 198200 12646 198228 15286
rect 201038 15286 201172 15314
rect 201038 15200 201094 15286
rect 200854 13288 200910 13297
rect 200854 13223 200910 13232
rect 200868 13190 200896 13223
rect 198556 13184 198608 13190
rect 198556 13126 198608 13132
rect 200488 13184 200540 13190
rect 200488 13126 200540 13132
rect 200856 13184 200908 13190
rect 200856 13126 200908 13132
rect 198372 12844 198424 12850
rect 198372 12786 198424 12792
rect 198188 12640 198240 12646
rect 198188 12582 198240 12588
rect 198384 12238 198412 12786
rect 198568 12782 198596 13126
rect 198556 12776 198608 12782
rect 198556 12718 198608 12724
rect 200396 12776 200448 12782
rect 200396 12718 200448 12724
rect 200408 12617 200436 12718
rect 200394 12608 200450 12617
rect 200394 12543 200450 12552
rect 200500 12306 200528 13126
rect 200672 12844 200724 12850
rect 200672 12786 200724 12792
rect 200684 12434 200712 12786
rect 201144 12646 201172 15286
rect 204074 15200 204130 16000
rect 207110 15314 207166 16000
rect 210238 15314 210294 16000
rect 213274 15314 213330 16000
rect 216310 15314 216366 16000
rect 207110 15286 207336 15314
rect 207110 15200 207166 15286
rect 201960 13456 202012 13462
rect 201960 13398 202012 13404
rect 203432 13456 203484 13462
rect 203432 13398 203484 13404
rect 201500 13320 201552 13326
rect 201500 13262 201552 13268
rect 201316 13184 201368 13190
rect 201316 13126 201368 13132
rect 201328 12850 201356 13126
rect 201316 12844 201368 12850
rect 201316 12786 201368 12792
rect 201132 12640 201184 12646
rect 201132 12582 201184 12588
rect 200592 12406 200712 12434
rect 200488 12300 200540 12306
rect 200488 12242 200540 12248
rect 200592 12238 200620 12406
rect 198372 12232 198424 12238
rect 198372 12174 198424 12180
rect 200580 12232 200632 12238
rect 200580 12174 200632 12180
rect 201040 12232 201092 12238
rect 201040 12174 201092 12180
rect 201052 11762 201080 12174
rect 197912 11756 197964 11762
rect 197912 11698 197964 11704
rect 201040 11756 201092 11762
rect 201040 11698 201092 11704
rect 197452 11620 197504 11626
rect 197452 11562 197504 11568
rect 196992 11552 197044 11558
rect 196992 11494 197044 11500
rect 201052 11218 201080 11698
rect 201328 11694 201356 12786
rect 201316 11688 201368 11694
rect 201316 11630 201368 11636
rect 201512 11558 201540 13262
rect 201972 12646 202000 13398
rect 202052 13388 202104 13394
rect 202052 13330 202104 13336
rect 201960 12640 202012 12646
rect 201960 12582 202012 12588
rect 202064 12306 202092 13330
rect 202144 13320 202196 13326
rect 203444 13297 203472 13398
rect 202144 13262 202196 13268
rect 203430 13288 203486 13297
rect 202156 12714 202184 13262
rect 202420 13252 202472 13258
rect 202420 13194 202472 13200
rect 203156 13252 203208 13258
rect 203430 13223 203486 13232
rect 203156 13194 203208 13200
rect 202144 12708 202196 12714
rect 202144 12650 202196 12656
rect 202432 12442 202460 13194
rect 202972 12912 203024 12918
rect 202972 12854 203024 12860
rect 202984 12782 203012 12854
rect 202880 12776 202932 12782
rect 202880 12718 202932 12724
rect 202972 12776 203024 12782
rect 202972 12718 203024 12724
rect 202420 12436 202472 12442
rect 202420 12378 202472 12384
rect 202052 12300 202104 12306
rect 202052 12242 202104 12248
rect 202892 11898 202920 12718
rect 203064 12096 203116 12102
rect 203064 12038 203116 12044
rect 202880 11892 202932 11898
rect 202880 11834 202932 11840
rect 203076 11762 203104 12038
rect 203168 11830 203196 13194
rect 203340 12912 203392 12918
rect 203340 12854 203392 12860
rect 203156 11824 203208 11830
rect 203156 11766 203208 11772
rect 203064 11756 203116 11762
rect 203064 11698 203116 11704
rect 202880 11688 202932 11694
rect 202880 11630 202932 11636
rect 201500 11552 201552 11558
rect 201500 11494 201552 11500
rect 196440 11212 196492 11218
rect 196440 11154 196492 11160
rect 201040 11212 201092 11218
rect 201040 11154 201092 11160
rect 201052 10606 201080 11154
rect 202696 11144 202748 11150
rect 202892 11098 202920 11630
rect 203352 11218 203380 12854
rect 203444 12102 203472 13223
rect 203524 12300 203576 12306
rect 203524 12242 203576 12248
rect 203432 12096 203484 12102
rect 203432 12038 203484 12044
rect 203444 11626 203472 12038
rect 203536 11694 203564 12242
rect 203524 11688 203576 11694
rect 203524 11630 203576 11636
rect 203432 11620 203484 11626
rect 203432 11562 203484 11568
rect 203340 11212 203392 11218
rect 203340 11154 203392 11160
rect 202748 11092 202920 11098
rect 202696 11086 202920 11092
rect 202708 11070 202920 11086
rect 201040 10600 201092 10606
rect 201040 10542 201092 10548
rect 203536 10470 203564 11630
rect 204088 11082 204116 15200
rect 207110 13560 207166 13569
rect 207110 13495 207112 13504
rect 207164 13495 207166 13504
rect 207112 13466 207164 13472
rect 206008 13456 206060 13462
rect 205652 13404 206008 13410
rect 205652 13398 206060 13404
rect 205652 13382 206048 13398
rect 205546 13288 205602 13297
rect 204260 13252 204312 13258
rect 204260 13194 204312 13200
rect 205456 13252 205508 13258
rect 205546 13223 205602 13232
rect 205456 13194 205508 13200
rect 204168 12776 204220 12782
rect 204168 12718 204220 12724
rect 204180 12434 204208 12718
rect 204272 12646 204300 13194
rect 205088 12776 205140 12782
rect 205088 12718 205140 12724
rect 205180 12776 205232 12782
rect 205180 12718 205232 12724
rect 204260 12640 204312 12646
rect 204260 12582 204312 12588
rect 204536 12640 204588 12646
rect 204536 12582 204588 12588
rect 204180 12406 204300 12434
rect 204272 12102 204300 12406
rect 204548 12238 204576 12582
rect 204536 12232 204588 12238
rect 204536 12174 204588 12180
rect 204260 12096 204312 12102
rect 204260 12038 204312 12044
rect 204548 11898 204576 12174
rect 204996 12164 205048 12170
rect 204996 12106 205048 12112
rect 204536 11892 204588 11898
rect 204536 11834 204588 11840
rect 204904 11620 204956 11626
rect 204904 11562 204956 11568
rect 204812 11552 204864 11558
rect 204812 11494 204864 11500
rect 204076 11076 204128 11082
rect 204076 11018 204128 11024
rect 204824 10674 204852 11494
rect 204916 11150 204944 11562
rect 205008 11218 205036 12106
rect 204996 11212 205048 11218
rect 204996 11154 205048 11160
rect 204904 11144 204956 11150
rect 204904 11086 204956 11092
rect 205100 10810 205128 12718
rect 205192 12646 205220 12718
rect 205180 12640 205232 12646
rect 205272 12640 205324 12646
rect 205180 12582 205232 12588
rect 205270 12608 205272 12617
rect 205324 12608 205326 12617
rect 205270 12543 205326 12552
rect 205468 11082 205496 13194
rect 205560 11830 205588 13223
rect 205652 13190 205680 13382
rect 207204 13320 207256 13326
rect 205730 13288 205786 13297
rect 207202 13288 207204 13297
rect 207256 13288 207258 13297
rect 205730 13223 205786 13232
rect 206376 13252 206428 13258
rect 205744 13190 205772 13223
rect 207202 13223 207258 13232
rect 206376 13194 206428 13200
rect 205640 13184 205692 13190
rect 205640 13126 205692 13132
rect 205732 13184 205784 13190
rect 205732 13126 205784 13132
rect 205640 12912 205692 12918
rect 205640 12854 205692 12860
rect 205652 12442 205680 12854
rect 205640 12436 205692 12442
rect 205640 12378 205692 12384
rect 205548 11824 205600 11830
rect 205548 11766 205600 11772
rect 206388 11762 206416 13194
rect 206560 12980 206612 12986
rect 206560 12922 206612 12928
rect 206572 11898 206600 12922
rect 207308 12714 207336 15286
rect 210238 15286 210372 15314
rect 210238 15200 210294 15286
rect 208030 13560 208086 13569
rect 210344 13530 210372 15286
rect 213274 15286 213408 15314
rect 213274 15200 213330 15286
rect 213380 13530 213408 15286
rect 216310 15286 216444 15314
rect 216310 15200 216366 15286
rect 208030 13495 208086 13504
rect 210332 13524 210384 13530
rect 208044 13462 208072 13495
rect 210332 13466 210384 13472
rect 213368 13524 213420 13530
rect 213368 13466 213420 13472
rect 216416 13462 216444 15286
rect 219438 15200 219494 16000
rect 222474 15314 222530 16000
rect 225602 15314 225658 16000
rect 228638 15314 228694 16000
rect 231674 15314 231730 16000
rect 234802 15314 234858 16000
rect 222474 15286 222792 15314
rect 222474 15200 222530 15286
rect 219452 13462 219480 15200
rect 207756 13456 207808 13462
rect 207756 13398 207808 13404
rect 208032 13456 208084 13462
rect 213276 13456 213328 13462
rect 208032 13398 208084 13404
rect 213274 13424 213276 13433
rect 216404 13456 216456 13462
rect 213328 13424 213330 13433
rect 207572 13252 207624 13258
rect 207624 13212 207704 13240
rect 207572 13194 207624 13200
rect 207388 13184 207440 13190
rect 207388 13126 207440 13132
rect 207400 12986 207428 13126
rect 207388 12980 207440 12986
rect 207388 12922 207440 12928
rect 207676 12850 207704 13212
rect 207664 12844 207716 12850
rect 207664 12786 207716 12792
rect 207296 12708 207348 12714
rect 207296 12650 207348 12656
rect 207676 12442 207704 12786
rect 207664 12436 207716 12442
rect 207768 12434 207796 13398
rect 216404 13398 216456 13404
rect 219440 13456 219492 13462
rect 219440 13398 219492 13404
rect 219806 13424 219862 13433
rect 213274 13359 213330 13368
rect 219806 13359 219862 13368
rect 207940 13320 207992 13326
rect 207938 13288 207940 13297
rect 213552 13320 213604 13326
rect 207992 13288 207994 13297
rect 213552 13262 213604 13268
rect 216588 13320 216640 13326
rect 216588 13262 216640 13268
rect 207938 13223 207994 13232
rect 213564 13190 213592 13262
rect 213552 13184 213604 13190
rect 213552 13126 213604 13132
rect 207848 12980 207900 12986
rect 207848 12922 207900 12928
rect 207860 12753 207888 12922
rect 210608 12912 210660 12918
rect 210608 12854 210660 12860
rect 207846 12744 207902 12753
rect 207846 12679 207902 12688
rect 210620 12646 210648 12854
rect 216600 12850 216628 13262
rect 219820 12986 219848 13359
rect 222764 13190 222792 15286
rect 225602 15286 225736 15314
rect 225602 15200 225658 15286
rect 224052 13518 224448 13546
rect 224052 13394 224080 13518
rect 224132 13456 224184 13462
rect 224132 13398 224184 13404
rect 224040 13388 224092 13394
rect 224040 13330 224092 13336
rect 224052 13190 224080 13330
rect 224144 13190 224172 13398
rect 224420 13394 224448 13518
rect 224408 13388 224460 13394
rect 224408 13330 224460 13336
rect 224236 13258 224448 13274
rect 224224 13252 224460 13258
rect 224276 13246 224408 13252
rect 224224 13194 224276 13200
rect 224408 13194 224460 13200
rect 225708 13190 225736 15286
rect 228638 15286 228864 15314
rect 228638 15200 228694 15286
rect 226444 13518 227208 13546
rect 226444 13462 226472 13518
rect 226432 13456 226484 13462
rect 226432 13398 226484 13404
rect 226616 13456 226668 13462
rect 226616 13398 226668 13404
rect 226892 13456 226944 13462
rect 226892 13398 226944 13404
rect 227074 13424 227130 13433
rect 222752 13184 222804 13190
rect 222752 13126 222804 13132
rect 223672 13184 223724 13190
rect 223672 13126 223724 13132
rect 224040 13184 224092 13190
rect 224040 13126 224092 13132
rect 224132 13184 224184 13190
rect 225420 13184 225472 13190
rect 224132 13126 224184 13132
rect 225418 13152 225420 13161
rect 225696 13184 225748 13190
rect 225472 13152 225474 13161
rect 219808 12980 219860 12986
rect 219808 12922 219860 12928
rect 223684 12850 223712 13126
rect 225696 13126 225748 13132
rect 225418 13087 225474 13096
rect 226628 12866 226656 13398
rect 226628 12850 226840 12866
rect 216588 12844 216640 12850
rect 216588 12786 216640 12792
rect 219808 12844 219860 12850
rect 219808 12786 219860 12792
rect 223672 12844 223724 12850
rect 226628 12844 226852 12850
rect 226628 12838 226800 12844
rect 223672 12786 223724 12792
rect 226800 12786 226852 12792
rect 219820 12714 219848 12786
rect 219808 12708 219860 12714
rect 219808 12650 219860 12656
rect 226904 12646 226932 13398
rect 227180 13394 227208 13518
rect 227904 13456 227956 13462
rect 227956 13404 228036 13410
rect 227904 13398 228036 13404
rect 227074 13359 227076 13368
rect 227128 13359 227130 13368
rect 227168 13388 227220 13394
rect 227076 13330 227128 13336
rect 227916 13382 228036 13398
rect 227168 13330 227220 13336
rect 227076 13184 227128 13190
rect 227074 13152 227076 13161
rect 227128 13152 227130 13161
rect 227180 13138 227208 13330
rect 227720 13320 227772 13326
rect 227720 13262 227772 13268
rect 228008 13274 228036 13382
rect 227628 13184 227680 13190
rect 227180 13110 227300 13138
rect 227628 13126 227680 13132
rect 227074 13087 227130 13096
rect 210608 12640 210660 12646
rect 210608 12582 210660 12588
rect 226892 12640 226944 12646
rect 226892 12582 226944 12588
rect 207768 12406 207888 12434
rect 207664 12378 207716 12384
rect 206560 11892 206612 11898
rect 206560 11834 206612 11840
rect 206376 11756 206428 11762
rect 206376 11698 206428 11704
rect 207860 11694 207888 12406
rect 227272 11694 227300 13110
rect 227640 12730 227668 13126
rect 227732 12866 227760 13262
rect 228008 13258 228128 13274
rect 228008 13252 228140 13258
rect 228008 13246 228088 13252
rect 228088 13194 228140 13200
rect 227904 13184 227956 13190
rect 227904 13126 227956 13132
rect 227732 12838 227852 12866
rect 227916 12850 227944 13126
rect 228272 12912 228324 12918
rect 228272 12854 228324 12860
rect 227640 12702 227760 12730
rect 227732 11830 227760 12702
rect 227824 11898 227852 12838
rect 227904 12844 227956 12850
rect 227904 12786 227956 12792
rect 228284 12782 228312 12854
rect 228272 12776 228324 12782
rect 228272 12718 228324 12724
rect 228836 12374 228864 15286
rect 231674 15286 231808 15314
rect 231674 15200 231730 15286
rect 231780 13682 231808 15286
rect 234802 15286 234936 15314
rect 234802 15200 234858 15286
rect 231780 13654 232084 13682
rect 229192 13456 229244 13462
rect 229190 13424 229192 13433
rect 229244 13424 229246 13433
rect 229190 13359 229246 13368
rect 231780 13394 231992 13410
rect 231780 13388 232004 13394
rect 231780 13382 231952 13388
rect 230388 13320 230440 13326
rect 230386 13288 230388 13297
rect 230440 13288 230442 13297
rect 230386 13223 230442 13232
rect 230756 13252 230808 13258
rect 230756 13194 230808 13200
rect 229544 13084 229852 13093
rect 229544 13082 229550 13084
rect 229606 13082 229630 13084
rect 229686 13082 229710 13084
rect 229766 13082 229790 13084
rect 229846 13082 229852 13084
rect 229606 13030 229608 13082
rect 229788 13030 229790 13082
rect 229544 13028 229550 13030
rect 229606 13028 229630 13030
rect 229686 13028 229710 13030
rect 229766 13028 229790 13030
rect 229846 13028 229852 13030
rect 229544 13019 229852 13028
rect 230388 12912 230440 12918
rect 230388 12854 230440 12860
rect 230296 12844 230348 12850
rect 230296 12786 230348 12792
rect 230204 12776 230256 12782
rect 230204 12718 230256 12724
rect 230216 12646 230244 12718
rect 229560 12640 229612 12646
rect 229560 12582 229612 12588
rect 230112 12640 230164 12646
rect 230112 12582 230164 12588
rect 230204 12640 230256 12646
rect 230204 12582 230256 12588
rect 228824 12368 228876 12374
rect 228824 12310 228876 12316
rect 228824 12096 228876 12102
rect 229572 12084 229600 12582
rect 230124 12442 230152 12582
rect 230112 12436 230164 12442
rect 230112 12378 230164 12384
rect 229928 12232 229980 12238
rect 229928 12174 229980 12180
rect 228824 12038 228876 12044
rect 229480 12056 229600 12084
rect 228836 11898 228864 12038
rect 227812 11892 227864 11898
rect 227812 11834 227864 11840
rect 228824 11892 228876 11898
rect 228824 11834 228876 11840
rect 227720 11824 227772 11830
rect 229480 11778 229508 12056
rect 229544 11996 229852 12005
rect 229544 11994 229550 11996
rect 229606 11994 229630 11996
rect 229686 11994 229710 11996
rect 229766 11994 229790 11996
rect 229846 11994 229852 11996
rect 229606 11942 229608 11994
rect 229788 11942 229790 11994
rect 229544 11940 229550 11942
rect 229606 11940 229630 11942
rect 229686 11940 229710 11942
rect 229766 11940 229790 11942
rect 229846 11940 229852 11942
rect 229544 11931 229852 11940
rect 229940 11898 229968 12174
rect 229928 11892 229980 11898
rect 229928 11834 229980 11840
rect 227720 11766 227772 11772
rect 229388 11762 229508 11778
rect 229376 11756 229508 11762
rect 229428 11750 229508 11756
rect 229376 11698 229428 11704
rect 207848 11688 207900 11694
rect 207848 11630 207900 11636
rect 227260 11688 227312 11694
rect 227260 11630 227312 11636
rect 230308 11626 230336 12786
rect 230400 11898 230428 12854
rect 230388 11892 230440 11898
rect 230388 11834 230440 11840
rect 230296 11620 230348 11626
rect 230296 11562 230348 11568
rect 229376 11552 229428 11558
rect 229376 11494 229428 11500
rect 229388 11150 229416 11494
rect 229376 11144 229428 11150
rect 229376 11086 229428 11092
rect 230768 11082 230796 13194
rect 231032 12912 231084 12918
rect 231032 12854 231084 12860
rect 230848 12164 230900 12170
rect 230848 12106 230900 12112
rect 230860 11830 230888 12106
rect 231044 11898 231072 12854
rect 231124 12368 231176 12374
rect 231124 12310 231176 12316
rect 231136 12170 231164 12310
rect 231676 12300 231728 12306
rect 231676 12242 231728 12248
rect 231308 12232 231360 12238
rect 231308 12174 231360 12180
rect 231124 12164 231176 12170
rect 231124 12106 231176 12112
rect 231216 12096 231268 12102
rect 231320 12084 231348 12174
rect 231400 12096 231452 12102
rect 231320 12056 231400 12084
rect 231216 12038 231268 12044
rect 231400 12038 231452 12044
rect 231032 11892 231084 11898
rect 231032 11834 231084 11840
rect 230848 11824 230900 11830
rect 230848 11766 230900 11772
rect 231228 11762 231256 12038
rect 231688 11898 231716 12242
rect 231780 12102 231808 13382
rect 231952 13330 232004 13336
rect 232056 13326 232084 13654
rect 233148 13388 233200 13394
rect 233148 13330 233200 13336
rect 233332 13388 233384 13394
rect 233332 13330 233384 13336
rect 231860 13320 231912 13326
rect 231860 13262 231912 13268
rect 232044 13320 232096 13326
rect 233056 13320 233108 13326
rect 232044 13262 232096 13268
rect 232134 13288 232190 13297
rect 231872 12442 231900 13262
rect 233056 13262 233108 13268
rect 232134 13223 232190 13232
rect 232148 13190 232176 13223
rect 232136 13184 232188 13190
rect 232136 13126 232188 13132
rect 232320 12912 232372 12918
rect 232320 12854 232372 12860
rect 232332 12646 232360 12854
rect 233068 12850 233096 13262
rect 233160 13172 233188 13330
rect 233240 13184 233292 13190
rect 233160 13144 233240 13172
rect 233240 13126 233292 13132
rect 233344 13002 233372 13330
rect 234908 13190 234936 15286
rect 237838 15200 237894 16000
rect 240874 15314 240930 16000
rect 244002 15314 244058 16000
rect 247038 15314 247094 16000
rect 250074 15314 250130 16000
rect 240874 15286 241284 15314
rect 240874 15200 240930 15286
rect 234896 13184 234948 13190
rect 234896 13126 234948 13132
rect 237012 13184 237064 13190
rect 237012 13126 237064 13132
rect 233160 12974 233372 13002
rect 233056 12844 233108 12850
rect 233056 12786 233108 12792
rect 232320 12640 232372 12646
rect 232320 12582 232372 12588
rect 232504 12640 232556 12646
rect 232504 12582 232556 12588
rect 231860 12436 231912 12442
rect 231860 12378 231912 12384
rect 232516 12374 232544 12582
rect 232504 12368 232556 12374
rect 232504 12310 232556 12316
rect 233068 12238 233096 12786
rect 233160 12646 233188 12974
rect 237024 12850 237052 13126
rect 237012 12844 237064 12850
rect 237012 12786 237064 12792
rect 237852 12714 237880 15200
rect 239496 13456 239548 13462
rect 238114 13424 238170 13433
rect 237932 13388 237984 13394
rect 238114 13359 238116 13368
rect 237932 13330 237984 13336
rect 238168 13359 238170 13368
rect 239494 13424 239496 13433
rect 239548 13424 239550 13433
rect 239494 13359 239550 13368
rect 238116 13330 238168 13336
rect 237944 12714 237972 13330
rect 238208 13320 238260 13326
rect 238208 13262 238260 13268
rect 238220 12986 238248 13262
rect 238484 13252 238536 13258
rect 238484 13194 238536 13200
rect 238208 12980 238260 12986
rect 238208 12922 238260 12928
rect 238300 12912 238352 12918
rect 238300 12854 238352 12860
rect 238312 12753 238340 12854
rect 238392 12844 238444 12850
rect 238392 12786 238444 12792
rect 238298 12744 238354 12753
rect 237840 12708 237892 12714
rect 237840 12650 237892 12656
rect 237932 12708 237984 12714
rect 238298 12679 238354 12688
rect 237932 12650 237984 12656
rect 233148 12640 233200 12646
rect 233148 12582 233200 12588
rect 238404 12238 238432 12786
rect 238496 12646 238524 13194
rect 239036 12912 239088 12918
rect 239036 12854 239088 12860
rect 238484 12640 238536 12646
rect 238484 12582 238536 12588
rect 238852 12640 238904 12646
rect 238852 12582 238904 12588
rect 238864 12306 238892 12582
rect 239048 12442 239076 12854
rect 239128 12640 239180 12646
rect 239128 12582 239180 12588
rect 239036 12436 239088 12442
rect 239036 12378 239088 12384
rect 238852 12300 238904 12306
rect 238852 12242 238904 12248
rect 239140 12238 239168 12582
rect 239312 12300 239364 12306
rect 239312 12242 239364 12248
rect 232136 12232 232188 12238
rect 232136 12174 232188 12180
rect 233056 12232 233108 12238
rect 233056 12174 233108 12180
rect 238024 12232 238076 12238
rect 238024 12174 238076 12180
rect 238392 12232 238444 12238
rect 238392 12174 238444 12180
rect 239128 12232 239180 12238
rect 239128 12174 239180 12180
rect 231768 12096 231820 12102
rect 231768 12038 231820 12044
rect 231676 11892 231728 11898
rect 231676 11834 231728 11840
rect 231216 11756 231268 11762
rect 231216 11698 231268 11704
rect 231688 11558 231716 11834
rect 232148 11626 232176 12174
rect 233068 12102 233096 12174
rect 233056 12096 233108 12102
rect 233056 12038 233108 12044
rect 232136 11620 232188 11626
rect 232136 11562 232188 11568
rect 231676 11552 231728 11558
rect 231676 11494 231728 11500
rect 238036 11218 238064 12174
rect 239324 11694 239352 12242
rect 239508 12238 239536 13359
rect 239772 13320 239824 13326
rect 239772 13262 239824 13268
rect 239496 12232 239548 12238
rect 239496 12174 239548 12180
rect 239312 11688 239364 11694
rect 239312 11630 239364 11636
rect 239404 11552 239456 11558
rect 239404 11494 239456 11500
rect 239416 11354 239444 11494
rect 239784 11354 239812 13262
rect 241060 13252 241112 13258
rect 241060 13194 241112 13200
rect 240048 12912 240100 12918
rect 240048 12854 240100 12860
rect 240968 12912 241020 12918
rect 240968 12854 241020 12860
rect 239956 12300 240008 12306
rect 239956 12242 240008 12248
rect 239968 11694 239996 12242
rect 239956 11688 240008 11694
rect 239956 11630 240008 11636
rect 240060 11354 240088 12854
rect 240324 12640 240376 12646
rect 240324 12582 240376 12588
rect 240140 12436 240192 12442
rect 240140 12378 240192 12384
rect 240152 11830 240180 12378
rect 240336 11898 240364 12582
rect 240876 12096 240928 12102
rect 240876 12038 240928 12044
rect 240324 11892 240376 11898
rect 240324 11834 240376 11840
rect 240140 11824 240192 11830
rect 240140 11766 240192 11772
rect 239404 11348 239456 11354
rect 239404 11290 239456 11296
rect 239772 11348 239824 11354
rect 239772 11290 239824 11296
rect 240048 11348 240100 11354
rect 240048 11290 240100 11296
rect 238024 11212 238076 11218
rect 238024 11154 238076 11160
rect 240888 11150 240916 12038
rect 240980 11354 241008 12854
rect 241072 11898 241100 13194
rect 241060 11892 241112 11898
rect 241060 11834 241112 11840
rect 241256 11558 241284 15286
rect 244002 15286 244228 15314
rect 244002 15200 244058 15286
rect 244096 13388 244148 13394
rect 244096 13330 244148 13336
rect 241796 13252 241848 13258
rect 241796 13194 241848 13200
rect 243636 13252 243688 13258
rect 243636 13194 243688 13200
rect 241520 12096 241572 12102
rect 241520 12038 241572 12044
rect 241532 11830 241560 12038
rect 241808 11898 241836 13194
rect 242532 13184 242584 13190
rect 242532 13126 242584 13132
rect 242072 12844 242124 12850
rect 242072 12786 242124 12792
rect 242256 12844 242308 12850
rect 242256 12786 242308 12792
rect 241796 11892 241848 11898
rect 241796 11834 241848 11840
rect 241520 11824 241572 11830
rect 241520 11766 241572 11772
rect 241980 11688 242032 11694
rect 241980 11630 242032 11636
rect 241244 11552 241296 11558
rect 241244 11494 241296 11500
rect 240968 11348 241020 11354
rect 240968 11290 241020 11296
rect 241992 11150 242020 11630
rect 242084 11354 242112 12786
rect 242162 12744 242218 12753
rect 242162 12679 242164 12688
rect 242216 12679 242218 12688
rect 242164 12650 242216 12656
rect 242268 12374 242296 12786
rect 242440 12640 242492 12646
rect 242440 12582 242492 12588
rect 242256 12368 242308 12374
rect 242256 12310 242308 12316
rect 242452 12306 242480 12582
rect 242440 12300 242492 12306
rect 242440 12242 242492 12248
rect 242164 12232 242216 12238
rect 242452 12186 242480 12242
rect 242216 12180 242480 12186
rect 242164 12174 242480 12180
rect 242176 12158 242480 12174
rect 242544 12102 242572 13126
rect 242900 12640 242952 12646
rect 242900 12582 242952 12588
rect 242912 12306 242940 12582
rect 243648 12442 243676 13194
rect 243636 12436 243688 12442
rect 243636 12378 243688 12384
rect 242992 12368 243044 12374
rect 243044 12316 243216 12322
rect 242992 12310 243216 12316
rect 243004 12306 243216 12310
rect 242900 12300 242952 12306
rect 243004 12300 243228 12306
rect 243004 12294 243176 12300
rect 242900 12242 242952 12248
rect 243176 12242 243228 12248
rect 244108 12102 244136 13330
rect 244200 12442 244228 15286
rect 247038 15286 247172 15314
rect 247038 15200 247094 15286
rect 247144 13462 247172 15286
rect 250074 15286 250208 15314
rect 250074 15200 250130 15286
rect 244648 13456 244700 13462
rect 244648 13398 244700 13404
rect 245384 13456 245436 13462
rect 245384 13398 245436 13404
rect 247132 13456 247184 13462
rect 247132 13398 247184 13404
rect 244660 13002 244688 13398
rect 244924 13252 244976 13258
rect 244924 13194 244976 13200
rect 244568 12974 244688 13002
rect 244568 12850 244596 12974
rect 244936 12918 244964 13194
rect 245396 12918 245424 13398
rect 244648 12912 244700 12918
rect 244648 12854 244700 12860
rect 244924 12912 244976 12918
rect 244924 12854 244976 12860
rect 245384 12912 245436 12918
rect 245384 12854 245436 12860
rect 244556 12844 244608 12850
rect 244556 12786 244608 12792
rect 244188 12436 244240 12442
rect 244188 12378 244240 12384
rect 242532 12096 242584 12102
rect 242532 12038 242584 12044
rect 244096 12096 244148 12102
rect 244096 12038 244148 12044
rect 242544 11762 242572 12038
rect 242532 11756 242584 11762
rect 242532 11698 242584 11704
rect 244568 11694 244596 12786
rect 244660 12714 244688 12854
rect 244832 12844 244884 12850
rect 244832 12786 244884 12792
rect 244648 12708 244700 12714
rect 244648 12650 244700 12656
rect 244844 11830 244872 12786
rect 250180 12714 250208 15286
rect 253202 15200 253258 16000
rect 256238 15200 256294 16000
rect 259366 15200 259422 16000
rect 262402 15314 262458 16000
rect 262402 15286 262536 15314
rect 262402 15200 262458 15286
rect 251008 13518 251496 13546
rect 251008 13394 251036 13518
rect 251088 13456 251140 13462
rect 251140 13404 251312 13410
rect 251088 13398 251312 13404
rect 250996 13388 251048 13394
rect 251100 13382 251312 13398
rect 250996 13330 251048 13336
rect 251088 13320 251140 13326
rect 251088 13262 251140 13268
rect 251100 12986 251128 13262
rect 251180 13184 251232 13190
rect 251180 13126 251232 13132
rect 251088 12980 251140 12986
rect 251088 12922 251140 12928
rect 251192 12850 251220 13126
rect 251180 12844 251232 12850
rect 251180 12786 251232 12792
rect 248328 12708 248380 12714
rect 248328 12650 248380 12656
rect 250168 12708 250220 12714
rect 250168 12650 250220 12656
rect 248340 12306 248368 12650
rect 248328 12300 248380 12306
rect 248328 12242 248380 12248
rect 249248 12300 249300 12306
rect 249248 12242 249300 12248
rect 249260 12170 249288 12242
rect 251284 12238 251312 13382
rect 251364 13252 251416 13258
rect 251364 13194 251416 13200
rect 251376 12442 251404 13194
rect 251364 12436 251416 12442
rect 251364 12378 251416 12384
rect 251468 12374 251496 13518
rect 252468 13456 252520 13462
rect 252468 13398 252520 13404
rect 252376 13252 252428 13258
rect 252376 13194 252428 13200
rect 251640 12912 251692 12918
rect 251640 12854 251692 12860
rect 251548 12844 251600 12850
rect 251548 12786 251600 12792
rect 251456 12368 251508 12374
rect 251456 12310 251508 12316
rect 251272 12232 251324 12238
rect 251272 12174 251324 12180
rect 249064 12164 249116 12170
rect 249064 12106 249116 12112
rect 249248 12164 249300 12170
rect 249248 12106 249300 12112
rect 244832 11824 244884 11830
rect 244832 11766 244884 11772
rect 242716 11688 242768 11694
rect 242716 11630 242768 11636
rect 244556 11688 244608 11694
rect 244556 11630 244608 11636
rect 242072 11348 242124 11354
rect 242072 11290 242124 11296
rect 242728 11218 242756 11630
rect 249076 11558 249104 12106
rect 249064 11552 249116 11558
rect 249064 11494 249116 11500
rect 242716 11212 242768 11218
rect 242716 11154 242768 11160
rect 240876 11144 240928 11150
rect 240876 11086 240928 11092
rect 241980 11144 242032 11150
rect 241980 11086 242032 11092
rect 205456 11076 205508 11082
rect 205456 11018 205508 11024
rect 230756 11076 230808 11082
rect 230756 11018 230808 11024
rect 229544 10908 229852 10917
rect 229544 10906 229550 10908
rect 229606 10906 229630 10908
rect 229686 10906 229710 10908
rect 229766 10906 229790 10908
rect 229846 10906 229852 10908
rect 229606 10854 229608 10906
rect 229788 10854 229790 10906
rect 229544 10852 229550 10854
rect 229606 10852 229630 10854
rect 229686 10852 229710 10854
rect 229766 10852 229790 10854
rect 229846 10852 229852 10854
rect 229544 10843 229852 10852
rect 205088 10804 205140 10810
rect 205088 10746 205140 10752
rect 204812 10668 204864 10674
rect 204812 10610 204864 10616
rect 203524 10464 203576 10470
rect 203524 10406 203576 10412
rect 229544 9820 229852 9829
rect 229544 9818 229550 9820
rect 229606 9818 229630 9820
rect 229686 9818 229710 9820
rect 229766 9818 229790 9820
rect 229846 9818 229852 9820
rect 229606 9766 229608 9818
rect 229788 9766 229790 9818
rect 229544 9764 229550 9766
rect 229606 9764 229630 9766
rect 229686 9764 229710 9766
rect 229766 9764 229790 9766
rect 229846 9764 229852 9766
rect 229544 9755 229852 9764
rect 195980 9512 196032 9518
rect 195980 9454 196032 9460
rect 194508 9444 194560 9450
rect 194508 9386 194560 9392
rect 191445 9276 191753 9285
rect 191445 9274 191451 9276
rect 191507 9274 191531 9276
rect 191587 9274 191611 9276
rect 191667 9274 191691 9276
rect 191747 9274 191753 9276
rect 191507 9222 191509 9274
rect 191689 9222 191691 9274
rect 191445 9220 191451 9222
rect 191507 9220 191531 9222
rect 191587 9220 191611 9222
rect 191667 9220 191691 9222
rect 191747 9220 191753 9222
rect 191445 9211 191753 9220
rect 229544 8732 229852 8741
rect 229544 8730 229550 8732
rect 229606 8730 229630 8732
rect 229686 8730 229710 8732
rect 229766 8730 229790 8732
rect 229846 8730 229852 8732
rect 229606 8678 229608 8730
rect 229788 8678 229790 8730
rect 229544 8676 229550 8678
rect 229606 8676 229630 8678
rect 229686 8676 229710 8678
rect 229766 8676 229790 8678
rect 229846 8676 229852 8678
rect 229544 8667 229852 8676
rect 187516 8356 187568 8362
rect 187516 8298 187568 8304
rect 191445 8188 191753 8197
rect 191445 8186 191451 8188
rect 191507 8186 191531 8188
rect 191587 8186 191611 8188
rect 191667 8186 191691 8188
rect 191747 8186 191753 8188
rect 191507 8134 191509 8186
rect 191689 8134 191691 8186
rect 191445 8132 191451 8134
rect 191507 8132 191531 8134
rect 191587 8132 191611 8134
rect 191667 8132 191691 8134
rect 191747 8132 191753 8134
rect 191445 8123 191753 8132
rect 153346 7644 153654 7653
rect 153346 7642 153352 7644
rect 153408 7642 153432 7644
rect 153488 7642 153512 7644
rect 153568 7642 153592 7644
rect 153648 7642 153654 7644
rect 153408 7590 153410 7642
rect 153590 7590 153592 7642
rect 153346 7588 153352 7590
rect 153408 7588 153432 7590
rect 153488 7588 153512 7590
rect 153568 7588 153592 7590
rect 153648 7588 153654 7590
rect 153346 7579 153654 7588
rect 229544 7644 229852 7653
rect 229544 7642 229550 7644
rect 229606 7642 229630 7644
rect 229686 7642 229710 7644
rect 229766 7642 229790 7644
rect 229846 7642 229852 7644
rect 229606 7590 229608 7642
rect 229788 7590 229790 7642
rect 229544 7588 229550 7590
rect 229606 7588 229630 7590
rect 229686 7588 229710 7590
rect 229766 7588 229790 7590
rect 229846 7588 229852 7590
rect 229544 7579 229852 7588
rect 191445 7100 191753 7109
rect 191445 7098 191451 7100
rect 191507 7098 191531 7100
rect 191587 7098 191611 7100
rect 191667 7098 191691 7100
rect 191747 7098 191753 7100
rect 191507 7046 191509 7098
rect 191689 7046 191691 7098
rect 191445 7044 191451 7046
rect 191507 7044 191531 7046
rect 191587 7044 191611 7046
rect 191667 7044 191691 7046
rect 191747 7044 191753 7046
rect 191445 7035 191753 7044
rect 153346 6556 153654 6565
rect 153346 6554 153352 6556
rect 153408 6554 153432 6556
rect 153488 6554 153512 6556
rect 153568 6554 153592 6556
rect 153648 6554 153654 6556
rect 153408 6502 153410 6554
rect 153590 6502 153592 6554
rect 153346 6500 153352 6502
rect 153408 6500 153432 6502
rect 153488 6500 153512 6502
rect 153568 6500 153592 6502
rect 153648 6500 153654 6502
rect 153346 6491 153654 6500
rect 229544 6556 229852 6565
rect 229544 6554 229550 6556
rect 229606 6554 229630 6556
rect 229686 6554 229710 6556
rect 229766 6554 229790 6556
rect 229846 6554 229852 6556
rect 229606 6502 229608 6554
rect 229788 6502 229790 6554
rect 229544 6500 229550 6502
rect 229606 6500 229630 6502
rect 229686 6500 229710 6502
rect 229766 6500 229790 6502
rect 229846 6500 229852 6502
rect 229544 6491 229852 6500
rect 249076 6254 249104 11494
rect 251560 11150 251588 12786
rect 251652 11626 251680 12854
rect 252100 12776 252152 12782
rect 252100 12718 252152 12724
rect 251824 12708 251876 12714
rect 251824 12650 251876 12656
rect 251836 12481 251864 12650
rect 251916 12640 251968 12646
rect 251914 12608 251916 12617
rect 252008 12640 252060 12646
rect 251968 12608 251970 12617
rect 252008 12582 252060 12588
rect 251914 12543 251970 12552
rect 251822 12472 251878 12481
rect 251822 12407 251878 12416
rect 251916 12436 251968 12442
rect 251916 12378 251968 12384
rect 251928 12238 251956 12378
rect 251916 12232 251968 12238
rect 251916 12174 251968 12180
rect 252020 11762 252048 12582
rect 252112 12374 252140 12718
rect 252388 12434 252416 13194
rect 252480 12918 252508 13398
rect 253020 13252 253072 13258
rect 253020 13194 253072 13200
rect 252468 12912 252520 12918
rect 252468 12854 252520 12860
rect 253032 12434 253060 13194
rect 252388 12406 252508 12434
rect 252100 12368 252152 12374
rect 252100 12310 252152 12316
rect 252008 11756 252060 11762
rect 252008 11698 252060 11704
rect 252112 11694 252140 12310
rect 252100 11688 252152 11694
rect 252100 11630 252152 11636
rect 251640 11620 251692 11626
rect 251640 11562 251692 11568
rect 252480 11354 252508 12406
rect 252940 12406 253060 12434
rect 252940 11898 252968 12406
rect 253112 12164 253164 12170
rect 253112 12106 253164 12112
rect 252928 11892 252980 11898
rect 252928 11834 252980 11840
rect 252744 11756 252796 11762
rect 252744 11698 252796 11704
rect 253020 11756 253072 11762
rect 253020 11698 253072 11704
rect 252468 11348 252520 11354
rect 252468 11290 252520 11296
rect 252756 11286 252784 11698
rect 252744 11280 252796 11286
rect 252744 11222 252796 11228
rect 251548 11144 251600 11150
rect 251548 11086 251600 11092
rect 252756 9994 252784 11222
rect 253032 11150 253060 11698
rect 253124 11354 253152 12106
rect 253112 11348 253164 11354
rect 253112 11290 253164 11296
rect 253216 11286 253244 15200
rect 254952 13456 255004 13462
rect 254688 13416 254952 13444
rect 253480 13184 253532 13190
rect 253480 13126 253532 13132
rect 253492 12764 253520 13126
rect 254688 12986 254716 13416
rect 254952 13398 255004 13404
rect 256252 13410 256280 15200
rect 259380 13682 259408 15200
rect 259380 13654 259500 13682
rect 259472 13462 259500 13654
rect 259460 13456 259512 13462
rect 256252 13382 256556 13410
rect 259460 13398 259512 13404
rect 256240 13320 256292 13326
rect 256240 13262 256292 13268
rect 254952 13252 255004 13258
rect 254952 13194 255004 13200
rect 255320 13252 255372 13258
rect 255320 13194 255372 13200
rect 254676 12980 254728 12986
rect 254676 12922 254728 12928
rect 253664 12776 253716 12782
rect 253492 12736 253664 12764
rect 253664 12718 253716 12724
rect 253940 12776 253992 12782
rect 253940 12718 253992 12724
rect 253952 12322 253980 12718
rect 254308 12368 254360 12374
rect 253952 12294 254072 12322
rect 254308 12310 254360 12316
rect 253296 11552 253348 11558
rect 253296 11494 253348 11500
rect 253204 11280 253256 11286
rect 253204 11222 253256 11228
rect 253308 11150 253336 11494
rect 254044 11354 254072 12294
rect 254320 11830 254348 12310
rect 254400 12096 254452 12102
rect 254400 12038 254452 12044
rect 254308 11824 254360 11830
rect 254308 11766 254360 11772
rect 254032 11348 254084 11354
rect 254032 11290 254084 11296
rect 254412 11150 254440 12038
rect 254688 11898 254716 12922
rect 254964 12434 254992 13194
rect 255332 13138 255360 13194
rect 255240 13110 255360 13138
rect 255136 12776 255188 12782
rect 255136 12718 255188 12724
rect 255044 12708 255096 12714
rect 255044 12650 255096 12656
rect 254780 12406 254992 12434
rect 254780 11898 254808 12406
rect 255056 12186 255084 12650
rect 255148 12238 255176 12718
rect 255240 12434 255268 13110
rect 256252 12986 256280 13262
rect 256332 13184 256384 13190
rect 256332 13126 256384 13132
rect 256240 12980 256292 12986
rect 256240 12922 256292 12928
rect 256344 12782 256372 13126
rect 256332 12776 256384 12782
rect 256332 12718 256384 12724
rect 256424 12776 256476 12782
rect 256424 12718 256476 12724
rect 255240 12406 255360 12434
rect 255228 12368 255280 12374
rect 255228 12310 255280 12316
rect 254964 12158 255084 12186
rect 255136 12232 255188 12238
rect 255136 12174 255188 12180
rect 254676 11892 254728 11898
rect 254676 11834 254728 11840
rect 254768 11892 254820 11898
rect 254768 11834 254820 11840
rect 254688 11150 254716 11834
rect 253020 11144 253072 11150
rect 253020 11086 253072 11092
rect 253296 11144 253348 11150
rect 253296 11086 253348 11092
rect 254400 11144 254452 11150
rect 254400 11086 254452 11092
rect 254676 11144 254728 11150
rect 254676 11086 254728 11092
rect 254964 10674 254992 12158
rect 255240 12102 255268 12310
rect 255044 12096 255096 12102
rect 255044 12038 255096 12044
rect 255228 12096 255280 12102
rect 255228 12038 255280 12044
rect 255056 11898 255084 12038
rect 255044 11892 255096 11898
rect 255044 11834 255096 11840
rect 255332 11676 255360 12406
rect 255596 12300 255648 12306
rect 255596 12242 255648 12248
rect 255608 11694 255636 12242
rect 256240 12232 256292 12238
rect 256240 12174 256292 12180
rect 256332 12232 256384 12238
rect 256332 12174 256384 12180
rect 256252 11762 256280 12174
rect 256344 12102 256372 12174
rect 256332 12096 256384 12102
rect 256332 12038 256384 12044
rect 256240 11756 256292 11762
rect 256240 11698 256292 11704
rect 256436 11694 256464 12718
rect 256528 12442 256556 13382
rect 256976 13252 257028 13258
rect 256976 13194 257028 13200
rect 261852 13252 261904 13258
rect 261852 13194 261904 13200
rect 256606 13016 256662 13025
rect 256606 12951 256662 12960
rect 256620 12850 256648 12951
rect 256608 12844 256660 12850
rect 256608 12786 256660 12792
rect 256516 12436 256568 12442
rect 256516 12378 256568 12384
rect 256988 12374 257016 13194
rect 257988 13184 258040 13190
rect 257988 13126 258040 13132
rect 258000 13025 258028 13126
rect 257986 13016 258042 13025
rect 257986 12951 258042 12960
rect 257252 12912 257304 12918
rect 257252 12854 257304 12860
rect 261760 12912 261812 12918
rect 261760 12854 261812 12860
rect 257160 12776 257212 12782
rect 257160 12718 257212 12724
rect 257068 12708 257120 12714
rect 257068 12650 257120 12656
rect 257080 12617 257108 12650
rect 257066 12608 257122 12617
rect 257066 12543 257122 12552
rect 257172 12481 257200 12718
rect 257158 12472 257214 12481
rect 257158 12407 257214 12416
rect 256976 12368 257028 12374
rect 256976 12310 257028 12316
rect 257264 11762 257292 12854
rect 257252 11756 257304 11762
rect 257252 11698 257304 11704
rect 255240 11648 255360 11676
rect 255596 11688 255648 11694
rect 255240 10810 255268 11648
rect 255596 11630 255648 11636
rect 256424 11688 256476 11694
rect 256424 11630 256476 11636
rect 261772 11558 261800 12854
rect 261864 12850 261892 13194
rect 261852 12844 261904 12850
rect 261852 12786 261904 12792
rect 261864 12306 261892 12786
rect 262312 12776 262364 12782
rect 262310 12744 262312 12753
rect 262364 12744 262366 12753
rect 262310 12679 262366 12688
rect 262220 12640 262272 12646
rect 262272 12600 262444 12628
rect 262220 12582 262272 12588
rect 262416 12306 262444 12600
rect 262508 12442 262536 15286
rect 265438 15200 265494 16000
rect 268566 15200 268622 16000
rect 271602 15314 271658 16000
rect 274638 15314 274694 16000
rect 277766 15314 277822 16000
rect 280802 15314 280858 16000
rect 283930 15314 283986 16000
rect 271602 15286 271828 15314
rect 271602 15200 271658 15286
rect 263508 13456 263560 13462
rect 263508 13398 263560 13404
rect 263414 13288 263470 13297
rect 263520 13258 263548 13398
rect 264152 13388 264204 13394
rect 264152 13330 264204 13336
rect 263414 13223 263416 13232
rect 263468 13223 263470 13232
rect 263508 13252 263560 13258
rect 263416 13194 263468 13200
rect 263508 13194 263560 13200
rect 262956 13184 263008 13190
rect 263324 13184 263376 13190
rect 263008 13144 263088 13172
rect 262956 13126 263008 13132
rect 262680 12708 262732 12714
rect 262680 12650 262732 12656
rect 262496 12436 262548 12442
rect 262496 12378 262548 12384
rect 261852 12300 261904 12306
rect 261852 12242 261904 12248
rect 262404 12300 262456 12306
rect 262404 12242 262456 12248
rect 262692 11558 262720 12650
rect 263060 12238 263088 13144
rect 263324 13126 263376 13132
rect 263336 12918 263364 13126
rect 263324 12912 263376 12918
rect 263324 12854 263376 12860
rect 263506 12744 263562 12753
rect 263506 12679 263508 12688
rect 263560 12679 263562 12688
rect 263508 12650 263560 12656
rect 263968 12640 264020 12646
rect 263968 12582 264020 12588
rect 263048 12232 263100 12238
rect 263048 12174 263100 12180
rect 263980 11694 264008 12582
rect 264164 12306 264192 13330
rect 264428 13252 264480 13258
rect 264428 13194 264480 13200
rect 264612 13252 264664 13258
rect 264612 13194 264664 13200
rect 264980 13252 265032 13258
rect 264980 13194 265032 13200
rect 264440 12850 264468 13194
rect 264624 12986 264652 13194
rect 264612 12980 264664 12986
rect 264612 12922 264664 12928
rect 264336 12844 264388 12850
rect 264336 12786 264388 12792
rect 264428 12844 264480 12850
rect 264428 12786 264480 12792
rect 264348 12753 264376 12786
rect 264334 12744 264390 12753
rect 264334 12679 264390 12688
rect 264992 12374 265020 13194
rect 264980 12368 265032 12374
rect 264980 12310 265032 12316
rect 264152 12300 264204 12306
rect 264152 12242 264204 12248
rect 265164 12300 265216 12306
rect 265164 12242 265216 12248
rect 264336 12232 264388 12238
rect 264336 12174 264388 12180
rect 264348 11762 264376 12174
rect 265176 12170 265204 12242
rect 265164 12164 265216 12170
rect 265164 12106 265216 12112
rect 265176 11914 265204 12106
rect 265176 11886 265296 11914
rect 265268 11762 265296 11886
rect 264336 11756 264388 11762
rect 264336 11698 264388 11704
rect 265164 11756 265216 11762
rect 265164 11698 265216 11704
rect 265256 11756 265308 11762
rect 265256 11698 265308 11704
rect 263968 11688 264020 11694
rect 263968 11630 264020 11636
rect 261760 11552 261812 11558
rect 261760 11494 261812 11500
rect 262680 11552 262732 11558
rect 262680 11494 262732 11500
rect 264348 11150 264376 11698
rect 265176 11286 265204 11698
rect 265452 11354 265480 15200
rect 267643 13628 267951 13637
rect 267643 13626 267649 13628
rect 267705 13626 267729 13628
rect 267785 13626 267809 13628
rect 267865 13626 267889 13628
rect 267945 13626 267951 13628
rect 267705 13574 267707 13626
rect 267887 13574 267889 13626
rect 267643 13572 267649 13574
rect 267705 13572 267729 13574
rect 267785 13572 267809 13574
rect 267865 13572 267889 13574
rect 267945 13572 267951 13574
rect 267643 13563 267951 13572
rect 265532 13456 265584 13462
rect 265532 13398 265584 13404
rect 265544 13297 265572 13398
rect 265530 13288 265586 13297
rect 265586 13246 265664 13274
rect 265530 13223 265586 13232
rect 265532 12912 265584 12918
rect 265532 12854 265584 12860
rect 265544 12442 265572 12854
rect 265532 12436 265584 12442
rect 265532 12378 265584 12384
rect 265636 12306 265664 13246
rect 266912 13252 266964 13258
rect 266912 13194 266964 13200
rect 266544 12912 266596 12918
rect 266544 12854 266596 12860
rect 265624 12300 265676 12306
rect 265624 12242 265676 12248
rect 265440 11348 265492 11354
rect 265440 11290 265492 11296
rect 265164 11280 265216 11286
rect 265164 11222 265216 11228
rect 265636 11150 265664 12242
rect 266268 11552 266320 11558
rect 266268 11494 266320 11500
rect 266360 11552 266412 11558
rect 266360 11494 266412 11500
rect 266280 11354 266308 11494
rect 266268 11348 266320 11354
rect 266268 11290 266320 11296
rect 264336 11144 264388 11150
rect 264336 11086 264388 11092
rect 264888 11144 264940 11150
rect 264888 11086 264940 11092
rect 265624 11144 265676 11150
rect 265624 11086 265676 11092
rect 255228 10804 255280 10810
rect 255228 10746 255280 10752
rect 264900 10742 264928 11086
rect 264888 10736 264940 10742
rect 264888 10678 264940 10684
rect 266372 10674 266400 11494
rect 266556 10810 266584 12854
rect 266820 12164 266872 12170
rect 266820 12106 266872 12112
rect 266832 11898 266860 12106
rect 266820 11892 266872 11898
rect 266820 11834 266872 11840
rect 266544 10804 266596 10810
rect 266544 10746 266596 10752
rect 254952 10668 255004 10674
rect 254952 10610 255004 10616
rect 266360 10668 266412 10674
rect 266360 10610 266412 10616
rect 266924 10266 266952 13194
rect 267648 13184 267700 13190
rect 267648 13126 267700 13132
rect 267004 12776 267056 12782
rect 267556 12776 267608 12782
rect 267004 12718 267056 12724
rect 267094 12744 267150 12753
rect 267016 12646 267044 12718
rect 267660 12753 267688 13126
rect 268384 12980 268436 12986
rect 268384 12922 268436 12928
rect 268292 12844 268344 12850
rect 268292 12786 268344 12792
rect 268016 12776 268068 12782
rect 267556 12718 267608 12724
rect 267646 12744 267702 12753
rect 267094 12679 267150 12688
rect 267108 12646 267136 12679
rect 267568 12646 267596 12718
rect 268016 12718 268068 12724
rect 268106 12744 268162 12753
rect 267646 12679 267702 12688
rect 267004 12640 267056 12646
rect 267004 12582 267056 12588
rect 267096 12640 267148 12646
rect 267096 12582 267148 12588
rect 267556 12640 267608 12646
rect 267556 12582 267608 12588
rect 267016 12102 267044 12582
rect 267643 12540 267951 12549
rect 267643 12538 267649 12540
rect 267705 12538 267729 12540
rect 267785 12538 267809 12540
rect 267865 12538 267889 12540
rect 267945 12538 267951 12540
rect 267705 12486 267707 12538
rect 267887 12486 267889 12538
rect 267643 12484 267649 12486
rect 267705 12484 267729 12486
rect 267785 12484 267809 12486
rect 267865 12484 267889 12486
rect 267945 12484 267951 12486
rect 267643 12475 267951 12484
rect 268028 12442 268056 12718
rect 268106 12679 268162 12688
rect 268016 12436 268068 12442
rect 268016 12378 268068 12384
rect 267280 12164 267332 12170
rect 267280 12106 267332 12112
rect 267004 12096 267056 12102
rect 267004 12038 267056 12044
rect 267292 11218 267320 12106
rect 268028 11626 268056 12378
rect 268120 12238 268148 12679
rect 268108 12232 268160 12238
rect 268108 12174 268160 12180
rect 268016 11620 268068 11626
rect 268016 11562 268068 11568
rect 267643 11452 267951 11461
rect 267643 11450 267649 11452
rect 267705 11450 267729 11452
rect 267785 11450 267809 11452
rect 267865 11450 267889 11452
rect 267945 11450 267951 11452
rect 267705 11398 267707 11450
rect 267887 11398 267889 11450
rect 267643 11396 267649 11398
rect 267705 11396 267729 11398
rect 267785 11396 267809 11398
rect 267865 11396 267889 11398
rect 267945 11396 267951 11398
rect 267643 11387 267951 11396
rect 268028 11218 268056 11562
rect 267280 11212 267332 11218
rect 267280 11154 267332 11160
rect 268016 11212 268068 11218
rect 268016 11154 268068 11160
rect 267643 10364 267951 10373
rect 267643 10362 267649 10364
rect 267705 10362 267729 10364
rect 267785 10362 267809 10364
rect 267865 10362 267889 10364
rect 267945 10362 267951 10364
rect 267705 10310 267707 10362
rect 267887 10310 267889 10362
rect 267643 10308 267649 10310
rect 267705 10308 267729 10310
rect 267785 10308 267809 10310
rect 267865 10308 267889 10310
rect 267945 10308 267951 10310
rect 267643 10299 267951 10308
rect 266912 10260 266964 10266
rect 266912 10202 266964 10208
rect 267740 10124 267792 10130
rect 267740 10066 267792 10072
rect 252744 9988 252796 9994
rect 252744 9930 252796 9936
rect 267752 9926 267780 10066
rect 268120 10062 268148 12174
rect 268200 12164 268252 12170
rect 268200 12106 268252 12112
rect 268212 10810 268240 12106
rect 268304 11830 268332 12786
rect 268396 12782 268424 12922
rect 268384 12776 268436 12782
rect 268384 12718 268436 12724
rect 268384 12436 268436 12442
rect 268384 12378 268436 12384
rect 268292 11824 268344 11830
rect 268292 11766 268344 11772
rect 268304 11082 268332 11766
rect 268292 11076 268344 11082
rect 268292 11018 268344 11024
rect 268200 10804 268252 10810
rect 268200 10746 268252 10752
rect 268396 10198 268424 12378
rect 268476 12096 268528 12102
rect 268476 12038 268528 12044
rect 268488 11762 268516 12038
rect 268476 11756 268528 11762
rect 268476 11698 268528 11704
rect 268488 11218 268516 11698
rect 268476 11212 268528 11218
rect 268476 11154 268528 11160
rect 268580 10266 268608 15200
rect 271800 13530 271828 15286
rect 274638 15286 274956 15314
rect 274638 15200 274694 15286
rect 274928 13530 274956 15286
rect 277766 15286 277900 15314
rect 277766 15200 277822 15286
rect 277872 13530 277900 15286
rect 280802 15286 280936 15314
rect 280802 15200 280858 15286
rect 280908 13530 280936 15286
rect 283930 15286 284248 15314
rect 283930 15200 283986 15286
rect 268936 13524 268988 13530
rect 268936 13466 268988 13472
rect 269580 13524 269632 13530
rect 269580 13466 269632 13472
rect 271788 13524 271840 13530
rect 271788 13466 271840 13472
rect 274916 13524 274968 13530
rect 274916 13466 274968 13472
rect 277860 13524 277912 13530
rect 277860 13466 277912 13472
rect 280896 13524 280948 13530
rect 284220 13512 284248 15286
rect 286966 15200 287022 16000
rect 290002 15314 290058 16000
rect 293130 15314 293186 16000
rect 296166 15314 296222 16000
rect 299202 15314 299258 16000
rect 302330 15314 302386 16000
rect 290002 15286 290136 15314
rect 290002 15200 290058 15286
rect 284300 13524 284352 13530
rect 284220 13484 284300 13512
rect 280896 13466 280948 13472
rect 286980 13512 287008 15200
rect 290108 13530 290136 15286
rect 293130 15286 293264 15314
rect 293130 15200 293186 15286
rect 293236 13530 293264 15286
rect 296166 15286 296300 15314
rect 296166 15200 296222 15286
rect 296272 13530 296300 15286
rect 299202 15286 299336 15314
rect 299202 15200 299258 15286
rect 299308 13530 299336 15286
rect 302330 15286 302648 15314
rect 302330 15200 302386 15286
rect 301412 13728 301464 13734
rect 301412 13670 301464 13676
rect 301424 13530 301452 13670
rect 287060 13524 287112 13530
rect 286980 13484 287060 13512
rect 284300 13466 284352 13472
rect 287060 13466 287112 13472
rect 290096 13524 290148 13530
rect 290096 13466 290148 13472
rect 293224 13524 293276 13530
rect 293224 13466 293276 13472
rect 296260 13524 296312 13530
rect 296260 13466 296312 13472
rect 299296 13524 299348 13530
rect 299296 13466 299348 13472
rect 301412 13524 301464 13530
rect 301412 13466 301464 13472
rect 268948 13433 268976 13466
rect 268934 13424 268990 13433
rect 268934 13359 268990 13368
rect 268948 13326 268976 13359
rect 268936 13320 268988 13326
rect 268936 13262 268988 13268
rect 269026 13288 269082 13297
rect 268752 13252 268804 13258
rect 268752 13194 268804 13200
rect 268660 12232 268712 12238
rect 268660 12174 268712 12180
rect 268672 12102 268700 12174
rect 268660 12096 268712 12102
rect 268660 12038 268712 12044
rect 268764 10538 268792 13194
rect 268948 11218 268976 13262
rect 269026 13223 269082 13232
rect 269040 12850 269068 13223
rect 269028 12844 269080 12850
rect 269028 12786 269080 12792
rect 269396 12776 269448 12782
rect 269316 12736 269396 12764
rect 269120 12640 269172 12646
rect 269172 12600 269252 12628
rect 269120 12582 269172 12588
rect 269120 12300 269172 12306
rect 269120 12242 269172 12248
rect 269132 11762 269160 12242
rect 269120 11756 269172 11762
rect 269120 11698 269172 11704
rect 268936 11212 268988 11218
rect 268936 11154 268988 11160
rect 268948 11082 268976 11154
rect 268936 11076 268988 11082
rect 268936 11018 268988 11024
rect 268844 11008 268896 11014
rect 268844 10950 268896 10956
rect 268752 10532 268804 10538
rect 268752 10474 268804 10480
rect 268568 10260 268620 10266
rect 268568 10202 268620 10208
rect 268384 10192 268436 10198
rect 268384 10134 268436 10140
rect 268856 10130 268884 10950
rect 269028 10668 269080 10674
rect 269028 10610 269080 10616
rect 268844 10124 268896 10130
rect 268844 10066 268896 10072
rect 269040 10062 269068 10610
rect 269224 10062 269252 12600
rect 269316 11354 269344 12736
rect 269396 12718 269448 12724
rect 269488 12164 269540 12170
rect 269488 12106 269540 12112
rect 269396 11688 269448 11694
rect 269396 11630 269448 11636
rect 269304 11348 269356 11354
rect 269304 11290 269356 11296
rect 269408 10810 269436 11630
rect 269396 10804 269448 10810
rect 269396 10746 269448 10752
rect 269500 10198 269528 12106
rect 269592 10470 269620 13466
rect 270408 13456 270460 13462
rect 272984 13456 273036 13462
rect 270408 13398 270460 13404
rect 272812 13404 272984 13410
rect 272812 13398 273036 13404
rect 273166 13424 273222 13433
rect 269672 12300 269724 12306
rect 269672 12242 269724 12248
rect 269684 11150 269712 12242
rect 270420 12186 270448 13398
rect 272812 13382 273024 13398
rect 270684 13252 270736 13258
rect 270684 13194 270736 13200
rect 270960 13252 271012 13258
rect 270960 13194 271012 13200
rect 270328 12158 270448 12186
rect 269856 11824 269908 11830
rect 269856 11766 269908 11772
rect 269672 11144 269724 11150
rect 269672 11086 269724 11092
rect 269580 10464 269632 10470
rect 269580 10406 269632 10412
rect 269488 10192 269540 10198
rect 269488 10134 269540 10140
rect 268108 10056 268160 10062
rect 268108 9998 268160 10004
rect 269028 10056 269080 10062
rect 269028 9998 269080 10004
rect 269212 10056 269264 10062
rect 269212 9998 269264 10004
rect 267740 9920 267792 9926
rect 267740 9862 267792 9868
rect 268120 9586 268148 9998
rect 269868 9654 269896 11766
rect 269948 11688 270000 11694
rect 269948 11630 270000 11636
rect 269960 11082 269988 11630
rect 269948 11076 270000 11082
rect 269948 11018 270000 11024
rect 270040 11008 270092 11014
rect 270040 10950 270092 10956
rect 270052 10742 270080 10950
rect 270040 10736 270092 10742
rect 270040 10678 270092 10684
rect 270328 10674 270356 12158
rect 270408 12096 270460 12102
rect 270408 12038 270460 12044
rect 270420 11150 270448 12038
rect 270696 11898 270724 13194
rect 270776 13184 270828 13190
rect 270776 13126 270828 13132
rect 270788 11898 270816 13126
rect 270868 12844 270920 12850
rect 270868 12786 270920 12792
rect 270880 12646 270908 12786
rect 270868 12640 270920 12646
rect 270868 12582 270920 12588
rect 270684 11892 270736 11898
rect 270684 11834 270736 11840
rect 270776 11892 270828 11898
rect 270776 11834 270828 11840
rect 270880 11150 270908 12582
rect 270408 11144 270460 11150
rect 270408 11086 270460 11092
rect 270868 11144 270920 11150
rect 270868 11086 270920 11092
rect 270316 10668 270368 10674
rect 270316 10610 270368 10616
rect 270972 9926 271000 13194
rect 271788 13184 271840 13190
rect 271788 13126 271840 13132
rect 271800 12918 271828 13126
rect 272812 12918 272840 13382
rect 273166 13359 273168 13368
rect 273220 13359 273222 13368
rect 273168 13330 273220 13336
rect 273260 13320 273312 13326
rect 273258 13288 273260 13297
rect 275100 13320 275152 13326
rect 273312 13288 273314 13297
rect 275100 13262 275152 13268
rect 281080 13320 281132 13326
rect 281080 13262 281132 13268
rect 284760 13320 284812 13326
rect 284760 13262 284812 13268
rect 290280 13320 290332 13326
rect 290280 13262 290332 13268
rect 299480 13320 299532 13326
rect 299480 13262 299532 13268
rect 273258 13223 273314 13232
rect 272892 13184 272944 13190
rect 272892 13126 272944 13132
rect 271052 12912 271104 12918
rect 271052 12854 271104 12860
rect 271788 12912 271840 12918
rect 271788 12854 271840 12860
rect 272800 12912 272852 12918
rect 272800 12854 272852 12860
rect 271064 12442 271092 12854
rect 272616 12844 272668 12850
rect 272616 12786 272668 12792
rect 272248 12776 272300 12782
rect 272248 12718 272300 12724
rect 271144 12640 271196 12646
rect 271144 12582 271196 12588
rect 271052 12436 271104 12442
rect 271052 12378 271104 12384
rect 271156 12306 271184 12582
rect 272260 12306 272288 12718
rect 272628 12646 272656 12786
rect 272904 12782 272932 13126
rect 273168 12912 273220 12918
rect 273168 12854 273220 12860
rect 273180 12782 273208 12854
rect 272892 12776 272944 12782
rect 272892 12718 272944 12724
rect 273168 12776 273220 12782
rect 273168 12718 273220 12724
rect 272800 12708 272852 12714
rect 272800 12650 272852 12656
rect 272524 12640 272576 12646
rect 272524 12582 272576 12588
rect 272616 12640 272668 12646
rect 272616 12582 272668 12588
rect 271144 12300 271196 12306
rect 271144 12242 271196 12248
rect 272248 12300 272300 12306
rect 272248 12242 272300 12248
rect 271328 12232 271380 12238
rect 271328 12174 271380 12180
rect 271340 11762 271368 12174
rect 271328 11756 271380 11762
rect 271328 11698 271380 11704
rect 272260 11218 272288 12242
rect 272248 11212 272300 11218
rect 272248 11154 272300 11160
rect 272536 10606 272564 12582
rect 272812 12306 272840 12650
rect 272800 12300 272852 12306
rect 272800 12242 272852 12248
rect 272904 12238 272932 12718
rect 272892 12232 272944 12238
rect 272892 12174 272944 12180
rect 273180 11694 273208 12718
rect 273168 11688 273220 11694
rect 273168 11630 273220 11636
rect 275112 11558 275140 13262
rect 281092 12646 281120 13262
rect 281080 12640 281132 12646
rect 281080 12582 281132 12588
rect 284772 12102 284800 13262
rect 290292 12850 290320 13262
rect 295892 13184 295944 13190
rect 295892 13126 295944 13132
rect 295904 12918 295932 13126
rect 295892 12912 295944 12918
rect 299492 12889 299520 13262
rect 302620 12986 302648 15286
rect 305366 15200 305422 16000
rect 303526 13968 303582 13977
rect 303526 13903 303582 13912
rect 302792 13796 302844 13802
rect 302792 13738 302844 13744
rect 302608 12980 302660 12986
rect 302608 12922 302660 12928
rect 295892 12854 295944 12860
rect 299478 12880 299534 12889
rect 290280 12844 290332 12850
rect 302804 12850 302832 13738
rect 303540 13326 303568 13903
rect 305000 13388 305052 13394
rect 305000 13330 305052 13336
rect 303528 13320 303580 13326
rect 303528 13262 303580 13268
rect 305012 12918 305040 13330
rect 305380 12986 305408 15200
rect 305368 12980 305420 12986
rect 305368 12922 305420 12928
rect 305000 12912 305052 12918
rect 305000 12854 305052 12860
rect 305460 12912 305512 12918
rect 305460 12854 305512 12860
rect 299478 12815 299534 12824
rect 302792 12844 302844 12850
rect 290280 12786 290332 12792
rect 302792 12786 302844 12792
rect 305472 12442 305500 12854
rect 305460 12436 305512 12442
rect 305460 12378 305512 12384
rect 284760 12096 284812 12102
rect 284760 12038 284812 12044
rect 275100 11552 275152 11558
rect 275100 11494 275152 11500
rect 272524 10600 272576 10606
rect 272524 10542 272576 10548
rect 304448 10056 304500 10062
rect 304446 10024 304448 10033
rect 304500 10024 304502 10033
rect 304446 9959 304502 9968
rect 270960 9920 271012 9926
rect 270960 9862 271012 9868
rect 269856 9648 269908 9654
rect 269856 9590 269908 9596
rect 268108 9580 268160 9586
rect 268108 9522 268160 9528
rect 267643 9276 267951 9285
rect 267643 9274 267649 9276
rect 267705 9274 267729 9276
rect 267785 9274 267809 9276
rect 267865 9274 267889 9276
rect 267945 9274 267951 9276
rect 267705 9222 267707 9274
rect 267887 9222 267889 9274
rect 267643 9220 267649 9222
rect 267705 9220 267729 9222
rect 267785 9220 267809 9222
rect 267865 9220 267889 9222
rect 267945 9220 267951 9222
rect 267643 9211 267951 9220
rect 267643 8188 267951 8197
rect 267643 8186 267649 8188
rect 267705 8186 267729 8188
rect 267785 8186 267809 8188
rect 267865 8186 267889 8188
rect 267945 8186 267951 8188
rect 267705 8134 267707 8186
rect 267887 8134 267889 8186
rect 267643 8132 267649 8134
rect 267705 8132 267729 8134
rect 267785 8132 267809 8134
rect 267865 8132 267889 8134
rect 267945 8132 267951 8134
rect 267643 8123 267951 8132
rect 267643 7100 267951 7109
rect 267643 7098 267649 7100
rect 267705 7098 267729 7100
rect 267785 7098 267809 7100
rect 267865 7098 267889 7100
rect 267945 7098 267951 7100
rect 267705 7046 267707 7098
rect 267887 7046 267889 7098
rect 267643 7044 267649 7046
rect 267705 7044 267729 7046
rect 267785 7044 267809 7046
rect 267865 7044 267889 7046
rect 267945 7044 267951 7046
rect 267643 7035 267951 7044
rect 303988 6316 304040 6322
rect 303988 6258 304040 6264
rect 249064 6248 249116 6254
rect 249064 6190 249116 6196
rect 191445 6012 191753 6021
rect 191445 6010 191451 6012
rect 191507 6010 191531 6012
rect 191587 6010 191611 6012
rect 191667 6010 191691 6012
rect 191747 6010 191753 6012
rect 191507 5958 191509 6010
rect 191689 5958 191691 6010
rect 191445 5956 191451 5958
rect 191507 5956 191531 5958
rect 191587 5956 191611 5958
rect 191667 5956 191691 5958
rect 191747 5956 191753 5958
rect 191445 5947 191753 5956
rect 267643 6012 267951 6021
rect 267643 6010 267649 6012
rect 267705 6010 267729 6012
rect 267785 6010 267809 6012
rect 267865 6010 267889 6012
rect 267945 6010 267951 6012
rect 267705 5958 267707 6010
rect 267887 5958 267889 6010
rect 267643 5956 267649 5958
rect 267705 5956 267729 5958
rect 267785 5956 267809 5958
rect 267865 5956 267889 5958
rect 267945 5956 267951 5958
rect 267643 5947 267951 5956
rect 304000 5953 304028 6258
rect 303986 5944 304042 5953
rect 303986 5879 304042 5888
rect 153346 5468 153654 5477
rect 153346 5466 153352 5468
rect 153408 5466 153432 5468
rect 153488 5466 153512 5468
rect 153568 5466 153592 5468
rect 153648 5466 153654 5468
rect 153408 5414 153410 5466
rect 153590 5414 153592 5466
rect 153346 5412 153352 5414
rect 153408 5412 153432 5414
rect 153488 5412 153512 5414
rect 153568 5412 153592 5414
rect 153648 5412 153654 5414
rect 153346 5403 153654 5412
rect 229544 5468 229852 5477
rect 229544 5466 229550 5468
rect 229606 5466 229630 5468
rect 229686 5466 229710 5468
rect 229766 5466 229790 5468
rect 229846 5466 229852 5468
rect 229606 5414 229608 5466
rect 229788 5414 229790 5466
rect 229544 5412 229550 5414
rect 229606 5412 229630 5414
rect 229686 5412 229710 5414
rect 229766 5412 229790 5414
rect 229846 5412 229852 5414
rect 229544 5403 229852 5412
rect 191445 4924 191753 4933
rect 191445 4922 191451 4924
rect 191507 4922 191531 4924
rect 191587 4922 191611 4924
rect 191667 4922 191691 4924
rect 191747 4922 191753 4924
rect 191507 4870 191509 4922
rect 191689 4870 191691 4922
rect 191445 4868 191451 4870
rect 191507 4868 191531 4870
rect 191587 4868 191611 4870
rect 191667 4868 191691 4870
rect 191747 4868 191753 4870
rect 191445 4859 191753 4868
rect 267643 4924 267951 4933
rect 267643 4922 267649 4924
rect 267705 4922 267729 4924
rect 267785 4922 267809 4924
rect 267865 4922 267889 4924
rect 267945 4922 267951 4924
rect 267705 4870 267707 4922
rect 267887 4870 267889 4922
rect 267643 4868 267649 4870
rect 267705 4868 267729 4870
rect 267785 4868 267809 4870
rect 267865 4868 267889 4870
rect 267945 4868 267951 4870
rect 267643 4859 267951 4868
rect 153346 4380 153654 4389
rect 153346 4378 153352 4380
rect 153408 4378 153432 4380
rect 153488 4378 153512 4380
rect 153568 4378 153592 4380
rect 153648 4378 153654 4380
rect 153408 4326 153410 4378
rect 153590 4326 153592 4378
rect 153346 4324 153352 4326
rect 153408 4324 153432 4326
rect 153488 4324 153512 4326
rect 153568 4324 153592 4326
rect 153648 4324 153654 4326
rect 153346 4315 153654 4324
rect 229544 4380 229852 4389
rect 229544 4378 229550 4380
rect 229606 4378 229630 4380
rect 229686 4378 229710 4380
rect 229766 4378 229790 4380
rect 229846 4378 229852 4380
rect 229606 4326 229608 4378
rect 229788 4326 229790 4378
rect 229544 4324 229550 4326
rect 229606 4324 229630 4326
rect 229686 4324 229710 4326
rect 229766 4324 229790 4326
rect 229846 4324 229852 4326
rect 229544 4315 229852 4324
rect 191445 3836 191753 3845
rect 191445 3834 191451 3836
rect 191507 3834 191531 3836
rect 191587 3834 191611 3836
rect 191667 3834 191691 3836
rect 191747 3834 191753 3836
rect 191507 3782 191509 3834
rect 191689 3782 191691 3834
rect 191445 3780 191451 3782
rect 191507 3780 191531 3782
rect 191587 3780 191611 3782
rect 191667 3780 191691 3782
rect 191747 3780 191753 3782
rect 191445 3771 191753 3780
rect 267643 3836 267951 3845
rect 267643 3834 267649 3836
rect 267705 3834 267729 3836
rect 267785 3834 267809 3836
rect 267865 3834 267889 3836
rect 267945 3834 267951 3836
rect 267705 3782 267707 3834
rect 267887 3782 267889 3834
rect 267643 3780 267649 3782
rect 267705 3780 267729 3782
rect 267785 3780 267809 3782
rect 267865 3780 267889 3782
rect 267945 3780 267951 3782
rect 267643 3771 267951 3780
rect 153346 3292 153654 3301
rect 153346 3290 153352 3292
rect 153408 3290 153432 3292
rect 153488 3290 153512 3292
rect 153568 3290 153592 3292
rect 153648 3290 153654 3292
rect 153408 3238 153410 3290
rect 153590 3238 153592 3290
rect 153346 3236 153352 3238
rect 153408 3236 153432 3238
rect 153488 3236 153512 3238
rect 153568 3236 153592 3238
rect 153648 3236 153654 3238
rect 153346 3227 153654 3236
rect 229544 3292 229852 3301
rect 229544 3290 229550 3292
rect 229606 3290 229630 3292
rect 229686 3290 229710 3292
rect 229766 3290 229790 3292
rect 229846 3290 229852 3292
rect 229606 3238 229608 3290
rect 229788 3238 229790 3290
rect 229544 3236 229550 3238
rect 229606 3236 229630 3238
rect 229686 3236 229710 3238
rect 229766 3236 229790 3238
rect 229846 3236 229852 3238
rect 229544 3227 229852 3236
rect 191445 2748 191753 2757
rect 191445 2746 191451 2748
rect 191507 2746 191531 2748
rect 191587 2746 191611 2748
rect 191667 2746 191691 2748
rect 191747 2746 191753 2748
rect 191507 2694 191509 2746
rect 191689 2694 191691 2746
rect 191445 2692 191451 2694
rect 191507 2692 191531 2694
rect 191587 2692 191611 2694
rect 191667 2692 191691 2694
rect 191747 2692 191753 2694
rect 191445 2683 191753 2692
rect 267643 2748 267951 2757
rect 267643 2746 267649 2748
rect 267705 2746 267729 2748
rect 267785 2746 267809 2748
rect 267865 2746 267889 2748
rect 267945 2746 267951 2748
rect 267705 2694 267707 2746
rect 267887 2694 267889 2746
rect 267643 2692 267649 2694
rect 267705 2692 267729 2694
rect 267785 2692 267809 2694
rect 267865 2692 267889 2694
rect 267945 2692 267951 2694
rect 267643 2683 267951 2692
rect 149428 2644 149480 2650
rect 149428 2586 149480 2592
rect 302240 2644 302292 2650
rect 302240 2586 302292 2592
rect 77148 2204 77456 2213
rect 77148 2202 77154 2204
rect 77210 2202 77234 2204
rect 77290 2202 77314 2204
rect 77370 2202 77394 2204
rect 77450 2202 77456 2204
rect 77210 2150 77212 2202
rect 77392 2150 77394 2202
rect 77148 2148 77154 2150
rect 77210 2148 77234 2150
rect 77290 2148 77314 2150
rect 77370 2148 77394 2150
rect 77450 2148 77456 2150
rect 77148 2139 77456 2148
rect 153346 2204 153654 2213
rect 153346 2202 153352 2204
rect 153408 2202 153432 2204
rect 153488 2202 153512 2204
rect 153568 2202 153592 2204
rect 153648 2202 153654 2204
rect 153408 2150 153410 2202
rect 153590 2150 153592 2202
rect 153346 2148 153352 2150
rect 153408 2148 153432 2150
rect 153488 2148 153512 2150
rect 153568 2148 153592 2150
rect 153648 2148 153654 2150
rect 153346 2139 153654 2148
rect 229544 2204 229852 2213
rect 229544 2202 229550 2204
rect 229606 2202 229630 2204
rect 229686 2202 229710 2204
rect 229766 2202 229790 2204
rect 229846 2202 229852 2204
rect 229606 2150 229608 2202
rect 229788 2150 229790 2202
rect 229544 2148 229550 2150
rect 229606 2148 229630 2150
rect 229686 2148 229710 2150
rect 229766 2148 229790 2150
rect 229846 2148 229852 2150
rect 229544 2139 229852 2148
rect 302252 2009 302280 2586
rect 302238 2000 302294 2009
rect 302238 1935 302294 1944
<< via2 >>
rect 29366 12180 29368 12200
rect 29368 12180 29420 12200
rect 29420 12180 29422 12200
rect 29366 12144 29422 12180
rect 30746 12144 30802 12200
rect 31390 12144 31446 12200
rect 39055 13626 39111 13628
rect 39135 13626 39191 13628
rect 39215 13626 39271 13628
rect 39295 13626 39351 13628
rect 39055 13574 39101 13626
rect 39101 13574 39111 13626
rect 39135 13574 39165 13626
rect 39165 13574 39177 13626
rect 39177 13574 39191 13626
rect 39215 13574 39229 13626
rect 39229 13574 39241 13626
rect 39241 13574 39271 13626
rect 39295 13574 39305 13626
rect 39305 13574 39351 13626
rect 39055 13572 39111 13574
rect 39135 13572 39191 13574
rect 39215 13572 39271 13574
rect 39295 13572 39351 13574
rect 39055 12538 39111 12540
rect 39135 12538 39191 12540
rect 39215 12538 39271 12540
rect 39295 12538 39351 12540
rect 39055 12486 39101 12538
rect 39101 12486 39111 12538
rect 39135 12486 39165 12538
rect 39165 12486 39177 12538
rect 39177 12486 39191 12538
rect 39215 12486 39229 12538
rect 39229 12486 39241 12538
rect 39241 12486 39271 12538
rect 39295 12486 39305 12538
rect 39305 12486 39351 12538
rect 39055 12484 39111 12486
rect 39135 12484 39191 12486
rect 39215 12484 39271 12486
rect 39295 12484 39351 12486
rect 39055 11450 39111 11452
rect 39135 11450 39191 11452
rect 39215 11450 39271 11452
rect 39295 11450 39351 11452
rect 39055 11398 39101 11450
rect 39101 11398 39111 11450
rect 39135 11398 39165 11450
rect 39165 11398 39177 11450
rect 39177 11398 39191 11450
rect 39215 11398 39229 11450
rect 39229 11398 39241 11450
rect 39241 11398 39271 11450
rect 39295 11398 39305 11450
rect 39305 11398 39351 11450
rect 39055 11396 39111 11398
rect 39135 11396 39191 11398
rect 39215 11396 39271 11398
rect 39295 11396 39351 11398
rect 40590 12180 40592 12200
rect 40592 12180 40644 12200
rect 40644 12180 40646 12200
rect 40590 12144 40646 12180
rect 42430 12144 42486 12200
rect 77154 13082 77210 13084
rect 77234 13082 77290 13084
rect 77314 13082 77370 13084
rect 77394 13082 77450 13084
rect 77154 13030 77200 13082
rect 77200 13030 77210 13082
rect 77234 13030 77264 13082
rect 77264 13030 77276 13082
rect 77276 13030 77290 13082
rect 77314 13030 77328 13082
rect 77328 13030 77340 13082
rect 77340 13030 77370 13082
rect 77394 13030 77404 13082
rect 77404 13030 77450 13082
rect 77154 13028 77210 13030
rect 77234 13028 77290 13030
rect 77314 13028 77370 13030
rect 77394 13028 77450 13030
rect 77154 11994 77210 11996
rect 77234 11994 77290 11996
rect 77314 11994 77370 11996
rect 77394 11994 77450 11996
rect 77154 11942 77200 11994
rect 77200 11942 77210 11994
rect 77234 11942 77264 11994
rect 77264 11942 77276 11994
rect 77276 11942 77290 11994
rect 77314 11942 77328 11994
rect 77328 11942 77340 11994
rect 77340 11942 77370 11994
rect 77394 11942 77404 11994
rect 77404 11942 77450 11994
rect 77154 11940 77210 11942
rect 77234 11940 77290 11942
rect 77314 11940 77370 11942
rect 77394 11940 77450 11942
rect 86958 13096 87014 13152
rect 87786 12688 87842 12744
rect 88154 12300 88210 12336
rect 88154 12280 88156 12300
rect 88156 12280 88208 12300
rect 88208 12280 88210 12300
rect 91834 13096 91890 13152
rect 89902 12280 89958 12336
rect 90730 12688 90786 12744
rect 77154 10906 77210 10908
rect 77234 10906 77290 10908
rect 77314 10906 77370 10908
rect 77394 10906 77450 10908
rect 77154 10854 77200 10906
rect 77200 10854 77210 10906
rect 77234 10854 77264 10906
rect 77264 10854 77276 10906
rect 77276 10854 77290 10906
rect 77314 10854 77328 10906
rect 77328 10854 77340 10906
rect 77340 10854 77370 10906
rect 77394 10854 77404 10906
rect 77404 10854 77450 10906
rect 77154 10852 77210 10854
rect 77234 10852 77290 10854
rect 77314 10852 77370 10854
rect 77394 10852 77450 10854
rect 39055 10362 39111 10364
rect 39135 10362 39191 10364
rect 39215 10362 39271 10364
rect 39295 10362 39351 10364
rect 39055 10310 39101 10362
rect 39101 10310 39111 10362
rect 39135 10310 39165 10362
rect 39165 10310 39177 10362
rect 39177 10310 39191 10362
rect 39215 10310 39229 10362
rect 39229 10310 39241 10362
rect 39241 10310 39271 10362
rect 39295 10310 39305 10362
rect 39305 10310 39351 10362
rect 39055 10308 39111 10310
rect 39135 10308 39191 10310
rect 39215 10308 39271 10310
rect 39295 10308 39351 10310
rect 77154 9818 77210 9820
rect 77234 9818 77290 9820
rect 77314 9818 77370 9820
rect 77394 9818 77450 9820
rect 77154 9766 77200 9818
rect 77200 9766 77210 9818
rect 77234 9766 77264 9818
rect 77264 9766 77276 9818
rect 77276 9766 77290 9818
rect 77314 9766 77328 9818
rect 77328 9766 77340 9818
rect 77340 9766 77370 9818
rect 77394 9766 77404 9818
rect 77404 9766 77450 9818
rect 77154 9764 77210 9766
rect 77234 9764 77290 9766
rect 77314 9764 77370 9766
rect 77394 9764 77450 9766
rect 115253 13626 115309 13628
rect 115333 13626 115389 13628
rect 115413 13626 115469 13628
rect 115493 13626 115549 13628
rect 115253 13574 115299 13626
rect 115299 13574 115309 13626
rect 115333 13574 115363 13626
rect 115363 13574 115375 13626
rect 115375 13574 115389 13626
rect 115413 13574 115427 13626
rect 115427 13574 115439 13626
rect 115439 13574 115469 13626
rect 115493 13574 115503 13626
rect 115503 13574 115549 13626
rect 115253 13572 115309 13574
rect 115333 13572 115389 13574
rect 115413 13572 115469 13574
rect 115493 13572 115549 13574
rect 115253 12538 115309 12540
rect 115333 12538 115389 12540
rect 115413 12538 115469 12540
rect 115493 12538 115549 12540
rect 115253 12486 115299 12538
rect 115299 12486 115309 12538
rect 115333 12486 115363 12538
rect 115363 12486 115375 12538
rect 115375 12486 115389 12538
rect 115413 12486 115427 12538
rect 115427 12486 115439 12538
rect 115439 12486 115469 12538
rect 115493 12486 115503 12538
rect 115503 12486 115549 12538
rect 115253 12484 115309 12486
rect 115333 12484 115389 12486
rect 115413 12484 115469 12486
rect 115493 12484 115549 12486
rect 115253 11450 115309 11452
rect 115333 11450 115389 11452
rect 115413 11450 115469 11452
rect 115493 11450 115549 11452
rect 115253 11398 115299 11450
rect 115299 11398 115309 11450
rect 115333 11398 115363 11450
rect 115363 11398 115375 11450
rect 115375 11398 115389 11450
rect 115413 11398 115427 11450
rect 115427 11398 115439 11450
rect 115439 11398 115469 11450
rect 115493 11398 115503 11450
rect 115503 11398 115549 11450
rect 115253 11396 115309 11398
rect 115333 11396 115389 11398
rect 115413 11396 115469 11398
rect 115493 11396 115549 11398
rect 115253 10362 115309 10364
rect 115333 10362 115389 10364
rect 115413 10362 115469 10364
rect 115493 10362 115549 10364
rect 115253 10310 115299 10362
rect 115299 10310 115309 10362
rect 115333 10310 115363 10362
rect 115363 10310 115375 10362
rect 115375 10310 115389 10362
rect 115413 10310 115427 10362
rect 115427 10310 115439 10362
rect 115439 10310 115469 10362
rect 115493 10310 115503 10362
rect 115503 10310 115549 10362
rect 115253 10308 115309 10310
rect 115333 10308 115389 10310
rect 115413 10308 115469 10310
rect 115493 10308 115549 10310
rect 39055 9274 39111 9276
rect 39135 9274 39191 9276
rect 39215 9274 39271 9276
rect 39295 9274 39351 9276
rect 39055 9222 39101 9274
rect 39101 9222 39111 9274
rect 39135 9222 39165 9274
rect 39165 9222 39177 9274
rect 39177 9222 39191 9274
rect 39215 9222 39229 9274
rect 39229 9222 39241 9274
rect 39241 9222 39271 9274
rect 39295 9222 39305 9274
rect 39305 9222 39351 9274
rect 39055 9220 39111 9222
rect 39135 9220 39191 9222
rect 39215 9220 39271 9222
rect 39295 9220 39351 9222
rect 115253 9274 115309 9276
rect 115333 9274 115389 9276
rect 115413 9274 115469 9276
rect 115493 9274 115549 9276
rect 115253 9222 115299 9274
rect 115299 9222 115309 9274
rect 115333 9222 115363 9274
rect 115363 9222 115375 9274
rect 115375 9222 115389 9274
rect 115413 9222 115427 9274
rect 115427 9222 115439 9274
rect 115439 9222 115469 9274
rect 115493 9222 115503 9274
rect 115503 9222 115549 9274
rect 115253 9220 115309 9222
rect 115333 9220 115389 9222
rect 115413 9220 115469 9222
rect 115493 9220 115549 9222
rect 77154 8730 77210 8732
rect 77234 8730 77290 8732
rect 77314 8730 77370 8732
rect 77394 8730 77450 8732
rect 77154 8678 77200 8730
rect 77200 8678 77210 8730
rect 77234 8678 77264 8730
rect 77264 8678 77276 8730
rect 77276 8678 77290 8730
rect 77314 8678 77328 8730
rect 77328 8678 77340 8730
rect 77340 8678 77370 8730
rect 77394 8678 77404 8730
rect 77404 8678 77450 8730
rect 77154 8676 77210 8678
rect 77234 8676 77290 8678
rect 77314 8676 77370 8678
rect 77394 8676 77450 8678
rect 39055 8186 39111 8188
rect 39135 8186 39191 8188
rect 39215 8186 39271 8188
rect 39295 8186 39351 8188
rect 39055 8134 39101 8186
rect 39101 8134 39111 8186
rect 39135 8134 39165 8186
rect 39165 8134 39177 8186
rect 39177 8134 39191 8186
rect 39215 8134 39229 8186
rect 39229 8134 39241 8186
rect 39241 8134 39271 8186
rect 39295 8134 39305 8186
rect 39305 8134 39351 8186
rect 39055 8132 39111 8134
rect 39135 8132 39191 8134
rect 39215 8132 39271 8134
rect 39295 8132 39351 8134
rect 115253 8186 115309 8188
rect 115333 8186 115389 8188
rect 115413 8186 115469 8188
rect 115493 8186 115549 8188
rect 115253 8134 115299 8186
rect 115299 8134 115309 8186
rect 115333 8134 115363 8186
rect 115363 8134 115375 8186
rect 115375 8134 115389 8186
rect 115413 8134 115427 8186
rect 115427 8134 115439 8186
rect 115439 8134 115469 8186
rect 115493 8134 115503 8186
rect 115503 8134 115549 8186
rect 115253 8132 115309 8134
rect 115333 8132 115389 8134
rect 115413 8132 115469 8134
rect 115493 8132 115549 8134
rect 1398 8064 1454 8120
rect 77154 7642 77210 7644
rect 77234 7642 77290 7644
rect 77314 7642 77370 7644
rect 77394 7642 77450 7644
rect 77154 7590 77200 7642
rect 77200 7590 77210 7642
rect 77234 7590 77264 7642
rect 77264 7590 77276 7642
rect 77276 7590 77290 7642
rect 77314 7590 77328 7642
rect 77328 7590 77340 7642
rect 77340 7590 77370 7642
rect 77394 7590 77404 7642
rect 77404 7590 77450 7642
rect 77154 7588 77210 7590
rect 77234 7588 77290 7590
rect 77314 7588 77370 7590
rect 77394 7588 77450 7590
rect 39055 7098 39111 7100
rect 39135 7098 39191 7100
rect 39215 7098 39271 7100
rect 39295 7098 39351 7100
rect 39055 7046 39101 7098
rect 39101 7046 39111 7098
rect 39135 7046 39165 7098
rect 39165 7046 39177 7098
rect 39177 7046 39191 7098
rect 39215 7046 39229 7098
rect 39229 7046 39241 7098
rect 39241 7046 39271 7098
rect 39295 7046 39305 7098
rect 39305 7046 39351 7098
rect 39055 7044 39111 7046
rect 39135 7044 39191 7046
rect 39215 7044 39271 7046
rect 39295 7044 39351 7046
rect 115253 7098 115309 7100
rect 115333 7098 115389 7100
rect 115413 7098 115469 7100
rect 115493 7098 115549 7100
rect 115253 7046 115299 7098
rect 115299 7046 115309 7098
rect 115333 7046 115363 7098
rect 115363 7046 115375 7098
rect 115375 7046 115389 7098
rect 115413 7046 115427 7098
rect 115427 7046 115439 7098
rect 115439 7046 115469 7098
rect 115493 7046 115503 7098
rect 115503 7046 115549 7098
rect 115253 7044 115309 7046
rect 115333 7044 115389 7046
rect 115413 7044 115469 7046
rect 115493 7044 115549 7046
rect 77154 6554 77210 6556
rect 77234 6554 77290 6556
rect 77314 6554 77370 6556
rect 77394 6554 77450 6556
rect 77154 6502 77200 6554
rect 77200 6502 77210 6554
rect 77234 6502 77264 6554
rect 77264 6502 77276 6554
rect 77276 6502 77290 6554
rect 77314 6502 77328 6554
rect 77328 6502 77340 6554
rect 77340 6502 77370 6554
rect 77394 6502 77404 6554
rect 77404 6502 77450 6554
rect 77154 6500 77210 6502
rect 77234 6500 77290 6502
rect 77314 6500 77370 6502
rect 77394 6500 77450 6502
rect 39055 6010 39111 6012
rect 39135 6010 39191 6012
rect 39215 6010 39271 6012
rect 39295 6010 39351 6012
rect 39055 5958 39101 6010
rect 39101 5958 39111 6010
rect 39135 5958 39165 6010
rect 39165 5958 39177 6010
rect 39177 5958 39191 6010
rect 39215 5958 39229 6010
rect 39229 5958 39241 6010
rect 39241 5958 39271 6010
rect 39295 5958 39305 6010
rect 39305 5958 39351 6010
rect 39055 5956 39111 5958
rect 39135 5956 39191 5958
rect 39215 5956 39271 5958
rect 39295 5956 39351 5958
rect 115253 6010 115309 6012
rect 115333 6010 115389 6012
rect 115413 6010 115469 6012
rect 115493 6010 115549 6012
rect 115253 5958 115299 6010
rect 115299 5958 115309 6010
rect 115333 5958 115363 6010
rect 115363 5958 115375 6010
rect 115375 5958 115389 6010
rect 115413 5958 115427 6010
rect 115427 5958 115439 6010
rect 115439 5958 115469 6010
rect 115493 5958 115503 6010
rect 115503 5958 115549 6010
rect 115253 5956 115309 5958
rect 115333 5956 115389 5958
rect 115413 5956 115469 5958
rect 115493 5956 115549 5958
rect 77154 5466 77210 5468
rect 77234 5466 77290 5468
rect 77314 5466 77370 5468
rect 77394 5466 77450 5468
rect 77154 5414 77200 5466
rect 77200 5414 77210 5466
rect 77234 5414 77264 5466
rect 77264 5414 77276 5466
rect 77276 5414 77290 5466
rect 77314 5414 77328 5466
rect 77328 5414 77340 5466
rect 77340 5414 77370 5466
rect 77394 5414 77404 5466
rect 77404 5414 77450 5466
rect 77154 5412 77210 5414
rect 77234 5412 77290 5414
rect 77314 5412 77370 5414
rect 77394 5412 77450 5414
rect 39055 4922 39111 4924
rect 39135 4922 39191 4924
rect 39215 4922 39271 4924
rect 39295 4922 39351 4924
rect 39055 4870 39101 4922
rect 39101 4870 39111 4922
rect 39135 4870 39165 4922
rect 39165 4870 39177 4922
rect 39177 4870 39191 4922
rect 39215 4870 39229 4922
rect 39229 4870 39241 4922
rect 39241 4870 39271 4922
rect 39295 4870 39305 4922
rect 39305 4870 39351 4922
rect 39055 4868 39111 4870
rect 39135 4868 39191 4870
rect 39215 4868 39271 4870
rect 39295 4868 39351 4870
rect 115253 4922 115309 4924
rect 115333 4922 115389 4924
rect 115413 4922 115469 4924
rect 115493 4922 115549 4924
rect 115253 4870 115299 4922
rect 115299 4870 115309 4922
rect 115333 4870 115363 4922
rect 115363 4870 115375 4922
rect 115375 4870 115389 4922
rect 115413 4870 115427 4922
rect 115427 4870 115439 4922
rect 115439 4870 115469 4922
rect 115493 4870 115503 4922
rect 115503 4870 115549 4922
rect 115253 4868 115309 4870
rect 115333 4868 115389 4870
rect 115413 4868 115469 4870
rect 115493 4868 115549 4870
rect 77154 4378 77210 4380
rect 77234 4378 77290 4380
rect 77314 4378 77370 4380
rect 77394 4378 77450 4380
rect 77154 4326 77200 4378
rect 77200 4326 77210 4378
rect 77234 4326 77264 4378
rect 77264 4326 77276 4378
rect 77276 4326 77290 4378
rect 77314 4326 77328 4378
rect 77328 4326 77340 4378
rect 77340 4326 77370 4378
rect 77394 4326 77404 4378
rect 77404 4326 77450 4378
rect 77154 4324 77210 4326
rect 77234 4324 77290 4326
rect 77314 4324 77370 4326
rect 77394 4324 77450 4326
rect 39055 3834 39111 3836
rect 39135 3834 39191 3836
rect 39215 3834 39271 3836
rect 39295 3834 39351 3836
rect 39055 3782 39101 3834
rect 39101 3782 39111 3834
rect 39135 3782 39165 3834
rect 39165 3782 39177 3834
rect 39177 3782 39191 3834
rect 39215 3782 39229 3834
rect 39229 3782 39241 3834
rect 39241 3782 39271 3834
rect 39295 3782 39305 3834
rect 39305 3782 39351 3834
rect 39055 3780 39111 3782
rect 39135 3780 39191 3782
rect 39215 3780 39271 3782
rect 39295 3780 39351 3782
rect 115253 3834 115309 3836
rect 115333 3834 115389 3836
rect 115413 3834 115469 3836
rect 115493 3834 115549 3836
rect 115253 3782 115299 3834
rect 115299 3782 115309 3834
rect 115333 3782 115363 3834
rect 115363 3782 115375 3834
rect 115375 3782 115389 3834
rect 115413 3782 115427 3834
rect 115427 3782 115439 3834
rect 115439 3782 115469 3834
rect 115493 3782 115503 3834
rect 115503 3782 115549 3834
rect 115253 3780 115309 3782
rect 115333 3780 115389 3782
rect 115413 3780 115469 3782
rect 115493 3780 115549 3782
rect 77154 3290 77210 3292
rect 77234 3290 77290 3292
rect 77314 3290 77370 3292
rect 77394 3290 77450 3292
rect 77154 3238 77200 3290
rect 77200 3238 77210 3290
rect 77234 3238 77264 3290
rect 77264 3238 77276 3290
rect 77276 3238 77290 3290
rect 77314 3238 77328 3290
rect 77328 3238 77340 3290
rect 77340 3238 77370 3290
rect 77394 3238 77404 3290
rect 77404 3238 77450 3290
rect 77154 3236 77210 3238
rect 77234 3236 77290 3238
rect 77314 3236 77370 3238
rect 77394 3236 77450 3238
rect 39055 2746 39111 2748
rect 39135 2746 39191 2748
rect 39215 2746 39271 2748
rect 39295 2746 39351 2748
rect 39055 2694 39101 2746
rect 39101 2694 39111 2746
rect 39135 2694 39165 2746
rect 39165 2694 39177 2746
rect 39177 2694 39191 2746
rect 39215 2694 39229 2746
rect 39229 2694 39241 2746
rect 39241 2694 39271 2746
rect 39295 2694 39305 2746
rect 39305 2694 39351 2746
rect 39055 2692 39111 2694
rect 39135 2692 39191 2694
rect 39215 2692 39271 2694
rect 39295 2692 39351 2694
rect 115253 2746 115309 2748
rect 115333 2746 115389 2748
rect 115413 2746 115469 2748
rect 115493 2746 115549 2748
rect 115253 2694 115299 2746
rect 115299 2694 115309 2746
rect 115333 2694 115363 2746
rect 115363 2694 115375 2746
rect 115375 2694 115389 2746
rect 115413 2694 115427 2746
rect 115427 2694 115439 2746
rect 115439 2694 115469 2746
rect 115493 2694 115503 2746
rect 115503 2694 115549 2746
rect 115253 2692 115309 2694
rect 115333 2692 115389 2694
rect 115413 2692 115469 2694
rect 115493 2692 115549 2694
rect 153352 13082 153408 13084
rect 153432 13082 153488 13084
rect 153512 13082 153568 13084
rect 153592 13082 153648 13084
rect 153352 13030 153398 13082
rect 153398 13030 153408 13082
rect 153432 13030 153462 13082
rect 153462 13030 153474 13082
rect 153474 13030 153488 13082
rect 153512 13030 153526 13082
rect 153526 13030 153538 13082
rect 153538 13030 153568 13082
rect 153592 13030 153602 13082
rect 153602 13030 153648 13082
rect 153352 13028 153408 13030
rect 153432 13028 153488 13030
rect 153512 13028 153568 13030
rect 153592 13028 153648 13030
rect 153352 11994 153408 11996
rect 153432 11994 153488 11996
rect 153512 11994 153568 11996
rect 153592 11994 153648 11996
rect 153352 11942 153398 11994
rect 153398 11942 153408 11994
rect 153432 11942 153462 11994
rect 153462 11942 153474 11994
rect 153474 11942 153488 11994
rect 153512 11942 153526 11994
rect 153526 11942 153538 11994
rect 153538 11942 153568 11994
rect 153592 11942 153602 11994
rect 153602 11942 153648 11994
rect 153352 11940 153408 11942
rect 153432 11940 153488 11942
rect 153512 11940 153568 11942
rect 153592 11940 153648 11942
rect 155038 12824 155094 12880
rect 157890 12588 157892 12608
rect 157892 12588 157944 12608
rect 157944 12588 157946 12608
rect 157890 12552 157946 12588
rect 153352 10906 153408 10908
rect 153432 10906 153488 10908
rect 153512 10906 153568 10908
rect 153592 10906 153648 10908
rect 153352 10854 153398 10906
rect 153398 10854 153408 10906
rect 153432 10854 153462 10906
rect 153462 10854 153474 10906
rect 153474 10854 153488 10906
rect 153512 10854 153526 10906
rect 153526 10854 153538 10906
rect 153538 10854 153568 10906
rect 153592 10854 153602 10906
rect 153602 10854 153648 10906
rect 153352 10852 153408 10854
rect 153432 10852 153488 10854
rect 153512 10852 153568 10854
rect 153592 10852 153648 10854
rect 153352 9818 153408 9820
rect 153432 9818 153488 9820
rect 153512 9818 153568 9820
rect 153592 9818 153648 9820
rect 153352 9766 153398 9818
rect 153398 9766 153408 9818
rect 153432 9766 153462 9818
rect 153462 9766 153474 9818
rect 153474 9766 153488 9818
rect 153512 9766 153526 9818
rect 153526 9766 153538 9818
rect 153538 9766 153568 9818
rect 153592 9766 153602 9818
rect 153602 9766 153648 9818
rect 153352 9764 153408 9766
rect 153432 9764 153488 9766
rect 153512 9764 153568 9766
rect 153592 9764 153648 9766
rect 160282 12588 160284 12608
rect 160284 12588 160336 12608
rect 160336 12588 160338 12608
rect 160282 12552 160338 12588
rect 163594 12300 163650 12336
rect 163594 12280 163596 12300
rect 163596 12280 163648 12300
rect 163648 12280 163650 12300
rect 189630 11756 189686 11792
rect 189630 11736 189632 11756
rect 189632 11736 189684 11756
rect 189684 11736 189686 11756
rect 153352 8730 153408 8732
rect 153432 8730 153488 8732
rect 153512 8730 153568 8732
rect 153592 8730 153648 8732
rect 153352 8678 153398 8730
rect 153398 8678 153408 8730
rect 153432 8678 153462 8730
rect 153462 8678 153474 8730
rect 153474 8678 153488 8730
rect 153512 8678 153526 8730
rect 153526 8678 153538 8730
rect 153538 8678 153568 8730
rect 153592 8678 153602 8730
rect 153602 8678 153648 8730
rect 153352 8676 153408 8678
rect 153432 8676 153488 8678
rect 153512 8676 153568 8678
rect 153592 8676 153648 8678
rect 191451 13626 191507 13628
rect 191531 13626 191587 13628
rect 191611 13626 191667 13628
rect 191691 13626 191747 13628
rect 191451 13574 191497 13626
rect 191497 13574 191507 13626
rect 191531 13574 191561 13626
rect 191561 13574 191573 13626
rect 191573 13574 191587 13626
rect 191611 13574 191625 13626
rect 191625 13574 191637 13626
rect 191637 13574 191667 13626
rect 191691 13574 191701 13626
rect 191701 13574 191747 13626
rect 191451 13572 191507 13574
rect 191531 13572 191587 13574
rect 191611 13572 191667 13574
rect 191691 13572 191747 13574
rect 191838 12552 191894 12608
rect 191451 12538 191507 12540
rect 191531 12538 191587 12540
rect 191611 12538 191667 12540
rect 191691 12538 191747 12540
rect 191451 12486 191497 12538
rect 191497 12486 191507 12538
rect 191531 12486 191561 12538
rect 191561 12486 191573 12538
rect 191573 12486 191587 12538
rect 191611 12486 191625 12538
rect 191625 12486 191637 12538
rect 191637 12486 191667 12538
rect 191691 12486 191701 12538
rect 191701 12486 191747 12538
rect 191451 12484 191507 12486
rect 191531 12484 191587 12486
rect 191611 12484 191667 12486
rect 191691 12484 191747 12486
rect 192206 12552 192262 12608
rect 191451 11450 191507 11452
rect 191531 11450 191587 11452
rect 191611 11450 191667 11452
rect 191691 11450 191747 11452
rect 191451 11398 191497 11450
rect 191497 11398 191507 11450
rect 191531 11398 191561 11450
rect 191561 11398 191573 11450
rect 191573 11398 191587 11450
rect 191611 11398 191625 11450
rect 191625 11398 191637 11450
rect 191637 11398 191667 11450
rect 191691 11398 191701 11450
rect 191701 11398 191747 11450
rect 191451 11396 191507 11398
rect 191531 11396 191587 11398
rect 191611 11396 191667 11398
rect 191691 11396 191747 11398
rect 191451 10362 191507 10364
rect 191531 10362 191587 10364
rect 191611 10362 191667 10364
rect 191691 10362 191747 10364
rect 191451 10310 191497 10362
rect 191497 10310 191507 10362
rect 191531 10310 191561 10362
rect 191561 10310 191573 10362
rect 191573 10310 191587 10362
rect 191611 10310 191625 10362
rect 191625 10310 191637 10362
rect 191637 10310 191667 10362
rect 191691 10310 191701 10362
rect 191701 10310 191747 10362
rect 191451 10308 191507 10310
rect 191531 10308 191587 10310
rect 191611 10308 191667 10310
rect 191691 10308 191747 10310
rect 193034 12280 193090 12336
rect 193034 11736 193090 11792
rect 194598 12824 194654 12880
rect 195058 12688 195114 12744
rect 195794 12824 195850 12880
rect 197358 12844 197414 12880
rect 197358 12824 197360 12844
rect 197360 12824 197412 12844
rect 197412 12824 197414 12844
rect 200854 13232 200910 13288
rect 200394 12552 200450 12608
rect 203430 13232 203486 13288
rect 207110 13524 207166 13560
rect 207110 13504 207112 13524
rect 207112 13504 207164 13524
rect 207164 13504 207166 13524
rect 205546 13232 205602 13288
rect 205270 12588 205272 12608
rect 205272 12588 205324 12608
rect 205324 12588 205326 12608
rect 205270 12552 205326 12588
rect 205730 13232 205786 13288
rect 207202 13268 207204 13288
rect 207204 13268 207256 13288
rect 207256 13268 207258 13288
rect 207202 13232 207258 13268
rect 208030 13504 208086 13560
rect 213274 13404 213276 13424
rect 213276 13404 213328 13424
rect 213328 13404 213330 13424
rect 213274 13368 213330 13404
rect 219806 13368 219862 13424
rect 207938 13268 207940 13288
rect 207940 13268 207992 13288
rect 207992 13268 207994 13288
rect 207938 13232 207994 13268
rect 207846 12688 207902 12744
rect 225418 13132 225420 13152
rect 225420 13132 225472 13152
rect 225472 13132 225474 13152
rect 225418 13096 225474 13132
rect 227074 13388 227130 13424
rect 227074 13368 227076 13388
rect 227076 13368 227128 13388
rect 227128 13368 227130 13388
rect 227074 13132 227076 13152
rect 227076 13132 227128 13152
rect 227128 13132 227130 13152
rect 227074 13096 227130 13132
rect 229190 13404 229192 13424
rect 229192 13404 229244 13424
rect 229244 13404 229246 13424
rect 229190 13368 229246 13404
rect 230386 13268 230388 13288
rect 230388 13268 230440 13288
rect 230440 13268 230442 13288
rect 230386 13232 230442 13268
rect 229550 13082 229606 13084
rect 229630 13082 229686 13084
rect 229710 13082 229766 13084
rect 229790 13082 229846 13084
rect 229550 13030 229596 13082
rect 229596 13030 229606 13082
rect 229630 13030 229660 13082
rect 229660 13030 229672 13082
rect 229672 13030 229686 13082
rect 229710 13030 229724 13082
rect 229724 13030 229736 13082
rect 229736 13030 229766 13082
rect 229790 13030 229800 13082
rect 229800 13030 229846 13082
rect 229550 13028 229606 13030
rect 229630 13028 229686 13030
rect 229710 13028 229766 13030
rect 229790 13028 229846 13030
rect 229550 11994 229606 11996
rect 229630 11994 229686 11996
rect 229710 11994 229766 11996
rect 229790 11994 229846 11996
rect 229550 11942 229596 11994
rect 229596 11942 229606 11994
rect 229630 11942 229660 11994
rect 229660 11942 229672 11994
rect 229672 11942 229686 11994
rect 229710 11942 229724 11994
rect 229724 11942 229736 11994
rect 229736 11942 229766 11994
rect 229790 11942 229800 11994
rect 229800 11942 229846 11994
rect 229550 11940 229606 11942
rect 229630 11940 229686 11942
rect 229710 11940 229766 11942
rect 229790 11940 229846 11942
rect 232134 13232 232190 13288
rect 238114 13388 238170 13424
rect 238114 13368 238116 13388
rect 238116 13368 238168 13388
rect 238168 13368 238170 13388
rect 239494 13404 239496 13424
rect 239496 13404 239548 13424
rect 239548 13404 239550 13424
rect 239494 13368 239550 13404
rect 238298 12688 238354 12744
rect 242162 12708 242218 12744
rect 242162 12688 242164 12708
rect 242164 12688 242216 12708
rect 242216 12688 242218 12708
rect 229550 10906 229606 10908
rect 229630 10906 229686 10908
rect 229710 10906 229766 10908
rect 229790 10906 229846 10908
rect 229550 10854 229596 10906
rect 229596 10854 229606 10906
rect 229630 10854 229660 10906
rect 229660 10854 229672 10906
rect 229672 10854 229686 10906
rect 229710 10854 229724 10906
rect 229724 10854 229736 10906
rect 229736 10854 229766 10906
rect 229790 10854 229800 10906
rect 229800 10854 229846 10906
rect 229550 10852 229606 10854
rect 229630 10852 229686 10854
rect 229710 10852 229766 10854
rect 229790 10852 229846 10854
rect 229550 9818 229606 9820
rect 229630 9818 229686 9820
rect 229710 9818 229766 9820
rect 229790 9818 229846 9820
rect 229550 9766 229596 9818
rect 229596 9766 229606 9818
rect 229630 9766 229660 9818
rect 229660 9766 229672 9818
rect 229672 9766 229686 9818
rect 229710 9766 229724 9818
rect 229724 9766 229736 9818
rect 229736 9766 229766 9818
rect 229790 9766 229800 9818
rect 229800 9766 229846 9818
rect 229550 9764 229606 9766
rect 229630 9764 229686 9766
rect 229710 9764 229766 9766
rect 229790 9764 229846 9766
rect 191451 9274 191507 9276
rect 191531 9274 191587 9276
rect 191611 9274 191667 9276
rect 191691 9274 191747 9276
rect 191451 9222 191497 9274
rect 191497 9222 191507 9274
rect 191531 9222 191561 9274
rect 191561 9222 191573 9274
rect 191573 9222 191587 9274
rect 191611 9222 191625 9274
rect 191625 9222 191637 9274
rect 191637 9222 191667 9274
rect 191691 9222 191701 9274
rect 191701 9222 191747 9274
rect 191451 9220 191507 9222
rect 191531 9220 191587 9222
rect 191611 9220 191667 9222
rect 191691 9220 191747 9222
rect 229550 8730 229606 8732
rect 229630 8730 229686 8732
rect 229710 8730 229766 8732
rect 229790 8730 229846 8732
rect 229550 8678 229596 8730
rect 229596 8678 229606 8730
rect 229630 8678 229660 8730
rect 229660 8678 229672 8730
rect 229672 8678 229686 8730
rect 229710 8678 229724 8730
rect 229724 8678 229736 8730
rect 229736 8678 229766 8730
rect 229790 8678 229800 8730
rect 229800 8678 229846 8730
rect 229550 8676 229606 8678
rect 229630 8676 229686 8678
rect 229710 8676 229766 8678
rect 229790 8676 229846 8678
rect 191451 8186 191507 8188
rect 191531 8186 191587 8188
rect 191611 8186 191667 8188
rect 191691 8186 191747 8188
rect 191451 8134 191497 8186
rect 191497 8134 191507 8186
rect 191531 8134 191561 8186
rect 191561 8134 191573 8186
rect 191573 8134 191587 8186
rect 191611 8134 191625 8186
rect 191625 8134 191637 8186
rect 191637 8134 191667 8186
rect 191691 8134 191701 8186
rect 191701 8134 191747 8186
rect 191451 8132 191507 8134
rect 191531 8132 191587 8134
rect 191611 8132 191667 8134
rect 191691 8132 191747 8134
rect 153352 7642 153408 7644
rect 153432 7642 153488 7644
rect 153512 7642 153568 7644
rect 153592 7642 153648 7644
rect 153352 7590 153398 7642
rect 153398 7590 153408 7642
rect 153432 7590 153462 7642
rect 153462 7590 153474 7642
rect 153474 7590 153488 7642
rect 153512 7590 153526 7642
rect 153526 7590 153538 7642
rect 153538 7590 153568 7642
rect 153592 7590 153602 7642
rect 153602 7590 153648 7642
rect 153352 7588 153408 7590
rect 153432 7588 153488 7590
rect 153512 7588 153568 7590
rect 153592 7588 153648 7590
rect 229550 7642 229606 7644
rect 229630 7642 229686 7644
rect 229710 7642 229766 7644
rect 229790 7642 229846 7644
rect 229550 7590 229596 7642
rect 229596 7590 229606 7642
rect 229630 7590 229660 7642
rect 229660 7590 229672 7642
rect 229672 7590 229686 7642
rect 229710 7590 229724 7642
rect 229724 7590 229736 7642
rect 229736 7590 229766 7642
rect 229790 7590 229800 7642
rect 229800 7590 229846 7642
rect 229550 7588 229606 7590
rect 229630 7588 229686 7590
rect 229710 7588 229766 7590
rect 229790 7588 229846 7590
rect 191451 7098 191507 7100
rect 191531 7098 191587 7100
rect 191611 7098 191667 7100
rect 191691 7098 191747 7100
rect 191451 7046 191497 7098
rect 191497 7046 191507 7098
rect 191531 7046 191561 7098
rect 191561 7046 191573 7098
rect 191573 7046 191587 7098
rect 191611 7046 191625 7098
rect 191625 7046 191637 7098
rect 191637 7046 191667 7098
rect 191691 7046 191701 7098
rect 191701 7046 191747 7098
rect 191451 7044 191507 7046
rect 191531 7044 191587 7046
rect 191611 7044 191667 7046
rect 191691 7044 191747 7046
rect 153352 6554 153408 6556
rect 153432 6554 153488 6556
rect 153512 6554 153568 6556
rect 153592 6554 153648 6556
rect 153352 6502 153398 6554
rect 153398 6502 153408 6554
rect 153432 6502 153462 6554
rect 153462 6502 153474 6554
rect 153474 6502 153488 6554
rect 153512 6502 153526 6554
rect 153526 6502 153538 6554
rect 153538 6502 153568 6554
rect 153592 6502 153602 6554
rect 153602 6502 153648 6554
rect 153352 6500 153408 6502
rect 153432 6500 153488 6502
rect 153512 6500 153568 6502
rect 153592 6500 153648 6502
rect 229550 6554 229606 6556
rect 229630 6554 229686 6556
rect 229710 6554 229766 6556
rect 229790 6554 229846 6556
rect 229550 6502 229596 6554
rect 229596 6502 229606 6554
rect 229630 6502 229660 6554
rect 229660 6502 229672 6554
rect 229672 6502 229686 6554
rect 229710 6502 229724 6554
rect 229724 6502 229736 6554
rect 229736 6502 229766 6554
rect 229790 6502 229800 6554
rect 229800 6502 229846 6554
rect 229550 6500 229606 6502
rect 229630 6500 229686 6502
rect 229710 6500 229766 6502
rect 229790 6500 229846 6502
rect 251914 12588 251916 12608
rect 251916 12588 251968 12608
rect 251968 12588 251970 12608
rect 251914 12552 251970 12588
rect 251822 12416 251878 12472
rect 256606 12960 256662 13016
rect 257986 12960 258042 13016
rect 257066 12552 257122 12608
rect 257158 12416 257214 12472
rect 262310 12724 262312 12744
rect 262312 12724 262364 12744
rect 262364 12724 262366 12744
rect 262310 12688 262366 12724
rect 263414 13252 263470 13288
rect 263414 13232 263416 13252
rect 263416 13232 263468 13252
rect 263468 13232 263470 13252
rect 263506 12708 263562 12744
rect 263506 12688 263508 12708
rect 263508 12688 263560 12708
rect 263560 12688 263562 12708
rect 264334 12688 264390 12744
rect 267649 13626 267705 13628
rect 267729 13626 267785 13628
rect 267809 13626 267865 13628
rect 267889 13626 267945 13628
rect 267649 13574 267695 13626
rect 267695 13574 267705 13626
rect 267729 13574 267759 13626
rect 267759 13574 267771 13626
rect 267771 13574 267785 13626
rect 267809 13574 267823 13626
rect 267823 13574 267835 13626
rect 267835 13574 267865 13626
rect 267889 13574 267899 13626
rect 267899 13574 267945 13626
rect 267649 13572 267705 13574
rect 267729 13572 267785 13574
rect 267809 13572 267865 13574
rect 267889 13572 267945 13574
rect 265530 13232 265586 13288
rect 267094 12688 267150 12744
rect 267646 12688 267702 12744
rect 267649 12538 267705 12540
rect 267729 12538 267785 12540
rect 267809 12538 267865 12540
rect 267889 12538 267945 12540
rect 267649 12486 267695 12538
rect 267695 12486 267705 12538
rect 267729 12486 267759 12538
rect 267759 12486 267771 12538
rect 267771 12486 267785 12538
rect 267809 12486 267823 12538
rect 267823 12486 267835 12538
rect 267835 12486 267865 12538
rect 267889 12486 267899 12538
rect 267899 12486 267945 12538
rect 267649 12484 267705 12486
rect 267729 12484 267785 12486
rect 267809 12484 267865 12486
rect 267889 12484 267945 12486
rect 268106 12688 268162 12744
rect 267649 11450 267705 11452
rect 267729 11450 267785 11452
rect 267809 11450 267865 11452
rect 267889 11450 267945 11452
rect 267649 11398 267695 11450
rect 267695 11398 267705 11450
rect 267729 11398 267759 11450
rect 267759 11398 267771 11450
rect 267771 11398 267785 11450
rect 267809 11398 267823 11450
rect 267823 11398 267835 11450
rect 267835 11398 267865 11450
rect 267889 11398 267899 11450
rect 267899 11398 267945 11450
rect 267649 11396 267705 11398
rect 267729 11396 267785 11398
rect 267809 11396 267865 11398
rect 267889 11396 267945 11398
rect 267649 10362 267705 10364
rect 267729 10362 267785 10364
rect 267809 10362 267865 10364
rect 267889 10362 267945 10364
rect 267649 10310 267695 10362
rect 267695 10310 267705 10362
rect 267729 10310 267759 10362
rect 267759 10310 267771 10362
rect 267771 10310 267785 10362
rect 267809 10310 267823 10362
rect 267823 10310 267835 10362
rect 267835 10310 267865 10362
rect 267889 10310 267899 10362
rect 267899 10310 267945 10362
rect 267649 10308 267705 10310
rect 267729 10308 267785 10310
rect 267809 10308 267865 10310
rect 267889 10308 267945 10310
rect 268934 13368 268990 13424
rect 269026 13232 269082 13288
rect 273166 13388 273222 13424
rect 273166 13368 273168 13388
rect 273168 13368 273220 13388
rect 273220 13368 273222 13388
rect 273258 13268 273260 13288
rect 273260 13268 273312 13288
rect 273312 13268 273314 13288
rect 273258 13232 273314 13268
rect 303526 13912 303582 13968
rect 299478 12824 299534 12880
rect 304446 10004 304448 10024
rect 304448 10004 304500 10024
rect 304500 10004 304502 10024
rect 304446 9968 304502 10004
rect 267649 9274 267705 9276
rect 267729 9274 267785 9276
rect 267809 9274 267865 9276
rect 267889 9274 267945 9276
rect 267649 9222 267695 9274
rect 267695 9222 267705 9274
rect 267729 9222 267759 9274
rect 267759 9222 267771 9274
rect 267771 9222 267785 9274
rect 267809 9222 267823 9274
rect 267823 9222 267835 9274
rect 267835 9222 267865 9274
rect 267889 9222 267899 9274
rect 267899 9222 267945 9274
rect 267649 9220 267705 9222
rect 267729 9220 267785 9222
rect 267809 9220 267865 9222
rect 267889 9220 267945 9222
rect 267649 8186 267705 8188
rect 267729 8186 267785 8188
rect 267809 8186 267865 8188
rect 267889 8186 267945 8188
rect 267649 8134 267695 8186
rect 267695 8134 267705 8186
rect 267729 8134 267759 8186
rect 267759 8134 267771 8186
rect 267771 8134 267785 8186
rect 267809 8134 267823 8186
rect 267823 8134 267835 8186
rect 267835 8134 267865 8186
rect 267889 8134 267899 8186
rect 267899 8134 267945 8186
rect 267649 8132 267705 8134
rect 267729 8132 267785 8134
rect 267809 8132 267865 8134
rect 267889 8132 267945 8134
rect 267649 7098 267705 7100
rect 267729 7098 267785 7100
rect 267809 7098 267865 7100
rect 267889 7098 267945 7100
rect 267649 7046 267695 7098
rect 267695 7046 267705 7098
rect 267729 7046 267759 7098
rect 267759 7046 267771 7098
rect 267771 7046 267785 7098
rect 267809 7046 267823 7098
rect 267823 7046 267835 7098
rect 267835 7046 267865 7098
rect 267889 7046 267899 7098
rect 267899 7046 267945 7098
rect 267649 7044 267705 7046
rect 267729 7044 267785 7046
rect 267809 7044 267865 7046
rect 267889 7044 267945 7046
rect 191451 6010 191507 6012
rect 191531 6010 191587 6012
rect 191611 6010 191667 6012
rect 191691 6010 191747 6012
rect 191451 5958 191497 6010
rect 191497 5958 191507 6010
rect 191531 5958 191561 6010
rect 191561 5958 191573 6010
rect 191573 5958 191587 6010
rect 191611 5958 191625 6010
rect 191625 5958 191637 6010
rect 191637 5958 191667 6010
rect 191691 5958 191701 6010
rect 191701 5958 191747 6010
rect 191451 5956 191507 5958
rect 191531 5956 191587 5958
rect 191611 5956 191667 5958
rect 191691 5956 191747 5958
rect 267649 6010 267705 6012
rect 267729 6010 267785 6012
rect 267809 6010 267865 6012
rect 267889 6010 267945 6012
rect 267649 5958 267695 6010
rect 267695 5958 267705 6010
rect 267729 5958 267759 6010
rect 267759 5958 267771 6010
rect 267771 5958 267785 6010
rect 267809 5958 267823 6010
rect 267823 5958 267835 6010
rect 267835 5958 267865 6010
rect 267889 5958 267899 6010
rect 267899 5958 267945 6010
rect 267649 5956 267705 5958
rect 267729 5956 267785 5958
rect 267809 5956 267865 5958
rect 267889 5956 267945 5958
rect 303986 5888 304042 5944
rect 153352 5466 153408 5468
rect 153432 5466 153488 5468
rect 153512 5466 153568 5468
rect 153592 5466 153648 5468
rect 153352 5414 153398 5466
rect 153398 5414 153408 5466
rect 153432 5414 153462 5466
rect 153462 5414 153474 5466
rect 153474 5414 153488 5466
rect 153512 5414 153526 5466
rect 153526 5414 153538 5466
rect 153538 5414 153568 5466
rect 153592 5414 153602 5466
rect 153602 5414 153648 5466
rect 153352 5412 153408 5414
rect 153432 5412 153488 5414
rect 153512 5412 153568 5414
rect 153592 5412 153648 5414
rect 229550 5466 229606 5468
rect 229630 5466 229686 5468
rect 229710 5466 229766 5468
rect 229790 5466 229846 5468
rect 229550 5414 229596 5466
rect 229596 5414 229606 5466
rect 229630 5414 229660 5466
rect 229660 5414 229672 5466
rect 229672 5414 229686 5466
rect 229710 5414 229724 5466
rect 229724 5414 229736 5466
rect 229736 5414 229766 5466
rect 229790 5414 229800 5466
rect 229800 5414 229846 5466
rect 229550 5412 229606 5414
rect 229630 5412 229686 5414
rect 229710 5412 229766 5414
rect 229790 5412 229846 5414
rect 191451 4922 191507 4924
rect 191531 4922 191587 4924
rect 191611 4922 191667 4924
rect 191691 4922 191747 4924
rect 191451 4870 191497 4922
rect 191497 4870 191507 4922
rect 191531 4870 191561 4922
rect 191561 4870 191573 4922
rect 191573 4870 191587 4922
rect 191611 4870 191625 4922
rect 191625 4870 191637 4922
rect 191637 4870 191667 4922
rect 191691 4870 191701 4922
rect 191701 4870 191747 4922
rect 191451 4868 191507 4870
rect 191531 4868 191587 4870
rect 191611 4868 191667 4870
rect 191691 4868 191747 4870
rect 267649 4922 267705 4924
rect 267729 4922 267785 4924
rect 267809 4922 267865 4924
rect 267889 4922 267945 4924
rect 267649 4870 267695 4922
rect 267695 4870 267705 4922
rect 267729 4870 267759 4922
rect 267759 4870 267771 4922
rect 267771 4870 267785 4922
rect 267809 4870 267823 4922
rect 267823 4870 267835 4922
rect 267835 4870 267865 4922
rect 267889 4870 267899 4922
rect 267899 4870 267945 4922
rect 267649 4868 267705 4870
rect 267729 4868 267785 4870
rect 267809 4868 267865 4870
rect 267889 4868 267945 4870
rect 153352 4378 153408 4380
rect 153432 4378 153488 4380
rect 153512 4378 153568 4380
rect 153592 4378 153648 4380
rect 153352 4326 153398 4378
rect 153398 4326 153408 4378
rect 153432 4326 153462 4378
rect 153462 4326 153474 4378
rect 153474 4326 153488 4378
rect 153512 4326 153526 4378
rect 153526 4326 153538 4378
rect 153538 4326 153568 4378
rect 153592 4326 153602 4378
rect 153602 4326 153648 4378
rect 153352 4324 153408 4326
rect 153432 4324 153488 4326
rect 153512 4324 153568 4326
rect 153592 4324 153648 4326
rect 229550 4378 229606 4380
rect 229630 4378 229686 4380
rect 229710 4378 229766 4380
rect 229790 4378 229846 4380
rect 229550 4326 229596 4378
rect 229596 4326 229606 4378
rect 229630 4326 229660 4378
rect 229660 4326 229672 4378
rect 229672 4326 229686 4378
rect 229710 4326 229724 4378
rect 229724 4326 229736 4378
rect 229736 4326 229766 4378
rect 229790 4326 229800 4378
rect 229800 4326 229846 4378
rect 229550 4324 229606 4326
rect 229630 4324 229686 4326
rect 229710 4324 229766 4326
rect 229790 4324 229846 4326
rect 191451 3834 191507 3836
rect 191531 3834 191587 3836
rect 191611 3834 191667 3836
rect 191691 3834 191747 3836
rect 191451 3782 191497 3834
rect 191497 3782 191507 3834
rect 191531 3782 191561 3834
rect 191561 3782 191573 3834
rect 191573 3782 191587 3834
rect 191611 3782 191625 3834
rect 191625 3782 191637 3834
rect 191637 3782 191667 3834
rect 191691 3782 191701 3834
rect 191701 3782 191747 3834
rect 191451 3780 191507 3782
rect 191531 3780 191587 3782
rect 191611 3780 191667 3782
rect 191691 3780 191747 3782
rect 267649 3834 267705 3836
rect 267729 3834 267785 3836
rect 267809 3834 267865 3836
rect 267889 3834 267945 3836
rect 267649 3782 267695 3834
rect 267695 3782 267705 3834
rect 267729 3782 267759 3834
rect 267759 3782 267771 3834
rect 267771 3782 267785 3834
rect 267809 3782 267823 3834
rect 267823 3782 267835 3834
rect 267835 3782 267865 3834
rect 267889 3782 267899 3834
rect 267899 3782 267945 3834
rect 267649 3780 267705 3782
rect 267729 3780 267785 3782
rect 267809 3780 267865 3782
rect 267889 3780 267945 3782
rect 153352 3290 153408 3292
rect 153432 3290 153488 3292
rect 153512 3290 153568 3292
rect 153592 3290 153648 3292
rect 153352 3238 153398 3290
rect 153398 3238 153408 3290
rect 153432 3238 153462 3290
rect 153462 3238 153474 3290
rect 153474 3238 153488 3290
rect 153512 3238 153526 3290
rect 153526 3238 153538 3290
rect 153538 3238 153568 3290
rect 153592 3238 153602 3290
rect 153602 3238 153648 3290
rect 153352 3236 153408 3238
rect 153432 3236 153488 3238
rect 153512 3236 153568 3238
rect 153592 3236 153648 3238
rect 229550 3290 229606 3292
rect 229630 3290 229686 3292
rect 229710 3290 229766 3292
rect 229790 3290 229846 3292
rect 229550 3238 229596 3290
rect 229596 3238 229606 3290
rect 229630 3238 229660 3290
rect 229660 3238 229672 3290
rect 229672 3238 229686 3290
rect 229710 3238 229724 3290
rect 229724 3238 229736 3290
rect 229736 3238 229766 3290
rect 229790 3238 229800 3290
rect 229800 3238 229846 3290
rect 229550 3236 229606 3238
rect 229630 3236 229686 3238
rect 229710 3236 229766 3238
rect 229790 3236 229846 3238
rect 191451 2746 191507 2748
rect 191531 2746 191587 2748
rect 191611 2746 191667 2748
rect 191691 2746 191747 2748
rect 191451 2694 191497 2746
rect 191497 2694 191507 2746
rect 191531 2694 191561 2746
rect 191561 2694 191573 2746
rect 191573 2694 191587 2746
rect 191611 2694 191625 2746
rect 191625 2694 191637 2746
rect 191637 2694 191667 2746
rect 191691 2694 191701 2746
rect 191701 2694 191747 2746
rect 191451 2692 191507 2694
rect 191531 2692 191587 2694
rect 191611 2692 191667 2694
rect 191691 2692 191747 2694
rect 267649 2746 267705 2748
rect 267729 2746 267785 2748
rect 267809 2746 267865 2748
rect 267889 2746 267945 2748
rect 267649 2694 267695 2746
rect 267695 2694 267705 2746
rect 267729 2694 267759 2746
rect 267759 2694 267771 2746
rect 267771 2694 267785 2746
rect 267809 2694 267823 2746
rect 267823 2694 267835 2746
rect 267835 2694 267865 2746
rect 267889 2694 267899 2746
rect 267899 2694 267945 2746
rect 267649 2692 267705 2694
rect 267729 2692 267785 2694
rect 267809 2692 267865 2694
rect 267889 2692 267945 2694
rect 77154 2202 77210 2204
rect 77234 2202 77290 2204
rect 77314 2202 77370 2204
rect 77394 2202 77450 2204
rect 77154 2150 77200 2202
rect 77200 2150 77210 2202
rect 77234 2150 77264 2202
rect 77264 2150 77276 2202
rect 77276 2150 77290 2202
rect 77314 2150 77328 2202
rect 77328 2150 77340 2202
rect 77340 2150 77370 2202
rect 77394 2150 77404 2202
rect 77404 2150 77450 2202
rect 77154 2148 77210 2150
rect 77234 2148 77290 2150
rect 77314 2148 77370 2150
rect 77394 2148 77450 2150
rect 153352 2202 153408 2204
rect 153432 2202 153488 2204
rect 153512 2202 153568 2204
rect 153592 2202 153648 2204
rect 153352 2150 153398 2202
rect 153398 2150 153408 2202
rect 153432 2150 153462 2202
rect 153462 2150 153474 2202
rect 153474 2150 153488 2202
rect 153512 2150 153526 2202
rect 153526 2150 153538 2202
rect 153538 2150 153568 2202
rect 153592 2150 153602 2202
rect 153602 2150 153648 2202
rect 153352 2148 153408 2150
rect 153432 2148 153488 2150
rect 153512 2148 153568 2150
rect 153592 2148 153648 2150
rect 229550 2202 229606 2204
rect 229630 2202 229686 2204
rect 229710 2202 229766 2204
rect 229790 2202 229846 2204
rect 229550 2150 229596 2202
rect 229596 2150 229606 2202
rect 229630 2150 229660 2202
rect 229660 2150 229672 2202
rect 229672 2150 229686 2202
rect 229710 2150 229724 2202
rect 229724 2150 229736 2202
rect 229736 2150 229766 2202
rect 229790 2150 229800 2202
rect 229800 2150 229846 2202
rect 229550 2148 229606 2150
rect 229630 2148 229686 2150
rect 229710 2148 229766 2150
rect 229790 2148 229846 2150
rect 302238 1944 302294 2000
<< metal3 >>
rect 303521 13970 303587 13973
rect 306200 13970 307000 14000
rect 303521 13968 307000 13970
rect 303521 13912 303526 13968
rect 303582 13912 307000 13968
rect 303521 13910 307000 13912
rect 303521 13907 303587 13910
rect 306200 13880 307000 13910
rect 39045 13632 39361 13633
rect 39045 13568 39051 13632
rect 39115 13568 39131 13632
rect 39195 13568 39211 13632
rect 39275 13568 39291 13632
rect 39355 13568 39361 13632
rect 39045 13567 39361 13568
rect 115243 13632 115559 13633
rect 115243 13568 115249 13632
rect 115313 13568 115329 13632
rect 115393 13568 115409 13632
rect 115473 13568 115489 13632
rect 115553 13568 115559 13632
rect 115243 13567 115559 13568
rect 191441 13632 191757 13633
rect 191441 13568 191447 13632
rect 191511 13568 191527 13632
rect 191591 13568 191607 13632
rect 191671 13568 191687 13632
rect 191751 13568 191757 13632
rect 191441 13567 191757 13568
rect 267639 13632 267955 13633
rect 267639 13568 267645 13632
rect 267709 13568 267725 13632
rect 267789 13568 267805 13632
rect 267869 13568 267885 13632
rect 267949 13568 267955 13632
rect 267639 13567 267955 13568
rect 207105 13562 207171 13565
rect 208025 13562 208091 13565
rect 207105 13560 208091 13562
rect 207105 13504 207110 13560
rect 207166 13504 208030 13560
rect 208086 13504 208091 13560
rect 207105 13502 208091 13504
rect 207105 13499 207171 13502
rect 208025 13499 208091 13502
rect 213269 13426 213335 13429
rect 219801 13426 219867 13429
rect 213269 13424 219867 13426
rect 213269 13368 213274 13424
rect 213330 13368 219806 13424
rect 219862 13368 219867 13424
rect 213269 13366 219867 13368
rect 213269 13363 213335 13366
rect 219801 13363 219867 13366
rect 227069 13426 227135 13429
rect 229185 13426 229251 13429
rect 227069 13424 229251 13426
rect 227069 13368 227074 13424
rect 227130 13368 229190 13424
rect 229246 13368 229251 13424
rect 227069 13366 229251 13368
rect 227069 13363 227135 13366
rect 229185 13363 229251 13366
rect 238109 13426 238175 13429
rect 239489 13426 239555 13429
rect 238109 13424 239555 13426
rect 238109 13368 238114 13424
rect 238170 13368 239494 13424
rect 239550 13368 239555 13424
rect 238109 13366 239555 13368
rect 238109 13363 238175 13366
rect 239489 13363 239555 13366
rect 268929 13426 268995 13429
rect 273161 13426 273227 13429
rect 268929 13424 273227 13426
rect 268929 13368 268934 13424
rect 268990 13368 273166 13424
rect 273222 13368 273227 13424
rect 268929 13366 273227 13368
rect 268929 13363 268995 13366
rect 273161 13363 273227 13366
rect 200849 13290 200915 13293
rect 203425 13290 203491 13293
rect 200849 13288 203491 13290
rect 200849 13232 200854 13288
rect 200910 13232 203430 13288
rect 203486 13232 203491 13288
rect 200849 13230 203491 13232
rect 200849 13227 200915 13230
rect 203425 13227 203491 13230
rect 205541 13290 205607 13293
rect 205725 13290 205791 13293
rect 205541 13288 205791 13290
rect 205541 13232 205546 13288
rect 205602 13232 205730 13288
rect 205786 13232 205791 13288
rect 205541 13230 205791 13232
rect 205541 13227 205607 13230
rect 205725 13227 205791 13230
rect 207197 13290 207263 13293
rect 207933 13290 207999 13293
rect 207197 13288 207999 13290
rect 207197 13232 207202 13288
rect 207258 13232 207938 13288
rect 207994 13232 207999 13288
rect 207197 13230 207999 13232
rect 207197 13227 207263 13230
rect 207933 13227 207999 13230
rect 230381 13290 230447 13293
rect 232129 13290 232195 13293
rect 230381 13288 232195 13290
rect 230381 13232 230386 13288
rect 230442 13232 232134 13288
rect 232190 13232 232195 13288
rect 230381 13230 232195 13232
rect 230381 13227 230447 13230
rect 232129 13227 232195 13230
rect 263409 13290 263475 13293
rect 265525 13290 265591 13293
rect 263409 13288 265591 13290
rect 263409 13232 263414 13288
rect 263470 13232 265530 13288
rect 265586 13232 265591 13288
rect 263409 13230 265591 13232
rect 263409 13227 263475 13230
rect 265525 13227 265591 13230
rect 269021 13290 269087 13293
rect 273253 13290 273319 13293
rect 269021 13288 273319 13290
rect 269021 13232 269026 13288
rect 269082 13232 273258 13288
rect 273314 13232 273319 13288
rect 269021 13230 273319 13232
rect 269021 13227 269087 13230
rect 273253 13227 273319 13230
rect 86953 13154 87019 13157
rect 91829 13154 91895 13157
rect 86953 13152 91895 13154
rect 86953 13096 86958 13152
rect 87014 13096 91834 13152
rect 91890 13096 91895 13152
rect 86953 13094 91895 13096
rect 86953 13091 87019 13094
rect 91829 13091 91895 13094
rect 225413 13154 225479 13157
rect 227069 13154 227135 13157
rect 225413 13152 227135 13154
rect 225413 13096 225418 13152
rect 225474 13096 227074 13152
rect 227130 13096 227135 13152
rect 225413 13094 227135 13096
rect 225413 13091 225479 13094
rect 227069 13091 227135 13094
rect 77144 13088 77460 13089
rect 77144 13024 77150 13088
rect 77214 13024 77230 13088
rect 77294 13024 77310 13088
rect 77374 13024 77390 13088
rect 77454 13024 77460 13088
rect 77144 13023 77460 13024
rect 153342 13088 153658 13089
rect 153342 13024 153348 13088
rect 153412 13024 153428 13088
rect 153492 13024 153508 13088
rect 153572 13024 153588 13088
rect 153652 13024 153658 13088
rect 153342 13023 153658 13024
rect 229540 13088 229856 13089
rect 229540 13024 229546 13088
rect 229610 13024 229626 13088
rect 229690 13024 229706 13088
rect 229770 13024 229786 13088
rect 229850 13024 229856 13088
rect 229540 13023 229856 13024
rect 256601 13018 256667 13021
rect 257981 13018 258047 13021
rect 256601 13016 258047 13018
rect 256601 12960 256606 13016
rect 256662 12960 257986 13016
rect 258042 12960 258047 13016
rect 256601 12958 258047 12960
rect 256601 12955 256667 12958
rect 257981 12955 258047 12958
rect 155033 12882 155099 12885
rect 194593 12882 194659 12885
rect 195789 12882 195855 12885
rect 155033 12880 195855 12882
rect 155033 12824 155038 12880
rect 155094 12824 194598 12880
rect 194654 12824 195794 12880
rect 195850 12824 195855 12880
rect 155033 12822 195855 12824
rect 155033 12819 155099 12822
rect 194593 12819 194659 12822
rect 195789 12819 195855 12822
rect 197353 12882 197419 12885
rect 299473 12882 299539 12885
rect 197353 12880 299539 12882
rect 197353 12824 197358 12880
rect 197414 12824 299478 12880
rect 299534 12824 299539 12880
rect 197353 12822 299539 12824
rect 197353 12819 197419 12822
rect 299473 12819 299539 12822
rect 87781 12746 87847 12749
rect 90725 12746 90791 12749
rect 87781 12744 90791 12746
rect 87781 12688 87786 12744
rect 87842 12688 90730 12744
rect 90786 12688 90791 12744
rect 87781 12686 90791 12688
rect 87781 12683 87847 12686
rect 90725 12683 90791 12686
rect 195053 12746 195119 12749
rect 207841 12746 207907 12749
rect 195053 12744 207907 12746
rect 195053 12688 195058 12744
rect 195114 12688 207846 12744
rect 207902 12688 207907 12744
rect 195053 12686 207907 12688
rect 195053 12683 195119 12686
rect 207841 12683 207907 12686
rect 238293 12746 238359 12749
rect 242157 12746 242223 12749
rect 238293 12744 242223 12746
rect 238293 12688 238298 12744
rect 238354 12688 242162 12744
rect 242218 12688 242223 12744
rect 238293 12686 242223 12688
rect 238293 12683 238359 12686
rect 242157 12683 242223 12686
rect 262305 12746 262371 12749
rect 263501 12746 263567 12749
rect 262305 12744 263567 12746
rect 262305 12688 262310 12744
rect 262366 12688 263506 12744
rect 263562 12688 263567 12744
rect 262305 12686 263567 12688
rect 262305 12683 262371 12686
rect 263501 12683 263567 12686
rect 264329 12746 264395 12749
rect 267089 12746 267155 12749
rect 264329 12744 267155 12746
rect 264329 12688 264334 12744
rect 264390 12688 267094 12744
rect 267150 12688 267155 12744
rect 264329 12686 267155 12688
rect 264329 12683 264395 12686
rect 267089 12683 267155 12686
rect 267641 12746 267707 12749
rect 268101 12746 268167 12749
rect 267641 12744 268167 12746
rect 267641 12688 267646 12744
rect 267702 12688 268106 12744
rect 268162 12688 268167 12744
rect 267641 12686 268167 12688
rect 267641 12683 267707 12686
rect 268101 12683 268167 12686
rect 157885 12610 157951 12613
rect 160277 12610 160343 12613
rect 157885 12608 160343 12610
rect 157885 12552 157890 12608
rect 157946 12552 160282 12608
rect 160338 12552 160343 12608
rect 157885 12550 160343 12552
rect 157885 12547 157951 12550
rect 160277 12547 160343 12550
rect 191833 12610 191899 12613
rect 192201 12610 192267 12613
rect 191833 12608 192267 12610
rect 191833 12552 191838 12608
rect 191894 12552 192206 12608
rect 192262 12552 192267 12608
rect 191833 12550 192267 12552
rect 191833 12547 191899 12550
rect 192201 12547 192267 12550
rect 200389 12610 200455 12613
rect 205265 12610 205331 12613
rect 200389 12608 205331 12610
rect 200389 12552 200394 12608
rect 200450 12552 205270 12608
rect 205326 12552 205331 12608
rect 200389 12550 205331 12552
rect 200389 12547 200455 12550
rect 205265 12547 205331 12550
rect 251909 12610 251975 12613
rect 257061 12610 257127 12613
rect 251909 12608 257127 12610
rect 251909 12552 251914 12608
rect 251970 12552 257066 12608
rect 257122 12552 257127 12608
rect 251909 12550 257127 12552
rect 251909 12547 251975 12550
rect 257061 12547 257127 12550
rect 39045 12544 39361 12545
rect 39045 12480 39051 12544
rect 39115 12480 39131 12544
rect 39195 12480 39211 12544
rect 39275 12480 39291 12544
rect 39355 12480 39361 12544
rect 39045 12479 39361 12480
rect 115243 12544 115559 12545
rect 115243 12480 115249 12544
rect 115313 12480 115329 12544
rect 115393 12480 115409 12544
rect 115473 12480 115489 12544
rect 115553 12480 115559 12544
rect 115243 12479 115559 12480
rect 191441 12544 191757 12545
rect 191441 12480 191447 12544
rect 191511 12480 191527 12544
rect 191591 12480 191607 12544
rect 191671 12480 191687 12544
rect 191751 12480 191757 12544
rect 191441 12479 191757 12480
rect 267639 12544 267955 12545
rect 267639 12480 267645 12544
rect 267709 12480 267725 12544
rect 267789 12480 267805 12544
rect 267869 12480 267885 12544
rect 267949 12480 267955 12544
rect 267639 12479 267955 12480
rect 251817 12474 251883 12477
rect 257153 12474 257219 12477
rect 251817 12472 257219 12474
rect 251817 12416 251822 12472
rect 251878 12416 257158 12472
rect 257214 12416 257219 12472
rect 251817 12414 257219 12416
rect 251817 12411 251883 12414
rect 257153 12411 257219 12414
rect 88149 12338 88215 12341
rect 89897 12338 89963 12341
rect 88149 12336 89963 12338
rect 88149 12280 88154 12336
rect 88210 12280 89902 12336
rect 89958 12280 89963 12336
rect 88149 12278 89963 12280
rect 88149 12275 88215 12278
rect 89897 12275 89963 12278
rect 163589 12338 163655 12341
rect 193029 12338 193095 12341
rect 163589 12336 193095 12338
rect 163589 12280 163594 12336
rect 163650 12280 193034 12336
rect 193090 12280 193095 12336
rect 163589 12278 193095 12280
rect 163589 12275 163655 12278
rect 193029 12275 193095 12278
rect 29361 12202 29427 12205
rect 30741 12202 30807 12205
rect 31385 12202 31451 12205
rect 29361 12200 31451 12202
rect 29361 12144 29366 12200
rect 29422 12144 30746 12200
rect 30802 12144 31390 12200
rect 31446 12144 31451 12200
rect 29361 12142 31451 12144
rect 29361 12139 29427 12142
rect 30741 12139 30807 12142
rect 31385 12139 31451 12142
rect 40585 12202 40651 12205
rect 42425 12202 42491 12205
rect 40585 12200 42491 12202
rect 40585 12144 40590 12200
rect 40646 12144 42430 12200
rect 42486 12144 42491 12200
rect 40585 12142 42491 12144
rect 40585 12139 40651 12142
rect 42425 12139 42491 12142
rect 77144 12000 77460 12001
rect 77144 11936 77150 12000
rect 77214 11936 77230 12000
rect 77294 11936 77310 12000
rect 77374 11936 77390 12000
rect 77454 11936 77460 12000
rect 77144 11935 77460 11936
rect 153342 12000 153658 12001
rect 153342 11936 153348 12000
rect 153412 11936 153428 12000
rect 153492 11936 153508 12000
rect 153572 11936 153588 12000
rect 153652 11936 153658 12000
rect 153342 11935 153658 11936
rect 229540 12000 229856 12001
rect 229540 11936 229546 12000
rect 229610 11936 229626 12000
rect 229690 11936 229706 12000
rect 229770 11936 229786 12000
rect 229850 11936 229856 12000
rect 229540 11935 229856 11936
rect 189625 11794 189691 11797
rect 193029 11794 193095 11797
rect 189625 11792 193095 11794
rect 189625 11736 189630 11792
rect 189686 11736 193034 11792
rect 193090 11736 193095 11792
rect 189625 11734 193095 11736
rect 189625 11731 189691 11734
rect 193029 11731 193095 11734
rect 39045 11456 39361 11457
rect 39045 11392 39051 11456
rect 39115 11392 39131 11456
rect 39195 11392 39211 11456
rect 39275 11392 39291 11456
rect 39355 11392 39361 11456
rect 39045 11391 39361 11392
rect 115243 11456 115559 11457
rect 115243 11392 115249 11456
rect 115313 11392 115329 11456
rect 115393 11392 115409 11456
rect 115473 11392 115489 11456
rect 115553 11392 115559 11456
rect 115243 11391 115559 11392
rect 191441 11456 191757 11457
rect 191441 11392 191447 11456
rect 191511 11392 191527 11456
rect 191591 11392 191607 11456
rect 191671 11392 191687 11456
rect 191751 11392 191757 11456
rect 191441 11391 191757 11392
rect 267639 11456 267955 11457
rect 267639 11392 267645 11456
rect 267709 11392 267725 11456
rect 267789 11392 267805 11456
rect 267869 11392 267885 11456
rect 267949 11392 267955 11456
rect 267639 11391 267955 11392
rect 77144 10912 77460 10913
rect 77144 10848 77150 10912
rect 77214 10848 77230 10912
rect 77294 10848 77310 10912
rect 77374 10848 77390 10912
rect 77454 10848 77460 10912
rect 77144 10847 77460 10848
rect 153342 10912 153658 10913
rect 153342 10848 153348 10912
rect 153412 10848 153428 10912
rect 153492 10848 153508 10912
rect 153572 10848 153588 10912
rect 153652 10848 153658 10912
rect 153342 10847 153658 10848
rect 229540 10912 229856 10913
rect 229540 10848 229546 10912
rect 229610 10848 229626 10912
rect 229690 10848 229706 10912
rect 229770 10848 229786 10912
rect 229850 10848 229856 10912
rect 229540 10847 229856 10848
rect 39045 10368 39361 10369
rect 39045 10304 39051 10368
rect 39115 10304 39131 10368
rect 39195 10304 39211 10368
rect 39275 10304 39291 10368
rect 39355 10304 39361 10368
rect 39045 10303 39361 10304
rect 115243 10368 115559 10369
rect 115243 10304 115249 10368
rect 115313 10304 115329 10368
rect 115393 10304 115409 10368
rect 115473 10304 115489 10368
rect 115553 10304 115559 10368
rect 115243 10303 115559 10304
rect 191441 10368 191757 10369
rect 191441 10304 191447 10368
rect 191511 10304 191527 10368
rect 191591 10304 191607 10368
rect 191671 10304 191687 10368
rect 191751 10304 191757 10368
rect 191441 10303 191757 10304
rect 267639 10368 267955 10369
rect 267639 10304 267645 10368
rect 267709 10304 267725 10368
rect 267789 10304 267805 10368
rect 267869 10304 267885 10368
rect 267949 10304 267955 10368
rect 267639 10303 267955 10304
rect 304441 10026 304507 10029
rect 306200 10026 307000 10056
rect 304441 10024 307000 10026
rect 304441 9968 304446 10024
rect 304502 9968 307000 10024
rect 304441 9966 307000 9968
rect 304441 9963 304507 9966
rect 306200 9936 307000 9966
rect 77144 9824 77460 9825
rect 77144 9760 77150 9824
rect 77214 9760 77230 9824
rect 77294 9760 77310 9824
rect 77374 9760 77390 9824
rect 77454 9760 77460 9824
rect 77144 9759 77460 9760
rect 153342 9824 153658 9825
rect 153342 9760 153348 9824
rect 153412 9760 153428 9824
rect 153492 9760 153508 9824
rect 153572 9760 153588 9824
rect 153652 9760 153658 9824
rect 153342 9759 153658 9760
rect 229540 9824 229856 9825
rect 229540 9760 229546 9824
rect 229610 9760 229626 9824
rect 229690 9760 229706 9824
rect 229770 9760 229786 9824
rect 229850 9760 229856 9824
rect 229540 9759 229856 9760
rect 39045 9280 39361 9281
rect 39045 9216 39051 9280
rect 39115 9216 39131 9280
rect 39195 9216 39211 9280
rect 39275 9216 39291 9280
rect 39355 9216 39361 9280
rect 39045 9215 39361 9216
rect 115243 9280 115559 9281
rect 115243 9216 115249 9280
rect 115313 9216 115329 9280
rect 115393 9216 115409 9280
rect 115473 9216 115489 9280
rect 115553 9216 115559 9280
rect 115243 9215 115559 9216
rect 191441 9280 191757 9281
rect 191441 9216 191447 9280
rect 191511 9216 191527 9280
rect 191591 9216 191607 9280
rect 191671 9216 191687 9280
rect 191751 9216 191757 9280
rect 191441 9215 191757 9216
rect 267639 9280 267955 9281
rect 267639 9216 267645 9280
rect 267709 9216 267725 9280
rect 267789 9216 267805 9280
rect 267869 9216 267885 9280
rect 267949 9216 267955 9280
rect 267639 9215 267955 9216
rect 77144 8736 77460 8737
rect 77144 8672 77150 8736
rect 77214 8672 77230 8736
rect 77294 8672 77310 8736
rect 77374 8672 77390 8736
rect 77454 8672 77460 8736
rect 77144 8671 77460 8672
rect 153342 8736 153658 8737
rect 153342 8672 153348 8736
rect 153412 8672 153428 8736
rect 153492 8672 153508 8736
rect 153572 8672 153588 8736
rect 153652 8672 153658 8736
rect 153342 8671 153658 8672
rect 229540 8736 229856 8737
rect 229540 8672 229546 8736
rect 229610 8672 229626 8736
rect 229690 8672 229706 8736
rect 229770 8672 229786 8736
rect 229850 8672 229856 8736
rect 229540 8671 229856 8672
rect 39045 8192 39361 8193
rect 0 8122 800 8152
rect 39045 8128 39051 8192
rect 39115 8128 39131 8192
rect 39195 8128 39211 8192
rect 39275 8128 39291 8192
rect 39355 8128 39361 8192
rect 39045 8127 39361 8128
rect 115243 8192 115559 8193
rect 115243 8128 115249 8192
rect 115313 8128 115329 8192
rect 115393 8128 115409 8192
rect 115473 8128 115489 8192
rect 115553 8128 115559 8192
rect 115243 8127 115559 8128
rect 191441 8192 191757 8193
rect 191441 8128 191447 8192
rect 191511 8128 191527 8192
rect 191591 8128 191607 8192
rect 191671 8128 191687 8192
rect 191751 8128 191757 8192
rect 191441 8127 191757 8128
rect 267639 8192 267955 8193
rect 267639 8128 267645 8192
rect 267709 8128 267725 8192
rect 267789 8128 267805 8192
rect 267869 8128 267885 8192
rect 267949 8128 267955 8192
rect 267639 8127 267955 8128
rect 1393 8122 1459 8125
rect 0 8120 1459 8122
rect 0 8064 1398 8120
rect 1454 8064 1459 8120
rect 0 8062 1459 8064
rect 0 8032 800 8062
rect 1393 8059 1459 8062
rect 77144 7648 77460 7649
rect 77144 7584 77150 7648
rect 77214 7584 77230 7648
rect 77294 7584 77310 7648
rect 77374 7584 77390 7648
rect 77454 7584 77460 7648
rect 77144 7583 77460 7584
rect 153342 7648 153658 7649
rect 153342 7584 153348 7648
rect 153412 7584 153428 7648
rect 153492 7584 153508 7648
rect 153572 7584 153588 7648
rect 153652 7584 153658 7648
rect 153342 7583 153658 7584
rect 229540 7648 229856 7649
rect 229540 7584 229546 7648
rect 229610 7584 229626 7648
rect 229690 7584 229706 7648
rect 229770 7584 229786 7648
rect 229850 7584 229856 7648
rect 229540 7583 229856 7584
rect 39045 7104 39361 7105
rect 39045 7040 39051 7104
rect 39115 7040 39131 7104
rect 39195 7040 39211 7104
rect 39275 7040 39291 7104
rect 39355 7040 39361 7104
rect 39045 7039 39361 7040
rect 115243 7104 115559 7105
rect 115243 7040 115249 7104
rect 115313 7040 115329 7104
rect 115393 7040 115409 7104
rect 115473 7040 115489 7104
rect 115553 7040 115559 7104
rect 115243 7039 115559 7040
rect 191441 7104 191757 7105
rect 191441 7040 191447 7104
rect 191511 7040 191527 7104
rect 191591 7040 191607 7104
rect 191671 7040 191687 7104
rect 191751 7040 191757 7104
rect 191441 7039 191757 7040
rect 267639 7104 267955 7105
rect 267639 7040 267645 7104
rect 267709 7040 267725 7104
rect 267789 7040 267805 7104
rect 267869 7040 267885 7104
rect 267949 7040 267955 7104
rect 267639 7039 267955 7040
rect 77144 6560 77460 6561
rect 77144 6496 77150 6560
rect 77214 6496 77230 6560
rect 77294 6496 77310 6560
rect 77374 6496 77390 6560
rect 77454 6496 77460 6560
rect 77144 6495 77460 6496
rect 153342 6560 153658 6561
rect 153342 6496 153348 6560
rect 153412 6496 153428 6560
rect 153492 6496 153508 6560
rect 153572 6496 153588 6560
rect 153652 6496 153658 6560
rect 153342 6495 153658 6496
rect 229540 6560 229856 6561
rect 229540 6496 229546 6560
rect 229610 6496 229626 6560
rect 229690 6496 229706 6560
rect 229770 6496 229786 6560
rect 229850 6496 229856 6560
rect 229540 6495 229856 6496
rect 39045 6016 39361 6017
rect 39045 5952 39051 6016
rect 39115 5952 39131 6016
rect 39195 5952 39211 6016
rect 39275 5952 39291 6016
rect 39355 5952 39361 6016
rect 39045 5951 39361 5952
rect 115243 6016 115559 6017
rect 115243 5952 115249 6016
rect 115313 5952 115329 6016
rect 115393 5952 115409 6016
rect 115473 5952 115489 6016
rect 115553 5952 115559 6016
rect 115243 5951 115559 5952
rect 191441 6016 191757 6017
rect 191441 5952 191447 6016
rect 191511 5952 191527 6016
rect 191591 5952 191607 6016
rect 191671 5952 191687 6016
rect 191751 5952 191757 6016
rect 191441 5951 191757 5952
rect 267639 6016 267955 6017
rect 267639 5952 267645 6016
rect 267709 5952 267725 6016
rect 267789 5952 267805 6016
rect 267869 5952 267885 6016
rect 267949 5952 267955 6016
rect 267639 5951 267955 5952
rect 303981 5946 304047 5949
rect 306200 5946 307000 5976
rect 303981 5944 307000 5946
rect 303981 5888 303986 5944
rect 304042 5888 307000 5944
rect 303981 5886 307000 5888
rect 303981 5883 304047 5886
rect 306200 5856 307000 5886
rect 77144 5472 77460 5473
rect 77144 5408 77150 5472
rect 77214 5408 77230 5472
rect 77294 5408 77310 5472
rect 77374 5408 77390 5472
rect 77454 5408 77460 5472
rect 77144 5407 77460 5408
rect 153342 5472 153658 5473
rect 153342 5408 153348 5472
rect 153412 5408 153428 5472
rect 153492 5408 153508 5472
rect 153572 5408 153588 5472
rect 153652 5408 153658 5472
rect 153342 5407 153658 5408
rect 229540 5472 229856 5473
rect 229540 5408 229546 5472
rect 229610 5408 229626 5472
rect 229690 5408 229706 5472
rect 229770 5408 229786 5472
rect 229850 5408 229856 5472
rect 229540 5407 229856 5408
rect 39045 4928 39361 4929
rect 39045 4864 39051 4928
rect 39115 4864 39131 4928
rect 39195 4864 39211 4928
rect 39275 4864 39291 4928
rect 39355 4864 39361 4928
rect 39045 4863 39361 4864
rect 115243 4928 115559 4929
rect 115243 4864 115249 4928
rect 115313 4864 115329 4928
rect 115393 4864 115409 4928
rect 115473 4864 115489 4928
rect 115553 4864 115559 4928
rect 115243 4863 115559 4864
rect 191441 4928 191757 4929
rect 191441 4864 191447 4928
rect 191511 4864 191527 4928
rect 191591 4864 191607 4928
rect 191671 4864 191687 4928
rect 191751 4864 191757 4928
rect 191441 4863 191757 4864
rect 267639 4928 267955 4929
rect 267639 4864 267645 4928
rect 267709 4864 267725 4928
rect 267789 4864 267805 4928
rect 267869 4864 267885 4928
rect 267949 4864 267955 4928
rect 267639 4863 267955 4864
rect 77144 4384 77460 4385
rect 77144 4320 77150 4384
rect 77214 4320 77230 4384
rect 77294 4320 77310 4384
rect 77374 4320 77390 4384
rect 77454 4320 77460 4384
rect 77144 4319 77460 4320
rect 153342 4384 153658 4385
rect 153342 4320 153348 4384
rect 153412 4320 153428 4384
rect 153492 4320 153508 4384
rect 153572 4320 153588 4384
rect 153652 4320 153658 4384
rect 153342 4319 153658 4320
rect 229540 4384 229856 4385
rect 229540 4320 229546 4384
rect 229610 4320 229626 4384
rect 229690 4320 229706 4384
rect 229770 4320 229786 4384
rect 229850 4320 229856 4384
rect 229540 4319 229856 4320
rect 39045 3840 39361 3841
rect 39045 3776 39051 3840
rect 39115 3776 39131 3840
rect 39195 3776 39211 3840
rect 39275 3776 39291 3840
rect 39355 3776 39361 3840
rect 39045 3775 39361 3776
rect 115243 3840 115559 3841
rect 115243 3776 115249 3840
rect 115313 3776 115329 3840
rect 115393 3776 115409 3840
rect 115473 3776 115489 3840
rect 115553 3776 115559 3840
rect 115243 3775 115559 3776
rect 191441 3840 191757 3841
rect 191441 3776 191447 3840
rect 191511 3776 191527 3840
rect 191591 3776 191607 3840
rect 191671 3776 191687 3840
rect 191751 3776 191757 3840
rect 191441 3775 191757 3776
rect 267639 3840 267955 3841
rect 267639 3776 267645 3840
rect 267709 3776 267725 3840
rect 267789 3776 267805 3840
rect 267869 3776 267885 3840
rect 267949 3776 267955 3840
rect 267639 3775 267955 3776
rect 77144 3296 77460 3297
rect 77144 3232 77150 3296
rect 77214 3232 77230 3296
rect 77294 3232 77310 3296
rect 77374 3232 77390 3296
rect 77454 3232 77460 3296
rect 77144 3231 77460 3232
rect 153342 3296 153658 3297
rect 153342 3232 153348 3296
rect 153412 3232 153428 3296
rect 153492 3232 153508 3296
rect 153572 3232 153588 3296
rect 153652 3232 153658 3296
rect 153342 3231 153658 3232
rect 229540 3296 229856 3297
rect 229540 3232 229546 3296
rect 229610 3232 229626 3296
rect 229690 3232 229706 3296
rect 229770 3232 229786 3296
rect 229850 3232 229856 3296
rect 229540 3231 229856 3232
rect 39045 2752 39361 2753
rect 39045 2688 39051 2752
rect 39115 2688 39131 2752
rect 39195 2688 39211 2752
rect 39275 2688 39291 2752
rect 39355 2688 39361 2752
rect 39045 2687 39361 2688
rect 115243 2752 115559 2753
rect 115243 2688 115249 2752
rect 115313 2688 115329 2752
rect 115393 2688 115409 2752
rect 115473 2688 115489 2752
rect 115553 2688 115559 2752
rect 115243 2687 115559 2688
rect 191441 2752 191757 2753
rect 191441 2688 191447 2752
rect 191511 2688 191527 2752
rect 191591 2688 191607 2752
rect 191671 2688 191687 2752
rect 191751 2688 191757 2752
rect 191441 2687 191757 2688
rect 267639 2752 267955 2753
rect 267639 2688 267645 2752
rect 267709 2688 267725 2752
rect 267789 2688 267805 2752
rect 267869 2688 267885 2752
rect 267949 2688 267955 2752
rect 267639 2687 267955 2688
rect 77144 2208 77460 2209
rect 77144 2144 77150 2208
rect 77214 2144 77230 2208
rect 77294 2144 77310 2208
rect 77374 2144 77390 2208
rect 77454 2144 77460 2208
rect 77144 2143 77460 2144
rect 153342 2208 153658 2209
rect 153342 2144 153348 2208
rect 153412 2144 153428 2208
rect 153492 2144 153508 2208
rect 153572 2144 153588 2208
rect 153652 2144 153658 2208
rect 153342 2143 153658 2144
rect 229540 2208 229856 2209
rect 229540 2144 229546 2208
rect 229610 2144 229626 2208
rect 229690 2144 229706 2208
rect 229770 2144 229786 2208
rect 229850 2144 229856 2208
rect 229540 2143 229856 2144
rect 302233 2002 302299 2005
rect 306200 2002 307000 2032
rect 302233 2000 307000 2002
rect 302233 1944 302238 2000
rect 302294 1944 307000 2000
rect 302233 1942 307000 1944
rect 302233 1939 302299 1942
rect 306200 1912 307000 1942
<< via3 >>
rect 39051 13628 39115 13632
rect 39051 13572 39055 13628
rect 39055 13572 39111 13628
rect 39111 13572 39115 13628
rect 39051 13568 39115 13572
rect 39131 13628 39195 13632
rect 39131 13572 39135 13628
rect 39135 13572 39191 13628
rect 39191 13572 39195 13628
rect 39131 13568 39195 13572
rect 39211 13628 39275 13632
rect 39211 13572 39215 13628
rect 39215 13572 39271 13628
rect 39271 13572 39275 13628
rect 39211 13568 39275 13572
rect 39291 13628 39355 13632
rect 39291 13572 39295 13628
rect 39295 13572 39351 13628
rect 39351 13572 39355 13628
rect 39291 13568 39355 13572
rect 115249 13628 115313 13632
rect 115249 13572 115253 13628
rect 115253 13572 115309 13628
rect 115309 13572 115313 13628
rect 115249 13568 115313 13572
rect 115329 13628 115393 13632
rect 115329 13572 115333 13628
rect 115333 13572 115389 13628
rect 115389 13572 115393 13628
rect 115329 13568 115393 13572
rect 115409 13628 115473 13632
rect 115409 13572 115413 13628
rect 115413 13572 115469 13628
rect 115469 13572 115473 13628
rect 115409 13568 115473 13572
rect 115489 13628 115553 13632
rect 115489 13572 115493 13628
rect 115493 13572 115549 13628
rect 115549 13572 115553 13628
rect 115489 13568 115553 13572
rect 191447 13628 191511 13632
rect 191447 13572 191451 13628
rect 191451 13572 191507 13628
rect 191507 13572 191511 13628
rect 191447 13568 191511 13572
rect 191527 13628 191591 13632
rect 191527 13572 191531 13628
rect 191531 13572 191587 13628
rect 191587 13572 191591 13628
rect 191527 13568 191591 13572
rect 191607 13628 191671 13632
rect 191607 13572 191611 13628
rect 191611 13572 191667 13628
rect 191667 13572 191671 13628
rect 191607 13568 191671 13572
rect 191687 13628 191751 13632
rect 191687 13572 191691 13628
rect 191691 13572 191747 13628
rect 191747 13572 191751 13628
rect 191687 13568 191751 13572
rect 267645 13628 267709 13632
rect 267645 13572 267649 13628
rect 267649 13572 267705 13628
rect 267705 13572 267709 13628
rect 267645 13568 267709 13572
rect 267725 13628 267789 13632
rect 267725 13572 267729 13628
rect 267729 13572 267785 13628
rect 267785 13572 267789 13628
rect 267725 13568 267789 13572
rect 267805 13628 267869 13632
rect 267805 13572 267809 13628
rect 267809 13572 267865 13628
rect 267865 13572 267869 13628
rect 267805 13568 267869 13572
rect 267885 13628 267949 13632
rect 267885 13572 267889 13628
rect 267889 13572 267945 13628
rect 267945 13572 267949 13628
rect 267885 13568 267949 13572
rect 77150 13084 77214 13088
rect 77150 13028 77154 13084
rect 77154 13028 77210 13084
rect 77210 13028 77214 13084
rect 77150 13024 77214 13028
rect 77230 13084 77294 13088
rect 77230 13028 77234 13084
rect 77234 13028 77290 13084
rect 77290 13028 77294 13084
rect 77230 13024 77294 13028
rect 77310 13084 77374 13088
rect 77310 13028 77314 13084
rect 77314 13028 77370 13084
rect 77370 13028 77374 13084
rect 77310 13024 77374 13028
rect 77390 13084 77454 13088
rect 77390 13028 77394 13084
rect 77394 13028 77450 13084
rect 77450 13028 77454 13084
rect 77390 13024 77454 13028
rect 153348 13084 153412 13088
rect 153348 13028 153352 13084
rect 153352 13028 153408 13084
rect 153408 13028 153412 13084
rect 153348 13024 153412 13028
rect 153428 13084 153492 13088
rect 153428 13028 153432 13084
rect 153432 13028 153488 13084
rect 153488 13028 153492 13084
rect 153428 13024 153492 13028
rect 153508 13084 153572 13088
rect 153508 13028 153512 13084
rect 153512 13028 153568 13084
rect 153568 13028 153572 13084
rect 153508 13024 153572 13028
rect 153588 13084 153652 13088
rect 153588 13028 153592 13084
rect 153592 13028 153648 13084
rect 153648 13028 153652 13084
rect 153588 13024 153652 13028
rect 229546 13084 229610 13088
rect 229546 13028 229550 13084
rect 229550 13028 229606 13084
rect 229606 13028 229610 13084
rect 229546 13024 229610 13028
rect 229626 13084 229690 13088
rect 229626 13028 229630 13084
rect 229630 13028 229686 13084
rect 229686 13028 229690 13084
rect 229626 13024 229690 13028
rect 229706 13084 229770 13088
rect 229706 13028 229710 13084
rect 229710 13028 229766 13084
rect 229766 13028 229770 13084
rect 229706 13024 229770 13028
rect 229786 13084 229850 13088
rect 229786 13028 229790 13084
rect 229790 13028 229846 13084
rect 229846 13028 229850 13084
rect 229786 13024 229850 13028
rect 39051 12540 39115 12544
rect 39051 12484 39055 12540
rect 39055 12484 39111 12540
rect 39111 12484 39115 12540
rect 39051 12480 39115 12484
rect 39131 12540 39195 12544
rect 39131 12484 39135 12540
rect 39135 12484 39191 12540
rect 39191 12484 39195 12540
rect 39131 12480 39195 12484
rect 39211 12540 39275 12544
rect 39211 12484 39215 12540
rect 39215 12484 39271 12540
rect 39271 12484 39275 12540
rect 39211 12480 39275 12484
rect 39291 12540 39355 12544
rect 39291 12484 39295 12540
rect 39295 12484 39351 12540
rect 39351 12484 39355 12540
rect 39291 12480 39355 12484
rect 115249 12540 115313 12544
rect 115249 12484 115253 12540
rect 115253 12484 115309 12540
rect 115309 12484 115313 12540
rect 115249 12480 115313 12484
rect 115329 12540 115393 12544
rect 115329 12484 115333 12540
rect 115333 12484 115389 12540
rect 115389 12484 115393 12540
rect 115329 12480 115393 12484
rect 115409 12540 115473 12544
rect 115409 12484 115413 12540
rect 115413 12484 115469 12540
rect 115469 12484 115473 12540
rect 115409 12480 115473 12484
rect 115489 12540 115553 12544
rect 115489 12484 115493 12540
rect 115493 12484 115549 12540
rect 115549 12484 115553 12540
rect 115489 12480 115553 12484
rect 191447 12540 191511 12544
rect 191447 12484 191451 12540
rect 191451 12484 191507 12540
rect 191507 12484 191511 12540
rect 191447 12480 191511 12484
rect 191527 12540 191591 12544
rect 191527 12484 191531 12540
rect 191531 12484 191587 12540
rect 191587 12484 191591 12540
rect 191527 12480 191591 12484
rect 191607 12540 191671 12544
rect 191607 12484 191611 12540
rect 191611 12484 191667 12540
rect 191667 12484 191671 12540
rect 191607 12480 191671 12484
rect 191687 12540 191751 12544
rect 191687 12484 191691 12540
rect 191691 12484 191747 12540
rect 191747 12484 191751 12540
rect 191687 12480 191751 12484
rect 267645 12540 267709 12544
rect 267645 12484 267649 12540
rect 267649 12484 267705 12540
rect 267705 12484 267709 12540
rect 267645 12480 267709 12484
rect 267725 12540 267789 12544
rect 267725 12484 267729 12540
rect 267729 12484 267785 12540
rect 267785 12484 267789 12540
rect 267725 12480 267789 12484
rect 267805 12540 267869 12544
rect 267805 12484 267809 12540
rect 267809 12484 267865 12540
rect 267865 12484 267869 12540
rect 267805 12480 267869 12484
rect 267885 12540 267949 12544
rect 267885 12484 267889 12540
rect 267889 12484 267945 12540
rect 267945 12484 267949 12540
rect 267885 12480 267949 12484
rect 77150 11996 77214 12000
rect 77150 11940 77154 11996
rect 77154 11940 77210 11996
rect 77210 11940 77214 11996
rect 77150 11936 77214 11940
rect 77230 11996 77294 12000
rect 77230 11940 77234 11996
rect 77234 11940 77290 11996
rect 77290 11940 77294 11996
rect 77230 11936 77294 11940
rect 77310 11996 77374 12000
rect 77310 11940 77314 11996
rect 77314 11940 77370 11996
rect 77370 11940 77374 11996
rect 77310 11936 77374 11940
rect 77390 11996 77454 12000
rect 77390 11940 77394 11996
rect 77394 11940 77450 11996
rect 77450 11940 77454 11996
rect 77390 11936 77454 11940
rect 153348 11996 153412 12000
rect 153348 11940 153352 11996
rect 153352 11940 153408 11996
rect 153408 11940 153412 11996
rect 153348 11936 153412 11940
rect 153428 11996 153492 12000
rect 153428 11940 153432 11996
rect 153432 11940 153488 11996
rect 153488 11940 153492 11996
rect 153428 11936 153492 11940
rect 153508 11996 153572 12000
rect 153508 11940 153512 11996
rect 153512 11940 153568 11996
rect 153568 11940 153572 11996
rect 153508 11936 153572 11940
rect 153588 11996 153652 12000
rect 153588 11940 153592 11996
rect 153592 11940 153648 11996
rect 153648 11940 153652 11996
rect 153588 11936 153652 11940
rect 229546 11996 229610 12000
rect 229546 11940 229550 11996
rect 229550 11940 229606 11996
rect 229606 11940 229610 11996
rect 229546 11936 229610 11940
rect 229626 11996 229690 12000
rect 229626 11940 229630 11996
rect 229630 11940 229686 11996
rect 229686 11940 229690 11996
rect 229626 11936 229690 11940
rect 229706 11996 229770 12000
rect 229706 11940 229710 11996
rect 229710 11940 229766 11996
rect 229766 11940 229770 11996
rect 229706 11936 229770 11940
rect 229786 11996 229850 12000
rect 229786 11940 229790 11996
rect 229790 11940 229846 11996
rect 229846 11940 229850 11996
rect 229786 11936 229850 11940
rect 39051 11452 39115 11456
rect 39051 11396 39055 11452
rect 39055 11396 39111 11452
rect 39111 11396 39115 11452
rect 39051 11392 39115 11396
rect 39131 11452 39195 11456
rect 39131 11396 39135 11452
rect 39135 11396 39191 11452
rect 39191 11396 39195 11452
rect 39131 11392 39195 11396
rect 39211 11452 39275 11456
rect 39211 11396 39215 11452
rect 39215 11396 39271 11452
rect 39271 11396 39275 11452
rect 39211 11392 39275 11396
rect 39291 11452 39355 11456
rect 39291 11396 39295 11452
rect 39295 11396 39351 11452
rect 39351 11396 39355 11452
rect 39291 11392 39355 11396
rect 115249 11452 115313 11456
rect 115249 11396 115253 11452
rect 115253 11396 115309 11452
rect 115309 11396 115313 11452
rect 115249 11392 115313 11396
rect 115329 11452 115393 11456
rect 115329 11396 115333 11452
rect 115333 11396 115389 11452
rect 115389 11396 115393 11452
rect 115329 11392 115393 11396
rect 115409 11452 115473 11456
rect 115409 11396 115413 11452
rect 115413 11396 115469 11452
rect 115469 11396 115473 11452
rect 115409 11392 115473 11396
rect 115489 11452 115553 11456
rect 115489 11396 115493 11452
rect 115493 11396 115549 11452
rect 115549 11396 115553 11452
rect 115489 11392 115553 11396
rect 191447 11452 191511 11456
rect 191447 11396 191451 11452
rect 191451 11396 191507 11452
rect 191507 11396 191511 11452
rect 191447 11392 191511 11396
rect 191527 11452 191591 11456
rect 191527 11396 191531 11452
rect 191531 11396 191587 11452
rect 191587 11396 191591 11452
rect 191527 11392 191591 11396
rect 191607 11452 191671 11456
rect 191607 11396 191611 11452
rect 191611 11396 191667 11452
rect 191667 11396 191671 11452
rect 191607 11392 191671 11396
rect 191687 11452 191751 11456
rect 191687 11396 191691 11452
rect 191691 11396 191747 11452
rect 191747 11396 191751 11452
rect 191687 11392 191751 11396
rect 267645 11452 267709 11456
rect 267645 11396 267649 11452
rect 267649 11396 267705 11452
rect 267705 11396 267709 11452
rect 267645 11392 267709 11396
rect 267725 11452 267789 11456
rect 267725 11396 267729 11452
rect 267729 11396 267785 11452
rect 267785 11396 267789 11452
rect 267725 11392 267789 11396
rect 267805 11452 267869 11456
rect 267805 11396 267809 11452
rect 267809 11396 267865 11452
rect 267865 11396 267869 11452
rect 267805 11392 267869 11396
rect 267885 11452 267949 11456
rect 267885 11396 267889 11452
rect 267889 11396 267945 11452
rect 267945 11396 267949 11452
rect 267885 11392 267949 11396
rect 77150 10908 77214 10912
rect 77150 10852 77154 10908
rect 77154 10852 77210 10908
rect 77210 10852 77214 10908
rect 77150 10848 77214 10852
rect 77230 10908 77294 10912
rect 77230 10852 77234 10908
rect 77234 10852 77290 10908
rect 77290 10852 77294 10908
rect 77230 10848 77294 10852
rect 77310 10908 77374 10912
rect 77310 10852 77314 10908
rect 77314 10852 77370 10908
rect 77370 10852 77374 10908
rect 77310 10848 77374 10852
rect 77390 10908 77454 10912
rect 77390 10852 77394 10908
rect 77394 10852 77450 10908
rect 77450 10852 77454 10908
rect 77390 10848 77454 10852
rect 153348 10908 153412 10912
rect 153348 10852 153352 10908
rect 153352 10852 153408 10908
rect 153408 10852 153412 10908
rect 153348 10848 153412 10852
rect 153428 10908 153492 10912
rect 153428 10852 153432 10908
rect 153432 10852 153488 10908
rect 153488 10852 153492 10908
rect 153428 10848 153492 10852
rect 153508 10908 153572 10912
rect 153508 10852 153512 10908
rect 153512 10852 153568 10908
rect 153568 10852 153572 10908
rect 153508 10848 153572 10852
rect 153588 10908 153652 10912
rect 153588 10852 153592 10908
rect 153592 10852 153648 10908
rect 153648 10852 153652 10908
rect 153588 10848 153652 10852
rect 229546 10908 229610 10912
rect 229546 10852 229550 10908
rect 229550 10852 229606 10908
rect 229606 10852 229610 10908
rect 229546 10848 229610 10852
rect 229626 10908 229690 10912
rect 229626 10852 229630 10908
rect 229630 10852 229686 10908
rect 229686 10852 229690 10908
rect 229626 10848 229690 10852
rect 229706 10908 229770 10912
rect 229706 10852 229710 10908
rect 229710 10852 229766 10908
rect 229766 10852 229770 10908
rect 229706 10848 229770 10852
rect 229786 10908 229850 10912
rect 229786 10852 229790 10908
rect 229790 10852 229846 10908
rect 229846 10852 229850 10908
rect 229786 10848 229850 10852
rect 39051 10364 39115 10368
rect 39051 10308 39055 10364
rect 39055 10308 39111 10364
rect 39111 10308 39115 10364
rect 39051 10304 39115 10308
rect 39131 10364 39195 10368
rect 39131 10308 39135 10364
rect 39135 10308 39191 10364
rect 39191 10308 39195 10364
rect 39131 10304 39195 10308
rect 39211 10364 39275 10368
rect 39211 10308 39215 10364
rect 39215 10308 39271 10364
rect 39271 10308 39275 10364
rect 39211 10304 39275 10308
rect 39291 10364 39355 10368
rect 39291 10308 39295 10364
rect 39295 10308 39351 10364
rect 39351 10308 39355 10364
rect 39291 10304 39355 10308
rect 115249 10364 115313 10368
rect 115249 10308 115253 10364
rect 115253 10308 115309 10364
rect 115309 10308 115313 10364
rect 115249 10304 115313 10308
rect 115329 10364 115393 10368
rect 115329 10308 115333 10364
rect 115333 10308 115389 10364
rect 115389 10308 115393 10364
rect 115329 10304 115393 10308
rect 115409 10364 115473 10368
rect 115409 10308 115413 10364
rect 115413 10308 115469 10364
rect 115469 10308 115473 10364
rect 115409 10304 115473 10308
rect 115489 10364 115553 10368
rect 115489 10308 115493 10364
rect 115493 10308 115549 10364
rect 115549 10308 115553 10364
rect 115489 10304 115553 10308
rect 191447 10364 191511 10368
rect 191447 10308 191451 10364
rect 191451 10308 191507 10364
rect 191507 10308 191511 10364
rect 191447 10304 191511 10308
rect 191527 10364 191591 10368
rect 191527 10308 191531 10364
rect 191531 10308 191587 10364
rect 191587 10308 191591 10364
rect 191527 10304 191591 10308
rect 191607 10364 191671 10368
rect 191607 10308 191611 10364
rect 191611 10308 191667 10364
rect 191667 10308 191671 10364
rect 191607 10304 191671 10308
rect 191687 10364 191751 10368
rect 191687 10308 191691 10364
rect 191691 10308 191747 10364
rect 191747 10308 191751 10364
rect 191687 10304 191751 10308
rect 267645 10364 267709 10368
rect 267645 10308 267649 10364
rect 267649 10308 267705 10364
rect 267705 10308 267709 10364
rect 267645 10304 267709 10308
rect 267725 10364 267789 10368
rect 267725 10308 267729 10364
rect 267729 10308 267785 10364
rect 267785 10308 267789 10364
rect 267725 10304 267789 10308
rect 267805 10364 267869 10368
rect 267805 10308 267809 10364
rect 267809 10308 267865 10364
rect 267865 10308 267869 10364
rect 267805 10304 267869 10308
rect 267885 10364 267949 10368
rect 267885 10308 267889 10364
rect 267889 10308 267945 10364
rect 267945 10308 267949 10364
rect 267885 10304 267949 10308
rect 77150 9820 77214 9824
rect 77150 9764 77154 9820
rect 77154 9764 77210 9820
rect 77210 9764 77214 9820
rect 77150 9760 77214 9764
rect 77230 9820 77294 9824
rect 77230 9764 77234 9820
rect 77234 9764 77290 9820
rect 77290 9764 77294 9820
rect 77230 9760 77294 9764
rect 77310 9820 77374 9824
rect 77310 9764 77314 9820
rect 77314 9764 77370 9820
rect 77370 9764 77374 9820
rect 77310 9760 77374 9764
rect 77390 9820 77454 9824
rect 77390 9764 77394 9820
rect 77394 9764 77450 9820
rect 77450 9764 77454 9820
rect 77390 9760 77454 9764
rect 153348 9820 153412 9824
rect 153348 9764 153352 9820
rect 153352 9764 153408 9820
rect 153408 9764 153412 9820
rect 153348 9760 153412 9764
rect 153428 9820 153492 9824
rect 153428 9764 153432 9820
rect 153432 9764 153488 9820
rect 153488 9764 153492 9820
rect 153428 9760 153492 9764
rect 153508 9820 153572 9824
rect 153508 9764 153512 9820
rect 153512 9764 153568 9820
rect 153568 9764 153572 9820
rect 153508 9760 153572 9764
rect 153588 9820 153652 9824
rect 153588 9764 153592 9820
rect 153592 9764 153648 9820
rect 153648 9764 153652 9820
rect 153588 9760 153652 9764
rect 229546 9820 229610 9824
rect 229546 9764 229550 9820
rect 229550 9764 229606 9820
rect 229606 9764 229610 9820
rect 229546 9760 229610 9764
rect 229626 9820 229690 9824
rect 229626 9764 229630 9820
rect 229630 9764 229686 9820
rect 229686 9764 229690 9820
rect 229626 9760 229690 9764
rect 229706 9820 229770 9824
rect 229706 9764 229710 9820
rect 229710 9764 229766 9820
rect 229766 9764 229770 9820
rect 229706 9760 229770 9764
rect 229786 9820 229850 9824
rect 229786 9764 229790 9820
rect 229790 9764 229846 9820
rect 229846 9764 229850 9820
rect 229786 9760 229850 9764
rect 39051 9276 39115 9280
rect 39051 9220 39055 9276
rect 39055 9220 39111 9276
rect 39111 9220 39115 9276
rect 39051 9216 39115 9220
rect 39131 9276 39195 9280
rect 39131 9220 39135 9276
rect 39135 9220 39191 9276
rect 39191 9220 39195 9276
rect 39131 9216 39195 9220
rect 39211 9276 39275 9280
rect 39211 9220 39215 9276
rect 39215 9220 39271 9276
rect 39271 9220 39275 9276
rect 39211 9216 39275 9220
rect 39291 9276 39355 9280
rect 39291 9220 39295 9276
rect 39295 9220 39351 9276
rect 39351 9220 39355 9276
rect 39291 9216 39355 9220
rect 115249 9276 115313 9280
rect 115249 9220 115253 9276
rect 115253 9220 115309 9276
rect 115309 9220 115313 9276
rect 115249 9216 115313 9220
rect 115329 9276 115393 9280
rect 115329 9220 115333 9276
rect 115333 9220 115389 9276
rect 115389 9220 115393 9276
rect 115329 9216 115393 9220
rect 115409 9276 115473 9280
rect 115409 9220 115413 9276
rect 115413 9220 115469 9276
rect 115469 9220 115473 9276
rect 115409 9216 115473 9220
rect 115489 9276 115553 9280
rect 115489 9220 115493 9276
rect 115493 9220 115549 9276
rect 115549 9220 115553 9276
rect 115489 9216 115553 9220
rect 191447 9276 191511 9280
rect 191447 9220 191451 9276
rect 191451 9220 191507 9276
rect 191507 9220 191511 9276
rect 191447 9216 191511 9220
rect 191527 9276 191591 9280
rect 191527 9220 191531 9276
rect 191531 9220 191587 9276
rect 191587 9220 191591 9276
rect 191527 9216 191591 9220
rect 191607 9276 191671 9280
rect 191607 9220 191611 9276
rect 191611 9220 191667 9276
rect 191667 9220 191671 9276
rect 191607 9216 191671 9220
rect 191687 9276 191751 9280
rect 191687 9220 191691 9276
rect 191691 9220 191747 9276
rect 191747 9220 191751 9276
rect 191687 9216 191751 9220
rect 267645 9276 267709 9280
rect 267645 9220 267649 9276
rect 267649 9220 267705 9276
rect 267705 9220 267709 9276
rect 267645 9216 267709 9220
rect 267725 9276 267789 9280
rect 267725 9220 267729 9276
rect 267729 9220 267785 9276
rect 267785 9220 267789 9276
rect 267725 9216 267789 9220
rect 267805 9276 267869 9280
rect 267805 9220 267809 9276
rect 267809 9220 267865 9276
rect 267865 9220 267869 9276
rect 267805 9216 267869 9220
rect 267885 9276 267949 9280
rect 267885 9220 267889 9276
rect 267889 9220 267945 9276
rect 267945 9220 267949 9276
rect 267885 9216 267949 9220
rect 77150 8732 77214 8736
rect 77150 8676 77154 8732
rect 77154 8676 77210 8732
rect 77210 8676 77214 8732
rect 77150 8672 77214 8676
rect 77230 8732 77294 8736
rect 77230 8676 77234 8732
rect 77234 8676 77290 8732
rect 77290 8676 77294 8732
rect 77230 8672 77294 8676
rect 77310 8732 77374 8736
rect 77310 8676 77314 8732
rect 77314 8676 77370 8732
rect 77370 8676 77374 8732
rect 77310 8672 77374 8676
rect 77390 8732 77454 8736
rect 77390 8676 77394 8732
rect 77394 8676 77450 8732
rect 77450 8676 77454 8732
rect 77390 8672 77454 8676
rect 153348 8732 153412 8736
rect 153348 8676 153352 8732
rect 153352 8676 153408 8732
rect 153408 8676 153412 8732
rect 153348 8672 153412 8676
rect 153428 8732 153492 8736
rect 153428 8676 153432 8732
rect 153432 8676 153488 8732
rect 153488 8676 153492 8732
rect 153428 8672 153492 8676
rect 153508 8732 153572 8736
rect 153508 8676 153512 8732
rect 153512 8676 153568 8732
rect 153568 8676 153572 8732
rect 153508 8672 153572 8676
rect 153588 8732 153652 8736
rect 153588 8676 153592 8732
rect 153592 8676 153648 8732
rect 153648 8676 153652 8732
rect 153588 8672 153652 8676
rect 229546 8732 229610 8736
rect 229546 8676 229550 8732
rect 229550 8676 229606 8732
rect 229606 8676 229610 8732
rect 229546 8672 229610 8676
rect 229626 8732 229690 8736
rect 229626 8676 229630 8732
rect 229630 8676 229686 8732
rect 229686 8676 229690 8732
rect 229626 8672 229690 8676
rect 229706 8732 229770 8736
rect 229706 8676 229710 8732
rect 229710 8676 229766 8732
rect 229766 8676 229770 8732
rect 229706 8672 229770 8676
rect 229786 8732 229850 8736
rect 229786 8676 229790 8732
rect 229790 8676 229846 8732
rect 229846 8676 229850 8732
rect 229786 8672 229850 8676
rect 39051 8188 39115 8192
rect 39051 8132 39055 8188
rect 39055 8132 39111 8188
rect 39111 8132 39115 8188
rect 39051 8128 39115 8132
rect 39131 8188 39195 8192
rect 39131 8132 39135 8188
rect 39135 8132 39191 8188
rect 39191 8132 39195 8188
rect 39131 8128 39195 8132
rect 39211 8188 39275 8192
rect 39211 8132 39215 8188
rect 39215 8132 39271 8188
rect 39271 8132 39275 8188
rect 39211 8128 39275 8132
rect 39291 8188 39355 8192
rect 39291 8132 39295 8188
rect 39295 8132 39351 8188
rect 39351 8132 39355 8188
rect 39291 8128 39355 8132
rect 115249 8188 115313 8192
rect 115249 8132 115253 8188
rect 115253 8132 115309 8188
rect 115309 8132 115313 8188
rect 115249 8128 115313 8132
rect 115329 8188 115393 8192
rect 115329 8132 115333 8188
rect 115333 8132 115389 8188
rect 115389 8132 115393 8188
rect 115329 8128 115393 8132
rect 115409 8188 115473 8192
rect 115409 8132 115413 8188
rect 115413 8132 115469 8188
rect 115469 8132 115473 8188
rect 115409 8128 115473 8132
rect 115489 8188 115553 8192
rect 115489 8132 115493 8188
rect 115493 8132 115549 8188
rect 115549 8132 115553 8188
rect 115489 8128 115553 8132
rect 191447 8188 191511 8192
rect 191447 8132 191451 8188
rect 191451 8132 191507 8188
rect 191507 8132 191511 8188
rect 191447 8128 191511 8132
rect 191527 8188 191591 8192
rect 191527 8132 191531 8188
rect 191531 8132 191587 8188
rect 191587 8132 191591 8188
rect 191527 8128 191591 8132
rect 191607 8188 191671 8192
rect 191607 8132 191611 8188
rect 191611 8132 191667 8188
rect 191667 8132 191671 8188
rect 191607 8128 191671 8132
rect 191687 8188 191751 8192
rect 191687 8132 191691 8188
rect 191691 8132 191747 8188
rect 191747 8132 191751 8188
rect 191687 8128 191751 8132
rect 267645 8188 267709 8192
rect 267645 8132 267649 8188
rect 267649 8132 267705 8188
rect 267705 8132 267709 8188
rect 267645 8128 267709 8132
rect 267725 8188 267789 8192
rect 267725 8132 267729 8188
rect 267729 8132 267785 8188
rect 267785 8132 267789 8188
rect 267725 8128 267789 8132
rect 267805 8188 267869 8192
rect 267805 8132 267809 8188
rect 267809 8132 267865 8188
rect 267865 8132 267869 8188
rect 267805 8128 267869 8132
rect 267885 8188 267949 8192
rect 267885 8132 267889 8188
rect 267889 8132 267945 8188
rect 267945 8132 267949 8188
rect 267885 8128 267949 8132
rect 77150 7644 77214 7648
rect 77150 7588 77154 7644
rect 77154 7588 77210 7644
rect 77210 7588 77214 7644
rect 77150 7584 77214 7588
rect 77230 7644 77294 7648
rect 77230 7588 77234 7644
rect 77234 7588 77290 7644
rect 77290 7588 77294 7644
rect 77230 7584 77294 7588
rect 77310 7644 77374 7648
rect 77310 7588 77314 7644
rect 77314 7588 77370 7644
rect 77370 7588 77374 7644
rect 77310 7584 77374 7588
rect 77390 7644 77454 7648
rect 77390 7588 77394 7644
rect 77394 7588 77450 7644
rect 77450 7588 77454 7644
rect 77390 7584 77454 7588
rect 153348 7644 153412 7648
rect 153348 7588 153352 7644
rect 153352 7588 153408 7644
rect 153408 7588 153412 7644
rect 153348 7584 153412 7588
rect 153428 7644 153492 7648
rect 153428 7588 153432 7644
rect 153432 7588 153488 7644
rect 153488 7588 153492 7644
rect 153428 7584 153492 7588
rect 153508 7644 153572 7648
rect 153508 7588 153512 7644
rect 153512 7588 153568 7644
rect 153568 7588 153572 7644
rect 153508 7584 153572 7588
rect 153588 7644 153652 7648
rect 153588 7588 153592 7644
rect 153592 7588 153648 7644
rect 153648 7588 153652 7644
rect 153588 7584 153652 7588
rect 229546 7644 229610 7648
rect 229546 7588 229550 7644
rect 229550 7588 229606 7644
rect 229606 7588 229610 7644
rect 229546 7584 229610 7588
rect 229626 7644 229690 7648
rect 229626 7588 229630 7644
rect 229630 7588 229686 7644
rect 229686 7588 229690 7644
rect 229626 7584 229690 7588
rect 229706 7644 229770 7648
rect 229706 7588 229710 7644
rect 229710 7588 229766 7644
rect 229766 7588 229770 7644
rect 229706 7584 229770 7588
rect 229786 7644 229850 7648
rect 229786 7588 229790 7644
rect 229790 7588 229846 7644
rect 229846 7588 229850 7644
rect 229786 7584 229850 7588
rect 39051 7100 39115 7104
rect 39051 7044 39055 7100
rect 39055 7044 39111 7100
rect 39111 7044 39115 7100
rect 39051 7040 39115 7044
rect 39131 7100 39195 7104
rect 39131 7044 39135 7100
rect 39135 7044 39191 7100
rect 39191 7044 39195 7100
rect 39131 7040 39195 7044
rect 39211 7100 39275 7104
rect 39211 7044 39215 7100
rect 39215 7044 39271 7100
rect 39271 7044 39275 7100
rect 39211 7040 39275 7044
rect 39291 7100 39355 7104
rect 39291 7044 39295 7100
rect 39295 7044 39351 7100
rect 39351 7044 39355 7100
rect 39291 7040 39355 7044
rect 115249 7100 115313 7104
rect 115249 7044 115253 7100
rect 115253 7044 115309 7100
rect 115309 7044 115313 7100
rect 115249 7040 115313 7044
rect 115329 7100 115393 7104
rect 115329 7044 115333 7100
rect 115333 7044 115389 7100
rect 115389 7044 115393 7100
rect 115329 7040 115393 7044
rect 115409 7100 115473 7104
rect 115409 7044 115413 7100
rect 115413 7044 115469 7100
rect 115469 7044 115473 7100
rect 115409 7040 115473 7044
rect 115489 7100 115553 7104
rect 115489 7044 115493 7100
rect 115493 7044 115549 7100
rect 115549 7044 115553 7100
rect 115489 7040 115553 7044
rect 191447 7100 191511 7104
rect 191447 7044 191451 7100
rect 191451 7044 191507 7100
rect 191507 7044 191511 7100
rect 191447 7040 191511 7044
rect 191527 7100 191591 7104
rect 191527 7044 191531 7100
rect 191531 7044 191587 7100
rect 191587 7044 191591 7100
rect 191527 7040 191591 7044
rect 191607 7100 191671 7104
rect 191607 7044 191611 7100
rect 191611 7044 191667 7100
rect 191667 7044 191671 7100
rect 191607 7040 191671 7044
rect 191687 7100 191751 7104
rect 191687 7044 191691 7100
rect 191691 7044 191747 7100
rect 191747 7044 191751 7100
rect 191687 7040 191751 7044
rect 267645 7100 267709 7104
rect 267645 7044 267649 7100
rect 267649 7044 267705 7100
rect 267705 7044 267709 7100
rect 267645 7040 267709 7044
rect 267725 7100 267789 7104
rect 267725 7044 267729 7100
rect 267729 7044 267785 7100
rect 267785 7044 267789 7100
rect 267725 7040 267789 7044
rect 267805 7100 267869 7104
rect 267805 7044 267809 7100
rect 267809 7044 267865 7100
rect 267865 7044 267869 7100
rect 267805 7040 267869 7044
rect 267885 7100 267949 7104
rect 267885 7044 267889 7100
rect 267889 7044 267945 7100
rect 267945 7044 267949 7100
rect 267885 7040 267949 7044
rect 77150 6556 77214 6560
rect 77150 6500 77154 6556
rect 77154 6500 77210 6556
rect 77210 6500 77214 6556
rect 77150 6496 77214 6500
rect 77230 6556 77294 6560
rect 77230 6500 77234 6556
rect 77234 6500 77290 6556
rect 77290 6500 77294 6556
rect 77230 6496 77294 6500
rect 77310 6556 77374 6560
rect 77310 6500 77314 6556
rect 77314 6500 77370 6556
rect 77370 6500 77374 6556
rect 77310 6496 77374 6500
rect 77390 6556 77454 6560
rect 77390 6500 77394 6556
rect 77394 6500 77450 6556
rect 77450 6500 77454 6556
rect 77390 6496 77454 6500
rect 153348 6556 153412 6560
rect 153348 6500 153352 6556
rect 153352 6500 153408 6556
rect 153408 6500 153412 6556
rect 153348 6496 153412 6500
rect 153428 6556 153492 6560
rect 153428 6500 153432 6556
rect 153432 6500 153488 6556
rect 153488 6500 153492 6556
rect 153428 6496 153492 6500
rect 153508 6556 153572 6560
rect 153508 6500 153512 6556
rect 153512 6500 153568 6556
rect 153568 6500 153572 6556
rect 153508 6496 153572 6500
rect 153588 6556 153652 6560
rect 153588 6500 153592 6556
rect 153592 6500 153648 6556
rect 153648 6500 153652 6556
rect 153588 6496 153652 6500
rect 229546 6556 229610 6560
rect 229546 6500 229550 6556
rect 229550 6500 229606 6556
rect 229606 6500 229610 6556
rect 229546 6496 229610 6500
rect 229626 6556 229690 6560
rect 229626 6500 229630 6556
rect 229630 6500 229686 6556
rect 229686 6500 229690 6556
rect 229626 6496 229690 6500
rect 229706 6556 229770 6560
rect 229706 6500 229710 6556
rect 229710 6500 229766 6556
rect 229766 6500 229770 6556
rect 229706 6496 229770 6500
rect 229786 6556 229850 6560
rect 229786 6500 229790 6556
rect 229790 6500 229846 6556
rect 229846 6500 229850 6556
rect 229786 6496 229850 6500
rect 39051 6012 39115 6016
rect 39051 5956 39055 6012
rect 39055 5956 39111 6012
rect 39111 5956 39115 6012
rect 39051 5952 39115 5956
rect 39131 6012 39195 6016
rect 39131 5956 39135 6012
rect 39135 5956 39191 6012
rect 39191 5956 39195 6012
rect 39131 5952 39195 5956
rect 39211 6012 39275 6016
rect 39211 5956 39215 6012
rect 39215 5956 39271 6012
rect 39271 5956 39275 6012
rect 39211 5952 39275 5956
rect 39291 6012 39355 6016
rect 39291 5956 39295 6012
rect 39295 5956 39351 6012
rect 39351 5956 39355 6012
rect 39291 5952 39355 5956
rect 115249 6012 115313 6016
rect 115249 5956 115253 6012
rect 115253 5956 115309 6012
rect 115309 5956 115313 6012
rect 115249 5952 115313 5956
rect 115329 6012 115393 6016
rect 115329 5956 115333 6012
rect 115333 5956 115389 6012
rect 115389 5956 115393 6012
rect 115329 5952 115393 5956
rect 115409 6012 115473 6016
rect 115409 5956 115413 6012
rect 115413 5956 115469 6012
rect 115469 5956 115473 6012
rect 115409 5952 115473 5956
rect 115489 6012 115553 6016
rect 115489 5956 115493 6012
rect 115493 5956 115549 6012
rect 115549 5956 115553 6012
rect 115489 5952 115553 5956
rect 191447 6012 191511 6016
rect 191447 5956 191451 6012
rect 191451 5956 191507 6012
rect 191507 5956 191511 6012
rect 191447 5952 191511 5956
rect 191527 6012 191591 6016
rect 191527 5956 191531 6012
rect 191531 5956 191587 6012
rect 191587 5956 191591 6012
rect 191527 5952 191591 5956
rect 191607 6012 191671 6016
rect 191607 5956 191611 6012
rect 191611 5956 191667 6012
rect 191667 5956 191671 6012
rect 191607 5952 191671 5956
rect 191687 6012 191751 6016
rect 191687 5956 191691 6012
rect 191691 5956 191747 6012
rect 191747 5956 191751 6012
rect 191687 5952 191751 5956
rect 267645 6012 267709 6016
rect 267645 5956 267649 6012
rect 267649 5956 267705 6012
rect 267705 5956 267709 6012
rect 267645 5952 267709 5956
rect 267725 6012 267789 6016
rect 267725 5956 267729 6012
rect 267729 5956 267785 6012
rect 267785 5956 267789 6012
rect 267725 5952 267789 5956
rect 267805 6012 267869 6016
rect 267805 5956 267809 6012
rect 267809 5956 267865 6012
rect 267865 5956 267869 6012
rect 267805 5952 267869 5956
rect 267885 6012 267949 6016
rect 267885 5956 267889 6012
rect 267889 5956 267945 6012
rect 267945 5956 267949 6012
rect 267885 5952 267949 5956
rect 77150 5468 77214 5472
rect 77150 5412 77154 5468
rect 77154 5412 77210 5468
rect 77210 5412 77214 5468
rect 77150 5408 77214 5412
rect 77230 5468 77294 5472
rect 77230 5412 77234 5468
rect 77234 5412 77290 5468
rect 77290 5412 77294 5468
rect 77230 5408 77294 5412
rect 77310 5468 77374 5472
rect 77310 5412 77314 5468
rect 77314 5412 77370 5468
rect 77370 5412 77374 5468
rect 77310 5408 77374 5412
rect 77390 5468 77454 5472
rect 77390 5412 77394 5468
rect 77394 5412 77450 5468
rect 77450 5412 77454 5468
rect 77390 5408 77454 5412
rect 153348 5468 153412 5472
rect 153348 5412 153352 5468
rect 153352 5412 153408 5468
rect 153408 5412 153412 5468
rect 153348 5408 153412 5412
rect 153428 5468 153492 5472
rect 153428 5412 153432 5468
rect 153432 5412 153488 5468
rect 153488 5412 153492 5468
rect 153428 5408 153492 5412
rect 153508 5468 153572 5472
rect 153508 5412 153512 5468
rect 153512 5412 153568 5468
rect 153568 5412 153572 5468
rect 153508 5408 153572 5412
rect 153588 5468 153652 5472
rect 153588 5412 153592 5468
rect 153592 5412 153648 5468
rect 153648 5412 153652 5468
rect 153588 5408 153652 5412
rect 229546 5468 229610 5472
rect 229546 5412 229550 5468
rect 229550 5412 229606 5468
rect 229606 5412 229610 5468
rect 229546 5408 229610 5412
rect 229626 5468 229690 5472
rect 229626 5412 229630 5468
rect 229630 5412 229686 5468
rect 229686 5412 229690 5468
rect 229626 5408 229690 5412
rect 229706 5468 229770 5472
rect 229706 5412 229710 5468
rect 229710 5412 229766 5468
rect 229766 5412 229770 5468
rect 229706 5408 229770 5412
rect 229786 5468 229850 5472
rect 229786 5412 229790 5468
rect 229790 5412 229846 5468
rect 229846 5412 229850 5468
rect 229786 5408 229850 5412
rect 39051 4924 39115 4928
rect 39051 4868 39055 4924
rect 39055 4868 39111 4924
rect 39111 4868 39115 4924
rect 39051 4864 39115 4868
rect 39131 4924 39195 4928
rect 39131 4868 39135 4924
rect 39135 4868 39191 4924
rect 39191 4868 39195 4924
rect 39131 4864 39195 4868
rect 39211 4924 39275 4928
rect 39211 4868 39215 4924
rect 39215 4868 39271 4924
rect 39271 4868 39275 4924
rect 39211 4864 39275 4868
rect 39291 4924 39355 4928
rect 39291 4868 39295 4924
rect 39295 4868 39351 4924
rect 39351 4868 39355 4924
rect 39291 4864 39355 4868
rect 115249 4924 115313 4928
rect 115249 4868 115253 4924
rect 115253 4868 115309 4924
rect 115309 4868 115313 4924
rect 115249 4864 115313 4868
rect 115329 4924 115393 4928
rect 115329 4868 115333 4924
rect 115333 4868 115389 4924
rect 115389 4868 115393 4924
rect 115329 4864 115393 4868
rect 115409 4924 115473 4928
rect 115409 4868 115413 4924
rect 115413 4868 115469 4924
rect 115469 4868 115473 4924
rect 115409 4864 115473 4868
rect 115489 4924 115553 4928
rect 115489 4868 115493 4924
rect 115493 4868 115549 4924
rect 115549 4868 115553 4924
rect 115489 4864 115553 4868
rect 191447 4924 191511 4928
rect 191447 4868 191451 4924
rect 191451 4868 191507 4924
rect 191507 4868 191511 4924
rect 191447 4864 191511 4868
rect 191527 4924 191591 4928
rect 191527 4868 191531 4924
rect 191531 4868 191587 4924
rect 191587 4868 191591 4924
rect 191527 4864 191591 4868
rect 191607 4924 191671 4928
rect 191607 4868 191611 4924
rect 191611 4868 191667 4924
rect 191667 4868 191671 4924
rect 191607 4864 191671 4868
rect 191687 4924 191751 4928
rect 191687 4868 191691 4924
rect 191691 4868 191747 4924
rect 191747 4868 191751 4924
rect 191687 4864 191751 4868
rect 267645 4924 267709 4928
rect 267645 4868 267649 4924
rect 267649 4868 267705 4924
rect 267705 4868 267709 4924
rect 267645 4864 267709 4868
rect 267725 4924 267789 4928
rect 267725 4868 267729 4924
rect 267729 4868 267785 4924
rect 267785 4868 267789 4924
rect 267725 4864 267789 4868
rect 267805 4924 267869 4928
rect 267805 4868 267809 4924
rect 267809 4868 267865 4924
rect 267865 4868 267869 4924
rect 267805 4864 267869 4868
rect 267885 4924 267949 4928
rect 267885 4868 267889 4924
rect 267889 4868 267945 4924
rect 267945 4868 267949 4924
rect 267885 4864 267949 4868
rect 77150 4380 77214 4384
rect 77150 4324 77154 4380
rect 77154 4324 77210 4380
rect 77210 4324 77214 4380
rect 77150 4320 77214 4324
rect 77230 4380 77294 4384
rect 77230 4324 77234 4380
rect 77234 4324 77290 4380
rect 77290 4324 77294 4380
rect 77230 4320 77294 4324
rect 77310 4380 77374 4384
rect 77310 4324 77314 4380
rect 77314 4324 77370 4380
rect 77370 4324 77374 4380
rect 77310 4320 77374 4324
rect 77390 4380 77454 4384
rect 77390 4324 77394 4380
rect 77394 4324 77450 4380
rect 77450 4324 77454 4380
rect 77390 4320 77454 4324
rect 153348 4380 153412 4384
rect 153348 4324 153352 4380
rect 153352 4324 153408 4380
rect 153408 4324 153412 4380
rect 153348 4320 153412 4324
rect 153428 4380 153492 4384
rect 153428 4324 153432 4380
rect 153432 4324 153488 4380
rect 153488 4324 153492 4380
rect 153428 4320 153492 4324
rect 153508 4380 153572 4384
rect 153508 4324 153512 4380
rect 153512 4324 153568 4380
rect 153568 4324 153572 4380
rect 153508 4320 153572 4324
rect 153588 4380 153652 4384
rect 153588 4324 153592 4380
rect 153592 4324 153648 4380
rect 153648 4324 153652 4380
rect 153588 4320 153652 4324
rect 229546 4380 229610 4384
rect 229546 4324 229550 4380
rect 229550 4324 229606 4380
rect 229606 4324 229610 4380
rect 229546 4320 229610 4324
rect 229626 4380 229690 4384
rect 229626 4324 229630 4380
rect 229630 4324 229686 4380
rect 229686 4324 229690 4380
rect 229626 4320 229690 4324
rect 229706 4380 229770 4384
rect 229706 4324 229710 4380
rect 229710 4324 229766 4380
rect 229766 4324 229770 4380
rect 229706 4320 229770 4324
rect 229786 4380 229850 4384
rect 229786 4324 229790 4380
rect 229790 4324 229846 4380
rect 229846 4324 229850 4380
rect 229786 4320 229850 4324
rect 39051 3836 39115 3840
rect 39051 3780 39055 3836
rect 39055 3780 39111 3836
rect 39111 3780 39115 3836
rect 39051 3776 39115 3780
rect 39131 3836 39195 3840
rect 39131 3780 39135 3836
rect 39135 3780 39191 3836
rect 39191 3780 39195 3836
rect 39131 3776 39195 3780
rect 39211 3836 39275 3840
rect 39211 3780 39215 3836
rect 39215 3780 39271 3836
rect 39271 3780 39275 3836
rect 39211 3776 39275 3780
rect 39291 3836 39355 3840
rect 39291 3780 39295 3836
rect 39295 3780 39351 3836
rect 39351 3780 39355 3836
rect 39291 3776 39355 3780
rect 115249 3836 115313 3840
rect 115249 3780 115253 3836
rect 115253 3780 115309 3836
rect 115309 3780 115313 3836
rect 115249 3776 115313 3780
rect 115329 3836 115393 3840
rect 115329 3780 115333 3836
rect 115333 3780 115389 3836
rect 115389 3780 115393 3836
rect 115329 3776 115393 3780
rect 115409 3836 115473 3840
rect 115409 3780 115413 3836
rect 115413 3780 115469 3836
rect 115469 3780 115473 3836
rect 115409 3776 115473 3780
rect 115489 3836 115553 3840
rect 115489 3780 115493 3836
rect 115493 3780 115549 3836
rect 115549 3780 115553 3836
rect 115489 3776 115553 3780
rect 191447 3836 191511 3840
rect 191447 3780 191451 3836
rect 191451 3780 191507 3836
rect 191507 3780 191511 3836
rect 191447 3776 191511 3780
rect 191527 3836 191591 3840
rect 191527 3780 191531 3836
rect 191531 3780 191587 3836
rect 191587 3780 191591 3836
rect 191527 3776 191591 3780
rect 191607 3836 191671 3840
rect 191607 3780 191611 3836
rect 191611 3780 191667 3836
rect 191667 3780 191671 3836
rect 191607 3776 191671 3780
rect 191687 3836 191751 3840
rect 191687 3780 191691 3836
rect 191691 3780 191747 3836
rect 191747 3780 191751 3836
rect 191687 3776 191751 3780
rect 267645 3836 267709 3840
rect 267645 3780 267649 3836
rect 267649 3780 267705 3836
rect 267705 3780 267709 3836
rect 267645 3776 267709 3780
rect 267725 3836 267789 3840
rect 267725 3780 267729 3836
rect 267729 3780 267785 3836
rect 267785 3780 267789 3836
rect 267725 3776 267789 3780
rect 267805 3836 267869 3840
rect 267805 3780 267809 3836
rect 267809 3780 267865 3836
rect 267865 3780 267869 3836
rect 267805 3776 267869 3780
rect 267885 3836 267949 3840
rect 267885 3780 267889 3836
rect 267889 3780 267945 3836
rect 267945 3780 267949 3836
rect 267885 3776 267949 3780
rect 77150 3292 77214 3296
rect 77150 3236 77154 3292
rect 77154 3236 77210 3292
rect 77210 3236 77214 3292
rect 77150 3232 77214 3236
rect 77230 3292 77294 3296
rect 77230 3236 77234 3292
rect 77234 3236 77290 3292
rect 77290 3236 77294 3292
rect 77230 3232 77294 3236
rect 77310 3292 77374 3296
rect 77310 3236 77314 3292
rect 77314 3236 77370 3292
rect 77370 3236 77374 3292
rect 77310 3232 77374 3236
rect 77390 3292 77454 3296
rect 77390 3236 77394 3292
rect 77394 3236 77450 3292
rect 77450 3236 77454 3292
rect 77390 3232 77454 3236
rect 153348 3292 153412 3296
rect 153348 3236 153352 3292
rect 153352 3236 153408 3292
rect 153408 3236 153412 3292
rect 153348 3232 153412 3236
rect 153428 3292 153492 3296
rect 153428 3236 153432 3292
rect 153432 3236 153488 3292
rect 153488 3236 153492 3292
rect 153428 3232 153492 3236
rect 153508 3292 153572 3296
rect 153508 3236 153512 3292
rect 153512 3236 153568 3292
rect 153568 3236 153572 3292
rect 153508 3232 153572 3236
rect 153588 3292 153652 3296
rect 153588 3236 153592 3292
rect 153592 3236 153648 3292
rect 153648 3236 153652 3292
rect 153588 3232 153652 3236
rect 229546 3292 229610 3296
rect 229546 3236 229550 3292
rect 229550 3236 229606 3292
rect 229606 3236 229610 3292
rect 229546 3232 229610 3236
rect 229626 3292 229690 3296
rect 229626 3236 229630 3292
rect 229630 3236 229686 3292
rect 229686 3236 229690 3292
rect 229626 3232 229690 3236
rect 229706 3292 229770 3296
rect 229706 3236 229710 3292
rect 229710 3236 229766 3292
rect 229766 3236 229770 3292
rect 229706 3232 229770 3236
rect 229786 3292 229850 3296
rect 229786 3236 229790 3292
rect 229790 3236 229846 3292
rect 229846 3236 229850 3292
rect 229786 3232 229850 3236
rect 39051 2748 39115 2752
rect 39051 2692 39055 2748
rect 39055 2692 39111 2748
rect 39111 2692 39115 2748
rect 39051 2688 39115 2692
rect 39131 2748 39195 2752
rect 39131 2692 39135 2748
rect 39135 2692 39191 2748
rect 39191 2692 39195 2748
rect 39131 2688 39195 2692
rect 39211 2748 39275 2752
rect 39211 2692 39215 2748
rect 39215 2692 39271 2748
rect 39271 2692 39275 2748
rect 39211 2688 39275 2692
rect 39291 2748 39355 2752
rect 39291 2692 39295 2748
rect 39295 2692 39351 2748
rect 39351 2692 39355 2748
rect 39291 2688 39355 2692
rect 115249 2748 115313 2752
rect 115249 2692 115253 2748
rect 115253 2692 115309 2748
rect 115309 2692 115313 2748
rect 115249 2688 115313 2692
rect 115329 2748 115393 2752
rect 115329 2692 115333 2748
rect 115333 2692 115389 2748
rect 115389 2692 115393 2748
rect 115329 2688 115393 2692
rect 115409 2748 115473 2752
rect 115409 2692 115413 2748
rect 115413 2692 115469 2748
rect 115469 2692 115473 2748
rect 115409 2688 115473 2692
rect 115489 2748 115553 2752
rect 115489 2692 115493 2748
rect 115493 2692 115549 2748
rect 115549 2692 115553 2748
rect 115489 2688 115553 2692
rect 191447 2748 191511 2752
rect 191447 2692 191451 2748
rect 191451 2692 191507 2748
rect 191507 2692 191511 2748
rect 191447 2688 191511 2692
rect 191527 2748 191591 2752
rect 191527 2692 191531 2748
rect 191531 2692 191587 2748
rect 191587 2692 191591 2748
rect 191527 2688 191591 2692
rect 191607 2748 191671 2752
rect 191607 2692 191611 2748
rect 191611 2692 191667 2748
rect 191667 2692 191671 2748
rect 191607 2688 191671 2692
rect 191687 2748 191751 2752
rect 191687 2692 191691 2748
rect 191691 2692 191747 2748
rect 191747 2692 191751 2748
rect 191687 2688 191751 2692
rect 267645 2748 267709 2752
rect 267645 2692 267649 2748
rect 267649 2692 267705 2748
rect 267705 2692 267709 2748
rect 267645 2688 267709 2692
rect 267725 2748 267789 2752
rect 267725 2692 267729 2748
rect 267729 2692 267785 2748
rect 267785 2692 267789 2748
rect 267725 2688 267789 2692
rect 267805 2748 267869 2752
rect 267805 2692 267809 2748
rect 267809 2692 267865 2748
rect 267865 2692 267869 2748
rect 267805 2688 267869 2692
rect 267885 2748 267949 2752
rect 267885 2692 267889 2748
rect 267889 2692 267945 2748
rect 267945 2692 267949 2748
rect 267885 2688 267949 2692
rect 77150 2204 77214 2208
rect 77150 2148 77154 2204
rect 77154 2148 77210 2204
rect 77210 2148 77214 2204
rect 77150 2144 77214 2148
rect 77230 2204 77294 2208
rect 77230 2148 77234 2204
rect 77234 2148 77290 2204
rect 77290 2148 77294 2204
rect 77230 2144 77294 2148
rect 77310 2204 77374 2208
rect 77310 2148 77314 2204
rect 77314 2148 77370 2204
rect 77370 2148 77374 2204
rect 77310 2144 77374 2148
rect 77390 2204 77454 2208
rect 77390 2148 77394 2204
rect 77394 2148 77450 2204
rect 77450 2148 77454 2204
rect 77390 2144 77454 2148
rect 153348 2204 153412 2208
rect 153348 2148 153352 2204
rect 153352 2148 153408 2204
rect 153408 2148 153412 2204
rect 153348 2144 153412 2148
rect 153428 2204 153492 2208
rect 153428 2148 153432 2204
rect 153432 2148 153488 2204
rect 153488 2148 153492 2204
rect 153428 2144 153492 2148
rect 153508 2204 153572 2208
rect 153508 2148 153512 2204
rect 153512 2148 153568 2204
rect 153568 2148 153572 2204
rect 153508 2144 153572 2148
rect 153588 2204 153652 2208
rect 153588 2148 153592 2204
rect 153592 2148 153648 2204
rect 153648 2148 153652 2204
rect 153588 2144 153652 2148
rect 229546 2204 229610 2208
rect 229546 2148 229550 2204
rect 229550 2148 229606 2204
rect 229606 2148 229610 2204
rect 229546 2144 229610 2148
rect 229626 2204 229690 2208
rect 229626 2148 229630 2204
rect 229630 2148 229686 2204
rect 229686 2148 229690 2204
rect 229626 2144 229690 2148
rect 229706 2204 229770 2208
rect 229706 2148 229710 2204
rect 229710 2148 229766 2204
rect 229766 2148 229770 2204
rect 229706 2144 229770 2148
rect 229786 2204 229850 2208
rect 229786 2148 229790 2204
rect 229790 2148 229846 2204
rect 229846 2148 229850 2204
rect 229786 2144 229850 2148
<< metal4 >>
rect -1076 15738 -756 15780
rect -1076 15502 -1034 15738
rect -798 15502 -756 15738
rect -1076 11030 -756 15502
rect -1076 10794 -1034 11030
rect -798 10794 -756 11030
rect -1076 8118 -756 10794
rect -1076 7882 -1034 8118
rect -798 7882 -756 8118
rect -1076 5206 -756 7882
rect -1076 4970 -1034 5206
rect -798 4970 -756 5206
rect -1076 274 -756 4970
rect -416 15078 -96 15120
rect -416 14842 -374 15078
rect -138 14842 -96 15078
rect -416 12486 -96 14842
rect -416 12250 -374 12486
rect -138 12250 -96 12486
rect -416 9574 -96 12250
rect -416 9338 -374 9574
rect -138 9338 -96 9574
rect -416 6662 -96 9338
rect -416 6426 -374 6662
rect -138 6426 -96 6662
rect -416 3750 -96 6426
rect -416 3514 -374 3750
rect -138 3514 -96 3750
rect -416 934 -96 3514
rect -416 698 -374 934
rect -138 698 -96 934
rect -416 656 -96 698
rect 39043 15078 39363 15780
rect 39043 14842 39085 15078
rect 39321 14842 39363 15078
rect 39043 13632 39363 14842
rect 39043 13568 39051 13632
rect 39115 13568 39131 13632
rect 39195 13568 39211 13632
rect 39275 13568 39291 13632
rect 39355 13568 39363 13632
rect 39043 12544 39363 13568
rect 39043 12480 39051 12544
rect 39115 12486 39131 12544
rect 39195 12486 39211 12544
rect 39275 12486 39291 12544
rect 39355 12480 39363 12544
rect 39043 12250 39085 12480
rect 39321 12250 39363 12480
rect 39043 11456 39363 12250
rect 39043 11392 39051 11456
rect 39115 11392 39131 11456
rect 39195 11392 39211 11456
rect 39275 11392 39291 11456
rect 39355 11392 39363 11456
rect 39043 10368 39363 11392
rect 39043 10304 39051 10368
rect 39115 10304 39131 10368
rect 39195 10304 39211 10368
rect 39275 10304 39291 10368
rect 39355 10304 39363 10368
rect 39043 9574 39363 10304
rect 39043 9338 39085 9574
rect 39321 9338 39363 9574
rect 39043 9280 39363 9338
rect 39043 9216 39051 9280
rect 39115 9216 39131 9280
rect 39195 9216 39211 9280
rect 39275 9216 39291 9280
rect 39355 9216 39363 9280
rect 39043 8192 39363 9216
rect 39043 8128 39051 8192
rect 39115 8128 39131 8192
rect 39195 8128 39211 8192
rect 39275 8128 39291 8192
rect 39355 8128 39363 8192
rect 39043 7104 39363 8128
rect 39043 7040 39051 7104
rect 39115 7040 39131 7104
rect 39195 7040 39211 7104
rect 39275 7040 39291 7104
rect 39355 7040 39363 7104
rect 39043 6662 39363 7040
rect 39043 6426 39085 6662
rect 39321 6426 39363 6662
rect 39043 6016 39363 6426
rect 39043 5952 39051 6016
rect 39115 5952 39131 6016
rect 39195 5952 39211 6016
rect 39275 5952 39291 6016
rect 39355 5952 39363 6016
rect 39043 4928 39363 5952
rect 39043 4864 39051 4928
rect 39115 4864 39131 4928
rect 39195 4864 39211 4928
rect 39275 4864 39291 4928
rect 39355 4864 39363 4928
rect 39043 3840 39363 4864
rect 39043 3776 39051 3840
rect 39115 3776 39131 3840
rect 39195 3776 39211 3840
rect 39275 3776 39291 3840
rect 39355 3776 39363 3840
rect 39043 3750 39363 3776
rect 39043 3514 39085 3750
rect 39321 3514 39363 3750
rect 39043 2752 39363 3514
rect 39043 2688 39051 2752
rect 39115 2688 39131 2752
rect 39195 2688 39211 2752
rect 39275 2688 39291 2752
rect 39355 2688 39363 2752
rect 39043 934 39363 2688
rect 39043 698 39085 934
rect 39321 698 39363 934
rect -1076 38 -1034 274
rect -798 38 -756 274
rect -1076 -4 -756 38
rect 39043 -4 39363 698
rect 77142 15738 77462 15780
rect 77142 15502 77184 15738
rect 77420 15502 77462 15738
rect 77142 13088 77462 15502
rect 77142 13024 77150 13088
rect 77214 13024 77230 13088
rect 77294 13024 77310 13088
rect 77374 13024 77390 13088
rect 77454 13024 77462 13088
rect 77142 12000 77462 13024
rect 77142 11936 77150 12000
rect 77214 11936 77230 12000
rect 77294 11936 77310 12000
rect 77374 11936 77390 12000
rect 77454 11936 77462 12000
rect 77142 11030 77462 11936
rect 77142 10912 77184 11030
rect 77420 10912 77462 11030
rect 77142 10848 77150 10912
rect 77454 10848 77462 10912
rect 77142 10794 77184 10848
rect 77420 10794 77462 10848
rect 77142 9824 77462 10794
rect 77142 9760 77150 9824
rect 77214 9760 77230 9824
rect 77294 9760 77310 9824
rect 77374 9760 77390 9824
rect 77454 9760 77462 9824
rect 77142 8736 77462 9760
rect 77142 8672 77150 8736
rect 77214 8672 77230 8736
rect 77294 8672 77310 8736
rect 77374 8672 77390 8736
rect 77454 8672 77462 8736
rect 77142 8118 77462 8672
rect 77142 7882 77184 8118
rect 77420 7882 77462 8118
rect 77142 7648 77462 7882
rect 77142 7584 77150 7648
rect 77214 7584 77230 7648
rect 77294 7584 77310 7648
rect 77374 7584 77390 7648
rect 77454 7584 77462 7648
rect 77142 6560 77462 7584
rect 77142 6496 77150 6560
rect 77214 6496 77230 6560
rect 77294 6496 77310 6560
rect 77374 6496 77390 6560
rect 77454 6496 77462 6560
rect 77142 5472 77462 6496
rect 77142 5408 77150 5472
rect 77214 5408 77230 5472
rect 77294 5408 77310 5472
rect 77374 5408 77390 5472
rect 77454 5408 77462 5472
rect 77142 5206 77462 5408
rect 77142 4970 77184 5206
rect 77420 4970 77462 5206
rect 77142 4384 77462 4970
rect 77142 4320 77150 4384
rect 77214 4320 77230 4384
rect 77294 4320 77310 4384
rect 77374 4320 77390 4384
rect 77454 4320 77462 4384
rect 77142 3296 77462 4320
rect 77142 3232 77150 3296
rect 77214 3232 77230 3296
rect 77294 3232 77310 3296
rect 77374 3232 77390 3296
rect 77454 3232 77462 3296
rect 77142 2208 77462 3232
rect 77142 2144 77150 2208
rect 77214 2144 77230 2208
rect 77294 2144 77310 2208
rect 77374 2144 77390 2208
rect 77454 2144 77462 2208
rect 77142 274 77462 2144
rect 77142 38 77184 274
rect 77420 38 77462 274
rect 77142 -4 77462 38
rect 115241 15078 115561 15780
rect 115241 14842 115283 15078
rect 115519 14842 115561 15078
rect 115241 13632 115561 14842
rect 115241 13568 115249 13632
rect 115313 13568 115329 13632
rect 115393 13568 115409 13632
rect 115473 13568 115489 13632
rect 115553 13568 115561 13632
rect 115241 12544 115561 13568
rect 115241 12480 115249 12544
rect 115313 12486 115329 12544
rect 115393 12486 115409 12544
rect 115473 12486 115489 12544
rect 115553 12480 115561 12544
rect 115241 12250 115283 12480
rect 115519 12250 115561 12480
rect 115241 11456 115561 12250
rect 115241 11392 115249 11456
rect 115313 11392 115329 11456
rect 115393 11392 115409 11456
rect 115473 11392 115489 11456
rect 115553 11392 115561 11456
rect 115241 10368 115561 11392
rect 115241 10304 115249 10368
rect 115313 10304 115329 10368
rect 115393 10304 115409 10368
rect 115473 10304 115489 10368
rect 115553 10304 115561 10368
rect 115241 9574 115561 10304
rect 115241 9338 115283 9574
rect 115519 9338 115561 9574
rect 115241 9280 115561 9338
rect 115241 9216 115249 9280
rect 115313 9216 115329 9280
rect 115393 9216 115409 9280
rect 115473 9216 115489 9280
rect 115553 9216 115561 9280
rect 115241 8192 115561 9216
rect 115241 8128 115249 8192
rect 115313 8128 115329 8192
rect 115393 8128 115409 8192
rect 115473 8128 115489 8192
rect 115553 8128 115561 8192
rect 115241 7104 115561 8128
rect 115241 7040 115249 7104
rect 115313 7040 115329 7104
rect 115393 7040 115409 7104
rect 115473 7040 115489 7104
rect 115553 7040 115561 7104
rect 115241 6662 115561 7040
rect 115241 6426 115283 6662
rect 115519 6426 115561 6662
rect 115241 6016 115561 6426
rect 115241 5952 115249 6016
rect 115313 5952 115329 6016
rect 115393 5952 115409 6016
rect 115473 5952 115489 6016
rect 115553 5952 115561 6016
rect 115241 4928 115561 5952
rect 115241 4864 115249 4928
rect 115313 4864 115329 4928
rect 115393 4864 115409 4928
rect 115473 4864 115489 4928
rect 115553 4864 115561 4928
rect 115241 3840 115561 4864
rect 115241 3776 115249 3840
rect 115313 3776 115329 3840
rect 115393 3776 115409 3840
rect 115473 3776 115489 3840
rect 115553 3776 115561 3840
rect 115241 3750 115561 3776
rect 115241 3514 115283 3750
rect 115519 3514 115561 3750
rect 115241 2752 115561 3514
rect 115241 2688 115249 2752
rect 115313 2688 115329 2752
rect 115393 2688 115409 2752
rect 115473 2688 115489 2752
rect 115553 2688 115561 2752
rect 115241 934 115561 2688
rect 115241 698 115283 934
rect 115519 698 115561 934
rect 115241 -4 115561 698
rect 153340 15738 153660 15780
rect 153340 15502 153382 15738
rect 153618 15502 153660 15738
rect 153340 13088 153660 15502
rect 153340 13024 153348 13088
rect 153412 13024 153428 13088
rect 153492 13024 153508 13088
rect 153572 13024 153588 13088
rect 153652 13024 153660 13088
rect 153340 12000 153660 13024
rect 153340 11936 153348 12000
rect 153412 11936 153428 12000
rect 153492 11936 153508 12000
rect 153572 11936 153588 12000
rect 153652 11936 153660 12000
rect 153340 11030 153660 11936
rect 153340 10912 153382 11030
rect 153618 10912 153660 11030
rect 153340 10848 153348 10912
rect 153652 10848 153660 10912
rect 153340 10794 153382 10848
rect 153618 10794 153660 10848
rect 153340 9824 153660 10794
rect 153340 9760 153348 9824
rect 153412 9760 153428 9824
rect 153492 9760 153508 9824
rect 153572 9760 153588 9824
rect 153652 9760 153660 9824
rect 153340 8736 153660 9760
rect 153340 8672 153348 8736
rect 153412 8672 153428 8736
rect 153492 8672 153508 8736
rect 153572 8672 153588 8736
rect 153652 8672 153660 8736
rect 153340 8118 153660 8672
rect 153340 7882 153382 8118
rect 153618 7882 153660 8118
rect 153340 7648 153660 7882
rect 153340 7584 153348 7648
rect 153412 7584 153428 7648
rect 153492 7584 153508 7648
rect 153572 7584 153588 7648
rect 153652 7584 153660 7648
rect 153340 6560 153660 7584
rect 153340 6496 153348 6560
rect 153412 6496 153428 6560
rect 153492 6496 153508 6560
rect 153572 6496 153588 6560
rect 153652 6496 153660 6560
rect 153340 5472 153660 6496
rect 153340 5408 153348 5472
rect 153412 5408 153428 5472
rect 153492 5408 153508 5472
rect 153572 5408 153588 5472
rect 153652 5408 153660 5472
rect 153340 5206 153660 5408
rect 153340 4970 153382 5206
rect 153618 4970 153660 5206
rect 153340 4384 153660 4970
rect 153340 4320 153348 4384
rect 153412 4320 153428 4384
rect 153492 4320 153508 4384
rect 153572 4320 153588 4384
rect 153652 4320 153660 4384
rect 153340 3296 153660 4320
rect 153340 3232 153348 3296
rect 153412 3232 153428 3296
rect 153492 3232 153508 3296
rect 153572 3232 153588 3296
rect 153652 3232 153660 3296
rect 153340 2208 153660 3232
rect 153340 2144 153348 2208
rect 153412 2144 153428 2208
rect 153492 2144 153508 2208
rect 153572 2144 153588 2208
rect 153652 2144 153660 2208
rect 153340 274 153660 2144
rect 153340 38 153382 274
rect 153618 38 153660 274
rect 153340 -4 153660 38
rect 191439 15078 191759 15780
rect 191439 14842 191481 15078
rect 191717 14842 191759 15078
rect 191439 13632 191759 14842
rect 191439 13568 191447 13632
rect 191511 13568 191527 13632
rect 191591 13568 191607 13632
rect 191671 13568 191687 13632
rect 191751 13568 191759 13632
rect 191439 12544 191759 13568
rect 191439 12480 191447 12544
rect 191511 12486 191527 12544
rect 191591 12486 191607 12544
rect 191671 12486 191687 12544
rect 191751 12480 191759 12544
rect 191439 12250 191481 12480
rect 191717 12250 191759 12480
rect 191439 11456 191759 12250
rect 191439 11392 191447 11456
rect 191511 11392 191527 11456
rect 191591 11392 191607 11456
rect 191671 11392 191687 11456
rect 191751 11392 191759 11456
rect 191439 10368 191759 11392
rect 191439 10304 191447 10368
rect 191511 10304 191527 10368
rect 191591 10304 191607 10368
rect 191671 10304 191687 10368
rect 191751 10304 191759 10368
rect 191439 9574 191759 10304
rect 191439 9338 191481 9574
rect 191717 9338 191759 9574
rect 191439 9280 191759 9338
rect 191439 9216 191447 9280
rect 191511 9216 191527 9280
rect 191591 9216 191607 9280
rect 191671 9216 191687 9280
rect 191751 9216 191759 9280
rect 191439 8192 191759 9216
rect 191439 8128 191447 8192
rect 191511 8128 191527 8192
rect 191591 8128 191607 8192
rect 191671 8128 191687 8192
rect 191751 8128 191759 8192
rect 191439 7104 191759 8128
rect 191439 7040 191447 7104
rect 191511 7040 191527 7104
rect 191591 7040 191607 7104
rect 191671 7040 191687 7104
rect 191751 7040 191759 7104
rect 191439 6662 191759 7040
rect 191439 6426 191481 6662
rect 191717 6426 191759 6662
rect 191439 6016 191759 6426
rect 191439 5952 191447 6016
rect 191511 5952 191527 6016
rect 191591 5952 191607 6016
rect 191671 5952 191687 6016
rect 191751 5952 191759 6016
rect 191439 4928 191759 5952
rect 191439 4864 191447 4928
rect 191511 4864 191527 4928
rect 191591 4864 191607 4928
rect 191671 4864 191687 4928
rect 191751 4864 191759 4928
rect 191439 3840 191759 4864
rect 191439 3776 191447 3840
rect 191511 3776 191527 3840
rect 191591 3776 191607 3840
rect 191671 3776 191687 3840
rect 191751 3776 191759 3840
rect 191439 3750 191759 3776
rect 191439 3514 191481 3750
rect 191717 3514 191759 3750
rect 191439 2752 191759 3514
rect 191439 2688 191447 2752
rect 191511 2688 191527 2752
rect 191591 2688 191607 2752
rect 191671 2688 191687 2752
rect 191751 2688 191759 2752
rect 191439 934 191759 2688
rect 191439 698 191481 934
rect 191717 698 191759 934
rect 191439 -4 191759 698
rect 229538 15738 229858 15780
rect 229538 15502 229580 15738
rect 229816 15502 229858 15738
rect 229538 13088 229858 15502
rect 229538 13024 229546 13088
rect 229610 13024 229626 13088
rect 229690 13024 229706 13088
rect 229770 13024 229786 13088
rect 229850 13024 229858 13088
rect 229538 12000 229858 13024
rect 229538 11936 229546 12000
rect 229610 11936 229626 12000
rect 229690 11936 229706 12000
rect 229770 11936 229786 12000
rect 229850 11936 229858 12000
rect 229538 11030 229858 11936
rect 229538 10912 229580 11030
rect 229816 10912 229858 11030
rect 229538 10848 229546 10912
rect 229850 10848 229858 10912
rect 229538 10794 229580 10848
rect 229816 10794 229858 10848
rect 229538 9824 229858 10794
rect 229538 9760 229546 9824
rect 229610 9760 229626 9824
rect 229690 9760 229706 9824
rect 229770 9760 229786 9824
rect 229850 9760 229858 9824
rect 229538 8736 229858 9760
rect 229538 8672 229546 8736
rect 229610 8672 229626 8736
rect 229690 8672 229706 8736
rect 229770 8672 229786 8736
rect 229850 8672 229858 8736
rect 229538 8118 229858 8672
rect 229538 7882 229580 8118
rect 229816 7882 229858 8118
rect 229538 7648 229858 7882
rect 229538 7584 229546 7648
rect 229610 7584 229626 7648
rect 229690 7584 229706 7648
rect 229770 7584 229786 7648
rect 229850 7584 229858 7648
rect 229538 6560 229858 7584
rect 229538 6496 229546 6560
rect 229610 6496 229626 6560
rect 229690 6496 229706 6560
rect 229770 6496 229786 6560
rect 229850 6496 229858 6560
rect 229538 5472 229858 6496
rect 229538 5408 229546 5472
rect 229610 5408 229626 5472
rect 229690 5408 229706 5472
rect 229770 5408 229786 5472
rect 229850 5408 229858 5472
rect 229538 5206 229858 5408
rect 229538 4970 229580 5206
rect 229816 4970 229858 5206
rect 229538 4384 229858 4970
rect 229538 4320 229546 4384
rect 229610 4320 229626 4384
rect 229690 4320 229706 4384
rect 229770 4320 229786 4384
rect 229850 4320 229858 4384
rect 229538 3296 229858 4320
rect 229538 3232 229546 3296
rect 229610 3232 229626 3296
rect 229690 3232 229706 3296
rect 229770 3232 229786 3296
rect 229850 3232 229858 3296
rect 229538 2208 229858 3232
rect 229538 2144 229546 2208
rect 229610 2144 229626 2208
rect 229690 2144 229706 2208
rect 229770 2144 229786 2208
rect 229850 2144 229858 2208
rect 229538 274 229858 2144
rect 229538 38 229580 274
rect 229816 38 229858 274
rect 229538 -4 229858 38
rect 267637 15078 267957 15780
rect 307668 15738 307988 15780
rect 307668 15502 307710 15738
rect 307946 15502 307988 15738
rect 267637 14842 267679 15078
rect 267915 14842 267957 15078
rect 267637 13632 267957 14842
rect 267637 13568 267645 13632
rect 267709 13568 267725 13632
rect 267789 13568 267805 13632
rect 267869 13568 267885 13632
rect 267949 13568 267957 13632
rect 267637 12544 267957 13568
rect 267637 12480 267645 12544
rect 267709 12486 267725 12544
rect 267789 12486 267805 12544
rect 267869 12486 267885 12544
rect 267949 12480 267957 12544
rect 267637 12250 267679 12480
rect 267915 12250 267957 12480
rect 267637 11456 267957 12250
rect 267637 11392 267645 11456
rect 267709 11392 267725 11456
rect 267789 11392 267805 11456
rect 267869 11392 267885 11456
rect 267949 11392 267957 11456
rect 267637 10368 267957 11392
rect 267637 10304 267645 10368
rect 267709 10304 267725 10368
rect 267789 10304 267805 10368
rect 267869 10304 267885 10368
rect 267949 10304 267957 10368
rect 267637 9574 267957 10304
rect 267637 9338 267679 9574
rect 267915 9338 267957 9574
rect 267637 9280 267957 9338
rect 267637 9216 267645 9280
rect 267709 9216 267725 9280
rect 267789 9216 267805 9280
rect 267869 9216 267885 9280
rect 267949 9216 267957 9280
rect 267637 8192 267957 9216
rect 267637 8128 267645 8192
rect 267709 8128 267725 8192
rect 267789 8128 267805 8192
rect 267869 8128 267885 8192
rect 267949 8128 267957 8192
rect 267637 7104 267957 8128
rect 267637 7040 267645 7104
rect 267709 7040 267725 7104
rect 267789 7040 267805 7104
rect 267869 7040 267885 7104
rect 267949 7040 267957 7104
rect 267637 6662 267957 7040
rect 267637 6426 267679 6662
rect 267915 6426 267957 6662
rect 267637 6016 267957 6426
rect 267637 5952 267645 6016
rect 267709 5952 267725 6016
rect 267789 5952 267805 6016
rect 267869 5952 267885 6016
rect 267949 5952 267957 6016
rect 267637 4928 267957 5952
rect 267637 4864 267645 4928
rect 267709 4864 267725 4928
rect 267789 4864 267805 4928
rect 267869 4864 267885 4928
rect 267949 4864 267957 4928
rect 267637 3840 267957 4864
rect 267637 3776 267645 3840
rect 267709 3776 267725 3840
rect 267789 3776 267805 3840
rect 267869 3776 267885 3840
rect 267949 3776 267957 3840
rect 267637 3750 267957 3776
rect 267637 3514 267679 3750
rect 267915 3514 267957 3750
rect 267637 2752 267957 3514
rect 267637 2688 267645 2752
rect 267709 2688 267725 2752
rect 267789 2688 267805 2752
rect 267869 2688 267885 2752
rect 267949 2688 267957 2752
rect 267637 934 267957 2688
rect 267637 698 267679 934
rect 267915 698 267957 934
rect 267637 -4 267957 698
rect 307008 15078 307328 15120
rect 307008 14842 307050 15078
rect 307286 14842 307328 15078
rect 307008 12486 307328 14842
rect 307008 12250 307050 12486
rect 307286 12250 307328 12486
rect 307008 9574 307328 12250
rect 307008 9338 307050 9574
rect 307286 9338 307328 9574
rect 307008 6662 307328 9338
rect 307008 6426 307050 6662
rect 307286 6426 307328 6662
rect 307008 3750 307328 6426
rect 307008 3514 307050 3750
rect 307286 3514 307328 3750
rect 307008 934 307328 3514
rect 307008 698 307050 934
rect 307286 698 307328 934
rect 307008 656 307328 698
rect 307668 11030 307988 15502
rect 307668 10794 307710 11030
rect 307946 10794 307988 11030
rect 307668 8118 307988 10794
rect 307668 7882 307710 8118
rect 307946 7882 307988 8118
rect 307668 5206 307988 7882
rect 307668 4970 307710 5206
rect 307946 4970 307988 5206
rect 307668 274 307988 4970
rect 307668 38 307710 274
rect 307946 38 307988 274
rect 307668 -4 307988 38
<< via4 >>
rect -1034 15502 -798 15738
rect -1034 10794 -798 11030
rect -1034 7882 -798 8118
rect -1034 4970 -798 5206
rect -374 14842 -138 15078
rect -374 12250 -138 12486
rect -374 9338 -138 9574
rect -374 6426 -138 6662
rect -374 3514 -138 3750
rect -374 698 -138 934
rect 39085 14842 39321 15078
rect 39085 12480 39115 12486
rect 39115 12480 39131 12486
rect 39131 12480 39195 12486
rect 39195 12480 39211 12486
rect 39211 12480 39275 12486
rect 39275 12480 39291 12486
rect 39291 12480 39321 12486
rect 39085 12250 39321 12480
rect 39085 9338 39321 9574
rect 39085 6426 39321 6662
rect 39085 3514 39321 3750
rect 39085 698 39321 934
rect -1034 38 -798 274
rect 77184 15502 77420 15738
rect 77184 10912 77420 11030
rect 77184 10848 77214 10912
rect 77214 10848 77230 10912
rect 77230 10848 77294 10912
rect 77294 10848 77310 10912
rect 77310 10848 77374 10912
rect 77374 10848 77390 10912
rect 77390 10848 77420 10912
rect 77184 10794 77420 10848
rect 77184 7882 77420 8118
rect 77184 4970 77420 5206
rect 77184 38 77420 274
rect 115283 14842 115519 15078
rect 115283 12480 115313 12486
rect 115313 12480 115329 12486
rect 115329 12480 115393 12486
rect 115393 12480 115409 12486
rect 115409 12480 115473 12486
rect 115473 12480 115489 12486
rect 115489 12480 115519 12486
rect 115283 12250 115519 12480
rect 115283 9338 115519 9574
rect 115283 6426 115519 6662
rect 115283 3514 115519 3750
rect 115283 698 115519 934
rect 153382 15502 153618 15738
rect 153382 10912 153618 11030
rect 153382 10848 153412 10912
rect 153412 10848 153428 10912
rect 153428 10848 153492 10912
rect 153492 10848 153508 10912
rect 153508 10848 153572 10912
rect 153572 10848 153588 10912
rect 153588 10848 153618 10912
rect 153382 10794 153618 10848
rect 153382 7882 153618 8118
rect 153382 4970 153618 5206
rect 153382 38 153618 274
rect 191481 14842 191717 15078
rect 191481 12480 191511 12486
rect 191511 12480 191527 12486
rect 191527 12480 191591 12486
rect 191591 12480 191607 12486
rect 191607 12480 191671 12486
rect 191671 12480 191687 12486
rect 191687 12480 191717 12486
rect 191481 12250 191717 12480
rect 191481 9338 191717 9574
rect 191481 6426 191717 6662
rect 191481 3514 191717 3750
rect 191481 698 191717 934
rect 229580 15502 229816 15738
rect 229580 10912 229816 11030
rect 229580 10848 229610 10912
rect 229610 10848 229626 10912
rect 229626 10848 229690 10912
rect 229690 10848 229706 10912
rect 229706 10848 229770 10912
rect 229770 10848 229786 10912
rect 229786 10848 229816 10912
rect 229580 10794 229816 10848
rect 229580 7882 229816 8118
rect 229580 4970 229816 5206
rect 229580 38 229816 274
rect 307710 15502 307946 15738
rect 267679 14842 267915 15078
rect 267679 12480 267709 12486
rect 267709 12480 267725 12486
rect 267725 12480 267789 12486
rect 267789 12480 267805 12486
rect 267805 12480 267869 12486
rect 267869 12480 267885 12486
rect 267885 12480 267915 12486
rect 267679 12250 267915 12480
rect 267679 9338 267915 9574
rect 267679 6426 267915 6662
rect 267679 3514 267915 3750
rect 267679 698 267915 934
rect 307050 14842 307286 15078
rect 307050 12250 307286 12486
rect 307050 9338 307286 9574
rect 307050 6426 307286 6662
rect 307050 3514 307286 3750
rect 307050 698 307286 934
rect 307710 10794 307946 11030
rect 307710 7882 307946 8118
rect 307710 4970 307946 5206
rect 307710 38 307946 274
<< metal5 >>
rect -1076 15738 307988 15780
rect -1076 15502 -1034 15738
rect -798 15502 77184 15738
rect 77420 15502 153382 15738
rect 153618 15502 229580 15738
rect 229816 15502 307710 15738
rect 307946 15502 307988 15738
rect -1076 15460 307988 15502
rect -416 15078 307328 15120
rect -416 14842 -374 15078
rect -138 14842 39085 15078
rect 39321 14842 115283 15078
rect 115519 14842 191481 15078
rect 191717 14842 267679 15078
rect 267915 14842 307050 15078
rect 307286 14842 307328 15078
rect -416 14800 307328 14842
rect -1076 12486 307988 12528
rect -1076 12250 -374 12486
rect -138 12250 39085 12486
rect 39321 12250 115283 12486
rect 115519 12250 191481 12486
rect 191717 12250 267679 12486
rect 267915 12250 307050 12486
rect 307286 12250 307988 12486
rect -1076 12208 307988 12250
rect -1076 11030 307988 11072
rect -1076 10794 -1034 11030
rect -798 10794 77184 11030
rect 77420 10794 153382 11030
rect 153618 10794 229580 11030
rect 229816 10794 307710 11030
rect 307946 10794 307988 11030
rect -1076 10752 307988 10794
rect -1076 9574 307988 9616
rect -1076 9338 -374 9574
rect -138 9338 39085 9574
rect 39321 9338 115283 9574
rect 115519 9338 191481 9574
rect 191717 9338 267679 9574
rect 267915 9338 307050 9574
rect 307286 9338 307988 9574
rect -1076 9296 307988 9338
rect -1076 8118 307988 8160
rect -1076 7882 -1034 8118
rect -798 7882 77184 8118
rect 77420 7882 153382 8118
rect 153618 7882 229580 8118
rect 229816 7882 307710 8118
rect 307946 7882 307988 8118
rect -1076 7840 307988 7882
rect -1076 6662 307988 6704
rect -1076 6426 -374 6662
rect -138 6426 39085 6662
rect 39321 6426 115283 6662
rect 115519 6426 191481 6662
rect 191717 6426 267679 6662
rect 267915 6426 307050 6662
rect 307286 6426 307988 6662
rect -1076 6384 307988 6426
rect -1076 5206 307988 5248
rect -1076 4970 -1034 5206
rect -798 4970 77184 5206
rect 77420 4970 153382 5206
rect 153618 4970 229580 5206
rect 229816 4970 307710 5206
rect 307946 4970 307988 5206
rect -1076 4928 307988 4970
rect -1076 3750 307988 3792
rect -1076 3514 -374 3750
rect -138 3514 39085 3750
rect 39321 3514 115283 3750
rect 115519 3514 191481 3750
rect 191717 3514 267679 3750
rect 267915 3514 307050 3750
rect 307286 3514 307988 3750
rect -1076 3472 307988 3514
rect -416 934 307328 976
rect -416 698 -374 934
rect -138 698 39085 934
rect 39321 698 115283 934
rect 115519 698 191481 934
rect 191717 698 267679 934
rect 267915 698 307050 934
rect 307286 698 307328 934
rect -416 656 307328 698
rect -1076 274 307988 316
rect -1076 38 -1034 274
rect -798 38 77184 274
rect 77420 38 153382 274
rect 153618 38 229580 274
rect 229816 38 307710 274
rect 307946 38 307988 274
rect -1076 -4 307988 38
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 43516 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1649977179
transform 1 0 55936 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1649977179
transform 1 0 154100 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1649977179
transform 1 0 153732 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1649977179
transform 1 0 155940 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1649977179
transform 1 0 153364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1649977179
transform 1 0 156308 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1649977179
transform 1 0 152996 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1649977179
transform 1 0 156676 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1649977179
transform 1 0 152628 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1649977179
transform 1 0 157044 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1649977179
transform 1 0 152260 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1649977179
transform -1 0 303508 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1649977179
transform -1 0 303140 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1649977179
transform -1 0 302312 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1649977179
transform -1 0 301944 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1649977179
transform -1 0 301576 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1649977179
transform 1 0 305348 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1649977179
transform 1 0 304888 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1649977179
transform 1 0 305348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1649977179
transform 1 0 304888 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1649977179
transform 1 0 305348 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1649977179
transform 1 0 1840 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1649977179
transform 1 0 2208 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1649977179
transform 1 0 2576 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1649977179
transform 1 0 2944 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1649977179
transform 1 0 268456 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1649977179
transform 1 0 252264 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1649977179
transform 1 0 197984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1649977179
transform 1 0 197800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1649977179
transform 1 0 295872 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1649977179
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1649977179
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1649977179
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1649977179
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1649977179
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1649977179
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1649977179
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1649977179
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1649977179
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1649977179
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1649977179
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1649977179
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1649977179
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1649977179
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1649977179
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1649977179
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1649977179
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1649977179
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1649977179
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1649977179
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1649977179
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1649977179
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1649977179
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1649977179
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1649977179
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1649977179
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_449
timestamp 1649977179
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_461
timestamp 1649977179
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1649977179
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1649977179
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1649977179
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1649977179
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_505
timestamp 1649977179
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_517
timestamp 1649977179
transform 1 0 48668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_529
timestamp 1649977179
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_533
timestamp 1649977179
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_545
timestamp 1649977179
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1649977179
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_561
timestamp 1649977179
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_573
timestamp 1649977179
transform 1 0 53820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_585
timestamp 1649977179
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_589
timestamp 1649977179
transform 1 0 55292 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_601
timestamp 1649977179
transform 1 0 56396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_613
timestamp 1649977179
transform 1 0 57500 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_617
timestamp 1649977179
transform 1 0 57868 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_629
timestamp 1649977179
transform 1 0 58972 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_641
timestamp 1649977179
transform 1 0 60076 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_645
timestamp 1649977179
transform 1 0 60444 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_657
timestamp 1649977179
transform 1 0 61548 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_669
timestamp 1649977179
transform 1 0 62652 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_673
timestamp 1649977179
transform 1 0 63020 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_685
timestamp 1649977179
transform 1 0 64124 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_697
timestamp 1649977179
transform 1 0 65228 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_701
timestamp 1649977179
transform 1 0 65596 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_713
timestamp 1649977179
transform 1 0 66700 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_725
timestamp 1649977179
transform 1 0 67804 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_729
timestamp 1649977179
transform 1 0 68172 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_741
timestamp 1649977179
transform 1 0 69276 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_753
timestamp 1649977179
transform 1 0 70380 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_757
timestamp 1649977179
transform 1 0 70748 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_769
timestamp 1649977179
transform 1 0 71852 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_781
timestamp 1649977179
transform 1 0 72956 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_785
timestamp 1649977179
transform 1 0 73324 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_797
timestamp 1649977179
transform 1 0 74428 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_809
timestamp 1649977179
transform 1 0 75532 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_813
timestamp 1649977179
transform 1 0 75900 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_825
timestamp 1649977179
transform 1 0 77004 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_837
timestamp 1649977179
transform 1 0 78108 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_841
timestamp 1649977179
transform 1 0 78476 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_853
timestamp 1649977179
transform 1 0 79580 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_865
timestamp 1649977179
transform 1 0 80684 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_869
timestamp 1649977179
transform 1 0 81052 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_881
timestamp 1649977179
transform 1 0 82156 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_893
timestamp 1649977179
transform 1 0 83260 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_897
timestamp 1649977179
transform 1 0 83628 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_909
timestamp 1649977179
transform 1 0 84732 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_921
timestamp 1649977179
transform 1 0 85836 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_925
timestamp 1649977179
transform 1 0 86204 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_937
timestamp 1649977179
transform 1 0 87308 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_949
timestamp 1649977179
transform 1 0 88412 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_953
timestamp 1649977179
transform 1 0 88780 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_965
timestamp 1649977179
transform 1 0 89884 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_977
timestamp 1649977179
transform 1 0 90988 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_981
timestamp 1649977179
transform 1 0 91356 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_993
timestamp 1649977179
transform 1 0 92460 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1005
timestamp 1649977179
transform 1 0 93564 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1009
timestamp 1649977179
transform 1 0 93932 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1021
timestamp 1649977179
transform 1 0 95036 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1033
timestamp 1649977179
transform 1 0 96140 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1037
timestamp 1649977179
transform 1 0 96508 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1049
timestamp 1649977179
transform 1 0 97612 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1061
timestamp 1649977179
transform 1 0 98716 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1065
timestamp 1649977179
transform 1 0 99084 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1077
timestamp 1649977179
transform 1 0 100188 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1089
timestamp 1649977179
transform 1 0 101292 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1093
timestamp 1649977179
transform 1 0 101660 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1105
timestamp 1649977179
transform 1 0 102764 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1117
timestamp 1649977179
transform 1 0 103868 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1121
timestamp 1649977179
transform 1 0 104236 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1133
timestamp 1649977179
transform 1 0 105340 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1145
timestamp 1649977179
transform 1 0 106444 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1149
timestamp 1649977179
transform 1 0 106812 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1161
timestamp 1649977179
transform 1 0 107916 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1173
timestamp 1649977179
transform 1 0 109020 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1177
timestamp 1649977179
transform 1 0 109388 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1189
timestamp 1649977179
transform 1 0 110492 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1201
timestamp 1649977179
transform 1 0 111596 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1205
timestamp 1649977179
transform 1 0 111964 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1217
timestamp 1649977179
transform 1 0 113068 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1229
timestamp 1649977179
transform 1 0 114172 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1233
timestamp 1649977179
transform 1 0 114540 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1245
timestamp 1649977179
transform 1 0 115644 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1257
timestamp 1649977179
transform 1 0 116748 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1261
timestamp 1649977179
transform 1 0 117116 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1273
timestamp 1649977179
transform 1 0 118220 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1285
timestamp 1649977179
transform 1 0 119324 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1289
timestamp 1649977179
transform 1 0 119692 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1301
timestamp 1649977179
transform 1 0 120796 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1313
timestamp 1649977179
transform 1 0 121900 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1317
timestamp 1649977179
transform 1 0 122268 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1329
timestamp 1649977179
transform 1 0 123372 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1341
timestamp 1649977179
transform 1 0 124476 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1345
timestamp 1649977179
transform 1 0 124844 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1357
timestamp 1649977179
transform 1 0 125948 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1369
timestamp 1649977179
transform 1 0 127052 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1373
timestamp 1649977179
transform 1 0 127420 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1385
timestamp 1649977179
transform 1 0 128524 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1397
timestamp 1649977179
transform 1 0 129628 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1401
timestamp 1649977179
transform 1 0 129996 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1413
timestamp 1649977179
transform 1 0 131100 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1425
timestamp 1649977179
transform 1 0 132204 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1429
timestamp 1649977179
transform 1 0 132572 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1441
timestamp 1649977179
transform 1 0 133676 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1453
timestamp 1649977179
transform 1 0 134780 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1457
timestamp 1649977179
transform 1 0 135148 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1469
timestamp 1649977179
transform 1 0 136252 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1481
timestamp 1649977179
transform 1 0 137356 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1485
timestamp 1649977179
transform 1 0 137724 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1497
timestamp 1649977179
transform 1 0 138828 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1509
timestamp 1649977179
transform 1 0 139932 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1513
timestamp 1649977179
transform 1 0 140300 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1525
timestamp 1649977179
transform 1 0 141404 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1537
timestamp 1649977179
transform 1 0 142508 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1541
timestamp 1649977179
transform 1 0 142876 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1553
timestamp 1649977179
transform 1 0 143980 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1565
timestamp 1649977179
transform 1 0 145084 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1569
timestamp 1649977179
transform 1 0 145452 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1581
timestamp 1649977179
transform 1 0 146556 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1593
timestamp 1649977179
transform 1 0 147660 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1597
timestamp 1649977179
transform 1 0 148028 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1609
timestamp 1649977179
transform 1 0 149132 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1621
timestamp 1649977179
transform 1 0 150236 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1625
timestamp 1649977179
transform 1 0 150604 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1637
timestamp 1649977179
transform 1 0 151708 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1649
timestamp 1649977179
transform 1 0 152812 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1653
timestamp 1649977179
transform 1 0 153180 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1665
timestamp 1649977179
transform 1 0 154284 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1677
timestamp 1649977179
transform 1 0 155388 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1681
timestamp 1649977179
transform 1 0 155756 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1693
timestamp 1649977179
transform 1 0 156860 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1705
timestamp 1649977179
transform 1 0 157964 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1709
timestamp 1649977179
transform 1 0 158332 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1721
timestamp 1649977179
transform 1 0 159436 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1733
timestamp 1649977179
transform 1 0 160540 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1737
timestamp 1649977179
transform 1 0 160908 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1749
timestamp 1649977179
transform 1 0 162012 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1761
timestamp 1649977179
transform 1 0 163116 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1765
timestamp 1649977179
transform 1 0 163484 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1777
timestamp 1649977179
transform 1 0 164588 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1789
timestamp 1649977179
transform 1 0 165692 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1793
timestamp 1649977179
transform 1 0 166060 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1805
timestamp 1649977179
transform 1 0 167164 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1817
timestamp 1649977179
transform 1 0 168268 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1821
timestamp 1649977179
transform 1 0 168636 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1833
timestamp 1649977179
transform 1 0 169740 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1845
timestamp 1649977179
transform 1 0 170844 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1849
timestamp 1649977179
transform 1 0 171212 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1861
timestamp 1649977179
transform 1 0 172316 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1873
timestamp 1649977179
transform 1 0 173420 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1877
timestamp 1649977179
transform 1 0 173788 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1889
timestamp 1649977179
transform 1 0 174892 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1901
timestamp 1649977179
transform 1 0 175996 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1905
timestamp 1649977179
transform 1 0 176364 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1917
timestamp 1649977179
transform 1 0 177468 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1929
timestamp 1649977179
transform 1 0 178572 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1933
timestamp 1649977179
transform 1 0 178940 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1945
timestamp 1649977179
transform 1 0 180044 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1957
timestamp 1649977179
transform 1 0 181148 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1961
timestamp 1649977179
transform 1 0 181516 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1973
timestamp 1649977179
transform 1 0 182620 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1985
timestamp 1649977179
transform 1 0 183724 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1989
timestamp 1649977179
transform 1 0 184092 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2001
timestamp 1649977179
transform 1 0 185196 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2013
timestamp 1649977179
transform 1 0 186300 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2017
timestamp 1649977179
transform 1 0 186668 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2029
timestamp 1649977179
transform 1 0 187772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2041
timestamp 1649977179
transform 1 0 188876 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2045
timestamp 1649977179
transform 1 0 189244 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2057
timestamp 1649977179
transform 1 0 190348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2069
timestamp 1649977179
transform 1 0 191452 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2073
timestamp 1649977179
transform 1 0 191820 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2085
timestamp 1649977179
transform 1 0 192924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2097
timestamp 1649977179
transform 1 0 194028 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2101
timestamp 1649977179
transform 1 0 194396 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2113
timestamp 1649977179
transform 1 0 195500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2125
timestamp 1649977179
transform 1 0 196604 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2129
timestamp 1649977179
transform 1 0 196972 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2141
timestamp 1649977179
transform 1 0 198076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2153
timestamp 1649977179
transform 1 0 199180 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2157
timestamp 1649977179
transform 1 0 199548 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2169
timestamp 1649977179
transform 1 0 200652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2181
timestamp 1649977179
transform 1 0 201756 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2185
timestamp 1649977179
transform 1 0 202124 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2197
timestamp 1649977179
transform 1 0 203228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2209
timestamp 1649977179
transform 1 0 204332 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2213
timestamp 1649977179
transform 1 0 204700 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2225
timestamp 1649977179
transform 1 0 205804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2237
timestamp 1649977179
transform 1 0 206908 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2241
timestamp 1649977179
transform 1 0 207276 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2253
timestamp 1649977179
transform 1 0 208380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2265
timestamp 1649977179
transform 1 0 209484 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2269
timestamp 1649977179
transform 1 0 209852 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2281
timestamp 1649977179
transform 1 0 210956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2293
timestamp 1649977179
transform 1 0 212060 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2297
timestamp 1649977179
transform 1 0 212428 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2309
timestamp 1649977179
transform 1 0 213532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2321
timestamp 1649977179
transform 1 0 214636 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2325
timestamp 1649977179
transform 1 0 215004 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2337
timestamp 1649977179
transform 1 0 216108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2349
timestamp 1649977179
transform 1 0 217212 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2353
timestamp 1649977179
transform 1 0 217580 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2365
timestamp 1649977179
transform 1 0 218684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2377
timestamp 1649977179
transform 1 0 219788 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2381
timestamp 1649977179
transform 1 0 220156 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2393
timestamp 1649977179
transform 1 0 221260 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2405
timestamp 1649977179
transform 1 0 222364 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2409
timestamp 1649977179
transform 1 0 222732 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2421
timestamp 1649977179
transform 1 0 223836 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2433
timestamp 1649977179
transform 1 0 224940 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2437
timestamp 1649977179
transform 1 0 225308 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2449
timestamp 1649977179
transform 1 0 226412 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2461
timestamp 1649977179
transform 1 0 227516 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2465
timestamp 1649977179
transform 1 0 227884 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2477
timestamp 1649977179
transform 1 0 228988 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2489
timestamp 1649977179
transform 1 0 230092 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2493
timestamp 1649977179
transform 1 0 230460 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2505
timestamp 1649977179
transform 1 0 231564 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2517
timestamp 1649977179
transform 1 0 232668 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2521
timestamp 1649977179
transform 1 0 233036 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2533
timestamp 1649977179
transform 1 0 234140 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2545
timestamp 1649977179
transform 1 0 235244 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2549
timestamp 1649977179
transform 1 0 235612 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2561
timestamp 1649977179
transform 1 0 236716 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2573
timestamp 1649977179
transform 1 0 237820 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2577
timestamp 1649977179
transform 1 0 238188 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2589
timestamp 1649977179
transform 1 0 239292 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2601
timestamp 1649977179
transform 1 0 240396 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2605
timestamp 1649977179
transform 1 0 240764 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2617
timestamp 1649977179
transform 1 0 241868 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2629
timestamp 1649977179
transform 1 0 242972 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2633
timestamp 1649977179
transform 1 0 243340 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2645
timestamp 1649977179
transform 1 0 244444 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2657
timestamp 1649977179
transform 1 0 245548 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2661
timestamp 1649977179
transform 1 0 245916 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2673
timestamp 1649977179
transform 1 0 247020 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2685
timestamp 1649977179
transform 1 0 248124 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2689
timestamp 1649977179
transform 1 0 248492 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2701
timestamp 1649977179
transform 1 0 249596 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2713
timestamp 1649977179
transform 1 0 250700 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2717
timestamp 1649977179
transform 1 0 251068 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2729
timestamp 1649977179
transform 1 0 252172 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2741
timestamp 1649977179
transform 1 0 253276 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2745
timestamp 1649977179
transform 1 0 253644 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2757
timestamp 1649977179
transform 1 0 254748 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2769
timestamp 1649977179
transform 1 0 255852 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2773
timestamp 1649977179
transform 1 0 256220 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2785
timestamp 1649977179
transform 1 0 257324 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2797
timestamp 1649977179
transform 1 0 258428 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2801
timestamp 1649977179
transform 1 0 258796 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2813
timestamp 1649977179
transform 1 0 259900 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2825
timestamp 1649977179
transform 1 0 261004 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2829
timestamp 1649977179
transform 1 0 261372 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2841
timestamp 1649977179
transform 1 0 262476 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2853
timestamp 1649977179
transform 1 0 263580 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2857
timestamp 1649977179
transform 1 0 263948 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2869
timestamp 1649977179
transform 1 0 265052 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2881
timestamp 1649977179
transform 1 0 266156 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2885
timestamp 1649977179
transform 1 0 266524 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2897
timestamp 1649977179
transform 1 0 267628 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2909
timestamp 1649977179
transform 1 0 268732 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2913
timestamp 1649977179
transform 1 0 269100 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2925
timestamp 1649977179
transform 1 0 270204 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2937
timestamp 1649977179
transform 1 0 271308 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2941
timestamp 1649977179
transform 1 0 271676 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2953
timestamp 1649977179
transform 1 0 272780 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2965
timestamp 1649977179
transform 1 0 273884 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2969
timestamp 1649977179
transform 1 0 274252 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2981
timestamp 1649977179
transform 1 0 275356 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2993
timestamp 1649977179
transform 1 0 276460 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2997
timestamp 1649977179
transform 1 0 276828 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3009
timestamp 1649977179
transform 1 0 277932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3021
timestamp 1649977179
transform 1 0 279036 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3025
timestamp 1649977179
transform 1 0 279404 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3037
timestamp 1649977179
transform 1 0 280508 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3049
timestamp 1649977179
transform 1 0 281612 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3053
timestamp 1649977179
transform 1 0 281980 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3065
timestamp 1649977179
transform 1 0 283084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3077
timestamp 1649977179
transform 1 0 284188 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3081
timestamp 1649977179
transform 1 0 284556 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3093
timestamp 1649977179
transform 1 0 285660 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3105
timestamp 1649977179
transform 1 0 286764 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3109
timestamp 1649977179
transform 1 0 287132 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3121
timestamp 1649977179
transform 1 0 288236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3133
timestamp 1649977179
transform 1 0 289340 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3137
timestamp 1649977179
transform 1 0 289708 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3149
timestamp 1649977179
transform 1 0 290812 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3161
timestamp 1649977179
transform 1 0 291916 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3165
timestamp 1649977179
transform 1 0 292284 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3177
timestamp 1649977179
transform 1 0 293388 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3189
timestamp 1649977179
transform 1 0 294492 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3193
timestamp 1649977179
transform 1 0 294860 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3205
timestamp 1649977179
transform 1 0 295964 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3217
timestamp 1649977179
transform 1 0 297068 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3221
timestamp 1649977179
transform 1 0 297436 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3233
timestamp 1649977179
transform 1 0 298540 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3245
timestamp 1649977179
transform 1 0 299644 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3249
timestamp 1649977179
transform 1 0 300012 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3261
timestamp 1649977179
transform 1 0 301116 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3273
timestamp 1649977179
transform 1 0 302220 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3277
timestamp 1649977179
transform 1 0 302588 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3289
timestamp 1649977179
transform 1 0 303692 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3301
timestamp 1649977179
transform 1 0 304796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3305 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 305164 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1649977179
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1649977179
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1649977179
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1649977179
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1649977179
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1649977179
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1649977179
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1649977179
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1649977179
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1649977179
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1649977179
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1649977179
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1649977179
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1649977179
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1649977179
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1649977179
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1649977179
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1649977179
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1649977179
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1649977179
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1649977179
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1649977179
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1649977179
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1649977179
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1649977179
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1649977179
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1649977179
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1649977179
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1649977179
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1649977179
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1649977179
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1649977179
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1649977179
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1649977179
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1649977179
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_517
timestamp 1649977179
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_529
timestamp 1649977179
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_541
timestamp 1649977179
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 1649977179
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1649977179
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_561
timestamp 1649977179
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_573
timestamp 1649977179
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_585
timestamp 1649977179
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_597
timestamp 1649977179
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 1649977179
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1649977179
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_617
timestamp 1649977179
transform 1 0 57868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_629
timestamp 1649977179
transform 1 0 58972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_641
timestamp 1649977179
transform 1 0 60076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_653
timestamp 1649977179
transform 1 0 61180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_665
timestamp 1649977179
transform 1 0 62284 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 1649977179
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_673
timestamp 1649977179
transform 1 0 63020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_685
timestamp 1649977179
transform 1 0 64124 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_697
timestamp 1649977179
transform 1 0 65228 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_709
timestamp 1649977179
transform 1 0 66332 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_721
timestamp 1649977179
transform 1 0 67436 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 1649977179
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_729
timestamp 1649977179
transform 1 0 68172 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_741
timestamp 1649977179
transform 1 0 69276 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_753
timestamp 1649977179
transform 1 0 70380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_765
timestamp 1649977179
transform 1 0 71484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_777
timestamp 1649977179
transform 1 0 72588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_783
timestamp 1649977179
transform 1 0 73140 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_785
timestamp 1649977179
transform 1 0 73324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_797
timestamp 1649977179
transform 1 0 74428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_809
timestamp 1649977179
transform 1 0 75532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_821
timestamp 1649977179
transform 1 0 76636 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_833
timestamp 1649977179
transform 1 0 77740 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_839
timestamp 1649977179
transform 1 0 78292 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_841
timestamp 1649977179
transform 1 0 78476 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_853
timestamp 1649977179
transform 1 0 79580 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_865
timestamp 1649977179
transform 1 0 80684 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_877
timestamp 1649977179
transform 1 0 81788 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_889
timestamp 1649977179
transform 1 0 82892 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_895
timestamp 1649977179
transform 1 0 83444 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_897
timestamp 1649977179
transform 1 0 83628 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_909
timestamp 1649977179
transform 1 0 84732 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_921
timestamp 1649977179
transform 1 0 85836 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_933
timestamp 1649977179
transform 1 0 86940 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_945
timestamp 1649977179
transform 1 0 88044 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_951
timestamp 1649977179
transform 1 0 88596 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_953
timestamp 1649977179
transform 1 0 88780 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_965
timestamp 1649977179
transform 1 0 89884 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_977
timestamp 1649977179
transform 1 0 90988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_989
timestamp 1649977179
transform 1 0 92092 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1001
timestamp 1649977179
transform 1 0 93196 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1007
timestamp 1649977179
transform 1 0 93748 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1009
timestamp 1649977179
transform 1 0 93932 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1021
timestamp 1649977179
transform 1 0 95036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1033
timestamp 1649977179
transform 1 0 96140 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1045
timestamp 1649977179
transform 1 0 97244 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1057
timestamp 1649977179
transform 1 0 98348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1063
timestamp 1649977179
transform 1 0 98900 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1065
timestamp 1649977179
transform 1 0 99084 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1077
timestamp 1649977179
transform 1 0 100188 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1089
timestamp 1649977179
transform 1 0 101292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1101
timestamp 1649977179
transform 1 0 102396 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1113
timestamp 1649977179
transform 1 0 103500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1119
timestamp 1649977179
transform 1 0 104052 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1121
timestamp 1649977179
transform 1 0 104236 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1133
timestamp 1649977179
transform 1 0 105340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1145
timestamp 1649977179
transform 1 0 106444 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1157
timestamp 1649977179
transform 1 0 107548 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1169
timestamp 1649977179
transform 1 0 108652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1175
timestamp 1649977179
transform 1 0 109204 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1177
timestamp 1649977179
transform 1 0 109388 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1189
timestamp 1649977179
transform 1 0 110492 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1201
timestamp 1649977179
transform 1 0 111596 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1213
timestamp 1649977179
transform 1 0 112700 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1225
timestamp 1649977179
transform 1 0 113804 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1231
timestamp 1649977179
transform 1 0 114356 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1233
timestamp 1649977179
transform 1 0 114540 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1245
timestamp 1649977179
transform 1 0 115644 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1257
timestamp 1649977179
transform 1 0 116748 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1269
timestamp 1649977179
transform 1 0 117852 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1281
timestamp 1649977179
transform 1 0 118956 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1287
timestamp 1649977179
transform 1 0 119508 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1289
timestamp 1649977179
transform 1 0 119692 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1301
timestamp 1649977179
transform 1 0 120796 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1313
timestamp 1649977179
transform 1 0 121900 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1325
timestamp 1649977179
transform 1 0 123004 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1337
timestamp 1649977179
transform 1 0 124108 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1343
timestamp 1649977179
transform 1 0 124660 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1345
timestamp 1649977179
transform 1 0 124844 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1357
timestamp 1649977179
transform 1 0 125948 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1369
timestamp 1649977179
transform 1 0 127052 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1381
timestamp 1649977179
transform 1 0 128156 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1393
timestamp 1649977179
transform 1 0 129260 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1399
timestamp 1649977179
transform 1 0 129812 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1401
timestamp 1649977179
transform 1 0 129996 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1413
timestamp 1649977179
transform 1 0 131100 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1425
timestamp 1649977179
transform 1 0 132204 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1437
timestamp 1649977179
transform 1 0 133308 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1449
timestamp 1649977179
transform 1 0 134412 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1455
timestamp 1649977179
transform 1 0 134964 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1457
timestamp 1649977179
transform 1 0 135148 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1469
timestamp 1649977179
transform 1 0 136252 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1481
timestamp 1649977179
transform 1 0 137356 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1493
timestamp 1649977179
transform 1 0 138460 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1505
timestamp 1649977179
transform 1 0 139564 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1511
timestamp 1649977179
transform 1 0 140116 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1513
timestamp 1649977179
transform 1 0 140300 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1525
timestamp 1649977179
transform 1 0 141404 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1537
timestamp 1649977179
transform 1 0 142508 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1549
timestamp 1649977179
transform 1 0 143612 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1561
timestamp 1649977179
transform 1 0 144716 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1567
timestamp 1649977179
transform 1 0 145268 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1569
timestamp 1649977179
transform 1 0 145452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1581
timestamp 1649977179
transform 1 0 146556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1593
timestamp 1649977179
transform 1 0 147660 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1605
timestamp 1649977179
transform 1 0 148764 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1617
timestamp 1649977179
transform 1 0 149868 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1623
timestamp 1649977179
transform 1 0 150420 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1625
timestamp 1649977179
transform 1 0 150604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1637
timestamp 1649977179
transform 1 0 151708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1649
timestamp 1649977179
transform 1 0 152812 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1661
timestamp 1649977179
transform 1 0 153916 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1673
timestamp 1649977179
transform 1 0 155020 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1679
timestamp 1649977179
transform 1 0 155572 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1681
timestamp 1649977179
transform 1 0 155756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1693
timestamp 1649977179
transform 1 0 156860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1705
timestamp 1649977179
transform 1 0 157964 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1717
timestamp 1649977179
transform 1 0 159068 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1729
timestamp 1649977179
transform 1 0 160172 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1735
timestamp 1649977179
transform 1 0 160724 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1737
timestamp 1649977179
transform 1 0 160908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1749
timestamp 1649977179
transform 1 0 162012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1761
timestamp 1649977179
transform 1 0 163116 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1773
timestamp 1649977179
transform 1 0 164220 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1785
timestamp 1649977179
transform 1 0 165324 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1791
timestamp 1649977179
transform 1 0 165876 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1793
timestamp 1649977179
transform 1 0 166060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1805
timestamp 1649977179
transform 1 0 167164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1817
timestamp 1649977179
transform 1 0 168268 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1829
timestamp 1649977179
transform 1 0 169372 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1841
timestamp 1649977179
transform 1 0 170476 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1847
timestamp 1649977179
transform 1 0 171028 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1849
timestamp 1649977179
transform 1 0 171212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1861
timestamp 1649977179
transform 1 0 172316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1873
timestamp 1649977179
transform 1 0 173420 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1885
timestamp 1649977179
transform 1 0 174524 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1897
timestamp 1649977179
transform 1 0 175628 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1903
timestamp 1649977179
transform 1 0 176180 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1905
timestamp 1649977179
transform 1 0 176364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1917
timestamp 1649977179
transform 1 0 177468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1929
timestamp 1649977179
transform 1 0 178572 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1941
timestamp 1649977179
transform 1 0 179676 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1953
timestamp 1649977179
transform 1 0 180780 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1959
timestamp 1649977179
transform 1 0 181332 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1961
timestamp 1649977179
transform 1 0 181516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1973
timestamp 1649977179
transform 1 0 182620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1985
timestamp 1649977179
transform 1 0 183724 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1997
timestamp 1649977179
transform 1 0 184828 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2009
timestamp 1649977179
transform 1 0 185932 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2015
timestamp 1649977179
transform 1 0 186484 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2017
timestamp 1649977179
transform 1 0 186668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2029
timestamp 1649977179
transform 1 0 187772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2041
timestamp 1649977179
transform 1 0 188876 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2053
timestamp 1649977179
transform 1 0 189980 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2065
timestamp 1649977179
transform 1 0 191084 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2071
timestamp 1649977179
transform 1 0 191636 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2073
timestamp 1649977179
transform 1 0 191820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2085
timestamp 1649977179
transform 1 0 192924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2097
timestamp 1649977179
transform 1 0 194028 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2109
timestamp 1649977179
transform 1 0 195132 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2121
timestamp 1649977179
transform 1 0 196236 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2127
timestamp 1649977179
transform 1 0 196788 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2129
timestamp 1649977179
transform 1 0 196972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2141
timestamp 1649977179
transform 1 0 198076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2153
timestamp 1649977179
transform 1 0 199180 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2165
timestamp 1649977179
transform 1 0 200284 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2177
timestamp 1649977179
transform 1 0 201388 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2183
timestamp 1649977179
transform 1 0 201940 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2185
timestamp 1649977179
transform 1 0 202124 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2197
timestamp 1649977179
transform 1 0 203228 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2209
timestamp 1649977179
transform 1 0 204332 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2221
timestamp 1649977179
transform 1 0 205436 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2233
timestamp 1649977179
transform 1 0 206540 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2239
timestamp 1649977179
transform 1 0 207092 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2241
timestamp 1649977179
transform 1 0 207276 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2253
timestamp 1649977179
transform 1 0 208380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2265
timestamp 1649977179
transform 1 0 209484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2277
timestamp 1649977179
transform 1 0 210588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2289
timestamp 1649977179
transform 1 0 211692 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2295
timestamp 1649977179
transform 1 0 212244 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2297
timestamp 1649977179
transform 1 0 212428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2309
timestamp 1649977179
transform 1 0 213532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2321
timestamp 1649977179
transform 1 0 214636 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2333
timestamp 1649977179
transform 1 0 215740 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2345
timestamp 1649977179
transform 1 0 216844 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2351
timestamp 1649977179
transform 1 0 217396 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2353
timestamp 1649977179
transform 1 0 217580 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2365
timestamp 1649977179
transform 1 0 218684 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2377
timestamp 1649977179
transform 1 0 219788 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2389
timestamp 1649977179
transform 1 0 220892 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2401
timestamp 1649977179
transform 1 0 221996 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2407
timestamp 1649977179
transform 1 0 222548 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2409
timestamp 1649977179
transform 1 0 222732 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2421
timestamp 1649977179
transform 1 0 223836 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2433
timestamp 1649977179
transform 1 0 224940 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2445
timestamp 1649977179
transform 1 0 226044 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2457
timestamp 1649977179
transform 1 0 227148 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2463
timestamp 1649977179
transform 1 0 227700 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2465
timestamp 1649977179
transform 1 0 227884 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2477
timestamp 1649977179
transform 1 0 228988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2489
timestamp 1649977179
transform 1 0 230092 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2501
timestamp 1649977179
transform 1 0 231196 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2513
timestamp 1649977179
transform 1 0 232300 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2519
timestamp 1649977179
transform 1 0 232852 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2521
timestamp 1649977179
transform 1 0 233036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2533
timestamp 1649977179
transform 1 0 234140 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2545
timestamp 1649977179
transform 1 0 235244 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2557
timestamp 1649977179
transform 1 0 236348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2569
timestamp 1649977179
transform 1 0 237452 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2575
timestamp 1649977179
transform 1 0 238004 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2577
timestamp 1649977179
transform 1 0 238188 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2589
timestamp 1649977179
transform 1 0 239292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2601
timestamp 1649977179
transform 1 0 240396 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2613
timestamp 1649977179
transform 1 0 241500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2625
timestamp 1649977179
transform 1 0 242604 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2631
timestamp 1649977179
transform 1 0 243156 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2633
timestamp 1649977179
transform 1 0 243340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2645
timestamp 1649977179
transform 1 0 244444 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2657
timestamp 1649977179
transform 1 0 245548 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2669
timestamp 1649977179
transform 1 0 246652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2681
timestamp 1649977179
transform 1 0 247756 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2687
timestamp 1649977179
transform 1 0 248308 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2689
timestamp 1649977179
transform 1 0 248492 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2701
timestamp 1649977179
transform 1 0 249596 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2713
timestamp 1649977179
transform 1 0 250700 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2725
timestamp 1649977179
transform 1 0 251804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2737
timestamp 1649977179
transform 1 0 252908 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2743
timestamp 1649977179
transform 1 0 253460 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2745
timestamp 1649977179
transform 1 0 253644 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2757
timestamp 1649977179
transform 1 0 254748 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2769
timestamp 1649977179
transform 1 0 255852 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2781
timestamp 1649977179
transform 1 0 256956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2793
timestamp 1649977179
transform 1 0 258060 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2799
timestamp 1649977179
transform 1 0 258612 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2801
timestamp 1649977179
transform 1 0 258796 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2813
timestamp 1649977179
transform 1 0 259900 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2825
timestamp 1649977179
transform 1 0 261004 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2837
timestamp 1649977179
transform 1 0 262108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2849
timestamp 1649977179
transform 1 0 263212 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2855
timestamp 1649977179
transform 1 0 263764 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2857
timestamp 1649977179
transform 1 0 263948 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2869
timestamp 1649977179
transform 1 0 265052 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2881
timestamp 1649977179
transform 1 0 266156 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2893
timestamp 1649977179
transform 1 0 267260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2905
timestamp 1649977179
transform 1 0 268364 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2911
timestamp 1649977179
transform 1 0 268916 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2913
timestamp 1649977179
transform 1 0 269100 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2925
timestamp 1649977179
transform 1 0 270204 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2937
timestamp 1649977179
transform 1 0 271308 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2949
timestamp 1649977179
transform 1 0 272412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2961
timestamp 1649977179
transform 1 0 273516 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2967
timestamp 1649977179
transform 1 0 274068 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2969
timestamp 1649977179
transform 1 0 274252 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2981
timestamp 1649977179
transform 1 0 275356 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2993
timestamp 1649977179
transform 1 0 276460 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3005
timestamp 1649977179
transform 1 0 277564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3017
timestamp 1649977179
transform 1 0 278668 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3023
timestamp 1649977179
transform 1 0 279220 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3025
timestamp 1649977179
transform 1 0 279404 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3037
timestamp 1649977179
transform 1 0 280508 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3049
timestamp 1649977179
transform 1 0 281612 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3061
timestamp 1649977179
transform 1 0 282716 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3073
timestamp 1649977179
transform 1 0 283820 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3079
timestamp 1649977179
transform 1 0 284372 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3081
timestamp 1649977179
transform 1 0 284556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3093
timestamp 1649977179
transform 1 0 285660 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3105
timestamp 1649977179
transform 1 0 286764 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3117
timestamp 1649977179
transform 1 0 287868 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3129
timestamp 1649977179
transform 1 0 288972 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3135
timestamp 1649977179
transform 1 0 289524 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3137
timestamp 1649977179
transform 1 0 289708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3149
timestamp 1649977179
transform 1 0 290812 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3161
timestamp 1649977179
transform 1 0 291916 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3173
timestamp 1649977179
transform 1 0 293020 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3185
timestamp 1649977179
transform 1 0 294124 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3191
timestamp 1649977179
transform 1 0 294676 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3193
timestamp 1649977179
transform 1 0 294860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3205
timestamp 1649977179
transform 1 0 295964 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3217
timestamp 1649977179
transform 1 0 297068 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3229
timestamp 1649977179
transform 1 0 298172 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3241
timestamp 1649977179
transform 1 0 299276 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3247
timestamp 1649977179
transform 1 0 299828 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3249
timestamp 1649977179
transform 1 0 300012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3261
timestamp 1649977179
transform 1 0 301116 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3273
timestamp 1649977179
transform 1 0 302220 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3285
timestamp 1649977179
transform 1 0 303324 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3297
timestamp 1649977179
transform 1 0 304428 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3303
timestamp 1649977179
transform 1 0 304980 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3305
timestamp 1649977179
transform 1 0 305164 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1649977179
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1649977179
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1649977179
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1649977179
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1649977179
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1649977179
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1649977179
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1649977179
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1649977179
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1649977179
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1649977179
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1649977179
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1649977179
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1649977179
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1649977179
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1649977179
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1649977179
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1649977179
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1649977179
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1649977179
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1649977179
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1649977179
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1649977179
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1649977179
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1649977179
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1649977179
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1649977179
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1649977179
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1649977179
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1649977179
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1649977179
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1649977179
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1649977179
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_557
timestamp 1649977179
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_569
timestamp 1649977179
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1649977179
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1649977179
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1649977179
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_601
timestamp 1649977179
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_613
timestamp 1649977179
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_625
timestamp 1649977179
transform 1 0 58604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_637
timestamp 1649977179
transform 1 0 59708 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 1649977179
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_645
timestamp 1649977179
transform 1 0 60444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_657
timestamp 1649977179
transform 1 0 61548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_669
timestamp 1649977179
transform 1 0 62652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_681
timestamp 1649977179
transform 1 0 63756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_693
timestamp 1649977179
transform 1 0 64860 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_699
timestamp 1649977179
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_701
timestamp 1649977179
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_713
timestamp 1649977179
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_725
timestamp 1649977179
transform 1 0 67804 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_737
timestamp 1649977179
transform 1 0 68908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_749
timestamp 1649977179
transform 1 0 70012 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_755
timestamp 1649977179
transform 1 0 70564 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_757
timestamp 1649977179
transform 1 0 70748 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_769
timestamp 1649977179
transform 1 0 71852 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_781
timestamp 1649977179
transform 1 0 72956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_793
timestamp 1649977179
transform 1 0 74060 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_805
timestamp 1649977179
transform 1 0 75164 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_811
timestamp 1649977179
transform 1 0 75716 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_813
timestamp 1649977179
transform 1 0 75900 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_825
timestamp 1649977179
transform 1 0 77004 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_837
timestamp 1649977179
transform 1 0 78108 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_849
timestamp 1649977179
transform 1 0 79212 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_861
timestamp 1649977179
transform 1 0 80316 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_867
timestamp 1649977179
transform 1 0 80868 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_869
timestamp 1649977179
transform 1 0 81052 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_881
timestamp 1649977179
transform 1 0 82156 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_893
timestamp 1649977179
transform 1 0 83260 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_905
timestamp 1649977179
transform 1 0 84364 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_917
timestamp 1649977179
transform 1 0 85468 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_923
timestamp 1649977179
transform 1 0 86020 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_925
timestamp 1649977179
transform 1 0 86204 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_937
timestamp 1649977179
transform 1 0 87308 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_949
timestamp 1649977179
transform 1 0 88412 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_961
timestamp 1649977179
transform 1 0 89516 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_973
timestamp 1649977179
transform 1 0 90620 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_979
timestamp 1649977179
transform 1 0 91172 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_981
timestamp 1649977179
transform 1 0 91356 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_993
timestamp 1649977179
transform 1 0 92460 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1005
timestamp 1649977179
transform 1 0 93564 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1017
timestamp 1649977179
transform 1 0 94668 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1029
timestamp 1649977179
transform 1 0 95772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1035
timestamp 1649977179
transform 1 0 96324 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1037
timestamp 1649977179
transform 1 0 96508 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1049
timestamp 1649977179
transform 1 0 97612 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1061
timestamp 1649977179
transform 1 0 98716 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1073
timestamp 1649977179
transform 1 0 99820 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1085
timestamp 1649977179
transform 1 0 100924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1091
timestamp 1649977179
transform 1 0 101476 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1093
timestamp 1649977179
transform 1 0 101660 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1105
timestamp 1649977179
transform 1 0 102764 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1117
timestamp 1649977179
transform 1 0 103868 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1129
timestamp 1649977179
transform 1 0 104972 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1141
timestamp 1649977179
transform 1 0 106076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1147
timestamp 1649977179
transform 1 0 106628 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1149
timestamp 1649977179
transform 1 0 106812 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1161
timestamp 1649977179
transform 1 0 107916 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1173
timestamp 1649977179
transform 1 0 109020 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1185
timestamp 1649977179
transform 1 0 110124 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1197
timestamp 1649977179
transform 1 0 111228 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1203
timestamp 1649977179
transform 1 0 111780 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1205
timestamp 1649977179
transform 1 0 111964 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1217
timestamp 1649977179
transform 1 0 113068 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1229
timestamp 1649977179
transform 1 0 114172 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1241
timestamp 1649977179
transform 1 0 115276 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1253
timestamp 1649977179
transform 1 0 116380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1259
timestamp 1649977179
transform 1 0 116932 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1261
timestamp 1649977179
transform 1 0 117116 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1273
timestamp 1649977179
transform 1 0 118220 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1285
timestamp 1649977179
transform 1 0 119324 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1297
timestamp 1649977179
transform 1 0 120428 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1309
timestamp 1649977179
transform 1 0 121532 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1315
timestamp 1649977179
transform 1 0 122084 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1317
timestamp 1649977179
transform 1 0 122268 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1329
timestamp 1649977179
transform 1 0 123372 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1341
timestamp 1649977179
transform 1 0 124476 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1353
timestamp 1649977179
transform 1 0 125580 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1365
timestamp 1649977179
transform 1 0 126684 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1371
timestamp 1649977179
transform 1 0 127236 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1373
timestamp 1649977179
transform 1 0 127420 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1385
timestamp 1649977179
transform 1 0 128524 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1397
timestamp 1649977179
transform 1 0 129628 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1409
timestamp 1649977179
transform 1 0 130732 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1421
timestamp 1649977179
transform 1 0 131836 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1427
timestamp 1649977179
transform 1 0 132388 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1429
timestamp 1649977179
transform 1 0 132572 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1441
timestamp 1649977179
transform 1 0 133676 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1453
timestamp 1649977179
transform 1 0 134780 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1465
timestamp 1649977179
transform 1 0 135884 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1477
timestamp 1649977179
transform 1 0 136988 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1483
timestamp 1649977179
transform 1 0 137540 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1485
timestamp 1649977179
transform 1 0 137724 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1497
timestamp 1649977179
transform 1 0 138828 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1509
timestamp 1649977179
transform 1 0 139932 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1521
timestamp 1649977179
transform 1 0 141036 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1533
timestamp 1649977179
transform 1 0 142140 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1539
timestamp 1649977179
transform 1 0 142692 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1541
timestamp 1649977179
transform 1 0 142876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1553
timestamp 1649977179
transform 1 0 143980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1565
timestamp 1649977179
transform 1 0 145084 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1577
timestamp 1649977179
transform 1 0 146188 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1589
timestamp 1649977179
transform 1 0 147292 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1595
timestamp 1649977179
transform 1 0 147844 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1597
timestamp 1649977179
transform 1 0 148028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1609
timestamp 1649977179
transform 1 0 149132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1621
timestamp 1649977179
transform 1 0 150236 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1633
timestamp 1649977179
transform 1 0 151340 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1645
timestamp 1649977179
transform 1 0 152444 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1651
timestamp 1649977179
transform 1 0 152996 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1653
timestamp 1649977179
transform 1 0 153180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1665
timestamp 1649977179
transform 1 0 154284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1677
timestamp 1649977179
transform 1 0 155388 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1689
timestamp 1649977179
transform 1 0 156492 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1701
timestamp 1649977179
transform 1 0 157596 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1707
timestamp 1649977179
transform 1 0 158148 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1709
timestamp 1649977179
transform 1 0 158332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1721
timestamp 1649977179
transform 1 0 159436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1733
timestamp 1649977179
transform 1 0 160540 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1745
timestamp 1649977179
transform 1 0 161644 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1757
timestamp 1649977179
transform 1 0 162748 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1763
timestamp 1649977179
transform 1 0 163300 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1765
timestamp 1649977179
transform 1 0 163484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1777
timestamp 1649977179
transform 1 0 164588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1789
timestamp 1649977179
transform 1 0 165692 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1801
timestamp 1649977179
transform 1 0 166796 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1813
timestamp 1649977179
transform 1 0 167900 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1819
timestamp 1649977179
transform 1 0 168452 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1821
timestamp 1649977179
transform 1 0 168636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1833
timestamp 1649977179
transform 1 0 169740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1845
timestamp 1649977179
transform 1 0 170844 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1857
timestamp 1649977179
transform 1 0 171948 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1869
timestamp 1649977179
transform 1 0 173052 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1875
timestamp 1649977179
transform 1 0 173604 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1877
timestamp 1649977179
transform 1 0 173788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1889
timestamp 1649977179
transform 1 0 174892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1901
timestamp 1649977179
transform 1 0 175996 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1913
timestamp 1649977179
transform 1 0 177100 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1925
timestamp 1649977179
transform 1 0 178204 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1931
timestamp 1649977179
transform 1 0 178756 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1933
timestamp 1649977179
transform 1 0 178940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1945
timestamp 1649977179
transform 1 0 180044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1957
timestamp 1649977179
transform 1 0 181148 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1969
timestamp 1649977179
transform 1 0 182252 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1981
timestamp 1649977179
transform 1 0 183356 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1987
timestamp 1649977179
transform 1 0 183908 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1989
timestamp 1649977179
transform 1 0 184092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2001
timestamp 1649977179
transform 1 0 185196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2013
timestamp 1649977179
transform 1 0 186300 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2025
timestamp 1649977179
transform 1 0 187404 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2037
timestamp 1649977179
transform 1 0 188508 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2043
timestamp 1649977179
transform 1 0 189060 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2045
timestamp 1649977179
transform 1 0 189244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2057
timestamp 1649977179
transform 1 0 190348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2069
timestamp 1649977179
transform 1 0 191452 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2081
timestamp 1649977179
transform 1 0 192556 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2093
timestamp 1649977179
transform 1 0 193660 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2099
timestamp 1649977179
transform 1 0 194212 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2101
timestamp 1649977179
transform 1 0 194396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2113
timestamp 1649977179
transform 1 0 195500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2125
timestamp 1649977179
transform 1 0 196604 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2137
timestamp 1649977179
transform 1 0 197708 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2149
timestamp 1649977179
transform 1 0 198812 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2155
timestamp 1649977179
transform 1 0 199364 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2157
timestamp 1649977179
transform 1 0 199548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2169
timestamp 1649977179
transform 1 0 200652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2181
timestamp 1649977179
transform 1 0 201756 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2193
timestamp 1649977179
transform 1 0 202860 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2205
timestamp 1649977179
transform 1 0 203964 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2211
timestamp 1649977179
transform 1 0 204516 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2213
timestamp 1649977179
transform 1 0 204700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2225
timestamp 1649977179
transform 1 0 205804 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2237
timestamp 1649977179
transform 1 0 206908 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2249
timestamp 1649977179
transform 1 0 208012 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2261
timestamp 1649977179
transform 1 0 209116 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2267
timestamp 1649977179
transform 1 0 209668 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2269
timestamp 1649977179
transform 1 0 209852 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2281
timestamp 1649977179
transform 1 0 210956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2293
timestamp 1649977179
transform 1 0 212060 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2305
timestamp 1649977179
transform 1 0 213164 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2317
timestamp 1649977179
transform 1 0 214268 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2323
timestamp 1649977179
transform 1 0 214820 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2325
timestamp 1649977179
transform 1 0 215004 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2337
timestamp 1649977179
transform 1 0 216108 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2349
timestamp 1649977179
transform 1 0 217212 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2361
timestamp 1649977179
transform 1 0 218316 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2373
timestamp 1649977179
transform 1 0 219420 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2379
timestamp 1649977179
transform 1 0 219972 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2381
timestamp 1649977179
transform 1 0 220156 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2393
timestamp 1649977179
transform 1 0 221260 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2405
timestamp 1649977179
transform 1 0 222364 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2417
timestamp 1649977179
transform 1 0 223468 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2429
timestamp 1649977179
transform 1 0 224572 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2435
timestamp 1649977179
transform 1 0 225124 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2437
timestamp 1649977179
transform 1 0 225308 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2449
timestamp 1649977179
transform 1 0 226412 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2461
timestamp 1649977179
transform 1 0 227516 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2473
timestamp 1649977179
transform 1 0 228620 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2485
timestamp 1649977179
transform 1 0 229724 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2491
timestamp 1649977179
transform 1 0 230276 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2493
timestamp 1649977179
transform 1 0 230460 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2505
timestamp 1649977179
transform 1 0 231564 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2517
timestamp 1649977179
transform 1 0 232668 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2529
timestamp 1649977179
transform 1 0 233772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2541
timestamp 1649977179
transform 1 0 234876 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2547
timestamp 1649977179
transform 1 0 235428 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2549
timestamp 1649977179
transform 1 0 235612 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2561
timestamp 1649977179
transform 1 0 236716 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2573
timestamp 1649977179
transform 1 0 237820 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2585
timestamp 1649977179
transform 1 0 238924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2597
timestamp 1649977179
transform 1 0 240028 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2603
timestamp 1649977179
transform 1 0 240580 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2605
timestamp 1649977179
transform 1 0 240764 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2617
timestamp 1649977179
transform 1 0 241868 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2629
timestamp 1649977179
transform 1 0 242972 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2641
timestamp 1649977179
transform 1 0 244076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2653
timestamp 1649977179
transform 1 0 245180 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2659
timestamp 1649977179
transform 1 0 245732 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2661
timestamp 1649977179
transform 1 0 245916 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2673
timestamp 1649977179
transform 1 0 247020 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2685
timestamp 1649977179
transform 1 0 248124 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2697
timestamp 1649977179
transform 1 0 249228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2709
timestamp 1649977179
transform 1 0 250332 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2715
timestamp 1649977179
transform 1 0 250884 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2717
timestamp 1649977179
transform 1 0 251068 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2729
timestamp 1649977179
transform 1 0 252172 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2741
timestamp 1649977179
transform 1 0 253276 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2753
timestamp 1649977179
transform 1 0 254380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2765
timestamp 1649977179
transform 1 0 255484 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2771
timestamp 1649977179
transform 1 0 256036 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2773
timestamp 1649977179
transform 1 0 256220 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2785
timestamp 1649977179
transform 1 0 257324 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2797
timestamp 1649977179
transform 1 0 258428 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2809
timestamp 1649977179
transform 1 0 259532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2821
timestamp 1649977179
transform 1 0 260636 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2827
timestamp 1649977179
transform 1 0 261188 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2829
timestamp 1649977179
transform 1 0 261372 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2841
timestamp 1649977179
transform 1 0 262476 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2853
timestamp 1649977179
transform 1 0 263580 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2865
timestamp 1649977179
transform 1 0 264684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2877
timestamp 1649977179
transform 1 0 265788 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2883
timestamp 1649977179
transform 1 0 266340 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2885
timestamp 1649977179
transform 1 0 266524 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2897
timestamp 1649977179
transform 1 0 267628 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2909
timestamp 1649977179
transform 1 0 268732 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2921
timestamp 1649977179
transform 1 0 269836 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2933
timestamp 1649977179
transform 1 0 270940 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2939
timestamp 1649977179
transform 1 0 271492 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2941
timestamp 1649977179
transform 1 0 271676 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2953
timestamp 1649977179
transform 1 0 272780 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2965
timestamp 1649977179
transform 1 0 273884 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2977
timestamp 1649977179
transform 1 0 274988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2989
timestamp 1649977179
transform 1 0 276092 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2995
timestamp 1649977179
transform 1 0 276644 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2997
timestamp 1649977179
transform 1 0 276828 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3009
timestamp 1649977179
transform 1 0 277932 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3021
timestamp 1649977179
transform 1 0 279036 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3033
timestamp 1649977179
transform 1 0 280140 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3045
timestamp 1649977179
transform 1 0 281244 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3051
timestamp 1649977179
transform 1 0 281796 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3053
timestamp 1649977179
transform 1 0 281980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3065
timestamp 1649977179
transform 1 0 283084 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3077
timestamp 1649977179
transform 1 0 284188 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3089
timestamp 1649977179
transform 1 0 285292 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3101
timestamp 1649977179
transform 1 0 286396 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3107
timestamp 1649977179
transform 1 0 286948 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3109
timestamp 1649977179
transform 1 0 287132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3121
timestamp 1649977179
transform 1 0 288236 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3133
timestamp 1649977179
transform 1 0 289340 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3145
timestamp 1649977179
transform 1 0 290444 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3157
timestamp 1649977179
transform 1 0 291548 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3163
timestamp 1649977179
transform 1 0 292100 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3165
timestamp 1649977179
transform 1 0 292284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3177
timestamp 1649977179
transform 1 0 293388 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3189
timestamp 1649977179
transform 1 0 294492 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3201
timestamp 1649977179
transform 1 0 295596 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3213
timestamp 1649977179
transform 1 0 296700 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3219
timestamp 1649977179
transform 1 0 297252 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3221
timestamp 1649977179
transform 1 0 297436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3233
timestamp 1649977179
transform 1 0 298540 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3245
timestamp 1649977179
transform 1 0 299644 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3257
timestamp 1649977179
transform 1 0 300748 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3269
timestamp 1649977179
transform 1 0 301852 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3275
timestamp 1649977179
transform 1 0 302404 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3277
timestamp 1649977179
transform 1 0 302588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3289
timestamp 1649977179
transform 1 0 303692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3301 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 304796 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1649977179
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1649977179
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1649977179
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1649977179
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1649977179
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1649977179
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1649977179
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1649977179
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1649977179
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1649977179
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1649977179
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1649977179
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1649977179
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1649977179
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1649977179
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1649977179
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1649977179
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1649977179
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1649977179
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1649977179
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1649977179
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1649977179
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1649977179
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1649977179
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1649977179
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1649977179
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1649977179
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1649977179
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1649977179
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1649977179
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1649977179
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1649977179
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1649977179
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1649977179
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1649977179
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1649977179
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1649977179
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1649977179
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1649977179
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1649977179
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1649977179
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1649977179
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_617
timestamp 1649977179
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_629
timestamp 1649977179
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_641
timestamp 1649977179
transform 1 0 60076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_653
timestamp 1649977179
transform 1 0 61180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 1649977179
transform 1 0 62284 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 1649977179
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1649977179
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1649977179
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1649977179
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_709
timestamp 1649977179
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 1649977179
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 1649977179
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_729
timestamp 1649977179
transform 1 0 68172 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_741
timestamp 1649977179
transform 1 0 69276 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_753
timestamp 1649977179
transform 1 0 70380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_765
timestamp 1649977179
transform 1 0 71484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_777
timestamp 1649977179
transform 1 0 72588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_783
timestamp 1649977179
transform 1 0 73140 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_785
timestamp 1649977179
transform 1 0 73324 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_797
timestamp 1649977179
transform 1 0 74428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_809
timestamp 1649977179
transform 1 0 75532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_821
timestamp 1649977179
transform 1 0 76636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_833
timestamp 1649977179
transform 1 0 77740 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_839
timestamp 1649977179
transform 1 0 78292 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_841
timestamp 1649977179
transform 1 0 78476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_853
timestamp 1649977179
transform 1 0 79580 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_865
timestamp 1649977179
transform 1 0 80684 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_877
timestamp 1649977179
transform 1 0 81788 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_889
timestamp 1649977179
transform 1 0 82892 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_895
timestamp 1649977179
transform 1 0 83444 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_897
timestamp 1649977179
transform 1 0 83628 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_909
timestamp 1649977179
transform 1 0 84732 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_921
timestamp 1649977179
transform 1 0 85836 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_933
timestamp 1649977179
transform 1 0 86940 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_945
timestamp 1649977179
transform 1 0 88044 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_951
timestamp 1649977179
transform 1 0 88596 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_953
timestamp 1649977179
transform 1 0 88780 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_965
timestamp 1649977179
transform 1 0 89884 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_977
timestamp 1649977179
transform 1 0 90988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_989
timestamp 1649977179
transform 1 0 92092 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1001
timestamp 1649977179
transform 1 0 93196 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1007
timestamp 1649977179
transform 1 0 93748 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1009
timestamp 1649977179
transform 1 0 93932 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1021
timestamp 1649977179
transform 1 0 95036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1033
timestamp 1649977179
transform 1 0 96140 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1045
timestamp 1649977179
transform 1 0 97244 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1057
timestamp 1649977179
transform 1 0 98348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1063
timestamp 1649977179
transform 1 0 98900 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1065
timestamp 1649977179
transform 1 0 99084 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1077
timestamp 1649977179
transform 1 0 100188 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1089
timestamp 1649977179
transform 1 0 101292 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1101
timestamp 1649977179
transform 1 0 102396 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1113
timestamp 1649977179
transform 1 0 103500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1119
timestamp 1649977179
transform 1 0 104052 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1121
timestamp 1649977179
transform 1 0 104236 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1133
timestamp 1649977179
transform 1 0 105340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1145
timestamp 1649977179
transform 1 0 106444 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1157
timestamp 1649977179
transform 1 0 107548 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1169
timestamp 1649977179
transform 1 0 108652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1175
timestamp 1649977179
transform 1 0 109204 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1177
timestamp 1649977179
transform 1 0 109388 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1189
timestamp 1649977179
transform 1 0 110492 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1201
timestamp 1649977179
transform 1 0 111596 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1213
timestamp 1649977179
transform 1 0 112700 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1225
timestamp 1649977179
transform 1 0 113804 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1231
timestamp 1649977179
transform 1 0 114356 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1233
timestamp 1649977179
transform 1 0 114540 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1245
timestamp 1649977179
transform 1 0 115644 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1257
timestamp 1649977179
transform 1 0 116748 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1269
timestamp 1649977179
transform 1 0 117852 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1281
timestamp 1649977179
transform 1 0 118956 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1287
timestamp 1649977179
transform 1 0 119508 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1289
timestamp 1649977179
transform 1 0 119692 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1301
timestamp 1649977179
transform 1 0 120796 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1313
timestamp 1649977179
transform 1 0 121900 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1325
timestamp 1649977179
transform 1 0 123004 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1337
timestamp 1649977179
transform 1 0 124108 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1343
timestamp 1649977179
transform 1 0 124660 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1345
timestamp 1649977179
transform 1 0 124844 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1357
timestamp 1649977179
transform 1 0 125948 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1369
timestamp 1649977179
transform 1 0 127052 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1381
timestamp 1649977179
transform 1 0 128156 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1393
timestamp 1649977179
transform 1 0 129260 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1399
timestamp 1649977179
transform 1 0 129812 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1401
timestamp 1649977179
transform 1 0 129996 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1413
timestamp 1649977179
transform 1 0 131100 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1425
timestamp 1649977179
transform 1 0 132204 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1437
timestamp 1649977179
transform 1 0 133308 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1449
timestamp 1649977179
transform 1 0 134412 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1455
timestamp 1649977179
transform 1 0 134964 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1457
timestamp 1649977179
transform 1 0 135148 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1469
timestamp 1649977179
transform 1 0 136252 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1481
timestamp 1649977179
transform 1 0 137356 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1493
timestamp 1649977179
transform 1 0 138460 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1505
timestamp 1649977179
transform 1 0 139564 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1511
timestamp 1649977179
transform 1 0 140116 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1513
timestamp 1649977179
transform 1 0 140300 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1525
timestamp 1649977179
transform 1 0 141404 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1537
timestamp 1649977179
transform 1 0 142508 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1549
timestamp 1649977179
transform 1 0 143612 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1561
timestamp 1649977179
transform 1 0 144716 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1567
timestamp 1649977179
transform 1 0 145268 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1569
timestamp 1649977179
transform 1 0 145452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1581
timestamp 1649977179
transform 1 0 146556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1593
timestamp 1649977179
transform 1 0 147660 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1605
timestamp 1649977179
transform 1 0 148764 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1617
timestamp 1649977179
transform 1 0 149868 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1623
timestamp 1649977179
transform 1 0 150420 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1625
timestamp 1649977179
transform 1 0 150604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1637
timestamp 1649977179
transform 1 0 151708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1649
timestamp 1649977179
transform 1 0 152812 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1661
timestamp 1649977179
transform 1 0 153916 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1673
timestamp 1649977179
transform 1 0 155020 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1679
timestamp 1649977179
transform 1 0 155572 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1681
timestamp 1649977179
transform 1 0 155756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1693
timestamp 1649977179
transform 1 0 156860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1705
timestamp 1649977179
transform 1 0 157964 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1717
timestamp 1649977179
transform 1 0 159068 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1729
timestamp 1649977179
transform 1 0 160172 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1735
timestamp 1649977179
transform 1 0 160724 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1737
timestamp 1649977179
transform 1 0 160908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1749
timestamp 1649977179
transform 1 0 162012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1761
timestamp 1649977179
transform 1 0 163116 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1773
timestamp 1649977179
transform 1 0 164220 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1785
timestamp 1649977179
transform 1 0 165324 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1791
timestamp 1649977179
transform 1 0 165876 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1793
timestamp 1649977179
transform 1 0 166060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1805
timestamp 1649977179
transform 1 0 167164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1817
timestamp 1649977179
transform 1 0 168268 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1829
timestamp 1649977179
transform 1 0 169372 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1841
timestamp 1649977179
transform 1 0 170476 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1847
timestamp 1649977179
transform 1 0 171028 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1849
timestamp 1649977179
transform 1 0 171212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1861
timestamp 1649977179
transform 1 0 172316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1873
timestamp 1649977179
transform 1 0 173420 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1885
timestamp 1649977179
transform 1 0 174524 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1897
timestamp 1649977179
transform 1 0 175628 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1903
timestamp 1649977179
transform 1 0 176180 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1905
timestamp 1649977179
transform 1 0 176364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1917
timestamp 1649977179
transform 1 0 177468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1929
timestamp 1649977179
transform 1 0 178572 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1941
timestamp 1649977179
transform 1 0 179676 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1953
timestamp 1649977179
transform 1 0 180780 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1959
timestamp 1649977179
transform 1 0 181332 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1961
timestamp 1649977179
transform 1 0 181516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1973
timestamp 1649977179
transform 1 0 182620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1985
timestamp 1649977179
transform 1 0 183724 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1997
timestamp 1649977179
transform 1 0 184828 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2009
timestamp 1649977179
transform 1 0 185932 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2015
timestamp 1649977179
transform 1 0 186484 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2017
timestamp 1649977179
transform 1 0 186668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2029
timestamp 1649977179
transform 1 0 187772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2041
timestamp 1649977179
transform 1 0 188876 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2053
timestamp 1649977179
transform 1 0 189980 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2065
timestamp 1649977179
transform 1 0 191084 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2071
timestamp 1649977179
transform 1 0 191636 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2073
timestamp 1649977179
transform 1 0 191820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2085
timestamp 1649977179
transform 1 0 192924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2097
timestamp 1649977179
transform 1 0 194028 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2109
timestamp 1649977179
transform 1 0 195132 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2121
timestamp 1649977179
transform 1 0 196236 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2127
timestamp 1649977179
transform 1 0 196788 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2129
timestamp 1649977179
transform 1 0 196972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2141
timestamp 1649977179
transform 1 0 198076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2153
timestamp 1649977179
transform 1 0 199180 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2165
timestamp 1649977179
transform 1 0 200284 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2177
timestamp 1649977179
transform 1 0 201388 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2183
timestamp 1649977179
transform 1 0 201940 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2185
timestamp 1649977179
transform 1 0 202124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2197
timestamp 1649977179
transform 1 0 203228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2209
timestamp 1649977179
transform 1 0 204332 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2221
timestamp 1649977179
transform 1 0 205436 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2233
timestamp 1649977179
transform 1 0 206540 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2239
timestamp 1649977179
transform 1 0 207092 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2241
timestamp 1649977179
transform 1 0 207276 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2253
timestamp 1649977179
transform 1 0 208380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2265
timestamp 1649977179
transform 1 0 209484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2277
timestamp 1649977179
transform 1 0 210588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2289
timestamp 1649977179
transform 1 0 211692 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2295
timestamp 1649977179
transform 1 0 212244 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2297
timestamp 1649977179
transform 1 0 212428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2309
timestamp 1649977179
transform 1 0 213532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2321
timestamp 1649977179
transform 1 0 214636 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2333
timestamp 1649977179
transform 1 0 215740 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2345
timestamp 1649977179
transform 1 0 216844 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2351
timestamp 1649977179
transform 1 0 217396 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2353
timestamp 1649977179
transform 1 0 217580 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2365
timestamp 1649977179
transform 1 0 218684 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2377
timestamp 1649977179
transform 1 0 219788 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2389
timestamp 1649977179
transform 1 0 220892 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2401
timestamp 1649977179
transform 1 0 221996 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2407
timestamp 1649977179
transform 1 0 222548 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2409
timestamp 1649977179
transform 1 0 222732 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2421
timestamp 1649977179
transform 1 0 223836 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2433
timestamp 1649977179
transform 1 0 224940 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2445
timestamp 1649977179
transform 1 0 226044 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2457
timestamp 1649977179
transform 1 0 227148 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2463
timestamp 1649977179
transform 1 0 227700 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2465
timestamp 1649977179
transform 1 0 227884 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2477
timestamp 1649977179
transform 1 0 228988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2489
timestamp 1649977179
transform 1 0 230092 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2501
timestamp 1649977179
transform 1 0 231196 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2513
timestamp 1649977179
transform 1 0 232300 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2519
timestamp 1649977179
transform 1 0 232852 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2521
timestamp 1649977179
transform 1 0 233036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2533
timestamp 1649977179
transform 1 0 234140 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2545
timestamp 1649977179
transform 1 0 235244 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2557
timestamp 1649977179
transform 1 0 236348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2569
timestamp 1649977179
transform 1 0 237452 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2575
timestamp 1649977179
transform 1 0 238004 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2577
timestamp 1649977179
transform 1 0 238188 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2589
timestamp 1649977179
transform 1 0 239292 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2601
timestamp 1649977179
transform 1 0 240396 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2613
timestamp 1649977179
transform 1 0 241500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2625
timestamp 1649977179
transform 1 0 242604 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2631
timestamp 1649977179
transform 1 0 243156 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2633
timestamp 1649977179
transform 1 0 243340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2645
timestamp 1649977179
transform 1 0 244444 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2657
timestamp 1649977179
transform 1 0 245548 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2669
timestamp 1649977179
transform 1 0 246652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2681
timestamp 1649977179
transform 1 0 247756 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2687
timestamp 1649977179
transform 1 0 248308 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2689
timestamp 1649977179
transform 1 0 248492 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2701
timestamp 1649977179
transform 1 0 249596 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2713
timestamp 1649977179
transform 1 0 250700 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2725
timestamp 1649977179
transform 1 0 251804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2737
timestamp 1649977179
transform 1 0 252908 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2743
timestamp 1649977179
transform 1 0 253460 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2745
timestamp 1649977179
transform 1 0 253644 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2757
timestamp 1649977179
transform 1 0 254748 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2769
timestamp 1649977179
transform 1 0 255852 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2781
timestamp 1649977179
transform 1 0 256956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2793
timestamp 1649977179
transform 1 0 258060 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2799
timestamp 1649977179
transform 1 0 258612 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2801
timestamp 1649977179
transform 1 0 258796 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2813
timestamp 1649977179
transform 1 0 259900 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2825
timestamp 1649977179
transform 1 0 261004 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2837
timestamp 1649977179
transform 1 0 262108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2849
timestamp 1649977179
transform 1 0 263212 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2855
timestamp 1649977179
transform 1 0 263764 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2857
timestamp 1649977179
transform 1 0 263948 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2869
timestamp 1649977179
transform 1 0 265052 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2881
timestamp 1649977179
transform 1 0 266156 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2893
timestamp 1649977179
transform 1 0 267260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2905
timestamp 1649977179
transform 1 0 268364 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2911
timestamp 1649977179
transform 1 0 268916 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2913
timestamp 1649977179
transform 1 0 269100 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2925
timestamp 1649977179
transform 1 0 270204 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2937
timestamp 1649977179
transform 1 0 271308 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2949
timestamp 1649977179
transform 1 0 272412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2961
timestamp 1649977179
transform 1 0 273516 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2967
timestamp 1649977179
transform 1 0 274068 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2969
timestamp 1649977179
transform 1 0 274252 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2981
timestamp 1649977179
transform 1 0 275356 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2993
timestamp 1649977179
transform 1 0 276460 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3005
timestamp 1649977179
transform 1 0 277564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3017
timestamp 1649977179
transform 1 0 278668 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3023
timestamp 1649977179
transform 1 0 279220 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3025
timestamp 1649977179
transform 1 0 279404 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3037
timestamp 1649977179
transform 1 0 280508 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3049
timestamp 1649977179
transform 1 0 281612 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3061
timestamp 1649977179
transform 1 0 282716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3073
timestamp 1649977179
transform 1 0 283820 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3079
timestamp 1649977179
transform 1 0 284372 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3081
timestamp 1649977179
transform 1 0 284556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3093
timestamp 1649977179
transform 1 0 285660 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3105
timestamp 1649977179
transform 1 0 286764 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3117
timestamp 1649977179
transform 1 0 287868 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3129
timestamp 1649977179
transform 1 0 288972 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3135
timestamp 1649977179
transform 1 0 289524 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3137
timestamp 1649977179
transform 1 0 289708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3149
timestamp 1649977179
transform 1 0 290812 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3161
timestamp 1649977179
transform 1 0 291916 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3173
timestamp 1649977179
transform 1 0 293020 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3185
timestamp 1649977179
transform 1 0 294124 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3191
timestamp 1649977179
transform 1 0 294676 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3193
timestamp 1649977179
transform 1 0 294860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3205
timestamp 1649977179
transform 1 0 295964 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3217
timestamp 1649977179
transform 1 0 297068 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3229
timestamp 1649977179
transform 1 0 298172 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3241
timestamp 1649977179
transform 1 0 299276 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3247
timestamp 1649977179
transform 1 0 299828 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3249
timestamp 1649977179
transform 1 0 300012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3261
timestamp 1649977179
transform 1 0 301116 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3273
timestamp 1649977179
transform 1 0 302220 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3285
timestamp 1649977179
transform 1 0 303324 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3297
timestamp 1649977179
transform 1 0 304428 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3303
timestamp 1649977179
transform 1 0 304980 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3305
timestamp 1649977179
transform 1 0 305164 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1649977179
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1649977179
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1649977179
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1649977179
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1649977179
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1649977179
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1649977179
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1649977179
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1649977179
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1649977179
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1649977179
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1649977179
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1649977179
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1649977179
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1649977179
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1649977179
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1649977179
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1649977179
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1649977179
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1649977179
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1649977179
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1649977179
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1649977179
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1649977179
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1649977179
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1649977179
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1649977179
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1649977179
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1649977179
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1649977179
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1649977179
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1649977179
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1649977179
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1649977179
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1649977179
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1649977179
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1649977179
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1649977179
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_613
timestamp 1649977179
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_625
timestamp 1649977179
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 1649977179
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 1649977179
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_645
timestamp 1649977179
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_657
timestamp 1649977179
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_669
timestamp 1649977179
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_681
timestamp 1649977179
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 1649977179
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 1649977179
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1649977179
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1649977179
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_725
timestamp 1649977179
transform 1 0 67804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_737
timestamp 1649977179
transform 1 0 68908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_749
timestamp 1649977179
transform 1 0 70012 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_755
timestamp 1649977179
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_757
timestamp 1649977179
transform 1 0 70748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_769
timestamp 1649977179
transform 1 0 71852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_781
timestamp 1649977179
transform 1 0 72956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_793
timestamp 1649977179
transform 1 0 74060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_805
timestamp 1649977179
transform 1 0 75164 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_811
timestamp 1649977179
transform 1 0 75716 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_813
timestamp 1649977179
transform 1 0 75900 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_825
timestamp 1649977179
transform 1 0 77004 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_837
timestamp 1649977179
transform 1 0 78108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_849
timestamp 1649977179
transform 1 0 79212 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_861
timestamp 1649977179
transform 1 0 80316 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_867
timestamp 1649977179
transform 1 0 80868 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_869
timestamp 1649977179
transform 1 0 81052 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_881
timestamp 1649977179
transform 1 0 82156 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_893
timestamp 1649977179
transform 1 0 83260 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_905
timestamp 1649977179
transform 1 0 84364 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_917
timestamp 1649977179
transform 1 0 85468 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_923
timestamp 1649977179
transform 1 0 86020 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_925
timestamp 1649977179
transform 1 0 86204 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_937
timestamp 1649977179
transform 1 0 87308 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_949
timestamp 1649977179
transform 1 0 88412 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_961
timestamp 1649977179
transform 1 0 89516 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_973
timestamp 1649977179
transform 1 0 90620 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_979
timestamp 1649977179
transform 1 0 91172 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_981
timestamp 1649977179
transform 1 0 91356 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_993
timestamp 1649977179
transform 1 0 92460 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1005
timestamp 1649977179
transform 1 0 93564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1017
timestamp 1649977179
transform 1 0 94668 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1029
timestamp 1649977179
transform 1 0 95772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1035
timestamp 1649977179
transform 1 0 96324 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1037
timestamp 1649977179
transform 1 0 96508 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1049
timestamp 1649977179
transform 1 0 97612 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1061
timestamp 1649977179
transform 1 0 98716 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1073
timestamp 1649977179
transform 1 0 99820 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1085
timestamp 1649977179
transform 1 0 100924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1091
timestamp 1649977179
transform 1 0 101476 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1093
timestamp 1649977179
transform 1 0 101660 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1105
timestamp 1649977179
transform 1 0 102764 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1117
timestamp 1649977179
transform 1 0 103868 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1129
timestamp 1649977179
transform 1 0 104972 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1141
timestamp 1649977179
transform 1 0 106076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1147
timestamp 1649977179
transform 1 0 106628 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1149
timestamp 1649977179
transform 1 0 106812 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1161
timestamp 1649977179
transform 1 0 107916 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1173
timestamp 1649977179
transform 1 0 109020 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1185
timestamp 1649977179
transform 1 0 110124 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1197
timestamp 1649977179
transform 1 0 111228 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1203
timestamp 1649977179
transform 1 0 111780 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1205
timestamp 1649977179
transform 1 0 111964 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1217
timestamp 1649977179
transform 1 0 113068 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1229
timestamp 1649977179
transform 1 0 114172 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1241
timestamp 1649977179
transform 1 0 115276 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1253
timestamp 1649977179
transform 1 0 116380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1259
timestamp 1649977179
transform 1 0 116932 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1261
timestamp 1649977179
transform 1 0 117116 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1273
timestamp 1649977179
transform 1 0 118220 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1285
timestamp 1649977179
transform 1 0 119324 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1297
timestamp 1649977179
transform 1 0 120428 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1309
timestamp 1649977179
transform 1 0 121532 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1315
timestamp 1649977179
transform 1 0 122084 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1317
timestamp 1649977179
transform 1 0 122268 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1329
timestamp 1649977179
transform 1 0 123372 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1341
timestamp 1649977179
transform 1 0 124476 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1353
timestamp 1649977179
transform 1 0 125580 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1365
timestamp 1649977179
transform 1 0 126684 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1371
timestamp 1649977179
transform 1 0 127236 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1373
timestamp 1649977179
transform 1 0 127420 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1385
timestamp 1649977179
transform 1 0 128524 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1397
timestamp 1649977179
transform 1 0 129628 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1409
timestamp 1649977179
transform 1 0 130732 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1421
timestamp 1649977179
transform 1 0 131836 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1427
timestamp 1649977179
transform 1 0 132388 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1429
timestamp 1649977179
transform 1 0 132572 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1441
timestamp 1649977179
transform 1 0 133676 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1453
timestamp 1649977179
transform 1 0 134780 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1465
timestamp 1649977179
transform 1 0 135884 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1477
timestamp 1649977179
transform 1 0 136988 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1483
timestamp 1649977179
transform 1 0 137540 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1485
timestamp 1649977179
transform 1 0 137724 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1497
timestamp 1649977179
transform 1 0 138828 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1509
timestamp 1649977179
transform 1 0 139932 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1521
timestamp 1649977179
transform 1 0 141036 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1533
timestamp 1649977179
transform 1 0 142140 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1539
timestamp 1649977179
transform 1 0 142692 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1541
timestamp 1649977179
transform 1 0 142876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1553
timestamp 1649977179
transform 1 0 143980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1565
timestamp 1649977179
transform 1 0 145084 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1577
timestamp 1649977179
transform 1 0 146188 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1589
timestamp 1649977179
transform 1 0 147292 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1595
timestamp 1649977179
transform 1 0 147844 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1597
timestamp 1649977179
transform 1 0 148028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1609
timestamp 1649977179
transform 1 0 149132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1621
timestamp 1649977179
transform 1 0 150236 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1633
timestamp 1649977179
transform 1 0 151340 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1645
timestamp 1649977179
transform 1 0 152444 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1651
timestamp 1649977179
transform 1 0 152996 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1653
timestamp 1649977179
transform 1 0 153180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1665
timestamp 1649977179
transform 1 0 154284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1677
timestamp 1649977179
transform 1 0 155388 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1689
timestamp 1649977179
transform 1 0 156492 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1701
timestamp 1649977179
transform 1 0 157596 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1707
timestamp 1649977179
transform 1 0 158148 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1709
timestamp 1649977179
transform 1 0 158332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1721
timestamp 1649977179
transform 1 0 159436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1733
timestamp 1649977179
transform 1 0 160540 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1745
timestamp 1649977179
transform 1 0 161644 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1757
timestamp 1649977179
transform 1 0 162748 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1763
timestamp 1649977179
transform 1 0 163300 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1765
timestamp 1649977179
transform 1 0 163484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1777
timestamp 1649977179
transform 1 0 164588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1789
timestamp 1649977179
transform 1 0 165692 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1801
timestamp 1649977179
transform 1 0 166796 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1813
timestamp 1649977179
transform 1 0 167900 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1819
timestamp 1649977179
transform 1 0 168452 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1821
timestamp 1649977179
transform 1 0 168636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1833
timestamp 1649977179
transform 1 0 169740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1845
timestamp 1649977179
transform 1 0 170844 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1857
timestamp 1649977179
transform 1 0 171948 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1869
timestamp 1649977179
transform 1 0 173052 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1875
timestamp 1649977179
transform 1 0 173604 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1877
timestamp 1649977179
transform 1 0 173788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1889
timestamp 1649977179
transform 1 0 174892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1901
timestamp 1649977179
transform 1 0 175996 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1913
timestamp 1649977179
transform 1 0 177100 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1925
timestamp 1649977179
transform 1 0 178204 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1931
timestamp 1649977179
transform 1 0 178756 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1933
timestamp 1649977179
transform 1 0 178940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1945
timestamp 1649977179
transform 1 0 180044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1957
timestamp 1649977179
transform 1 0 181148 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1969
timestamp 1649977179
transform 1 0 182252 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1981
timestamp 1649977179
transform 1 0 183356 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1987
timestamp 1649977179
transform 1 0 183908 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1989
timestamp 1649977179
transform 1 0 184092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2001
timestamp 1649977179
transform 1 0 185196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2013
timestamp 1649977179
transform 1 0 186300 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2025
timestamp 1649977179
transform 1 0 187404 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2037
timestamp 1649977179
transform 1 0 188508 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2043
timestamp 1649977179
transform 1 0 189060 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2045
timestamp 1649977179
transform 1 0 189244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2057
timestamp 1649977179
transform 1 0 190348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2069
timestamp 1649977179
transform 1 0 191452 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2081
timestamp 1649977179
transform 1 0 192556 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2093
timestamp 1649977179
transform 1 0 193660 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2099
timestamp 1649977179
transform 1 0 194212 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2101
timestamp 1649977179
transform 1 0 194396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2113
timestamp 1649977179
transform 1 0 195500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2125
timestamp 1649977179
transform 1 0 196604 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2137
timestamp 1649977179
transform 1 0 197708 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2149
timestamp 1649977179
transform 1 0 198812 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2155
timestamp 1649977179
transform 1 0 199364 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2157
timestamp 1649977179
transform 1 0 199548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2169
timestamp 1649977179
transform 1 0 200652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2181
timestamp 1649977179
transform 1 0 201756 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2193
timestamp 1649977179
transform 1 0 202860 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2205
timestamp 1649977179
transform 1 0 203964 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2211
timestamp 1649977179
transform 1 0 204516 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2213
timestamp 1649977179
transform 1 0 204700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2225
timestamp 1649977179
transform 1 0 205804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2237
timestamp 1649977179
transform 1 0 206908 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2249
timestamp 1649977179
transform 1 0 208012 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2261
timestamp 1649977179
transform 1 0 209116 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2267
timestamp 1649977179
transform 1 0 209668 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2269
timestamp 1649977179
transform 1 0 209852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2281
timestamp 1649977179
transform 1 0 210956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2293
timestamp 1649977179
transform 1 0 212060 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2305
timestamp 1649977179
transform 1 0 213164 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2317
timestamp 1649977179
transform 1 0 214268 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2323
timestamp 1649977179
transform 1 0 214820 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2325
timestamp 1649977179
transform 1 0 215004 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2337
timestamp 1649977179
transform 1 0 216108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2349
timestamp 1649977179
transform 1 0 217212 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2361
timestamp 1649977179
transform 1 0 218316 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2373
timestamp 1649977179
transform 1 0 219420 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2379
timestamp 1649977179
transform 1 0 219972 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2381
timestamp 1649977179
transform 1 0 220156 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2393
timestamp 1649977179
transform 1 0 221260 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2405
timestamp 1649977179
transform 1 0 222364 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2417
timestamp 1649977179
transform 1 0 223468 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2429
timestamp 1649977179
transform 1 0 224572 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2435
timestamp 1649977179
transform 1 0 225124 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2437
timestamp 1649977179
transform 1 0 225308 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2449
timestamp 1649977179
transform 1 0 226412 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2461
timestamp 1649977179
transform 1 0 227516 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2473
timestamp 1649977179
transform 1 0 228620 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2485
timestamp 1649977179
transform 1 0 229724 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2491
timestamp 1649977179
transform 1 0 230276 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2493
timestamp 1649977179
transform 1 0 230460 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2505
timestamp 1649977179
transform 1 0 231564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2517
timestamp 1649977179
transform 1 0 232668 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2529
timestamp 1649977179
transform 1 0 233772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2541
timestamp 1649977179
transform 1 0 234876 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2547
timestamp 1649977179
transform 1 0 235428 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2549
timestamp 1649977179
transform 1 0 235612 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2561
timestamp 1649977179
transform 1 0 236716 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2573
timestamp 1649977179
transform 1 0 237820 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2585
timestamp 1649977179
transform 1 0 238924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2597
timestamp 1649977179
transform 1 0 240028 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2603
timestamp 1649977179
transform 1 0 240580 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2605
timestamp 1649977179
transform 1 0 240764 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2617
timestamp 1649977179
transform 1 0 241868 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2629
timestamp 1649977179
transform 1 0 242972 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2641
timestamp 1649977179
transform 1 0 244076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2653
timestamp 1649977179
transform 1 0 245180 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2659
timestamp 1649977179
transform 1 0 245732 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2661
timestamp 1649977179
transform 1 0 245916 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2673
timestamp 1649977179
transform 1 0 247020 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2685
timestamp 1649977179
transform 1 0 248124 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2697
timestamp 1649977179
transform 1 0 249228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2709
timestamp 1649977179
transform 1 0 250332 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2715
timestamp 1649977179
transform 1 0 250884 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2717
timestamp 1649977179
transform 1 0 251068 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2729
timestamp 1649977179
transform 1 0 252172 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2741
timestamp 1649977179
transform 1 0 253276 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2753
timestamp 1649977179
transform 1 0 254380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2765
timestamp 1649977179
transform 1 0 255484 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2771
timestamp 1649977179
transform 1 0 256036 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2773
timestamp 1649977179
transform 1 0 256220 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2785
timestamp 1649977179
transform 1 0 257324 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2797
timestamp 1649977179
transform 1 0 258428 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2809
timestamp 1649977179
transform 1 0 259532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2821
timestamp 1649977179
transform 1 0 260636 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2827
timestamp 1649977179
transform 1 0 261188 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2829
timestamp 1649977179
transform 1 0 261372 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2841
timestamp 1649977179
transform 1 0 262476 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2853
timestamp 1649977179
transform 1 0 263580 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2865
timestamp 1649977179
transform 1 0 264684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2877
timestamp 1649977179
transform 1 0 265788 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2883
timestamp 1649977179
transform 1 0 266340 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2885
timestamp 1649977179
transform 1 0 266524 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2897
timestamp 1649977179
transform 1 0 267628 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2909
timestamp 1649977179
transform 1 0 268732 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2921
timestamp 1649977179
transform 1 0 269836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2933
timestamp 1649977179
transform 1 0 270940 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2939
timestamp 1649977179
transform 1 0 271492 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2941
timestamp 1649977179
transform 1 0 271676 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2953
timestamp 1649977179
transform 1 0 272780 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2965
timestamp 1649977179
transform 1 0 273884 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2977
timestamp 1649977179
transform 1 0 274988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2989
timestamp 1649977179
transform 1 0 276092 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2995
timestamp 1649977179
transform 1 0 276644 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2997
timestamp 1649977179
transform 1 0 276828 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3009
timestamp 1649977179
transform 1 0 277932 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3021
timestamp 1649977179
transform 1 0 279036 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3033
timestamp 1649977179
transform 1 0 280140 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3045
timestamp 1649977179
transform 1 0 281244 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3051
timestamp 1649977179
transform 1 0 281796 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3053
timestamp 1649977179
transform 1 0 281980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3065
timestamp 1649977179
transform 1 0 283084 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3077
timestamp 1649977179
transform 1 0 284188 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3089
timestamp 1649977179
transform 1 0 285292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3101
timestamp 1649977179
transform 1 0 286396 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3107
timestamp 1649977179
transform 1 0 286948 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3109
timestamp 1649977179
transform 1 0 287132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3121
timestamp 1649977179
transform 1 0 288236 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3133
timestamp 1649977179
transform 1 0 289340 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3145
timestamp 1649977179
transform 1 0 290444 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3157
timestamp 1649977179
transform 1 0 291548 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3163
timestamp 1649977179
transform 1 0 292100 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3165
timestamp 1649977179
transform 1 0 292284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3177
timestamp 1649977179
transform 1 0 293388 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3189
timestamp 1649977179
transform 1 0 294492 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3201
timestamp 1649977179
transform 1 0 295596 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3213
timestamp 1649977179
transform 1 0 296700 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3219
timestamp 1649977179
transform 1 0 297252 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3221
timestamp 1649977179
transform 1 0 297436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3233
timestamp 1649977179
transform 1 0 298540 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3245
timestamp 1649977179
transform 1 0 299644 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3257
timestamp 1649977179
transform 1 0 300748 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3269
timestamp 1649977179
transform 1 0 301852 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3275
timestamp 1649977179
transform 1 0 302404 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3277
timestamp 1649977179
transform 1 0 302588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3289
timestamp 1649977179
transform 1 0 303692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3301
timestamp 1649977179
transform 1 0 304796 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1649977179
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1649977179
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1649977179
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1649977179
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1649977179
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1649977179
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1649977179
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1649977179
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1649977179
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1649977179
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1649977179
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1649977179
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1649977179
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1649977179
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1649977179
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1649977179
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1649977179
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1649977179
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1649977179
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1649977179
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1649977179
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1649977179
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1649977179
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1649977179
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1649977179
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1649977179
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1649977179
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1649977179
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1649977179
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1649977179
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1649977179
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1649977179
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1649977179
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1649977179
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1649977179
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1649977179
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1649977179
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1649977179
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1649977179
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1649977179
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1649977179
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1649977179
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_617
timestamp 1649977179
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_629
timestamp 1649977179
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_641
timestamp 1649977179
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_653
timestamp 1649977179
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 1649977179
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 1649977179
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_673
timestamp 1649977179
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_685
timestamp 1649977179
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_697
timestamp 1649977179
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_709
timestamp 1649977179
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 1649977179
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 1649977179
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_729
timestamp 1649977179
transform 1 0 68172 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_741
timestamp 1649977179
transform 1 0 69276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_753
timestamp 1649977179
transform 1 0 70380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_765
timestamp 1649977179
transform 1 0 71484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_777
timestamp 1649977179
transform 1 0 72588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_783
timestamp 1649977179
transform 1 0 73140 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_785
timestamp 1649977179
transform 1 0 73324 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_797
timestamp 1649977179
transform 1 0 74428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_809
timestamp 1649977179
transform 1 0 75532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_821
timestamp 1649977179
transform 1 0 76636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_833
timestamp 1649977179
transform 1 0 77740 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_839
timestamp 1649977179
transform 1 0 78292 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_841
timestamp 1649977179
transform 1 0 78476 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_853
timestamp 1649977179
transform 1 0 79580 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_865
timestamp 1649977179
transform 1 0 80684 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_877
timestamp 1649977179
transform 1 0 81788 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_889
timestamp 1649977179
transform 1 0 82892 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_895
timestamp 1649977179
transform 1 0 83444 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_897
timestamp 1649977179
transform 1 0 83628 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_909
timestamp 1649977179
transform 1 0 84732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_921
timestamp 1649977179
transform 1 0 85836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_933
timestamp 1649977179
transform 1 0 86940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_945
timestamp 1649977179
transform 1 0 88044 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_951
timestamp 1649977179
transform 1 0 88596 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_953
timestamp 1649977179
transform 1 0 88780 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_965
timestamp 1649977179
transform 1 0 89884 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_977
timestamp 1649977179
transform 1 0 90988 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_989
timestamp 1649977179
transform 1 0 92092 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1001
timestamp 1649977179
transform 1 0 93196 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1007
timestamp 1649977179
transform 1 0 93748 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1009
timestamp 1649977179
transform 1 0 93932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1021
timestamp 1649977179
transform 1 0 95036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1033
timestamp 1649977179
transform 1 0 96140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1045
timestamp 1649977179
transform 1 0 97244 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1057
timestamp 1649977179
transform 1 0 98348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1063
timestamp 1649977179
transform 1 0 98900 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1065
timestamp 1649977179
transform 1 0 99084 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1077
timestamp 1649977179
transform 1 0 100188 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1089
timestamp 1649977179
transform 1 0 101292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1101
timestamp 1649977179
transform 1 0 102396 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1113
timestamp 1649977179
transform 1 0 103500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1119
timestamp 1649977179
transform 1 0 104052 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1121
timestamp 1649977179
transform 1 0 104236 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1133
timestamp 1649977179
transform 1 0 105340 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1145
timestamp 1649977179
transform 1 0 106444 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1157
timestamp 1649977179
transform 1 0 107548 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1169
timestamp 1649977179
transform 1 0 108652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1175
timestamp 1649977179
transform 1 0 109204 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1177
timestamp 1649977179
transform 1 0 109388 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1189
timestamp 1649977179
transform 1 0 110492 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1201
timestamp 1649977179
transform 1 0 111596 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1213
timestamp 1649977179
transform 1 0 112700 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1225
timestamp 1649977179
transform 1 0 113804 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1231
timestamp 1649977179
transform 1 0 114356 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1233
timestamp 1649977179
transform 1 0 114540 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1245
timestamp 1649977179
transform 1 0 115644 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1257
timestamp 1649977179
transform 1 0 116748 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1269
timestamp 1649977179
transform 1 0 117852 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1281
timestamp 1649977179
transform 1 0 118956 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1287
timestamp 1649977179
transform 1 0 119508 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1289
timestamp 1649977179
transform 1 0 119692 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1301
timestamp 1649977179
transform 1 0 120796 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1313
timestamp 1649977179
transform 1 0 121900 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1325
timestamp 1649977179
transform 1 0 123004 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1337
timestamp 1649977179
transform 1 0 124108 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1343
timestamp 1649977179
transform 1 0 124660 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1345
timestamp 1649977179
transform 1 0 124844 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1357
timestamp 1649977179
transform 1 0 125948 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1369
timestamp 1649977179
transform 1 0 127052 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1381
timestamp 1649977179
transform 1 0 128156 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1393
timestamp 1649977179
transform 1 0 129260 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1399
timestamp 1649977179
transform 1 0 129812 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1401
timestamp 1649977179
transform 1 0 129996 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1413
timestamp 1649977179
transform 1 0 131100 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1425
timestamp 1649977179
transform 1 0 132204 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1437
timestamp 1649977179
transform 1 0 133308 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1449
timestamp 1649977179
transform 1 0 134412 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1455
timestamp 1649977179
transform 1 0 134964 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1457
timestamp 1649977179
transform 1 0 135148 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1469
timestamp 1649977179
transform 1 0 136252 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1481
timestamp 1649977179
transform 1 0 137356 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1493
timestamp 1649977179
transform 1 0 138460 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1505
timestamp 1649977179
transform 1 0 139564 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1511
timestamp 1649977179
transform 1 0 140116 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1513
timestamp 1649977179
transform 1 0 140300 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1525
timestamp 1649977179
transform 1 0 141404 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1537
timestamp 1649977179
transform 1 0 142508 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1549
timestamp 1649977179
transform 1 0 143612 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1561
timestamp 1649977179
transform 1 0 144716 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1567
timestamp 1649977179
transform 1 0 145268 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1569
timestamp 1649977179
transform 1 0 145452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1581
timestamp 1649977179
transform 1 0 146556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1593
timestamp 1649977179
transform 1 0 147660 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1605
timestamp 1649977179
transform 1 0 148764 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1617
timestamp 1649977179
transform 1 0 149868 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1623
timestamp 1649977179
transform 1 0 150420 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1625
timestamp 1649977179
transform 1 0 150604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1637
timestamp 1649977179
transform 1 0 151708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1649
timestamp 1649977179
transform 1 0 152812 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1661
timestamp 1649977179
transform 1 0 153916 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1673
timestamp 1649977179
transform 1 0 155020 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1679
timestamp 1649977179
transform 1 0 155572 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1681
timestamp 1649977179
transform 1 0 155756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1693
timestamp 1649977179
transform 1 0 156860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1705
timestamp 1649977179
transform 1 0 157964 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1717
timestamp 1649977179
transform 1 0 159068 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1729
timestamp 1649977179
transform 1 0 160172 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1735
timestamp 1649977179
transform 1 0 160724 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1737
timestamp 1649977179
transform 1 0 160908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1749
timestamp 1649977179
transform 1 0 162012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1761
timestamp 1649977179
transform 1 0 163116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1773
timestamp 1649977179
transform 1 0 164220 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1785
timestamp 1649977179
transform 1 0 165324 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1791
timestamp 1649977179
transform 1 0 165876 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1793
timestamp 1649977179
transform 1 0 166060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1805
timestamp 1649977179
transform 1 0 167164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1817
timestamp 1649977179
transform 1 0 168268 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1829
timestamp 1649977179
transform 1 0 169372 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1841
timestamp 1649977179
transform 1 0 170476 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1847
timestamp 1649977179
transform 1 0 171028 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1849
timestamp 1649977179
transform 1 0 171212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1861
timestamp 1649977179
transform 1 0 172316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1873
timestamp 1649977179
transform 1 0 173420 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1885
timestamp 1649977179
transform 1 0 174524 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1897
timestamp 1649977179
transform 1 0 175628 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1903
timestamp 1649977179
transform 1 0 176180 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1905
timestamp 1649977179
transform 1 0 176364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1917
timestamp 1649977179
transform 1 0 177468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1929
timestamp 1649977179
transform 1 0 178572 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1941
timestamp 1649977179
transform 1 0 179676 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1953
timestamp 1649977179
transform 1 0 180780 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1959
timestamp 1649977179
transform 1 0 181332 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1961
timestamp 1649977179
transform 1 0 181516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1973
timestamp 1649977179
transform 1 0 182620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1985
timestamp 1649977179
transform 1 0 183724 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1997
timestamp 1649977179
transform 1 0 184828 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2009
timestamp 1649977179
transform 1 0 185932 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2015
timestamp 1649977179
transform 1 0 186484 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2017
timestamp 1649977179
transform 1 0 186668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2029
timestamp 1649977179
transform 1 0 187772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2041
timestamp 1649977179
transform 1 0 188876 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2053
timestamp 1649977179
transform 1 0 189980 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2065
timestamp 1649977179
transform 1 0 191084 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2071
timestamp 1649977179
transform 1 0 191636 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2073
timestamp 1649977179
transform 1 0 191820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2085
timestamp 1649977179
transform 1 0 192924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2097
timestamp 1649977179
transform 1 0 194028 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2109
timestamp 1649977179
transform 1 0 195132 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2121
timestamp 1649977179
transform 1 0 196236 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2127
timestamp 1649977179
transform 1 0 196788 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2129
timestamp 1649977179
transform 1 0 196972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2141
timestamp 1649977179
transform 1 0 198076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2153
timestamp 1649977179
transform 1 0 199180 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2165
timestamp 1649977179
transform 1 0 200284 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2177
timestamp 1649977179
transform 1 0 201388 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2183
timestamp 1649977179
transform 1 0 201940 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2185
timestamp 1649977179
transform 1 0 202124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2197
timestamp 1649977179
transform 1 0 203228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2209
timestamp 1649977179
transform 1 0 204332 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2221
timestamp 1649977179
transform 1 0 205436 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2233
timestamp 1649977179
transform 1 0 206540 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2239
timestamp 1649977179
transform 1 0 207092 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2241
timestamp 1649977179
transform 1 0 207276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2253
timestamp 1649977179
transform 1 0 208380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2265
timestamp 1649977179
transform 1 0 209484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2277
timestamp 1649977179
transform 1 0 210588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2289
timestamp 1649977179
transform 1 0 211692 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2295
timestamp 1649977179
transform 1 0 212244 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2297
timestamp 1649977179
transform 1 0 212428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2309
timestamp 1649977179
transform 1 0 213532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2321
timestamp 1649977179
transform 1 0 214636 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2333
timestamp 1649977179
transform 1 0 215740 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2345
timestamp 1649977179
transform 1 0 216844 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2351
timestamp 1649977179
transform 1 0 217396 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2353
timestamp 1649977179
transform 1 0 217580 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2365
timestamp 1649977179
transform 1 0 218684 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2377
timestamp 1649977179
transform 1 0 219788 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2389
timestamp 1649977179
transform 1 0 220892 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2401
timestamp 1649977179
transform 1 0 221996 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2407
timestamp 1649977179
transform 1 0 222548 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2409
timestamp 1649977179
transform 1 0 222732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2421
timestamp 1649977179
transform 1 0 223836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2433
timestamp 1649977179
transform 1 0 224940 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2445
timestamp 1649977179
transform 1 0 226044 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2457
timestamp 1649977179
transform 1 0 227148 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2463
timestamp 1649977179
transform 1 0 227700 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2465
timestamp 1649977179
transform 1 0 227884 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2477
timestamp 1649977179
transform 1 0 228988 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2489
timestamp 1649977179
transform 1 0 230092 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2501
timestamp 1649977179
transform 1 0 231196 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2513
timestamp 1649977179
transform 1 0 232300 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2519
timestamp 1649977179
transform 1 0 232852 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2521
timestamp 1649977179
transform 1 0 233036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2533
timestamp 1649977179
transform 1 0 234140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2545
timestamp 1649977179
transform 1 0 235244 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2557
timestamp 1649977179
transform 1 0 236348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2569
timestamp 1649977179
transform 1 0 237452 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2575
timestamp 1649977179
transform 1 0 238004 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2577
timestamp 1649977179
transform 1 0 238188 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2589
timestamp 1649977179
transform 1 0 239292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2601
timestamp 1649977179
transform 1 0 240396 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2613
timestamp 1649977179
transform 1 0 241500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2625
timestamp 1649977179
transform 1 0 242604 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2631
timestamp 1649977179
transform 1 0 243156 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2633
timestamp 1649977179
transform 1 0 243340 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2645
timestamp 1649977179
transform 1 0 244444 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2657
timestamp 1649977179
transform 1 0 245548 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2669
timestamp 1649977179
transform 1 0 246652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2681
timestamp 1649977179
transform 1 0 247756 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2687
timestamp 1649977179
transform 1 0 248308 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2689
timestamp 1649977179
transform 1 0 248492 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2701
timestamp 1649977179
transform 1 0 249596 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2713
timestamp 1649977179
transform 1 0 250700 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2725
timestamp 1649977179
transform 1 0 251804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2737
timestamp 1649977179
transform 1 0 252908 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2743
timestamp 1649977179
transform 1 0 253460 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2745
timestamp 1649977179
transform 1 0 253644 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2757
timestamp 1649977179
transform 1 0 254748 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2769
timestamp 1649977179
transform 1 0 255852 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2781
timestamp 1649977179
transform 1 0 256956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2793
timestamp 1649977179
transform 1 0 258060 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2799
timestamp 1649977179
transform 1 0 258612 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2801
timestamp 1649977179
transform 1 0 258796 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2813
timestamp 1649977179
transform 1 0 259900 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2825
timestamp 1649977179
transform 1 0 261004 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2837
timestamp 1649977179
transform 1 0 262108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2849
timestamp 1649977179
transform 1 0 263212 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2855
timestamp 1649977179
transform 1 0 263764 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2857
timestamp 1649977179
transform 1 0 263948 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2869
timestamp 1649977179
transform 1 0 265052 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2881
timestamp 1649977179
transform 1 0 266156 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2893
timestamp 1649977179
transform 1 0 267260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2905
timestamp 1649977179
transform 1 0 268364 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2911
timestamp 1649977179
transform 1 0 268916 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2913
timestamp 1649977179
transform 1 0 269100 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2925
timestamp 1649977179
transform 1 0 270204 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2937
timestamp 1649977179
transform 1 0 271308 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2949
timestamp 1649977179
transform 1 0 272412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2961
timestamp 1649977179
transform 1 0 273516 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2967
timestamp 1649977179
transform 1 0 274068 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2969
timestamp 1649977179
transform 1 0 274252 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2981
timestamp 1649977179
transform 1 0 275356 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2993
timestamp 1649977179
transform 1 0 276460 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3005
timestamp 1649977179
transform 1 0 277564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3017
timestamp 1649977179
transform 1 0 278668 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3023
timestamp 1649977179
transform 1 0 279220 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3025
timestamp 1649977179
transform 1 0 279404 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3037
timestamp 1649977179
transform 1 0 280508 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3049
timestamp 1649977179
transform 1 0 281612 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3061
timestamp 1649977179
transform 1 0 282716 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3073
timestamp 1649977179
transform 1 0 283820 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3079
timestamp 1649977179
transform 1 0 284372 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3081
timestamp 1649977179
transform 1 0 284556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3093
timestamp 1649977179
transform 1 0 285660 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3105
timestamp 1649977179
transform 1 0 286764 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3117
timestamp 1649977179
transform 1 0 287868 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3129
timestamp 1649977179
transform 1 0 288972 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3135
timestamp 1649977179
transform 1 0 289524 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3137
timestamp 1649977179
transform 1 0 289708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3149
timestamp 1649977179
transform 1 0 290812 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3161
timestamp 1649977179
transform 1 0 291916 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3173
timestamp 1649977179
transform 1 0 293020 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3185
timestamp 1649977179
transform 1 0 294124 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3191
timestamp 1649977179
transform 1 0 294676 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3193
timestamp 1649977179
transform 1 0 294860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3205
timestamp 1649977179
transform 1 0 295964 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3217
timestamp 1649977179
transform 1 0 297068 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3229
timestamp 1649977179
transform 1 0 298172 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3241
timestamp 1649977179
transform 1 0 299276 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3247
timestamp 1649977179
transform 1 0 299828 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3249
timestamp 1649977179
transform 1 0 300012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3261
timestamp 1649977179
transform 1 0 301116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3273
timestamp 1649977179
transform 1 0 302220 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3285
timestamp 1649977179
transform 1 0 303324 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3297
timestamp 1649977179
transform 1 0 304428 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3303
timestamp 1649977179
transform 1 0 304980 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3305
timestamp 1649977179
transform 1 0 305164 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1649977179
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1649977179
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1649977179
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1649977179
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1649977179
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1649977179
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1649977179
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1649977179
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1649977179
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1649977179
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1649977179
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1649977179
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1649977179
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1649977179
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1649977179
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1649977179
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1649977179
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1649977179
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1649977179
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1649977179
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1649977179
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1649977179
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1649977179
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1649977179
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1649977179
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1649977179
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1649977179
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1649977179
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1649977179
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1649977179
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1649977179
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1649977179
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1649977179
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1649977179
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1649977179
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1649977179
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1649977179
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1649977179
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1649977179
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1649977179
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1649977179
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_625
timestamp 1649977179
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1649977179
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1649977179
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1649977179
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1649977179
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_669
timestamp 1649977179
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_681
timestamp 1649977179
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1649977179
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1649977179
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_701
timestamp 1649977179
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_713
timestamp 1649977179
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_725
timestamp 1649977179
transform 1 0 67804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_737
timestamp 1649977179
transform 1 0 68908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_749
timestamp 1649977179
transform 1 0 70012 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_755
timestamp 1649977179
transform 1 0 70564 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_757
timestamp 1649977179
transform 1 0 70748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_769
timestamp 1649977179
transform 1 0 71852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_781
timestamp 1649977179
transform 1 0 72956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_793
timestamp 1649977179
transform 1 0 74060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_805
timestamp 1649977179
transform 1 0 75164 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_811
timestamp 1649977179
transform 1 0 75716 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_813
timestamp 1649977179
transform 1 0 75900 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_825
timestamp 1649977179
transform 1 0 77004 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_837
timestamp 1649977179
transform 1 0 78108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_849
timestamp 1649977179
transform 1 0 79212 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_861
timestamp 1649977179
transform 1 0 80316 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_867
timestamp 1649977179
transform 1 0 80868 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_869
timestamp 1649977179
transform 1 0 81052 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_881
timestamp 1649977179
transform 1 0 82156 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_893
timestamp 1649977179
transform 1 0 83260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_905
timestamp 1649977179
transform 1 0 84364 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_917
timestamp 1649977179
transform 1 0 85468 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_923
timestamp 1649977179
transform 1 0 86020 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_925
timestamp 1649977179
transform 1 0 86204 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_937
timestamp 1649977179
transform 1 0 87308 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_949
timestamp 1649977179
transform 1 0 88412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_961
timestamp 1649977179
transform 1 0 89516 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_973
timestamp 1649977179
transform 1 0 90620 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_979
timestamp 1649977179
transform 1 0 91172 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_981
timestamp 1649977179
transform 1 0 91356 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_993
timestamp 1649977179
transform 1 0 92460 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1005
timestamp 1649977179
transform 1 0 93564 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1017
timestamp 1649977179
transform 1 0 94668 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1029
timestamp 1649977179
transform 1 0 95772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1035
timestamp 1649977179
transform 1 0 96324 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1037
timestamp 1649977179
transform 1 0 96508 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1049
timestamp 1649977179
transform 1 0 97612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1061
timestamp 1649977179
transform 1 0 98716 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1073
timestamp 1649977179
transform 1 0 99820 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1085
timestamp 1649977179
transform 1 0 100924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1091
timestamp 1649977179
transform 1 0 101476 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1093
timestamp 1649977179
transform 1 0 101660 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1105
timestamp 1649977179
transform 1 0 102764 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1117
timestamp 1649977179
transform 1 0 103868 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1129
timestamp 1649977179
transform 1 0 104972 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1141
timestamp 1649977179
transform 1 0 106076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1147
timestamp 1649977179
transform 1 0 106628 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1149
timestamp 1649977179
transform 1 0 106812 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1161
timestamp 1649977179
transform 1 0 107916 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1173
timestamp 1649977179
transform 1 0 109020 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1185
timestamp 1649977179
transform 1 0 110124 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1197
timestamp 1649977179
transform 1 0 111228 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1203
timestamp 1649977179
transform 1 0 111780 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1205
timestamp 1649977179
transform 1 0 111964 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1217
timestamp 1649977179
transform 1 0 113068 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1229
timestamp 1649977179
transform 1 0 114172 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1241
timestamp 1649977179
transform 1 0 115276 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1253
timestamp 1649977179
transform 1 0 116380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1259
timestamp 1649977179
transform 1 0 116932 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1261
timestamp 1649977179
transform 1 0 117116 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1273
timestamp 1649977179
transform 1 0 118220 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1285
timestamp 1649977179
transform 1 0 119324 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1297
timestamp 1649977179
transform 1 0 120428 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1309
timestamp 1649977179
transform 1 0 121532 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1315
timestamp 1649977179
transform 1 0 122084 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1317
timestamp 1649977179
transform 1 0 122268 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1329
timestamp 1649977179
transform 1 0 123372 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1341
timestamp 1649977179
transform 1 0 124476 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1353
timestamp 1649977179
transform 1 0 125580 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1365
timestamp 1649977179
transform 1 0 126684 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1371
timestamp 1649977179
transform 1 0 127236 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1373
timestamp 1649977179
transform 1 0 127420 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1385
timestamp 1649977179
transform 1 0 128524 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1397
timestamp 1649977179
transform 1 0 129628 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1409
timestamp 1649977179
transform 1 0 130732 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1421
timestamp 1649977179
transform 1 0 131836 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1427
timestamp 1649977179
transform 1 0 132388 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1429
timestamp 1649977179
transform 1 0 132572 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1441
timestamp 1649977179
transform 1 0 133676 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1453
timestamp 1649977179
transform 1 0 134780 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1465
timestamp 1649977179
transform 1 0 135884 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1477
timestamp 1649977179
transform 1 0 136988 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1483
timestamp 1649977179
transform 1 0 137540 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1485
timestamp 1649977179
transform 1 0 137724 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1497
timestamp 1649977179
transform 1 0 138828 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1509
timestamp 1649977179
transform 1 0 139932 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1521
timestamp 1649977179
transform 1 0 141036 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1533
timestamp 1649977179
transform 1 0 142140 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1539
timestamp 1649977179
transform 1 0 142692 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1541
timestamp 1649977179
transform 1 0 142876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1553
timestamp 1649977179
transform 1 0 143980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1565
timestamp 1649977179
transform 1 0 145084 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1577
timestamp 1649977179
transform 1 0 146188 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1589
timestamp 1649977179
transform 1 0 147292 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1595
timestamp 1649977179
transform 1 0 147844 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1597
timestamp 1649977179
transform 1 0 148028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1609
timestamp 1649977179
transform 1 0 149132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1621
timestamp 1649977179
transform 1 0 150236 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1633
timestamp 1649977179
transform 1 0 151340 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1645
timestamp 1649977179
transform 1 0 152444 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1651
timestamp 1649977179
transform 1 0 152996 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1653
timestamp 1649977179
transform 1 0 153180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1665
timestamp 1649977179
transform 1 0 154284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1677
timestamp 1649977179
transform 1 0 155388 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1689
timestamp 1649977179
transform 1 0 156492 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1701
timestamp 1649977179
transform 1 0 157596 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1707
timestamp 1649977179
transform 1 0 158148 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1709
timestamp 1649977179
transform 1 0 158332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1721
timestamp 1649977179
transform 1 0 159436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1733
timestamp 1649977179
transform 1 0 160540 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1745
timestamp 1649977179
transform 1 0 161644 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1757
timestamp 1649977179
transform 1 0 162748 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1763
timestamp 1649977179
transform 1 0 163300 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1765
timestamp 1649977179
transform 1 0 163484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1777
timestamp 1649977179
transform 1 0 164588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1789
timestamp 1649977179
transform 1 0 165692 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1801
timestamp 1649977179
transform 1 0 166796 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1813
timestamp 1649977179
transform 1 0 167900 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1819
timestamp 1649977179
transform 1 0 168452 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1821
timestamp 1649977179
transform 1 0 168636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1833
timestamp 1649977179
transform 1 0 169740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1845
timestamp 1649977179
transform 1 0 170844 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1857
timestamp 1649977179
transform 1 0 171948 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1869
timestamp 1649977179
transform 1 0 173052 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1875
timestamp 1649977179
transform 1 0 173604 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1877
timestamp 1649977179
transform 1 0 173788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1889
timestamp 1649977179
transform 1 0 174892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1901
timestamp 1649977179
transform 1 0 175996 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1913
timestamp 1649977179
transform 1 0 177100 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1925
timestamp 1649977179
transform 1 0 178204 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1931
timestamp 1649977179
transform 1 0 178756 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1933
timestamp 1649977179
transform 1 0 178940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1945
timestamp 1649977179
transform 1 0 180044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1957
timestamp 1649977179
transform 1 0 181148 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1969
timestamp 1649977179
transform 1 0 182252 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1981
timestamp 1649977179
transform 1 0 183356 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1987
timestamp 1649977179
transform 1 0 183908 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1989
timestamp 1649977179
transform 1 0 184092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2001
timestamp 1649977179
transform 1 0 185196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2013
timestamp 1649977179
transform 1 0 186300 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2025
timestamp 1649977179
transform 1 0 187404 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2037
timestamp 1649977179
transform 1 0 188508 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2043
timestamp 1649977179
transform 1 0 189060 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2045
timestamp 1649977179
transform 1 0 189244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2057
timestamp 1649977179
transform 1 0 190348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2069
timestamp 1649977179
transform 1 0 191452 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2081
timestamp 1649977179
transform 1 0 192556 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2093
timestamp 1649977179
transform 1 0 193660 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2099
timestamp 1649977179
transform 1 0 194212 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2101
timestamp 1649977179
transform 1 0 194396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2113
timestamp 1649977179
transform 1 0 195500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2125
timestamp 1649977179
transform 1 0 196604 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2137
timestamp 1649977179
transform 1 0 197708 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2149
timestamp 1649977179
transform 1 0 198812 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2155
timestamp 1649977179
transform 1 0 199364 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2157
timestamp 1649977179
transform 1 0 199548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2169
timestamp 1649977179
transform 1 0 200652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2181
timestamp 1649977179
transform 1 0 201756 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2193
timestamp 1649977179
transform 1 0 202860 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2205
timestamp 1649977179
transform 1 0 203964 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2211
timestamp 1649977179
transform 1 0 204516 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2213
timestamp 1649977179
transform 1 0 204700 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2225
timestamp 1649977179
transform 1 0 205804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2237
timestamp 1649977179
transform 1 0 206908 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2249
timestamp 1649977179
transform 1 0 208012 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2261
timestamp 1649977179
transform 1 0 209116 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2267
timestamp 1649977179
transform 1 0 209668 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2269
timestamp 1649977179
transform 1 0 209852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2281
timestamp 1649977179
transform 1 0 210956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2293
timestamp 1649977179
transform 1 0 212060 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2305
timestamp 1649977179
transform 1 0 213164 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2317
timestamp 1649977179
transform 1 0 214268 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2323
timestamp 1649977179
transform 1 0 214820 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2325
timestamp 1649977179
transform 1 0 215004 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2337
timestamp 1649977179
transform 1 0 216108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2349
timestamp 1649977179
transform 1 0 217212 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2361
timestamp 1649977179
transform 1 0 218316 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2373
timestamp 1649977179
transform 1 0 219420 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2379
timestamp 1649977179
transform 1 0 219972 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2381
timestamp 1649977179
transform 1 0 220156 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2393
timestamp 1649977179
transform 1 0 221260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2405
timestamp 1649977179
transform 1 0 222364 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2417
timestamp 1649977179
transform 1 0 223468 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2429
timestamp 1649977179
transform 1 0 224572 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2435
timestamp 1649977179
transform 1 0 225124 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2437
timestamp 1649977179
transform 1 0 225308 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2449
timestamp 1649977179
transform 1 0 226412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2461
timestamp 1649977179
transform 1 0 227516 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2473
timestamp 1649977179
transform 1 0 228620 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2485
timestamp 1649977179
transform 1 0 229724 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2491
timestamp 1649977179
transform 1 0 230276 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2493
timestamp 1649977179
transform 1 0 230460 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2505
timestamp 1649977179
transform 1 0 231564 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2517
timestamp 1649977179
transform 1 0 232668 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2529
timestamp 1649977179
transform 1 0 233772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2541
timestamp 1649977179
transform 1 0 234876 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2547
timestamp 1649977179
transform 1 0 235428 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2549
timestamp 1649977179
transform 1 0 235612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2561
timestamp 1649977179
transform 1 0 236716 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2573
timestamp 1649977179
transform 1 0 237820 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2585
timestamp 1649977179
transform 1 0 238924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2597
timestamp 1649977179
transform 1 0 240028 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2603
timestamp 1649977179
transform 1 0 240580 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2605
timestamp 1649977179
transform 1 0 240764 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2617
timestamp 1649977179
transform 1 0 241868 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2629
timestamp 1649977179
transform 1 0 242972 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2641
timestamp 1649977179
transform 1 0 244076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2653
timestamp 1649977179
transform 1 0 245180 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2659
timestamp 1649977179
transform 1 0 245732 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2661
timestamp 1649977179
transform 1 0 245916 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2673
timestamp 1649977179
transform 1 0 247020 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2685
timestamp 1649977179
transform 1 0 248124 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2697
timestamp 1649977179
transform 1 0 249228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2709
timestamp 1649977179
transform 1 0 250332 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2715
timestamp 1649977179
transform 1 0 250884 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2717
timestamp 1649977179
transform 1 0 251068 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2729
timestamp 1649977179
transform 1 0 252172 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2741
timestamp 1649977179
transform 1 0 253276 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2753
timestamp 1649977179
transform 1 0 254380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2765
timestamp 1649977179
transform 1 0 255484 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2771
timestamp 1649977179
transform 1 0 256036 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2773
timestamp 1649977179
transform 1 0 256220 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2785
timestamp 1649977179
transform 1 0 257324 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2797
timestamp 1649977179
transform 1 0 258428 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2809
timestamp 1649977179
transform 1 0 259532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2821
timestamp 1649977179
transform 1 0 260636 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2827
timestamp 1649977179
transform 1 0 261188 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2829
timestamp 1649977179
transform 1 0 261372 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2841
timestamp 1649977179
transform 1 0 262476 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2853
timestamp 1649977179
transform 1 0 263580 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2865
timestamp 1649977179
transform 1 0 264684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2877
timestamp 1649977179
transform 1 0 265788 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2883
timestamp 1649977179
transform 1 0 266340 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2885
timestamp 1649977179
transform 1 0 266524 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2897
timestamp 1649977179
transform 1 0 267628 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2909
timestamp 1649977179
transform 1 0 268732 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2921
timestamp 1649977179
transform 1 0 269836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2933
timestamp 1649977179
transform 1 0 270940 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2939
timestamp 1649977179
transform 1 0 271492 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2941
timestamp 1649977179
transform 1 0 271676 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2953
timestamp 1649977179
transform 1 0 272780 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2965
timestamp 1649977179
transform 1 0 273884 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2977
timestamp 1649977179
transform 1 0 274988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2989
timestamp 1649977179
transform 1 0 276092 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2995
timestamp 1649977179
transform 1 0 276644 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2997
timestamp 1649977179
transform 1 0 276828 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3009
timestamp 1649977179
transform 1 0 277932 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3021
timestamp 1649977179
transform 1 0 279036 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3033
timestamp 1649977179
transform 1 0 280140 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3045
timestamp 1649977179
transform 1 0 281244 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3051
timestamp 1649977179
transform 1 0 281796 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3053
timestamp 1649977179
transform 1 0 281980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3065
timestamp 1649977179
transform 1 0 283084 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3077
timestamp 1649977179
transform 1 0 284188 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3089
timestamp 1649977179
transform 1 0 285292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3101
timestamp 1649977179
transform 1 0 286396 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3107
timestamp 1649977179
transform 1 0 286948 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3109
timestamp 1649977179
transform 1 0 287132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3121
timestamp 1649977179
transform 1 0 288236 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3133
timestamp 1649977179
transform 1 0 289340 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3145
timestamp 1649977179
transform 1 0 290444 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3157
timestamp 1649977179
transform 1 0 291548 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3163
timestamp 1649977179
transform 1 0 292100 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3165
timestamp 1649977179
transform 1 0 292284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3177
timestamp 1649977179
transform 1 0 293388 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3189
timestamp 1649977179
transform 1 0 294492 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3201
timestamp 1649977179
transform 1 0 295596 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3213
timestamp 1649977179
transform 1 0 296700 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3219
timestamp 1649977179
transform 1 0 297252 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3221
timestamp 1649977179
transform 1 0 297436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3233
timestamp 1649977179
transform 1 0 298540 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3245
timestamp 1649977179
transform 1 0 299644 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3257
timestamp 1649977179
transform 1 0 300748 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3269
timestamp 1649977179
transform 1 0 301852 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3275
timestamp 1649977179
transform 1 0 302404 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3277
timestamp 1649977179
transform 1 0 302588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3289
timestamp 1649977179
transform 1 0 303692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3301
timestamp 1649977179
transform 1 0 304796 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1649977179
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1649977179
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1649977179
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1649977179
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1649977179
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1649977179
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1649977179
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1649977179
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1649977179
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1649977179
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1649977179
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1649977179
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1649977179
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1649977179
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1649977179
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1649977179
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1649977179
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1649977179
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1649977179
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1649977179
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1649977179
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1649977179
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1649977179
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1649977179
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1649977179
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1649977179
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1649977179
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1649977179
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1649977179
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1649977179
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1649977179
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1649977179
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1649977179
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1649977179
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1649977179
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1649977179
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1649977179
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1649977179
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1649977179
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1649977179
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_617
timestamp 1649977179
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_629
timestamp 1649977179
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_641
timestamp 1649977179
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_653
timestamp 1649977179
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1649977179
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1649977179
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_673
timestamp 1649977179
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_685
timestamp 1649977179
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_697
timestamp 1649977179
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_709
timestamp 1649977179
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 1649977179
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1649977179
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_729
timestamp 1649977179
transform 1 0 68172 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_741
timestamp 1649977179
transform 1 0 69276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_753
timestamp 1649977179
transform 1 0 70380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_765
timestamp 1649977179
transform 1 0 71484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_777
timestamp 1649977179
transform 1 0 72588 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_783
timestamp 1649977179
transform 1 0 73140 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_785
timestamp 1649977179
transform 1 0 73324 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_797
timestamp 1649977179
transform 1 0 74428 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_809
timestamp 1649977179
transform 1 0 75532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_821
timestamp 1649977179
transform 1 0 76636 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_833
timestamp 1649977179
transform 1 0 77740 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_839
timestamp 1649977179
transform 1 0 78292 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_841
timestamp 1649977179
transform 1 0 78476 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_853
timestamp 1649977179
transform 1 0 79580 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_865
timestamp 1649977179
transform 1 0 80684 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_877
timestamp 1649977179
transform 1 0 81788 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_889
timestamp 1649977179
transform 1 0 82892 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_895
timestamp 1649977179
transform 1 0 83444 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_897
timestamp 1649977179
transform 1 0 83628 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_909
timestamp 1649977179
transform 1 0 84732 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_921
timestamp 1649977179
transform 1 0 85836 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_933
timestamp 1649977179
transform 1 0 86940 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_945
timestamp 1649977179
transform 1 0 88044 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_951
timestamp 1649977179
transform 1 0 88596 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_953
timestamp 1649977179
transform 1 0 88780 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_965
timestamp 1649977179
transform 1 0 89884 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_977
timestamp 1649977179
transform 1 0 90988 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_989
timestamp 1649977179
transform 1 0 92092 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1001
timestamp 1649977179
transform 1 0 93196 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1007
timestamp 1649977179
transform 1 0 93748 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1009
timestamp 1649977179
transform 1 0 93932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1021
timestamp 1649977179
transform 1 0 95036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1033
timestamp 1649977179
transform 1 0 96140 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1045
timestamp 1649977179
transform 1 0 97244 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1057
timestamp 1649977179
transform 1 0 98348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1063
timestamp 1649977179
transform 1 0 98900 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1065
timestamp 1649977179
transform 1 0 99084 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1077
timestamp 1649977179
transform 1 0 100188 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1089
timestamp 1649977179
transform 1 0 101292 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1101
timestamp 1649977179
transform 1 0 102396 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1113
timestamp 1649977179
transform 1 0 103500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1119
timestamp 1649977179
transform 1 0 104052 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1121
timestamp 1649977179
transform 1 0 104236 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1133
timestamp 1649977179
transform 1 0 105340 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1145
timestamp 1649977179
transform 1 0 106444 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1157
timestamp 1649977179
transform 1 0 107548 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1169
timestamp 1649977179
transform 1 0 108652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1175
timestamp 1649977179
transform 1 0 109204 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1177
timestamp 1649977179
transform 1 0 109388 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1189
timestamp 1649977179
transform 1 0 110492 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1201
timestamp 1649977179
transform 1 0 111596 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1213
timestamp 1649977179
transform 1 0 112700 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1225
timestamp 1649977179
transform 1 0 113804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1231
timestamp 1649977179
transform 1 0 114356 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1233
timestamp 1649977179
transform 1 0 114540 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1245
timestamp 1649977179
transform 1 0 115644 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1257
timestamp 1649977179
transform 1 0 116748 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1269
timestamp 1649977179
transform 1 0 117852 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1281
timestamp 1649977179
transform 1 0 118956 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1287
timestamp 1649977179
transform 1 0 119508 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1289
timestamp 1649977179
transform 1 0 119692 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1301
timestamp 1649977179
transform 1 0 120796 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1313
timestamp 1649977179
transform 1 0 121900 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1325
timestamp 1649977179
transform 1 0 123004 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1337
timestamp 1649977179
transform 1 0 124108 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1343
timestamp 1649977179
transform 1 0 124660 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1345
timestamp 1649977179
transform 1 0 124844 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1357
timestamp 1649977179
transform 1 0 125948 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1369
timestamp 1649977179
transform 1 0 127052 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1381
timestamp 1649977179
transform 1 0 128156 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1393
timestamp 1649977179
transform 1 0 129260 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1399
timestamp 1649977179
transform 1 0 129812 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1401
timestamp 1649977179
transform 1 0 129996 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1413
timestamp 1649977179
transform 1 0 131100 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1425
timestamp 1649977179
transform 1 0 132204 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1437
timestamp 1649977179
transform 1 0 133308 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1449
timestamp 1649977179
transform 1 0 134412 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1455
timestamp 1649977179
transform 1 0 134964 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1457
timestamp 1649977179
transform 1 0 135148 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1469
timestamp 1649977179
transform 1 0 136252 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1481
timestamp 1649977179
transform 1 0 137356 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1493
timestamp 1649977179
transform 1 0 138460 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1505
timestamp 1649977179
transform 1 0 139564 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1511
timestamp 1649977179
transform 1 0 140116 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1513
timestamp 1649977179
transform 1 0 140300 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1525
timestamp 1649977179
transform 1 0 141404 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1537
timestamp 1649977179
transform 1 0 142508 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1549
timestamp 1649977179
transform 1 0 143612 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1561
timestamp 1649977179
transform 1 0 144716 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1567
timestamp 1649977179
transform 1 0 145268 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1569
timestamp 1649977179
transform 1 0 145452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1581
timestamp 1649977179
transform 1 0 146556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1593
timestamp 1649977179
transform 1 0 147660 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1605
timestamp 1649977179
transform 1 0 148764 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1617
timestamp 1649977179
transform 1 0 149868 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1623
timestamp 1649977179
transform 1 0 150420 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1625
timestamp 1649977179
transform 1 0 150604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1637
timestamp 1649977179
transform 1 0 151708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1649
timestamp 1649977179
transform 1 0 152812 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1661
timestamp 1649977179
transform 1 0 153916 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1673
timestamp 1649977179
transform 1 0 155020 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1679
timestamp 1649977179
transform 1 0 155572 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1681
timestamp 1649977179
transform 1 0 155756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1693
timestamp 1649977179
transform 1 0 156860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1705
timestamp 1649977179
transform 1 0 157964 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1717
timestamp 1649977179
transform 1 0 159068 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1729
timestamp 1649977179
transform 1 0 160172 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1735
timestamp 1649977179
transform 1 0 160724 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1737
timestamp 1649977179
transform 1 0 160908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1749
timestamp 1649977179
transform 1 0 162012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1761
timestamp 1649977179
transform 1 0 163116 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1773
timestamp 1649977179
transform 1 0 164220 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1785
timestamp 1649977179
transform 1 0 165324 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1791
timestamp 1649977179
transform 1 0 165876 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1793
timestamp 1649977179
transform 1 0 166060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1805
timestamp 1649977179
transform 1 0 167164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1817
timestamp 1649977179
transform 1 0 168268 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1829
timestamp 1649977179
transform 1 0 169372 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1841
timestamp 1649977179
transform 1 0 170476 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1847
timestamp 1649977179
transform 1 0 171028 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1849
timestamp 1649977179
transform 1 0 171212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1861
timestamp 1649977179
transform 1 0 172316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1873
timestamp 1649977179
transform 1 0 173420 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1885
timestamp 1649977179
transform 1 0 174524 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1897
timestamp 1649977179
transform 1 0 175628 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1903
timestamp 1649977179
transform 1 0 176180 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1905
timestamp 1649977179
transform 1 0 176364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1917
timestamp 1649977179
transform 1 0 177468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1929
timestamp 1649977179
transform 1 0 178572 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1941
timestamp 1649977179
transform 1 0 179676 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1953
timestamp 1649977179
transform 1 0 180780 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1959
timestamp 1649977179
transform 1 0 181332 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1961
timestamp 1649977179
transform 1 0 181516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1973
timestamp 1649977179
transform 1 0 182620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1985
timestamp 1649977179
transform 1 0 183724 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1997
timestamp 1649977179
transform 1 0 184828 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2009
timestamp 1649977179
transform 1 0 185932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2015
timestamp 1649977179
transform 1 0 186484 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2017
timestamp 1649977179
transform 1 0 186668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2029
timestamp 1649977179
transform 1 0 187772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2041
timestamp 1649977179
transform 1 0 188876 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2053
timestamp 1649977179
transform 1 0 189980 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2065
timestamp 1649977179
transform 1 0 191084 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2071
timestamp 1649977179
transform 1 0 191636 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2073
timestamp 1649977179
transform 1 0 191820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2085
timestamp 1649977179
transform 1 0 192924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2097
timestamp 1649977179
transform 1 0 194028 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2109
timestamp 1649977179
transform 1 0 195132 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2121
timestamp 1649977179
transform 1 0 196236 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2127
timestamp 1649977179
transform 1 0 196788 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2129
timestamp 1649977179
transform 1 0 196972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2141
timestamp 1649977179
transform 1 0 198076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2153
timestamp 1649977179
transform 1 0 199180 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2165
timestamp 1649977179
transform 1 0 200284 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2177
timestamp 1649977179
transform 1 0 201388 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2183
timestamp 1649977179
transform 1 0 201940 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2185
timestamp 1649977179
transform 1 0 202124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2197
timestamp 1649977179
transform 1 0 203228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2209
timestamp 1649977179
transform 1 0 204332 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2221
timestamp 1649977179
transform 1 0 205436 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2233
timestamp 1649977179
transform 1 0 206540 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2239
timestamp 1649977179
transform 1 0 207092 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2241
timestamp 1649977179
transform 1 0 207276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2253
timestamp 1649977179
transform 1 0 208380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2265
timestamp 1649977179
transform 1 0 209484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2277
timestamp 1649977179
transform 1 0 210588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2289
timestamp 1649977179
transform 1 0 211692 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2295
timestamp 1649977179
transform 1 0 212244 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2297
timestamp 1649977179
transform 1 0 212428 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2309
timestamp 1649977179
transform 1 0 213532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2321
timestamp 1649977179
transform 1 0 214636 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2333
timestamp 1649977179
transform 1 0 215740 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2345
timestamp 1649977179
transform 1 0 216844 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2351
timestamp 1649977179
transform 1 0 217396 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2353
timestamp 1649977179
transform 1 0 217580 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2365
timestamp 1649977179
transform 1 0 218684 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2377
timestamp 1649977179
transform 1 0 219788 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2389
timestamp 1649977179
transform 1 0 220892 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2401
timestamp 1649977179
transform 1 0 221996 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2407
timestamp 1649977179
transform 1 0 222548 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2409
timestamp 1649977179
transform 1 0 222732 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2421
timestamp 1649977179
transform 1 0 223836 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2433
timestamp 1649977179
transform 1 0 224940 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2445
timestamp 1649977179
transform 1 0 226044 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2457
timestamp 1649977179
transform 1 0 227148 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2463
timestamp 1649977179
transform 1 0 227700 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2465
timestamp 1649977179
transform 1 0 227884 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2477
timestamp 1649977179
transform 1 0 228988 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2489
timestamp 1649977179
transform 1 0 230092 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2501
timestamp 1649977179
transform 1 0 231196 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2513
timestamp 1649977179
transform 1 0 232300 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2519
timestamp 1649977179
transform 1 0 232852 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2521
timestamp 1649977179
transform 1 0 233036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2533
timestamp 1649977179
transform 1 0 234140 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2545
timestamp 1649977179
transform 1 0 235244 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2557
timestamp 1649977179
transform 1 0 236348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2569
timestamp 1649977179
transform 1 0 237452 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2575
timestamp 1649977179
transform 1 0 238004 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2577
timestamp 1649977179
transform 1 0 238188 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2589
timestamp 1649977179
transform 1 0 239292 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2601
timestamp 1649977179
transform 1 0 240396 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2613
timestamp 1649977179
transform 1 0 241500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2625
timestamp 1649977179
transform 1 0 242604 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2631
timestamp 1649977179
transform 1 0 243156 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2633
timestamp 1649977179
transform 1 0 243340 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2645
timestamp 1649977179
transform 1 0 244444 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2657
timestamp 1649977179
transform 1 0 245548 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2669
timestamp 1649977179
transform 1 0 246652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2681
timestamp 1649977179
transform 1 0 247756 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2687
timestamp 1649977179
transform 1 0 248308 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2689
timestamp 1649977179
transform 1 0 248492 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2701
timestamp 1649977179
transform 1 0 249596 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2713
timestamp 1649977179
transform 1 0 250700 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2725
timestamp 1649977179
transform 1 0 251804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2737
timestamp 1649977179
transform 1 0 252908 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2743
timestamp 1649977179
transform 1 0 253460 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2745
timestamp 1649977179
transform 1 0 253644 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2757
timestamp 1649977179
transform 1 0 254748 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2769
timestamp 1649977179
transform 1 0 255852 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2781
timestamp 1649977179
transform 1 0 256956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2793
timestamp 1649977179
transform 1 0 258060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2799
timestamp 1649977179
transform 1 0 258612 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2801
timestamp 1649977179
transform 1 0 258796 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2813
timestamp 1649977179
transform 1 0 259900 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2825
timestamp 1649977179
transform 1 0 261004 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2837
timestamp 1649977179
transform 1 0 262108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2849
timestamp 1649977179
transform 1 0 263212 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2855
timestamp 1649977179
transform 1 0 263764 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2857
timestamp 1649977179
transform 1 0 263948 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2869
timestamp 1649977179
transform 1 0 265052 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2881
timestamp 1649977179
transform 1 0 266156 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2893
timestamp 1649977179
transform 1 0 267260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2905
timestamp 1649977179
transform 1 0 268364 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2911
timestamp 1649977179
transform 1 0 268916 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2913
timestamp 1649977179
transform 1 0 269100 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2925
timestamp 1649977179
transform 1 0 270204 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2937
timestamp 1649977179
transform 1 0 271308 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2949
timestamp 1649977179
transform 1 0 272412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2961
timestamp 1649977179
transform 1 0 273516 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2967
timestamp 1649977179
transform 1 0 274068 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2969
timestamp 1649977179
transform 1 0 274252 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2981
timestamp 1649977179
transform 1 0 275356 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2993
timestamp 1649977179
transform 1 0 276460 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3005
timestamp 1649977179
transform 1 0 277564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3017
timestamp 1649977179
transform 1 0 278668 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3023
timestamp 1649977179
transform 1 0 279220 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3025
timestamp 1649977179
transform 1 0 279404 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3037
timestamp 1649977179
transform 1 0 280508 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3049
timestamp 1649977179
transform 1 0 281612 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3061
timestamp 1649977179
transform 1 0 282716 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3073
timestamp 1649977179
transform 1 0 283820 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3079
timestamp 1649977179
transform 1 0 284372 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3081
timestamp 1649977179
transform 1 0 284556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3093
timestamp 1649977179
transform 1 0 285660 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3105
timestamp 1649977179
transform 1 0 286764 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3117
timestamp 1649977179
transform 1 0 287868 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3129
timestamp 1649977179
transform 1 0 288972 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3135
timestamp 1649977179
transform 1 0 289524 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3137
timestamp 1649977179
transform 1 0 289708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3149
timestamp 1649977179
transform 1 0 290812 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3161
timestamp 1649977179
transform 1 0 291916 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3173
timestamp 1649977179
transform 1 0 293020 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3185
timestamp 1649977179
transform 1 0 294124 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3191
timestamp 1649977179
transform 1 0 294676 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3193
timestamp 1649977179
transform 1 0 294860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3205
timestamp 1649977179
transform 1 0 295964 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3217
timestamp 1649977179
transform 1 0 297068 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3229
timestamp 1649977179
transform 1 0 298172 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3241
timestamp 1649977179
transform 1 0 299276 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3247
timestamp 1649977179
transform 1 0 299828 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3249
timestamp 1649977179
transform 1 0 300012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3261
timestamp 1649977179
transform 1 0 301116 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3273
timestamp 1649977179
transform 1 0 302220 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3285
timestamp 1649977179
transform 1 0 303324 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3300
timestamp 1649977179
transform 1 0 304704 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3305
timestamp 1649977179
transform 1 0 305164 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1649977179
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1649977179
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1649977179
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1649977179
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1649977179
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1649977179
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1649977179
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1649977179
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1649977179
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1649977179
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1649977179
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1649977179
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1649977179
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1649977179
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1649977179
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1649977179
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1649977179
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1649977179
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1649977179
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1649977179
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1649977179
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1649977179
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1649977179
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1649977179
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1649977179
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1649977179
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1649977179
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1649977179
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1649977179
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1649977179
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1649977179
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1649977179
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1649977179
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1649977179
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1649977179
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1649977179
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1649977179
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1649977179
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1649977179
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1649977179
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1649977179
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_625
timestamp 1649977179
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1649977179
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1649977179
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_645
timestamp 1649977179
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_657
timestamp 1649977179
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_669
timestamp 1649977179
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_681
timestamp 1649977179
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1649977179
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1649977179
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_701
timestamp 1649977179
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_713
timestamp 1649977179
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_725
timestamp 1649977179
transform 1 0 67804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_737
timestamp 1649977179
transform 1 0 68908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_749
timestamp 1649977179
transform 1 0 70012 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_755
timestamp 1649977179
transform 1 0 70564 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_757
timestamp 1649977179
transform 1 0 70748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_769
timestamp 1649977179
transform 1 0 71852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_781
timestamp 1649977179
transform 1 0 72956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_793
timestamp 1649977179
transform 1 0 74060 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_805
timestamp 1649977179
transform 1 0 75164 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_811
timestamp 1649977179
transform 1 0 75716 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_813
timestamp 1649977179
transform 1 0 75900 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_825
timestamp 1649977179
transform 1 0 77004 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_837
timestamp 1649977179
transform 1 0 78108 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_849
timestamp 1649977179
transform 1 0 79212 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_861
timestamp 1649977179
transform 1 0 80316 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_867
timestamp 1649977179
transform 1 0 80868 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_869
timestamp 1649977179
transform 1 0 81052 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_881
timestamp 1649977179
transform 1 0 82156 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_893
timestamp 1649977179
transform 1 0 83260 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_905
timestamp 1649977179
transform 1 0 84364 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_917
timestamp 1649977179
transform 1 0 85468 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_923
timestamp 1649977179
transform 1 0 86020 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_925
timestamp 1649977179
transform 1 0 86204 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_937
timestamp 1649977179
transform 1 0 87308 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_949
timestamp 1649977179
transform 1 0 88412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_961
timestamp 1649977179
transform 1 0 89516 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_973
timestamp 1649977179
transform 1 0 90620 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_979
timestamp 1649977179
transform 1 0 91172 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_981
timestamp 1649977179
transform 1 0 91356 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_993
timestamp 1649977179
transform 1 0 92460 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1005
timestamp 1649977179
transform 1 0 93564 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1017
timestamp 1649977179
transform 1 0 94668 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1029
timestamp 1649977179
transform 1 0 95772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1035
timestamp 1649977179
transform 1 0 96324 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1037
timestamp 1649977179
transform 1 0 96508 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1049
timestamp 1649977179
transform 1 0 97612 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1061
timestamp 1649977179
transform 1 0 98716 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1073
timestamp 1649977179
transform 1 0 99820 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1085
timestamp 1649977179
transform 1 0 100924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1091
timestamp 1649977179
transform 1 0 101476 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1093
timestamp 1649977179
transform 1 0 101660 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1105
timestamp 1649977179
transform 1 0 102764 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1117
timestamp 1649977179
transform 1 0 103868 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1129
timestamp 1649977179
transform 1 0 104972 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1141
timestamp 1649977179
transform 1 0 106076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1147
timestamp 1649977179
transform 1 0 106628 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1149
timestamp 1649977179
transform 1 0 106812 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1161
timestamp 1649977179
transform 1 0 107916 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1173
timestamp 1649977179
transform 1 0 109020 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1185
timestamp 1649977179
transform 1 0 110124 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1197
timestamp 1649977179
transform 1 0 111228 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1203
timestamp 1649977179
transform 1 0 111780 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1205
timestamp 1649977179
transform 1 0 111964 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1217
timestamp 1649977179
transform 1 0 113068 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1229
timestamp 1649977179
transform 1 0 114172 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1241
timestamp 1649977179
transform 1 0 115276 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1253
timestamp 1649977179
transform 1 0 116380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1259
timestamp 1649977179
transform 1 0 116932 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1261
timestamp 1649977179
transform 1 0 117116 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1273
timestamp 1649977179
transform 1 0 118220 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1285
timestamp 1649977179
transform 1 0 119324 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1297
timestamp 1649977179
transform 1 0 120428 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1309
timestamp 1649977179
transform 1 0 121532 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1315
timestamp 1649977179
transform 1 0 122084 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1317
timestamp 1649977179
transform 1 0 122268 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1329
timestamp 1649977179
transform 1 0 123372 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1341
timestamp 1649977179
transform 1 0 124476 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1353
timestamp 1649977179
transform 1 0 125580 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1365
timestamp 1649977179
transform 1 0 126684 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1371
timestamp 1649977179
transform 1 0 127236 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1373
timestamp 1649977179
transform 1 0 127420 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1385
timestamp 1649977179
transform 1 0 128524 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1397
timestamp 1649977179
transform 1 0 129628 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1409
timestamp 1649977179
transform 1 0 130732 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1421
timestamp 1649977179
transform 1 0 131836 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1427
timestamp 1649977179
transform 1 0 132388 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1429
timestamp 1649977179
transform 1 0 132572 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1441
timestamp 1649977179
transform 1 0 133676 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1453
timestamp 1649977179
transform 1 0 134780 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1465
timestamp 1649977179
transform 1 0 135884 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1477
timestamp 1649977179
transform 1 0 136988 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1483
timestamp 1649977179
transform 1 0 137540 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1485
timestamp 1649977179
transform 1 0 137724 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1497
timestamp 1649977179
transform 1 0 138828 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1509
timestamp 1649977179
transform 1 0 139932 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1521
timestamp 1649977179
transform 1 0 141036 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1533
timestamp 1649977179
transform 1 0 142140 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1539
timestamp 1649977179
transform 1 0 142692 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1541
timestamp 1649977179
transform 1 0 142876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1553
timestamp 1649977179
transform 1 0 143980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1565
timestamp 1649977179
transform 1 0 145084 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1577
timestamp 1649977179
transform 1 0 146188 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1589
timestamp 1649977179
transform 1 0 147292 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1595
timestamp 1649977179
transform 1 0 147844 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1597
timestamp 1649977179
transform 1 0 148028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1609
timestamp 1649977179
transform 1 0 149132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1621
timestamp 1649977179
transform 1 0 150236 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1633
timestamp 1649977179
transform 1 0 151340 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1645
timestamp 1649977179
transform 1 0 152444 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1651
timestamp 1649977179
transform 1 0 152996 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1653
timestamp 1649977179
transform 1 0 153180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1665
timestamp 1649977179
transform 1 0 154284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1677
timestamp 1649977179
transform 1 0 155388 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1689
timestamp 1649977179
transform 1 0 156492 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1701
timestamp 1649977179
transform 1 0 157596 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1707
timestamp 1649977179
transform 1 0 158148 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1709
timestamp 1649977179
transform 1 0 158332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1721
timestamp 1649977179
transform 1 0 159436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1733
timestamp 1649977179
transform 1 0 160540 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1745
timestamp 1649977179
transform 1 0 161644 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1757
timestamp 1649977179
transform 1 0 162748 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1763
timestamp 1649977179
transform 1 0 163300 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1765
timestamp 1649977179
transform 1 0 163484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1777
timestamp 1649977179
transform 1 0 164588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1789
timestamp 1649977179
transform 1 0 165692 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1801
timestamp 1649977179
transform 1 0 166796 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1813
timestamp 1649977179
transform 1 0 167900 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1819
timestamp 1649977179
transform 1 0 168452 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1821
timestamp 1649977179
transform 1 0 168636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1833
timestamp 1649977179
transform 1 0 169740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1845
timestamp 1649977179
transform 1 0 170844 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1857
timestamp 1649977179
transform 1 0 171948 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1869
timestamp 1649977179
transform 1 0 173052 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1875
timestamp 1649977179
transform 1 0 173604 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1877
timestamp 1649977179
transform 1 0 173788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1889
timestamp 1649977179
transform 1 0 174892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1901
timestamp 1649977179
transform 1 0 175996 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1913
timestamp 1649977179
transform 1 0 177100 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1925
timestamp 1649977179
transform 1 0 178204 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1931
timestamp 1649977179
transform 1 0 178756 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1933
timestamp 1649977179
transform 1 0 178940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1945
timestamp 1649977179
transform 1 0 180044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1957
timestamp 1649977179
transform 1 0 181148 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1969
timestamp 1649977179
transform 1 0 182252 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1981
timestamp 1649977179
transform 1 0 183356 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1987
timestamp 1649977179
transform 1 0 183908 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1989
timestamp 1649977179
transform 1 0 184092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2001
timestamp 1649977179
transform 1 0 185196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2013
timestamp 1649977179
transform 1 0 186300 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2025
timestamp 1649977179
transform 1 0 187404 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2037
timestamp 1649977179
transform 1 0 188508 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2043
timestamp 1649977179
transform 1 0 189060 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2045
timestamp 1649977179
transform 1 0 189244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2057
timestamp 1649977179
transform 1 0 190348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2069
timestamp 1649977179
transform 1 0 191452 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2081
timestamp 1649977179
transform 1 0 192556 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2093
timestamp 1649977179
transform 1 0 193660 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2099
timestamp 1649977179
transform 1 0 194212 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2101
timestamp 1649977179
transform 1 0 194396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2113
timestamp 1649977179
transform 1 0 195500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2125
timestamp 1649977179
transform 1 0 196604 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2137
timestamp 1649977179
transform 1 0 197708 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2149
timestamp 1649977179
transform 1 0 198812 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2155
timestamp 1649977179
transform 1 0 199364 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2157
timestamp 1649977179
transform 1 0 199548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2169
timestamp 1649977179
transform 1 0 200652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2181
timestamp 1649977179
transform 1 0 201756 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2193
timestamp 1649977179
transform 1 0 202860 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2205
timestamp 1649977179
transform 1 0 203964 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2211
timestamp 1649977179
transform 1 0 204516 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2213
timestamp 1649977179
transform 1 0 204700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2225
timestamp 1649977179
transform 1 0 205804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2237
timestamp 1649977179
transform 1 0 206908 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2249
timestamp 1649977179
transform 1 0 208012 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2261
timestamp 1649977179
transform 1 0 209116 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2267
timestamp 1649977179
transform 1 0 209668 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2269
timestamp 1649977179
transform 1 0 209852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2281
timestamp 1649977179
transform 1 0 210956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2293
timestamp 1649977179
transform 1 0 212060 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2305
timestamp 1649977179
transform 1 0 213164 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2317
timestamp 1649977179
transform 1 0 214268 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2323
timestamp 1649977179
transform 1 0 214820 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2325
timestamp 1649977179
transform 1 0 215004 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2337
timestamp 1649977179
transform 1 0 216108 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2349
timestamp 1649977179
transform 1 0 217212 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2361
timestamp 1649977179
transform 1 0 218316 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2373
timestamp 1649977179
transform 1 0 219420 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2379
timestamp 1649977179
transform 1 0 219972 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2381
timestamp 1649977179
transform 1 0 220156 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2393
timestamp 1649977179
transform 1 0 221260 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2405
timestamp 1649977179
transform 1 0 222364 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2417
timestamp 1649977179
transform 1 0 223468 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2429
timestamp 1649977179
transform 1 0 224572 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2435
timestamp 1649977179
transform 1 0 225124 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2437
timestamp 1649977179
transform 1 0 225308 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2449
timestamp 1649977179
transform 1 0 226412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2461
timestamp 1649977179
transform 1 0 227516 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2473
timestamp 1649977179
transform 1 0 228620 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2485
timestamp 1649977179
transform 1 0 229724 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2491
timestamp 1649977179
transform 1 0 230276 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2493
timestamp 1649977179
transform 1 0 230460 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2505
timestamp 1649977179
transform 1 0 231564 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2517
timestamp 1649977179
transform 1 0 232668 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2529
timestamp 1649977179
transform 1 0 233772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2541
timestamp 1649977179
transform 1 0 234876 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2547
timestamp 1649977179
transform 1 0 235428 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2549
timestamp 1649977179
transform 1 0 235612 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2561
timestamp 1649977179
transform 1 0 236716 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2573
timestamp 1649977179
transform 1 0 237820 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2585
timestamp 1649977179
transform 1 0 238924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2597
timestamp 1649977179
transform 1 0 240028 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2603
timestamp 1649977179
transform 1 0 240580 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2605
timestamp 1649977179
transform 1 0 240764 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2617
timestamp 1649977179
transform 1 0 241868 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2629
timestamp 1649977179
transform 1 0 242972 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2641
timestamp 1649977179
transform 1 0 244076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2653
timestamp 1649977179
transform 1 0 245180 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2659
timestamp 1649977179
transform 1 0 245732 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2661
timestamp 1649977179
transform 1 0 245916 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2673
timestamp 1649977179
transform 1 0 247020 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2685
timestamp 1649977179
transform 1 0 248124 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2697
timestamp 1649977179
transform 1 0 249228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2709
timestamp 1649977179
transform 1 0 250332 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2715
timestamp 1649977179
transform 1 0 250884 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2717
timestamp 1649977179
transform 1 0 251068 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2729
timestamp 1649977179
transform 1 0 252172 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2741
timestamp 1649977179
transform 1 0 253276 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2753
timestamp 1649977179
transform 1 0 254380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2765
timestamp 1649977179
transform 1 0 255484 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2771
timestamp 1649977179
transform 1 0 256036 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2773
timestamp 1649977179
transform 1 0 256220 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2785
timestamp 1649977179
transform 1 0 257324 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2797
timestamp 1649977179
transform 1 0 258428 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2809
timestamp 1649977179
transform 1 0 259532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2821
timestamp 1649977179
transform 1 0 260636 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2827
timestamp 1649977179
transform 1 0 261188 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2829
timestamp 1649977179
transform 1 0 261372 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2841
timestamp 1649977179
transform 1 0 262476 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2853
timestamp 1649977179
transform 1 0 263580 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2865
timestamp 1649977179
transform 1 0 264684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2877
timestamp 1649977179
transform 1 0 265788 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2883
timestamp 1649977179
transform 1 0 266340 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2885
timestamp 1649977179
transform 1 0 266524 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2897
timestamp 1649977179
transform 1 0 267628 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2909
timestamp 1649977179
transform 1 0 268732 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2921
timestamp 1649977179
transform 1 0 269836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2933
timestamp 1649977179
transform 1 0 270940 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2939
timestamp 1649977179
transform 1 0 271492 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2941
timestamp 1649977179
transform 1 0 271676 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2953
timestamp 1649977179
transform 1 0 272780 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2965
timestamp 1649977179
transform 1 0 273884 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2977
timestamp 1649977179
transform 1 0 274988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2989
timestamp 1649977179
transform 1 0 276092 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2995
timestamp 1649977179
transform 1 0 276644 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2997
timestamp 1649977179
transform 1 0 276828 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3009
timestamp 1649977179
transform 1 0 277932 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3021
timestamp 1649977179
transform 1 0 279036 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3033
timestamp 1649977179
transform 1 0 280140 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3045
timestamp 1649977179
transform 1 0 281244 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3051
timestamp 1649977179
transform 1 0 281796 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3053
timestamp 1649977179
transform 1 0 281980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3065
timestamp 1649977179
transform 1 0 283084 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3077
timestamp 1649977179
transform 1 0 284188 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3089
timestamp 1649977179
transform 1 0 285292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3101
timestamp 1649977179
transform 1 0 286396 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3107
timestamp 1649977179
transform 1 0 286948 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3109
timestamp 1649977179
transform 1 0 287132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3121
timestamp 1649977179
transform 1 0 288236 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3133
timestamp 1649977179
transform 1 0 289340 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3145
timestamp 1649977179
transform 1 0 290444 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3157
timestamp 1649977179
transform 1 0 291548 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3163
timestamp 1649977179
transform 1 0 292100 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3165
timestamp 1649977179
transform 1 0 292284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3177
timestamp 1649977179
transform 1 0 293388 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3189
timestamp 1649977179
transform 1 0 294492 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3201
timestamp 1649977179
transform 1 0 295596 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3213
timestamp 1649977179
transform 1 0 296700 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3219
timestamp 1649977179
transform 1 0 297252 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3221
timestamp 1649977179
transform 1 0 297436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3233
timestamp 1649977179
transform 1 0 298540 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3245
timestamp 1649977179
transform 1 0 299644 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3257
timestamp 1649977179
transform 1 0 300748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3269
timestamp 1649977179
transform 1 0 301852 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3275
timestamp 1649977179
transform 1 0 302404 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3277
timestamp 1649977179
transform 1 0 302588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3289
timestamp 1649977179
transform 1 0 303692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_3301
timestamp 1649977179
transform 1 0 304796 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1649977179
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1649977179
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1649977179
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1649977179
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1649977179
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1649977179
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1649977179
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1649977179
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1649977179
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1649977179
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1649977179
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1649977179
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1649977179
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1649977179
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1649977179
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1649977179
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1649977179
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1649977179
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1649977179
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1649977179
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1649977179
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1649977179
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1649977179
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1649977179
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1649977179
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1649977179
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1649977179
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1649977179
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1649977179
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1649977179
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1649977179
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1649977179
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1649977179
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1649977179
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1649977179
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1649977179
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1649977179
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1649977179
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1649977179
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1649977179
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_597
timestamp 1649977179
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1649977179
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1649977179
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_617
timestamp 1649977179
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_629
timestamp 1649977179
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_641
timestamp 1649977179
transform 1 0 60076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_653
timestamp 1649977179
transform 1 0 61180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_665
timestamp 1649977179
transform 1 0 62284 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_671
timestamp 1649977179
transform 1 0 62836 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_673
timestamp 1649977179
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_685
timestamp 1649977179
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_697
timestamp 1649977179
transform 1 0 65228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_709
timestamp 1649977179
transform 1 0 66332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_721
timestamp 1649977179
transform 1 0 67436 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_727
timestamp 1649977179
transform 1 0 67988 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_729
timestamp 1649977179
transform 1 0 68172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_741
timestamp 1649977179
transform 1 0 69276 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_753
timestamp 1649977179
transform 1 0 70380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_765
timestamp 1649977179
transform 1 0 71484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_777
timestamp 1649977179
transform 1 0 72588 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_783
timestamp 1649977179
transform 1 0 73140 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_785
timestamp 1649977179
transform 1 0 73324 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_797
timestamp 1649977179
transform 1 0 74428 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_809
timestamp 1649977179
transform 1 0 75532 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_821
timestamp 1649977179
transform 1 0 76636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_833
timestamp 1649977179
transform 1 0 77740 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_839
timestamp 1649977179
transform 1 0 78292 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_841
timestamp 1649977179
transform 1 0 78476 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_853
timestamp 1649977179
transform 1 0 79580 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_865
timestamp 1649977179
transform 1 0 80684 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_877
timestamp 1649977179
transform 1 0 81788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_889
timestamp 1649977179
transform 1 0 82892 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_895
timestamp 1649977179
transform 1 0 83444 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_897
timestamp 1649977179
transform 1 0 83628 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_909
timestamp 1649977179
transform 1 0 84732 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_921
timestamp 1649977179
transform 1 0 85836 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_933
timestamp 1649977179
transform 1 0 86940 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_945
timestamp 1649977179
transform 1 0 88044 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_951
timestamp 1649977179
transform 1 0 88596 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_953
timestamp 1649977179
transform 1 0 88780 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_965
timestamp 1649977179
transform 1 0 89884 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_977
timestamp 1649977179
transform 1 0 90988 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_989
timestamp 1649977179
transform 1 0 92092 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1001
timestamp 1649977179
transform 1 0 93196 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1007
timestamp 1649977179
transform 1 0 93748 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1009
timestamp 1649977179
transform 1 0 93932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1021
timestamp 1649977179
transform 1 0 95036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1033
timestamp 1649977179
transform 1 0 96140 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1045
timestamp 1649977179
transform 1 0 97244 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1057
timestamp 1649977179
transform 1 0 98348 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1063
timestamp 1649977179
transform 1 0 98900 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1065
timestamp 1649977179
transform 1 0 99084 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1077
timestamp 1649977179
transform 1 0 100188 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1089
timestamp 1649977179
transform 1 0 101292 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1101
timestamp 1649977179
transform 1 0 102396 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1113
timestamp 1649977179
transform 1 0 103500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1119
timestamp 1649977179
transform 1 0 104052 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1121
timestamp 1649977179
transform 1 0 104236 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1133
timestamp 1649977179
transform 1 0 105340 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1145
timestamp 1649977179
transform 1 0 106444 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1157
timestamp 1649977179
transform 1 0 107548 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1169
timestamp 1649977179
transform 1 0 108652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1175
timestamp 1649977179
transform 1 0 109204 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1177
timestamp 1649977179
transform 1 0 109388 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1189
timestamp 1649977179
transform 1 0 110492 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1201
timestamp 1649977179
transform 1 0 111596 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1213
timestamp 1649977179
transform 1 0 112700 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1225
timestamp 1649977179
transform 1 0 113804 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1231
timestamp 1649977179
transform 1 0 114356 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1233
timestamp 1649977179
transform 1 0 114540 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1245
timestamp 1649977179
transform 1 0 115644 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1257
timestamp 1649977179
transform 1 0 116748 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1269
timestamp 1649977179
transform 1 0 117852 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1281
timestamp 1649977179
transform 1 0 118956 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1287
timestamp 1649977179
transform 1 0 119508 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1289
timestamp 1649977179
transform 1 0 119692 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1301
timestamp 1649977179
transform 1 0 120796 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1313
timestamp 1649977179
transform 1 0 121900 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1325
timestamp 1649977179
transform 1 0 123004 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1337
timestamp 1649977179
transform 1 0 124108 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1343
timestamp 1649977179
transform 1 0 124660 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1345
timestamp 1649977179
transform 1 0 124844 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1357
timestamp 1649977179
transform 1 0 125948 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1369
timestamp 1649977179
transform 1 0 127052 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1381
timestamp 1649977179
transform 1 0 128156 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1393
timestamp 1649977179
transform 1 0 129260 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1399
timestamp 1649977179
transform 1 0 129812 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1401
timestamp 1649977179
transform 1 0 129996 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1413
timestamp 1649977179
transform 1 0 131100 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1425
timestamp 1649977179
transform 1 0 132204 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1437
timestamp 1649977179
transform 1 0 133308 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1449
timestamp 1649977179
transform 1 0 134412 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1455
timestamp 1649977179
transform 1 0 134964 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1457
timestamp 1649977179
transform 1 0 135148 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1469
timestamp 1649977179
transform 1 0 136252 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1481
timestamp 1649977179
transform 1 0 137356 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1493
timestamp 1649977179
transform 1 0 138460 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1505
timestamp 1649977179
transform 1 0 139564 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1511
timestamp 1649977179
transform 1 0 140116 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1513
timestamp 1649977179
transform 1 0 140300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1525
timestamp 1649977179
transform 1 0 141404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1537
timestamp 1649977179
transform 1 0 142508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1549
timestamp 1649977179
transform 1 0 143612 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1561
timestamp 1649977179
transform 1 0 144716 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1567
timestamp 1649977179
transform 1 0 145268 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1569
timestamp 1649977179
transform 1 0 145452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1581
timestamp 1649977179
transform 1 0 146556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1593
timestamp 1649977179
transform 1 0 147660 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1605
timestamp 1649977179
transform 1 0 148764 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1617
timestamp 1649977179
transform 1 0 149868 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1623
timestamp 1649977179
transform 1 0 150420 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1625
timestamp 1649977179
transform 1 0 150604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1637
timestamp 1649977179
transform 1 0 151708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1649
timestamp 1649977179
transform 1 0 152812 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1661
timestamp 1649977179
transform 1 0 153916 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1673
timestamp 1649977179
transform 1 0 155020 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1679
timestamp 1649977179
transform 1 0 155572 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1681
timestamp 1649977179
transform 1 0 155756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1693
timestamp 1649977179
transform 1 0 156860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1705
timestamp 1649977179
transform 1 0 157964 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1717
timestamp 1649977179
transform 1 0 159068 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1729
timestamp 1649977179
transform 1 0 160172 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1735
timestamp 1649977179
transform 1 0 160724 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1737
timestamp 1649977179
transform 1 0 160908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1749
timestamp 1649977179
transform 1 0 162012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1761
timestamp 1649977179
transform 1 0 163116 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1773
timestamp 1649977179
transform 1 0 164220 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1785
timestamp 1649977179
transform 1 0 165324 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1791
timestamp 1649977179
transform 1 0 165876 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1793
timestamp 1649977179
transform 1 0 166060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1805
timestamp 1649977179
transform 1 0 167164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1817
timestamp 1649977179
transform 1 0 168268 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1829
timestamp 1649977179
transform 1 0 169372 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1841
timestamp 1649977179
transform 1 0 170476 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1847
timestamp 1649977179
transform 1 0 171028 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1849
timestamp 1649977179
transform 1 0 171212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1861
timestamp 1649977179
transform 1 0 172316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1873
timestamp 1649977179
transform 1 0 173420 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1885
timestamp 1649977179
transform 1 0 174524 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1897
timestamp 1649977179
transform 1 0 175628 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1903
timestamp 1649977179
transform 1 0 176180 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1905
timestamp 1649977179
transform 1 0 176364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1917
timestamp 1649977179
transform 1 0 177468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1929
timestamp 1649977179
transform 1 0 178572 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1941
timestamp 1649977179
transform 1 0 179676 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1953
timestamp 1649977179
transform 1 0 180780 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1959
timestamp 1649977179
transform 1 0 181332 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1961
timestamp 1649977179
transform 1 0 181516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1973
timestamp 1649977179
transform 1 0 182620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1985
timestamp 1649977179
transform 1 0 183724 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1997
timestamp 1649977179
transform 1 0 184828 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2009
timestamp 1649977179
transform 1 0 185932 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2015
timestamp 1649977179
transform 1 0 186484 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2017
timestamp 1649977179
transform 1 0 186668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2029
timestamp 1649977179
transform 1 0 187772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2041
timestamp 1649977179
transform 1 0 188876 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2053
timestamp 1649977179
transform 1 0 189980 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2065
timestamp 1649977179
transform 1 0 191084 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2071
timestamp 1649977179
transform 1 0 191636 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2073
timestamp 1649977179
transform 1 0 191820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2085
timestamp 1649977179
transform 1 0 192924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2097
timestamp 1649977179
transform 1 0 194028 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2109
timestamp 1649977179
transform 1 0 195132 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2121
timestamp 1649977179
transform 1 0 196236 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2127
timestamp 1649977179
transform 1 0 196788 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2129
timestamp 1649977179
transform 1 0 196972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2141
timestamp 1649977179
transform 1 0 198076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2153
timestamp 1649977179
transform 1 0 199180 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2165
timestamp 1649977179
transform 1 0 200284 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2177
timestamp 1649977179
transform 1 0 201388 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2183
timestamp 1649977179
transform 1 0 201940 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2185
timestamp 1649977179
transform 1 0 202124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2197
timestamp 1649977179
transform 1 0 203228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2209
timestamp 1649977179
transform 1 0 204332 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2221
timestamp 1649977179
transform 1 0 205436 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2233
timestamp 1649977179
transform 1 0 206540 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2239
timestamp 1649977179
transform 1 0 207092 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2241
timestamp 1649977179
transform 1 0 207276 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2253
timestamp 1649977179
transform 1 0 208380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2265
timestamp 1649977179
transform 1 0 209484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2277
timestamp 1649977179
transform 1 0 210588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2289
timestamp 1649977179
transform 1 0 211692 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2295
timestamp 1649977179
transform 1 0 212244 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2297
timestamp 1649977179
transform 1 0 212428 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2309
timestamp 1649977179
transform 1 0 213532 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2321
timestamp 1649977179
transform 1 0 214636 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2333
timestamp 1649977179
transform 1 0 215740 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2345
timestamp 1649977179
transform 1 0 216844 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2351
timestamp 1649977179
transform 1 0 217396 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2353
timestamp 1649977179
transform 1 0 217580 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2365
timestamp 1649977179
transform 1 0 218684 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2377
timestamp 1649977179
transform 1 0 219788 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2389
timestamp 1649977179
transform 1 0 220892 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2401
timestamp 1649977179
transform 1 0 221996 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2407
timestamp 1649977179
transform 1 0 222548 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2409
timestamp 1649977179
transform 1 0 222732 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2421
timestamp 1649977179
transform 1 0 223836 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2433
timestamp 1649977179
transform 1 0 224940 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2445
timestamp 1649977179
transform 1 0 226044 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2457
timestamp 1649977179
transform 1 0 227148 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2463
timestamp 1649977179
transform 1 0 227700 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2465
timestamp 1649977179
transform 1 0 227884 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2477
timestamp 1649977179
transform 1 0 228988 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2489
timestamp 1649977179
transform 1 0 230092 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2501
timestamp 1649977179
transform 1 0 231196 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2513
timestamp 1649977179
transform 1 0 232300 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2519
timestamp 1649977179
transform 1 0 232852 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2521
timestamp 1649977179
transform 1 0 233036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2533
timestamp 1649977179
transform 1 0 234140 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2545
timestamp 1649977179
transform 1 0 235244 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2557
timestamp 1649977179
transform 1 0 236348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2569
timestamp 1649977179
transform 1 0 237452 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2575
timestamp 1649977179
transform 1 0 238004 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2577
timestamp 1649977179
transform 1 0 238188 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2589
timestamp 1649977179
transform 1 0 239292 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2601
timestamp 1649977179
transform 1 0 240396 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2613
timestamp 1649977179
transform 1 0 241500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2625
timestamp 1649977179
transform 1 0 242604 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2631
timestamp 1649977179
transform 1 0 243156 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2633
timestamp 1649977179
transform 1 0 243340 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2645
timestamp 1649977179
transform 1 0 244444 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2657
timestamp 1649977179
transform 1 0 245548 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2669
timestamp 1649977179
transform 1 0 246652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2681
timestamp 1649977179
transform 1 0 247756 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2687
timestamp 1649977179
transform 1 0 248308 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2689
timestamp 1649977179
transform 1 0 248492 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2701
timestamp 1649977179
transform 1 0 249596 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2713
timestamp 1649977179
transform 1 0 250700 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2725
timestamp 1649977179
transform 1 0 251804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2737
timestamp 1649977179
transform 1 0 252908 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2743
timestamp 1649977179
transform 1 0 253460 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2745
timestamp 1649977179
transform 1 0 253644 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2757
timestamp 1649977179
transform 1 0 254748 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2769
timestamp 1649977179
transform 1 0 255852 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2781
timestamp 1649977179
transform 1 0 256956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2793
timestamp 1649977179
transform 1 0 258060 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2799
timestamp 1649977179
transform 1 0 258612 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2801
timestamp 1649977179
transform 1 0 258796 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2813
timestamp 1649977179
transform 1 0 259900 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2825
timestamp 1649977179
transform 1 0 261004 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2837
timestamp 1649977179
transform 1 0 262108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2849
timestamp 1649977179
transform 1 0 263212 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2855
timestamp 1649977179
transform 1 0 263764 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2857
timestamp 1649977179
transform 1 0 263948 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2869
timestamp 1649977179
transform 1 0 265052 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2881
timestamp 1649977179
transform 1 0 266156 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2893
timestamp 1649977179
transform 1 0 267260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2905
timestamp 1649977179
transform 1 0 268364 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2911
timestamp 1649977179
transform 1 0 268916 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2913
timestamp 1649977179
transform 1 0 269100 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2925
timestamp 1649977179
transform 1 0 270204 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2937
timestamp 1649977179
transform 1 0 271308 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2949
timestamp 1649977179
transform 1 0 272412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2961
timestamp 1649977179
transform 1 0 273516 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2967
timestamp 1649977179
transform 1 0 274068 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2969
timestamp 1649977179
transform 1 0 274252 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2981
timestamp 1649977179
transform 1 0 275356 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2993
timestamp 1649977179
transform 1 0 276460 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3005
timestamp 1649977179
transform 1 0 277564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3017
timestamp 1649977179
transform 1 0 278668 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3023
timestamp 1649977179
transform 1 0 279220 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3025
timestamp 1649977179
transform 1 0 279404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3037
timestamp 1649977179
transform 1 0 280508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3049
timestamp 1649977179
transform 1 0 281612 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3061
timestamp 1649977179
transform 1 0 282716 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3073
timestamp 1649977179
transform 1 0 283820 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3079
timestamp 1649977179
transform 1 0 284372 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3081
timestamp 1649977179
transform 1 0 284556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3093
timestamp 1649977179
transform 1 0 285660 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3105
timestamp 1649977179
transform 1 0 286764 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3117
timestamp 1649977179
transform 1 0 287868 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3129
timestamp 1649977179
transform 1 0 288972 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3135
timestamp 1649977179
transform 1 0 289524 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3137
timestamp 1649977179
transform 1 0 289708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3149
timestamp 1649977179
transform 1 0 290812 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3161
timestamp 1649977179
transform 1 0 291916 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3173
timestamp 1649977179
transform 1 0 293020 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3185
timestamp 1649977179
transform 1 0 294124 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3191
timestamp 1649977179
transform 1 0 294676 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3193
timestamp 1649977179
transform 1 0 294860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3205
timestamp 1649977179
transform 1 0 295964 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3217
timestamp 1649977179
transform 1 0 297068 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3229
timestamp 1649977179
transform 1 0 298172 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3241
timestamp 1649977179
transform 1 0 299276 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3247
timestamp 1649977179
transform 1 0 299828 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3249
timestamp 1649977179
transform 1 0 300012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3261
timestamp 1649977179
transform 1 0 301116 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3273
timestamp 1649977179
transform 1 0 302220 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3285
timestamp 1649977179
transform 1 0 303324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3297
timestamp 1649977179
transform 1 0 304428 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3303
timestamp 1649977179
transform 1 0 304980 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3305
timestamp 1649977179
transform 1 0 305164 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1649977179
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1649977179
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1649977179
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1649977179
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1649977179
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1649977179
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1649977179
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1649977179
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1649977179
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1649977179
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1649977179
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1649977179
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1649977179
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1649977179
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1649977179
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1649977179
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1649977179
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1649977179
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1649977179
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1649977179
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1649977179
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1649977179
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1649977179
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1649977179
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1649977179
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1649977179
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1649977179
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1649977179
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1649977179
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1649977179
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1649977179
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1649977179
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1649977179
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1649977179
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1649977179
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1649977179
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1649977179
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1649977179
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1649977179
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1649977179
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1649977179
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1649977179
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_601
timestamp 1649977179
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_613
timestamp 1649977179
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_625
timestamp 1649977179
transform 1 0 58604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_637
timestamp 1649977179
transform 1 0 59708 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_643
timestamp 1649977179
transform 1 0 60260 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_645
timestamp 1649977179
transform 1 0 60444 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_657
timestamp 1649977179
transform 1 0 61548 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_669
timestamp 1649977179
transform 1 0 62652 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_681
timestamp 1649977179
transform 1 0 63756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_693
timestamp 1649977179
transform 1 0 64860 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_699
timestamp 1649977179
transform 1 0 65412 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_701
timestamp 1649977179
transform 1 0 65596 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_713
timestamp 1649977179
transform 1 0 66700 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_725
timestamp 1649977179
transform 1 0 67804 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_737
timestamp 1649977179
transform 1 0 68908 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_749
timestamp 1649977179
transform 1 0 70012 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_755
timestamp 1649977179
transform 1 0 70564 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_757
timestamp 1649977179
transform 1 0 70748 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_769
timestamp 1649977179
transform 1 0 71852 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_781
timestamp 1649977179
transform 1 0 72956 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_793
timestamp 1649977179
transform 1 0 74060 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_805
timestamp 1649977179
transform 1 0 75164 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_811
timestamp 1649977179
transform 1 0 75716 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_813
timestamp 1649977179
transform 1 0 75900 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_825
timestamp 1649977179
transform 1 0 77004 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_837
timestamp 1649977179
transform 1 0 78108 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_849
timestamp 1649977179
transform 1 0 79212 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_861
timestamp 1649977179
transform 1 0 80316 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_867
timestamp 1649977179
transform 1 0 80868 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_869
timestamp 1649977179
transform 1 0 81052 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_881
timestamp 1649977179
transform 1 0 82156 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_893
timestamp 1649977179
transform 1 0 83260 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_905
timestamp 1649977179
transform 1 0 84364 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_917
timestamp 1649977179
transform 1 0 85468 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_923
timestamp 1649977179
transform 1 0 86020 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_925
timestamp 1649977179
transform 1 0 86204 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_937
timestamp 1649977179
transform 1 0 87308 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_949
timestamp 1649977179
transform 1 0 88412 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_961
timestamp 1649977179
transform 1 0 89516 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_973
timestamp 1649977179
transform 1 0 90620 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_979
timestamp 1649977179
transform 1 0 91172 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_981
timestamp 1649977179
transform 1 0 91356 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_993
timestamp 1649977179
transform 1 0 92460 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1005
timestamp 1649977179
transform 1 0 93564 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1017
timestamp 1649977179
transform 1 0 94668 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1029
timestamp 1649977179
transform 1 0 95772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1035
timestamp 1649977179
transform 1 0 96324 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1037
timestamp 1649977179
transform 1 0 96508 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1049
timestamp 1649977179
transform 1 0 97612 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1061
timestamp 1649977179
transform 1 0 98716 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1073
timestamp 1649977179
transform 1 0 99820 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1085
timestamp 1649977179
transform 1 0 100924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1091
timestamp 1649977179
transform 1 0 101476 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1093
timestamp 1649977179
transform 1 0 101660 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1105
timestamp 1649977179
transform 1 0 102764 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1117
timestamp 1649977179
transform 1 0 103868 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1129
timestamp 1649977179
transform 1 0 104972 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1141
timestamp 1649977179
transform 1 0 106076 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1147
timestamp 1649977179
transform 1 0 106628 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1149
timestamp 1649977179
transform 1 0 106812 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1161
timestamp 1649977179
transform 1 0 107916 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1173
timestamp 1649977179
transform 1 0 109020 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1185
timestamp 1649977179
transform 1 0 110124 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1197
timestamp 1649977179
transform 1 0 111228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1203
timestamp 1649977179
transform 1 0 111780 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1205
timestamp 1649977179
transform 1 0 111964 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1217
timestamp 1649977179
transform 1 0 113068 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1229
timestamp 1649977179
transform 1 0 114172 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1241
timestamp 1649977179
transform 1 0 115276 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1253
timestamp 1649977179
transform 1 0 116380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1259
timestamp 1649977179
transform 1 0 116932 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1261
timestamp 1649977179
transform 1 0 117116 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1273
timestamp 1649977179
transform 1 0 118220 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1285
timestamp 1649977179
transform 1 0 119324 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1297
timestamp 1649977179
transform 1 0 120428 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1309
timestamp 1649977179
transform 1 0 121532 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1315
timestamp 1649977179
transform 1 0 122084 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1317
timestamp 1649977179
transform 1 0 122268 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1329
timestamp 1649977179
transform 1 0 123372 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1341
timestamp 1649977179
transform 1 0 124476 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1353
timestamp 1649977179
transform 1 0 125580 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1365
timestamp 1649977179
transform 1 0 126684 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1371
timestamp 1649977179
transform 1 0 127236 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1373
timestamp 1649977179
transform 1 0 127420 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1385
timestamp 1649977179
transform 1 0 128524 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1397
timestamp 1649977179
transform 1 0 129628 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1409
timestamp 1649977179
transform 1 0 130732 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1421
timestamp 1649977179
transform 1 0 131836 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1427
timestamp 1649977179
transform 1 0 132388 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1429
timestamp 1649977179
transform 1 0 132572 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1441
timestamp 1649977179
transform 1 0 133676 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1453
timestamp 1649977179
transform 1 0 134780 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1465
timestamp 1649977179
transform 1 0 135884 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1477
timestamp 1649977179
transform 1 0 136988 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1483
timestamp 1649977179
transform 1 0 137540 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1485
timestamp 1649977179
transform 1 0 137724 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1497
timestamp 1649977179
transform 1 0 138828 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1509
timestamp 1649977179
transform 1 0 139932 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1521
timestamp 1649977179
transform 1 0 141036 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1533
timestamp 1649977179
transform 1 0 142140 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1539
timestamp 1649977179
transform 1 0 142692 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1541
timestamp 1649977179
transform 1 0 142876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1553
timestamp 1649977179
transform 1 0 143980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1565
timestamp 1649977179
transform 1 0 145084 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1577
timestamp 1649977179
transform 1 0 146188 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1589
timestamp 1649977179
transform 1 0 147292 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1595
timestamp 1649977179
transform 1 0 147844 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1597
timestamp 1649977179
transform 1 0 148028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1609
timestamp 1649977179
transform 1 0 149132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1621
timestamp 1649977179
transform 1 0 150236 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1633
timestamp 1649977179
transform 1 0 151340 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1645
timestamp 1649977179
transform 1 0 152444 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1651
timestamp 1649977179
transform 1 0 152996 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1653
timestamp 1649977179
transform 1 0 153180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1665
timestamp 1649977179
transform 1 0 154284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1677
timestamp 1649977179
transform 1 0 155388 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1689
timestamp 1649977179
transform 1 0 156492 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1701
timestamp 1649977179
transform 1 0 157596 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1707
timestamp 1649977179
transform 1 0 158148 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1709
timestamp 1649977179
transform 1 0 158332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1721
timestamp 1649977179
transform 1 0 159436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1733
timestamp 1649977179
transform 1 0 160540 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1745
timestamp 1649977179
transform 1 0 161644 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1757
timestamp 1649977179
transform 1 0 162748 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1763
timestamp 1649977179
transform 1 0 163300 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1765
timestamp 1649977179
transform 1 0 163484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1777
timestamp 1649977179
transform 1 0 164588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1789
timestamp 1649977179
transform 1 0 165692 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1801
timestamp 1649977179
transform 1 0 166796 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1813
timestamp 1649977179
transform 1 0 167900 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1819
timestamp 1649977179
transform 1 0 168452 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1821
timestamp 1649977179
transform 1 0 168636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1833
timestamp 1649977179
transform 1 0 169740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1845
timestamp 1649977179
transform 1 0 170844 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1857
timestamp 1649977179
transform 1 0 171948 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1869
timestamp 1649977179
transform 1 0 173052 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1875
timestamp 1649977179
transform 1 0 173604 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1877
timestamp 1649977179
transform 1 0 173788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1889
timestamp 1649977179
transform 1 0 174892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1901
timestamp 1649977179
transform 1 0 175996 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1913
timestamp 1649977179
transform 1 0 177100 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1925
timestamp 1649977179
transform 1 0 178204 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1931
timestamp 1649977179
transform 1 0 178756 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1933
timestamp 1649977179
transform 1 0 178940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1945
timestamp 1649977179
transform 1 0 180044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1957
timestamp 1649977179
transform 1 0 181148 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1969
timestamp 1649977179
transform 1 0 182252 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1981
timestamp 1649977179
transform 1 0 183356 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1987
timestamp 1649977179
transform 1 0 183908 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1989
timestamp 1649977179
transform 1 0 184092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2001
timestamp 1649977179
transform 1 0 185196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2013
timestamp 1649977179
transform 1 0 186300 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2025
timestamp 1649977179
transform 1 0 187404 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2037
timestamp 1649977179
transform 1 0 188508 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2043
timestamp 1649977179
transform 1 0 189060 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2045
timestamp 1649977179
transform 1 0 189244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2057
timestamp 1649977179
transform 1 0 190348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2069
timestamp 1649977179
transform 1 0 191452 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2081
timestamp 1649977179
transform 1 0 192556 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2093
timestamp 1649977179
transform 1 0 193660 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2099
timestamp 1649977179
transform 1 0 194212 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2101
timestamp 1649977179
transform 1 0 194396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2113
timestamp 1649977179
transform 1 0 195500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2125
timestamp 1649977179
transform 1 0 196604 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2137
timestamp 1649977179
transform 1 0 197708 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2149
timestamp 1649977179
transform 1 0 198812 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2155
timestamp 1649977179
transform 1 0 199364 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2157
timestamp 1649977179
transform 1 0 199548 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2169
timestamp 1649977179
transform 1 0 200652 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2181
timestamp 1649977179
transform 1 0 201756 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2193
timestamp 1649977179
transform 1 0 202860 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2205
timestamp 1649977179
transform 1 0 203964 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2211
timestamp 1649977179
transform 1 0 204516 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2213
timestamp 1649977179
transform 1 0 204700 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2225
timestamp 1649977179
transform 1 0 205804 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2237
timestamp 1649977179
transform 1 0 206908 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2249
timestamp 1649977179
transform 1 0 208012 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2261
timestamp 1649977179
transform 1 0 209116 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2267
timestamp 1649977179
transform 1 0 209668 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2269
timestamp 1649977179
transform 1 0 209852 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2281
timestamp 1649977179
transform 1 0 210956 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2293
timestamp 1649977179
transform 1 0 212060 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2305
timestamp 1649977179
transform 1 0 213164 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2317
timestamp 1649977179
transform 1 0 214268 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2323
timestamp 1649977179
transform 1 0 214820 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2325
timestamp 1649977179
transform 1 0 215004 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2337
timestamp 1649977179
transform 1 0 216108 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2349
timestamp 1649977179
transform 1 0 217212 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2361
timestamp 1649977179
transform 1 0 218316 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2373
timestamp 1649977179
transform 1 0 219420 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2379
timestamp 1649977179
transform 1 0 219972 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2381
timestamp 1649977179
transform 1 0 220156 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2393
timestamp 1649977179
transform 1 0 221260 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2405
timestamp 1649977179
transform 1 0 222364 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2417
timestamp 1649977179
transform 1 0 223468 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2429
timestamp 1649977179
transform 1 0 224572 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2435
timestamp 1649977179
transform 1 0 225124 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2437
timestamp 1649977179
transform 1 0 225308 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2449
timestamp 1649977179
transform 1 0 226412 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2461
timestamp 1649977179
transform 1 0 227516 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2473
timestamp 1649977179
transform 1 0 228620 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2485
timestamp 1649977179
transform 1 0 229724 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2491
timestamp 1649977179
transform 1 0 230276 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2493
timestamp 1649977179
transform 1 0 230460 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2505
timestamp 1649977179
transform 1 0 231564 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2517
timestamp 1649977179
transform 1 0 232668 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2529
timestamp 1649977179
transform 1 0 233772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2541
timestamp 1649977179
transform 1 0 234876 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2547
timestamp 1649977179
transform 1 0 235428 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2549
timestamp 1649977179
transform 1 0 235612 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2561
timestamp 1649977179
transform 1 0 236716 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2573
timestamp 1649977179
transform 1 0 237820 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2585
timestamp 1649977179
transform 1 0 238924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2597
timestamp 1649977179
transform 1 0 240028 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2603
timestamp 1649977179
transform 1 0 240580 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2605
timestamp 1649977179
transform 1 0 240764 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2617
timestamp 1649977179
transform 1 0 241868 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2629
timestamp 1649977179
transform 1 0 242972 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2641
timestamp 1649977179
transform 1 0 244076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2653
timestamp 1649977179
transform 1 0 245180 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2659
timestamp 1649977179
transform 1 0 245732 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2661
timestamp 1649977179
transform 1 0 245916 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2673
timestamp 1649977179
transform 1 0 247020 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2685
timestamp 1649977179
transform 1 0 248124 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2697
timestamp 1649977179
transform 1 0 249228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2709
timestamp 1649977179
transform 1 0 250332 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2715
timestamp 1649977179
transform 1 0 250884 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2717
timestamp 1649977179
transform 1 0 251068 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2729
timestamp 1649977179
transform 1 0 252172 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2741
timestamp 1649977179
transform 1 0 253276 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2753
timestamp 1649977179
transform 1 0 254380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2765
timestamp 1649977179
transform 1 0 255484 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2771
timestamp 1649977179
transform 1 0 256036 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2773
timestamp 1649977179
transform 1 0 256220 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2785
timestamp 1649977179
transform 1 0 257324 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2797
timestamp 1649977179
transform 1 0 258428 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2809
timestamp 1649977179
transform 1 0 259532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2821
timestamp 1649977179
transform 1 0 260636 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2827
timestamp 1649977179
transform 1 0 261188 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2829
timestamp 1649977179
transform 1 0 261372 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2841
timestamp 1649977179
transform 1 0 262476 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2853
timestamp 1649977179
transform 1 0 263580 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2865
timestamp 1649977179
transform 1 0 264684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2877
timestamp 1649977179
transform 1 0 265788 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2883
timestamp 1649977179
transform 1 0 266340 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2885
timestamp 1649977179
transform 1 0 266524 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2897
timestamp 1649977179
transform 1 0 267628 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2909
timestamp 1649977179
transform 1 0 268732 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2921
timestamp 1649977179
transform 1 0 269836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2933
timestamp 1649977179
transform 1 0 270940 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2939
timestamp 1649977179
transform 1 0 271492 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2941
timestamp 1649977179
transform 1 0 271676 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2953
timestamp 1649977179
transform 1 0 272780 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2965
timestamp 1649977179
transform 1 0 273884 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2977
timestamp 1649977179
transform 1 0 274988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2989
timestamp 1649977179
transform 1 0 276092 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2995
timestamp 1649977179
transform 1 0 276644 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2997
timestamp 1649977179
transform 1 0 276828 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3009
timestamp 1649977179
transform 1 0 277932 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3021
timestamp 1649977179
transform 1 0 279036 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3033
timestamp 1649977179
transform 1 0 280140 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3045
timestamp 1649977179
transform 1 0 281244 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3051
timestamp 1649977179
transform 1 0 281796 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3053
timestamp 1649977179
transform 1 0 281980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3065
timestamp 1649977179
transform 1 0 283084 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3077
timestamp 1649977179
transform 1 0 284188 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3089
timestamp 1649977179
transform 1 0 285292 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3101
timestamp 1649977179
transform 1 0 286396 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3107
timestamp 1649977179
transform 1 0 286948 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3109
timestamp 1649977179
transform 1 0 287132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3121
timestamp 1649977179
transform 1 0 288236 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3133
timestamp 1649977179
transform 1 0 289340 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3145
timestamp 1649977179
transform 1 0 290444 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3157
timestamp 1649977179
transform 1 0 291548 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3163
timestamp 1649977179
transform 1 0 292100 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3165
timestamp 1649977179
transform 1 0 292284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3177
timestamp 1649977179
transform 1 0 293388 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3189
timestamp 1649977179
transform 1 0 294492 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3201
timestamp 1649977179
transform 1 0 295596 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3213
timestamp 1649977179
transform 1 0 296700 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3219
timestamp 1649977179
transform 1 0 297252 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3221
timestamp 1649977179
transform 1 0 297436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3233
timestamp 1649977179
transform 1 0 298540 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3245
timestamp 1649977179
transform 1 0 299644 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3257
timestamp 1649977179
transform 1 0 300748 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3269
timestamp 1649977179
transform 1 0 301852 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3275
timestamp 1649977179
transform 1 0 302404 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3277
timestamp 1649977179
transform 1 0 302588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3289
timestamp 1649977179
transform 1 0 303692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3301
timestamp 1649977179
transform 1 0 304796 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1656 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_10
timestamp 1649977179
transform 1 0 2024 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_14
timestamp 1649977179
transform 1 0 2392 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_18
timestamp 1649977179
transform 1 0 2760 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_22
timestamp 1649977179
transform 1 0 3128 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_34
timestamp 1649977179
transform 1 0 4232 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_46
timestamp 1649977179
transform 1 0 5336 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1649977179
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1649977179
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1649977179
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1649977179
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1649977179
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1649977179
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1649977179
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1649977179
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1649977179
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1649977179
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1649977179
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1649977179
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1649977179
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1649977179
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1649977179
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1649977179
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1649977179
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1649977179
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1649977179
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1649977179
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1649977179
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1649977179
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1649977179
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1649977179
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1649977179
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1649977179
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1649977179
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1649977179
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1649977179
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1649977179
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1649977179
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1649977179
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1649977179
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1649977179
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1649977179
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1649977179
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1649977179
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1649977179
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1649977179
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1649977179
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1649977179
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1649977179
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1649977179
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1649977179
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_597
timestamp 1649977179
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1649977179
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1649977179
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_617
timestamp 1649977179
transform 1 0 57868 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_629
timestamp 1649977179
transform 1 0 58972 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_641
timestamp 1649977179
transform 1 0 60076 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_653
timestamp 1649977179
transform 1 0 61180 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_665
timestamp 1649977179
transform 1 0 62284 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_671
timestamp 1649977179
transform 1 0 62836 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_673
timestamp 1649977179
transform 1 0 63020 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_685
timestamp 1649977179
transform 1 0 64124 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_697
timestamp 1649977179
transform 1 0 65228 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_709
timestamp 1649977179
transform 1 0 66332 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_721
timestamp 1649977179
transform 1 0 67436 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_727
timestamp 1649977179
transform 1 0 67988 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_729
timestamp 1649977179
transform 1 0 68172 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_741
timestamp 1649977179
transform 1 0 69276 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_753
timestamp 1649977179
transform 1 0 70380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_765
timestamp 1649977179
transform 1 0 71484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_777
timestamp 1649977179
transform 1 0 72588 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_783
timestamp 1649977179
transform 1 0 73140 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_785
timestamp 1649977179
transform 1 0 73324 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_797
timestamp 1649977179
transform 1 0 74428 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_809
timestamp 1649977179
transform 1 0 75532 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_821
timestamp 1649977179
transform 1 0 76636 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_833
timestamp 1649977179
transform 1 0 77740 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_839
timestamp 1649977179
transform 1 0 78292 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_841
timestamp 1649977179
transform 1 0 78476 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_853
timestamp 1649977179
transform 1 0 79580 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_865
timestamp 1649977179
transform 1 0 80684 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_877
timestamp 1649977179
transform 1 0 81788 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_889
timestamp 1649977179
transform 1 0 82892 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_895
timestamp 1649977179
transform 1 0 83444 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_897
timestamp 1649977179
transform 1 0 83628 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_909
timestamp 1649977179
transform 1 0 84732 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_921
timestamp 1649977179
transform 1 0 85836 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_933
timestamp 1649977179
transform 1 0 86940 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_945
timestamp 1649977179
transform 1 0 88044 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_951
timestamp 1649977179
transform 1 0 88596 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_953
timestamp 1649977179
transform 1 0 88780 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_965
timestamp 1649977179
transform 1 0 89884 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_977
timestamp 1649977179
transform 1 0 90988 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_989
timestamp 1649977179
transform 1 0 92092 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1001
timestamp 1649977179
transform 1 0 93196 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1007
timestamp 1649977179
transform 1 0 93748 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1009
timestamp 1649977179
transform 1 0 93932 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1021
timestamp 1649977179
transform 1 0 95036 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1033
timestamp 1649977179
transform 1 0 96140 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1045
timestamp 1649977179
transform 1 0 97244 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1057
timestamp 1649977179
transform 1 0 98348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1063
timestamp 1649977179
transform 1 0 98900 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1065
timestamp 1649977179
transform 1 0 99084 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1077
timestamp 1649977179
transform 1 0 100188 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1089
timestamp 1649977179
transform 1 0 101292 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1101
timestamp 1649977179
transform 1 0 102396 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1113
timestamp 1649977179
transform 1 0 103500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1119
timestamp 1649977179
transform 1 0 104052 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1121
timestamp 1649977179
transform 1 0 104236 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1133
timestamp 1649977179
transform 1 0 105340 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1145
timestamp 1649977179
transform 1 0 106444 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1157
timestamp 1649977179
transform 1 0 107548 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1169
timestamp 1649977179
transform 1 0 108652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1175
timestamp 1649977179
transform 1 0 109204 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1177
timestamp 1649977179
transform 1 0 109388 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1189
timestamp 1649977179
transform 1 0 110492 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1201
timestamp 1649977179
transform 1 0 111596 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1213
timestamp 1649977179
transform 1 0 112700 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1225
timestamp 1649977179
transform 1 0 113804 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1231
timestamp 1649977179
transform 1 0 114356 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1233
timestamp 1649977179
transform 1 0 114540 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1245
timestamp 1649977179
transform 1 0 115644 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1257
timestamp 1649977179
transform 1 0 116748 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1269
timestamp 1649977179
transform 1 0 117852 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1281
timestamp 1649977179
transform 1 0 118956 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1287
timestamp 1649977179
transform 1 0 119508 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1289
timestamp 1649977179
transform 1 0 119692 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1301
timestamp 1649977179
transform 1 0 120796 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1313
timestamp 1649977179
transform 1 0 121900 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1325
timestamp 1649977179
transform 1 0 123004 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1337
timestamp 1649977179
transform 1 0 124108 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1343
timestamp 1649977179
transform 1 0 124660 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1345
timestamp 1649977179
transform 1 0 124844 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1357
timestamp 1649977179
transform 1 0 125948 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1369
timestamp 1649977179
transform 1 0 127052 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1381
timestamp 1649977179
transform 1 0 128156 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1393
timestamp 1649977179
transform 1 0 129260 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1399
timestamp 1649977179
transform 1 0 129812 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1401
timestamp 1649977179
transform 1 0 129996 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1413
timestamp 1649977179
transform 1 0 131100 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1425
timestamp 1649977179
transform 1 0 132204 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1437
timestamp 1649977179
transform 1 0 133308 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1449
timestamp 1649977179
transform 1 0 134412 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1455
timestamp 1649977179
transform 1 0 134964 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1457
timestamp 1649977179
transform 1 0 135148 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1469
timestamp 1649977179
transform 1 0 136252 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1481
timestamp 1649977179
transform 1 0 137356 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1493
timestamp 1649977179
transform 1 0 138460 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1505
timestamp 1649977179
transform 1 0 139564 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1511
timestamp 1649977179
transform 1 0 140116 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1513
timestamp 1649977179
transform 1 0 140300 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1525
timestamp 1649977179
transform 1 0 141404 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1537
timestamp 1649977179
transform 1 0 142508 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1549
timestamp 1649977179
transform 1 0 143612 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1561
timestamp 1649977179
transform 1 0 144716 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1567
timestamp 1649977179
transform 1 0 145268 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1569
timestamp 1649977179
transform 1 0 145452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1581
timestamp 1649977179
transform 1 0 146556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1593
timestamp 1649977179
transform 1 0 147660 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1605
timestamp 1649977179
transform 1 0 148764 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1617
timestamp 1649977179
transform 1 0 149868 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1623
timestamp 1649977179
transform 1 0 150420 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1625
timestamp 1649977179
transform 1 0 150604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1637
timestamp 1649977179
transform 1 0 151708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1649
timestamp 1649977179
transform 1 0 152812 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1661
timestamp 1649977179
transform 1 0 153916 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1673
timestamp 1649977179
transform 1 0 155020 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1679
timestamp 1649977179
transform 1 0 155572 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1681
timestamp 1649977179
transform 1 0 155756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1693
timestamp 1649977179
transform 1 0 156860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1705
timestamp 1649977179
transform 1 0 157964 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1717
timestamp 1649977179
transform 1 0 159068 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1729
timestamp 1649977179
transform 1 0 160172 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1735
timestamp 1649977179
transform 1 0 160724 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1737
timestamp 1649977179
transform 1 0 160908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1749
timestamp 1649977179
transform 1 0 162012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1761
timestamp 1649977179
transform 1 0 163116 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1773
timestamp 1649977179
transform 1 0 164220 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1785
timestamp 1649977179
transform 1 0 165324 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1791
timestamp 1649977179
transform 1 0 165876 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1793
timestamp 1649977179
transform 1 0 166060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1805
timestamp 1649977179
transform 1 0 167164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1817
timestamp 1649977179
transform 1 0 168268 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1829
timestamp 1649977179
transform 1 0 169372 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1841
timestamp 1649977179
transform 1 0 170476 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1847
timestamp 1649977179
transform 1 0 171028 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1849
timestamp 1649977179
transform 1 0 171212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1861
timestamp 1649977179
transform 1 0 172316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1873
timestamp 1649977179
transform 1 0 173420 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1885
timestamp 1649977179
transform 1 0 174524 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1897
timestamp 1649977179
transform 1 0 175628 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1903
timestamp 1649977179
transform 1 0 176180 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1905
timestamp 1649977179
transform 1 0 176364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1917
timestamp 1649977179
transform 1 0 177468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1929
timestamp 1649977179
transform 1 0 178572 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1941
timestamp 1649977179
transform 1 0 179676 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1953
timestamp 1649977179
transform 1 0 180780 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1959
timestamp 1649977179
transform 1 0 181332 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1961
timestamp 1649977179
transform 1 0 181516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1973
timestamp 1649977179
transform 1 0 182620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1985
timestamp 1649977179
transform 1 0 183724 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1997
timestamp 1649977179
transform 1 0 184828 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2009
timestamp 1649977179
transform 1 0 185932 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2015
timestamp 1649977179
transform 1 0 186484 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2017
timestamp 1649977179
transform 1 0 186668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2029
timestamp 1649977179
transform 1 0 187772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2041
timestamp 1649977179
transform 1 0 188876 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2053
timestamp 1649977179
transform 1 0 189980 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2065
timestamp 1649977179
transform 1 0 191084 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2071
timestamp 1649977179
transform 1 0 191636 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2073
timestamp 1649977179
transform 1 0 191820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2085
timestamp 1649977179
transform 1 0 192924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2097
timestamp 1649977179
transform 1 0 194028 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2109
timestamp 1649977179
transform 1 0 195132 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2121
timestamp 1649977179
transform 1 0 196236 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2127
timestamp 1649977179
transform 1 0 196788 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2129
timestamp 1649977179
transform 1 0 196972 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2141
timestamp 1649977179
transform 1 0 198076 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2153
timestamp 1649977179
transform 1 0 199180 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2165
timestamp 1649977179
transform 1 0 200284 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2177
timestamp 1649977179
transform 1 0 201388 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2183
timestamp 1649977179
transform 1 0 201940 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2185
timestamp 1649977179
transform 1 0 202124 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2197
timestamp 1649977179
transform 1 0 203228 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2209
timestamp 1649977179
transform 1 0 204332 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2221
timestamp 1649977179
transform 1 0 205436 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2233
timestamp 1649977179
transform 1 0 206540 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2239
timestamp 1649977179
transform 1 0 207092 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2241
timestamp 1649977179
transform 1 0 207276 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2253
timestamp 1649977179
transform 1 0 208380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2265
timestamp 1649977179
transform 1 0 209484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2277
timestamp 1649977179
transform 1 0 210588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2289
timestamp 1649977179
transform 1 0 211692 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2295
timestamp 1649977179
transform 1 0 212244 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2297
timestamp 1649977179
transform 1 0 212428 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2309
timestamp 1649977179
transform 1 0 213532 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2321
timestamp 1649977179
transform 1 0 214636 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2333
timestamp 1649977179
transform 1 0 215740 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2345
timestamp 1649977179
transform 1 0 216844 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2351
timestamp 1649977179
transform 1 0 217396 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2353
timestamp 1649977179
transform 1 0 217580 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2365
timestamp 1649977179
transform 1 0 218684 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2377
timestamp 1649977179
transform 1 0 219788 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2389
timestamp 1649977179
transform 1 0 220892 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2401
timestamp 1649977179
transform 1 0 221996 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2407
timestamp 1649977179
transform 1 0 222548 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2409
timestamp 1649977179
transform 1 0 222732 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2421
timestamp 1649977179
transform 1 0 223836 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2433
timestamp 1649977179
transform 1 0 224940 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2445
timestamp 1649977179
transform 1 0 226044 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2457
timestamp 1649977179
transform 1 0 227148 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2463
timestamp 1649977179
transform 1 0 227700 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2465
timestamp 1649977179
transform 1 0 227884 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2477
timestamp 1649977179
transform 1 0 228988 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2489
timestamp 1649977179
transform 1 0 230092 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2501
timestamp 1649977179
transform 1 0 231196 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2513
timestamp 1649977179
transform 1 0 232300 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2519
timestamp 1649977179
transform 1 0 232852 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2521
timestamp 1649977179
transform 1 0 233036 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2533
timestamp 1649977179
transform 1 0 234140 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2545
timestamp 1649977179
transform 1 0 235244 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2557
timestamp 1649977179
transform 1 0 236348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2569
timestamp 1649977179
transform 1 0 237452 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2575
timestamp 1649977179
transform 1 0 238004 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2577
timestamp 1649977179
transform 1 0 238188 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2589
timestamp 1649977179
transform 1 0 239292 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2601
timestamp 1649977179
transform 1 0 240396 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2613
timestamp 1649977179
transform 1 0 241500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2625
timestamp 1649977179
transform 1 0 242604 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2631
timestamp 1649977179
transform 1 0 243156 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2633
timestamp 1649977179
transform 1 0 243340 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2645
timestamp 1649977179
transform 1 0 244444 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2657
timestamp 1649977179
transform 1 0 245548 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2669
timestamp 1649977179
transform 1 0 246652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2681
timestamp 1649977179
transform 1 0 247756 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2687
timestamp 1649977179
transform 1 0 248308 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2689
timestamp 1649977179
transform 1 0 248492 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2701
timestamp 1649977179
transform 1 0 249596 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2713
timestamp 1649977179
transform 1 0 250700 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2725
timestamp 1649977179
transform 1 0 251804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2737
timestamp 1649977179
transform 1 0 252908 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2743
timestamp 1649977179
transform 1 0 253460 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2745
timestamp 1649977179
transform 1 0 253644 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2757
timestamp 1649977179
transform 1 0 254748 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2769
timestamp 1649977179
transform 1 0 255852 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2781
timestamp 1649977179
transform 1 0 256956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2793
timestamp 1649977179
transform 1 0 258060 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2799
timestamp 1649977179
transform 1 0 258612 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2801
timestamp 1649977179
transform 1 0 258796 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2813
timestamp 1649977179
transform 1 0 259900 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2825
timestamp 1649977179
transform 1 0 261004 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2837
timestamp 1649977179
transform 1 0 262108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2849
timestamp 1649977179
transform 1 0 263212 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2855
timestamp 1649977179
transform 1 0 263764 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2857
timestamp 1649977179
transform 1 0 263948 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2869
timestamp 1649977179
transform 1 0 265052 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2881
timestamp 1649977179
transform 1 0 266156 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2893
timestamp 1649977179
transform 1 0 267260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2905
timestamp 1649977179
transform 1 0 268364 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2911
timestamp 1649977179
transform 1 0 268916 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2913
timestamp 1649977179
transform 1 0 269100 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2925
timestamp 1649977179
transform 1 0 270204 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2937
timestamp 1649977179
transform 1 0 271308 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2949
timestamp 1649977179
transform 1 0 272412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2961
timestamp 1649977179
transform 1 0 273516 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2967
timestamp 1649977179
transform 1 0 274068 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2969
timestamp 1649977179
transform 1 0 274252 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2981
timestamp 1649977179
transform 1 0 275356 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2993
timestamp 1649977179
transform 1 0 276460 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3005
timestamp 1649977179
transform 1 0 277564 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3017
timestamp 1649977179
transform 1 0 278668 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3023
timestamp 1649977179
transform 1 0 279220 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3025
timestamp 1649977179
transform 1 0 279404 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3037
timestamp 1649977179
transform 1 0 280508 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3049
timestamp 1649977179
transform 1 0 281612 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3061
timestamp 1649977179
transform 1 0 282716 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3073
timestamp 1649977179
transform 1 0 283820 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3079
timestamp 1649977179
transform 1 0 284372 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3081
timestamp 1649977179
transform 1 0 284556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3093
timestamp 1649977179
transform 1 0 285660 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3105
timestamp 1649977179
transform 1 0 286764 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3117
timestamp 1649977179
transform 1 0 287868 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3129
timestamp 1649977179
transform 1 0 288972 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3135
timestamp 1649977179
transform 1 0 289524 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3137
timestamp 1649977179
transform 1 0 289708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3149
timestamp 1649977179
transform 1 0 290812 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3161
timestamp 1649977179
transform 1 0 291916 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3173
timestamp 1649977179
transform 1 0 293020 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3185
timestamp 1649977179
transform 1 0 294124 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3191
timestamp 1649977179
transform 1 0 294676 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3193
timestamp 1649977179
transform 1 0 294860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3205
timestamp 1649977179
transform 1 0 295964 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3217
timestamp 1649977179
transform 1 0 297068 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3229
timestamp 1649977179
transform 1 0 298172 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3241
timestamp 1649977179
transform 1 0 299276 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3247
timestamp 1649977179
transform 1 0 299828 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3249
timestamp 1649977179
transform 1 0 300012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3261
timestamp 1649977179
transform 1 0 301116 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3273
timestamp 1649977179
transform 1 0 302220 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3285
timestamp 1649977179
transform 1 0 303324 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3297
timestamp 1649977179
transform 1 0 304428 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3303
timestamp 1649977179
transform 1 0 304980 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3305
timestamp 1649977179
transform 1 0 305164 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1649977179
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1649977179
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1649977179
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1649977179
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1649977179
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1649977179
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1649977179
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1649977179
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1649977179
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1649977179
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1649977179
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1649977179
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1649977179
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1649977179
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1649977179
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1649977179
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1649977179
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1649977179
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1649977179
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1649977179
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1649977179
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1649977179
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1649977179
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1649977179
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1649977179
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1649977179
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1649977179
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1649977179
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1649977179
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1649977179
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1649977179
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1649977179
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1649977179
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1649977179
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1649977179
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1649977179
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1649977179
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1649977179
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1649977179
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1649977179
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1649977179
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_601
timestamp 1649977179
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_613
timestamp 1649977179
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_625
timestamp 1649977179
transform 1 0 58604 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_637
timestamp 1649977179
transform 1 0 59708 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_643
timestamp 1649977179
transform 1 0 60260 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_645
timestamp 1649977179
transform 1 0 60444 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_657
timestamp 1649977179
transform 1 0 61548 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_669
timestamp 1649977179
transform 1 0 62652 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_681
timestamp 1649977179
transform 1 0 63756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_693
timestamp 1649977179
transform 1 0 64860 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_699
timestamp 1649977179
transform 1 0 65412 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_701
timestamp 1649977179
transform 1 0 65596 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_713
timestamp 1649977179
transform 1 0 66700 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_725
timestamp 1649977179
transform 1 0 67804 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_737
timestamp 1649977179
transform 1 0 68908 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_749
timestamp 1649977179
transform 1 0 70012 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_755
timestamp 1649977179
transform 1 0 70564 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_757
timestamp 1649977179
transform 1 0 70748 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_769
timestamp 1649977179
transform 1 0 71852 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_781
timestamp 1649977179
transform 1 0 72956 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_793
timestamp 1649977179
transform 1 0 74060 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_805
timestamp 1649977179
transform 1 0 75164 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_811
timestamp 1649977179
transform 1 0 75716 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_813
timestamp 1649977179
transform 1 0 75900 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_825
timestamp 1649977179
transform 1 0 77004 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_837
timestamp 1649977179
transform 1 0 78108 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_849
timestamp 1649977179
transform 1 0 79212 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_861
timestamp 1649977179
transform 1 0 80316 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_867
timestamp 1649977179
transform 1 0 80868 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_869
timestamp 1649977179
transform 1 0 81052 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_881
timestamp 1649977179
transform 1 0 82156 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_893
timestamp 1649977179
transform 1 0 83260 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_905
timestamp 1649977179
transform 1 0 84364 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_917
timestamp 1649977179
transform 1 0 85468 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_923
timestamp 1649977179
transform 1 0 86020 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_925
timestamp 1649977179
transform 1 0 86204 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_937
timestamp 1649977179
transform 1 0 87308 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_949
timestamp 1649977179
transform 1 0 88412 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_961
timestamp 1649977179
transform 1 0 89516 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_973
timestamp 1649977179
transform 1 0 90620 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_979
timestamp 1649977179
transform 1 0 91172 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_981
timestamp 1649977179
transform 1 0 91356 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_993
timestamp 1649977179
transform 1 0 92460 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1005
timestamp 1649977179
transform 1 0 93564 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1017
timestamp 1649977179
transform 1 0 94668 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1029
timestamp 1649977179
transform 1 0 95772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1035
timestamp 1649977179
transform 1 0 96324 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1037
timestamp 1649977179
transform 1 0 96508 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1049
timestamp 1649977179
transform 1 0 97612 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1061
timestamp 1649977179
transform 1 0 98716 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1073
timestamp 1649977179
transform 1 0 99820 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1085
timestamp 1649977179
transform 1 0 100924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1091
timestamp 1649977179
transform 1 0 101476 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1093
timestamp 1649977179
transform 1 0 101660 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1105
timestamp 1649977179
transform 1 0 102764 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1117
timestamp 1649977179
transform 1 0 103868 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1129
timestamp 1649977179
transform 1 0 104972 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1141
timestamp 1649977179
transform 1 0 106076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1147
timestamp 1649977179
transform 1 0 106628 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1149
timestamp 1649977179
transform 1 0 106812 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1161
timestamp 1649977179
transform 1 0 107916 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1173
timestamp 1649977179
transform 1 0 109020 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1185
timestamp 1649977179
transform 1 0 110124 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1197
timestamp 1649977179
transform 1 0 111228 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1203
timestamp 1649977179
transform 1 0 111780 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1205
timestamp 1649977179
transform 1 0 111964 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1217
timestamp 1649977179
transform 1 0 113068 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1229
timestamp 1649977179
transform 1 0 114172 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1241
timestamp 1649977179
transform 1 0 115276 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1253
timestamp 1649977179
transform 1 0 116380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1259
timestamp 1649977179
transform 1 0 116932 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1261
timestamp 1649977179
transform 1 0 117116 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1273
timestamp 1649977179
transform 1 0 118220 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1285
timestamp 1649977179
transform 1 0 119324 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1297
timestamp 1649977179
transform 1 0 120428 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1309
timestamp 1649977179
transform 1 0 121532 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1315
timestamp 1649977179
transform 1 0 122084 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1317
timestamp 1649977179
transform 1 0 122268 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1329
timestamp 1649977179
transform 1 0 123372 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1341
timestamp 1649977179
transform 1 0 124476 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1353
timestamp 1649977179
transform 1 0 125580 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1365
timestamp 1649977179
transform 1 0 126684 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1371
timestamp 1649977179
transform 1 0 127236 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1373
timestamp 1649977179
transform 1 0 127420 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1385
timestamp 1649977179
transform 1 0 128524 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1397
timestamp 1649977179
transform 1 0 129628 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1409
timestamp 1649977179
transform 1 0 130732 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1421
timestamp 1649977179
transform 1 0 131836 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1427
timestamp 1649977179
transform 1 0 132388 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1429
timestamp 1649977179
transform 1 0 132572 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1441
timestamp 1649977179
transform 1 0 133676 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1453
timestamp 1649977179
transform 1 0 134780 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1465
timestamp 1649977179
transform 1 0 135884 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1477
timestamp 1649977179
transform 1 0 136988 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1483
timestamp 1649977179
transform 1 0 137540 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1485
timestamp 1649977179
transform 1 0 137724 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1497
timestamp 1649977179
transform 1 0 138828 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1509
timestamp 1649977179
transform 1 0 139932 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1521
timestamp 1649977179
transform 1 0 141036 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1533
timestamp 1649977179
transform 1 0 142140 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1539
timestamp 1649977179
transform 1 0 142692 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1541
timestamp 1649977179
transform 1 0 142876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1553
timestamp 1649977179
transform 1 0 143980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1565
timestamp 1649977179
transform 1 0 145084 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1577
timestamp 1649977179
transform 1 0 146188 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1589
timestamp 1649977179
transform 1 0 147292 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1595
timestamp 1649977179
transform 1 0 147844 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1597
timestamp 1649977179
transform 1 0 148028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1609
timestamp 1649977179
transform 1 0 149132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1621
timestamp 1649977179
transform 1 0 150236 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1633
timestamp 1649977179
transform 1 0 151340 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1645
timestamp 1649977179
transform 1 0 152444 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1651
timestamp 1649977179
transform 1 0 152996 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1653
timestamp 1649977179
transform 1 0 153180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1665
timestamp 1649977179
transform 1 0 154284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1677
timestamp 1649977179
transform 1 0 155388 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1689
timestamp 1649977179
transform 1 0 156492 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1701
timestamp 1649977179
transform 1 0 157596 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1707
timestamp 1649977179
transform 1 0 158148 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1709
timestamp 1649977179
transform 1 0 158332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1721
timestamp 1649977179
transform 1 0 159436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1733
timestamp 1649977179
transform 1 0 160540 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1745
timestamp 1649977179
transform 1 0 161644 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1757
timestamp 1649977179
transform 1 0 162748 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1763
timestamp 1649977179
transform 1 0 163300 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1765
timestamp 1649977179
transform 1 0 163484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1777
timestamp 1649977179
transform 1 0 164588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1789
timestamp 1649977179
transform 1 0 165692 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1801
timestamp 1649977179
transform 1 0 166796 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1813
timestamp 1649977179
transform 1 0 167900 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1819
timestamp 1649977179
transform 1 0 168452 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1821
timestamp 1649977179
transform 1 0 168636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1833
timestamp 1649977179
transform 1 0 169740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1845
timestamp 1649977179
transform 1 0 170844 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1857
timestamp 1649977179
transform 1 0 171948 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1869
timestamp 1649977179
transform 1 0 173052 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1875
timestamp 1649977179
transform 1 0 173604 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1877
timestamp 1649977179
transform 1 0 173788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1889
timestamp 1649977179
transform 1 0 174892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1901
timestamp 1649977179
transform 1 0 175996 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1913
timestamp 1649977179
transform 1 0 177100 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1925
timestamp 1649977179
transform 1 0 178204 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1931
timestamp 1649977179
transform 1 0 178756 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1933
timestamp 1649977179
transform 1 0 178940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1945
timestamp 1649977179
transform 1 0 180044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1957
timestamp 1649977179
transform 1 0 181148 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1969
timestamp 1649977179
transform 1 0 182252 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1981
timestamp 1649977179
transform 1 0 183356 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1987
timestamp 1649977179
transform 1 0 183908 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1989
timestamp 1649977179
transform 1 0 184092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2001
timestamp 1649977179
transform 1 0 185196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2013
timestamp 1649977179
transform 1 0 186300 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2025
timestamp 1649977179
transform 1 0 187404 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2037
timestamp 1649977179
transform 1 0 188508 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2043
timestamp 1649977179
transform 1 0 189060 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2045
timestamp 1649977179
transform 1 0 189244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2057
timestamp 1649977179
transform 1 0 190348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2069
timestamp 1649977179
transform 1 0 191452 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2081
timestamp 1649977179
transform 1 0 192556 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2093
timestamp 1649977179
transform 1 0 193660 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2099
timestamp 1649977179
transform 1 0 194212 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2101
timestamp 1649977179
transform 1 0 194396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2113
timestamp 1649977179
transform 1 0 195500 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2125
timestamp 1649977179
transform 1 0 196604 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2137
timestamp 1649977179
transform 1 0 197708 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2149
timestamp 1649977179
transform 1 0 198812 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2155
timestamp 1649977179
transform 1 0 199364 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2157
timestamp 1649977179
transform 1 0 199548 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2169
timestamp 1649977179
transform 1 0 200652 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2181
timestamp 1649977179
transform 1 0 201756 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2193
timestamp 1649977179
transform 1 0 202860 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2205
timestamp 1649977179
transform 1 0 203964 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2211
timestamp 1649977179
transform 1 0 204516 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2213
timestamp 1649977179
transform 1 0 204700 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2225
timestamp 1649977179
transform 1 0 205804 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2237
timestamp 1649977179
transform 1 0 206908 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2249
timestamp 1649977179
transform 1 0 208012 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2261
timestamp 1649977179
transform 1 0 209116 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2267
timestamp 1649977179
transform 1 0 209668 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2269
timestamp 1649977179
transform 1 0 209852 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2281
timestamp 1649977179
transform 1 0 210956 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2293
timestamp 1649977179
transform 1 0 212060 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2305
timestamp 1649977179
transform 1 0 213164 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2317
timestamp 1649977179
transform 1 0 214268 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2323
timestamp 1649977179
transform 1 0 214820 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2325
timestamp 1649977179
transform 1 0 215004 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2337
timestamp 1649977179
transform 1 0 216108 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2349
timestamp 1649977179
transform 1 0 217212 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2361
timestamp 1649977179
transform 1 0 218316 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2373
timestamp 1649977179
transform 1 0 219420 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2379
timestamp 1649977179
transform 1 0 219972 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2381
timestamp 1649977179
transform 1 0 220156 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2393
timestamp 1649977179
transform 1 0 221260 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2405
timestamp 1649977179
transform 1 0 222364 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2417
timestamp 1649977179
transform 1 0 223468 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2429
timestamp 1649977179
transform 1 0 224572 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2435
timestamp 1649977179
transform 1 0 225124 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2437
timestamp 1649977179
transform 1 0 225308 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2449
timestamp 1649977179
transform 1 0 226412 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2461
timestamp 1649977179
transform 1 0 227516 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2473
timestamp 1649977179
transform 1 0 228620 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2485
timestamp 1649977179
transform 1 0 229724 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2491
timestamp 1649977179
transform 1 0 230276 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2493
timestamp 1649977179
transform 1 0 230460 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2505
timestamp 1649977179
transform 1 0 231564 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2517
timestamp 1649977179
transform 1 0 232668 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2529
timestamp 1649977179
transform 1 0 233772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2541
timestamp 1649977179
transform 1 0 234876 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2547
timestamp 1649977179
transform 1 0 235428 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2549
timestamp 1649977179
transform 1 0 235612 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2561
timestamp 1649977179
transform 1 0 236716 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2573
timestamp 1649977179
transform 1 0 237820 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2585
timestamp 1649977179
transform 1 0 238924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2597
timestamp 1649977179
transform 1 0 240028 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2603
timestamp 1649977179
transform 1 0 240580 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2605
timestamp 1649977179
transform 1 0 240764 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2617
timestamp 1649977179
transform 1 0 241868 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2629
timestamp 1649977179
transform 1 0 242972 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2641
timestamp 1649977179
transform 1 0 244076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2653
timestamp 1649977179
transform 1 0 245180 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2659
timestamp 1649977179
transform 1 0 245732 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2661
timestamp 1649977179
transform 1 0 245916 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2673
timestamp 1649977179
transform 1 0 247020 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2685
timestamp 1649977179
transform 1 0 248124 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2697
timestamp 1649977179
transform 1 0 249228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2709
timestamp 1649977179
transform 1 0 250332 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2715
timestamp 1649977179
transform 1 0 250884 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2717
timestamp 1649977179
transform 1 0 251068 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2729
timestamp 1649977179
transform 1 0 252172 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2741
timestamp 1649977179
transform 1 0 253276 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2753
timestamp 1649977179
transform 1 0 254380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2765
timestamp 1649977179
transform 1 0 255484 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2771
timestamp 1649977179
transform 1 0 256036 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2773
timestamp 1649977179
transform 1 0 256220 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2785
timestamp 1649977179
transform 1 0 257324 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2797
timestamp 1649977179
transform 1 0 258428 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2809
timestamp 1649977179
transform 1 0 259532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2821
timestamp 1649977179
transform 1 0 260636 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2827
timestamp 1649977179
transform 1 0 261188 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2829
timestamp 1649977179
transform 1 0 261372 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2841
timestamp 1649977179
transform 1 0 262476 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2853
timestamp 1649977179
transform 1 0 263580 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2865
timestamp 1649977179
transform 1 0 264684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2877
timestamp 1649977179
transform 1 0 265788 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2883
timestamp 1649977179
transform 1 0 266340 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2885
timestamp 1649977179
transform 1 0 266524 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2897
timestamp 1649977179
transform 1 0 267628 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2909
timestamp 1649977179
transform 1 0 268732 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2921
timestamp 1649977179
transform 1 0 269836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2933
timestamp 1649977179
transform 1 0 270940 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2939
timestamp 1649977179
transform 1 0 271492 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2941
timestamp 1649977179
transform 1 0 271676 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2953
timestamp 1649977179
transform 1 0 272780 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2965
timestamp 1649977179
transform 1 0 273884 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2977
timestamp 1649977179
transform 1 0 274988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2989
timestamp 1649977179
transform 1 0 276092 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2995
timestamp 1649977179
transform 1 0 276644 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2997
timestamp 1649977179
transform 1 0 276828 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3009
timestamp 1649977179
transform 1 0 277932 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3021
timestamp 1649977179
transform 1 0 279036 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3033
timestamp 1649977179
transform 1 0 280140 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3045
timestamp 1649977179
transform 1 0 281244 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3051
timestamp 1649977179
transform 1 0 281796 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3053
timestamp 1649977179
transform 1 0 281980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3065
timestamp 1649977179
transform 1 0 283084 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3077
timestamp 1649977179
transform 1 0 284188 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3089
timestamp 1649977179
transform 1 0 285292 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3101
timestamp 1649977179
transform 1 0 286396 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3107
timestamp 1649977179
transform 1 0 286948 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3109
timestamp 1649977179
transform 1 0 287132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3121
timestamp 1649977179
transform 1 0 288236 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3133
timestamp 1649977179
transform 1 0 289340 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3145
timestamp 1649977179
transform 1 0 290444 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3157
timestamp 1649977179
transform 1 0 291548 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3163
timestamp 1649977179
transform 1 0 292100 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3165
timestamp 1649977179
transform 1 0 292284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3177
timestamp 1649977179
transform 1 0 293388 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3189
timestamp 1649977179
transform 1 0 294492 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3201
timestamp 1649977179
transform 1 0 295596 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3213
timestamp 1649977179
transform 1 0 296700 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3219
timestamp 1649977179
transform 1 0 297252 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3221
timestamp 1649977179
transform 1 0 297436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3233
timestamp 1649977179
transform 1 0 298540 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3245
timestamp 1649977179
transform 1 0 299644 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3257
timestamp 1649977179
transform 1 0 300748 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3269
timestamp 1649977179
transform 1 0 301852 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3275
timestamp 1649977179
transform 1 0 302404 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3277
timestamp 1649977179
transform 1 0 302588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3289
timestamp 1649977179
transform 1 0 303692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3301
timestamp 1649977179
transform 1 0 304796 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1649977179
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1649977179
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1649977179
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1649977179
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1649977179
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1649977179
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1649977179
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1649977179
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1649977179
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1649977179
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1649977179
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1649977179
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1649977179
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_317
timestamp 1649977179
transform 1 0 30268 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_325
timestamp 1649977179
transform 1 0 31004 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1649977179
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1649977179
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_340
timestamp 1649977179
transform 1 0 32384 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_347
timestamp 1649977179
transform 1 0 33028 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_359
timestamp 1649977179
transform 1 0 34132 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_371
timestamp 1649977179
transform 1 0 35236 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_383
timestamp 1649977179
transform 1 0 36340 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1649977179
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1649977179
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1649977179
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1649977179
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1649977179
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1649977179
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1649977179
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1649977179
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1649977179
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1649977179
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1649977179
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1649977179
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1649977179
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1649977179
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1649977179
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1649977179
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1649977179
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1649977179
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1649977179
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1649977179
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1649977179
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1649977179
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_597
timestamp 1649977179
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1649977179
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1649977179
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_617
timestamp 1649977179
transform 1 0 57868 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_629
timestamp 1649977179
transform 1 0 58972 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_641
timestamp 1649977179
transform 1 0 60076 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_653
timestamp 1649977179
transform 1 0 61180 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_665
timestamp 1649977179
transform 1 0 62284 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_671
timestamp 1649977179
transform 1 0 62836 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_673
timestamp 1649977179
transform 1 0 63020 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_685
timestamp 1649977179
transform 1 0 64124 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_697
timestamp 1649977179
transform 1 0 65228 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_709
timestamp 1649977179
transform 1 0 66332 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_721
timestamp 1649977179
transform 1 0 67436 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_727
timestamp 1649977179
transform 1 0 67988 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_729
timestamp 1649977179
transform 1 0 68172 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_741
timestamp 1649977179
transform 1 0 69276 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_753
timestamp 1649977179
transform 1 0 70380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_765
timestamp 1649977179
transform 1 0 71484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_777
timestamp 1649977179
transform 1 0 72588 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_783
timestamp 1649977179
transform 1 0 73140 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_785
timestamp 1649977179
transform 1 0 73324 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_797
timestamp 1649977179
transform 1 0 74428 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_809
timestamp 1649977179
transform 1 0 75532 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_821
timestamp 1649977179
transform 1 0 76636 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_833
timestamp 1649977179
transform 1 0 77740 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_839
timestamp 1649977179
transform 1 0 78292 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_841
timestamp 1649977179
transform 1 0 78476 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_853
timestamp 1649977179
transform 1 0 79580 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_865
timestamp 1649977179
transform 1 0 80684 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_877
timestamp 1649977179
transform 1 0 81788 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_889
timestamp 1649977179
transform 1 0 82892 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_895
timestamp 1649977179
transform 1 0 83444 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_897
timestamp 1649977179
transform 1 0 83628 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_909
timestamp 1649977179
transform 1 0 84732 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_921
timestamp 1649977179
transform 1 0 85836 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_933
timestamp 1649977179
transform 1 0 86940 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_945
timestamp 1649977179
transform 1 0 88044 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_951
timestamp 1649977179
transform 1 0 88596 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_953
timestamp 1649977179
transform 1 0 88780 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_965
timestamp 1649977179
transform 1 0 89884 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_977
timestamp 1649977179
transform 1 0 90988 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_989
timestamp 1649977179
transform 1 0 92092 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1001
timestamp 1649977179
transform 1 0 93196 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1007
timestamp 1649977179
transform 1 0 93748 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1009
timestamp 1649977179
transform 1 0 93932 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1021
timestamp 1649977179
transform 1 0 95036 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1033
timestamp 1649977179
transform 1 0 96140 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1045
timestamp 1649977179
transform 1 0 97244 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1057
timestamp 1649977179
transform 1 0 98348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1063
timestamp 1649977179
transform 1 0 98900 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1065
timestamp 1649977179
transform 1 0 99084 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1077
timestamp 1649977179
transform 1 0 100188 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1089
timestamp 1649977179
transform 1 0 101292 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1101
timestamp 1649977179
transform 1 0 102396 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1113
timestamp 1649977179
transform 1 0 103500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1119
timestamp 1649977179
transform 1 0 104052 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1121
timestamp 1649977179
transform 1 0 104236 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1133
timestamp 1649977179
transform 1 0 105340 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1145
timestamp 1649977179
transform 1 0 106444 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1157
timestamp 1649977179
transform 1 0 107548 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1169
timestamp 1649977179
transform 1 0 108652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1175
timestamp 1649977179
transform 1 0 109204 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1177
timestamp 1649977179
transform 1 0 109388 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1189
timestamp 1649977179
transform 1 0 110492 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1201
timestamp 1649977179
transform 1 0 111596 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1213
timestamp 1649977179
transform 1 0 112700 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1225
timestamp 1649977179
transform 1 0 113804 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1231
timestamp 1649977179
transform 1 0 114356 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1233
timestamp 1649977179
transform 1 0 114540 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1245
timestamp 1649977179
transform 1 0 115644 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1257
timestamp 1649977179
transform 1 0 116748 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1269
timestamp 1649977179
transform 1 0 117852 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1281
timestamp 1649977179
transform 1 0 118956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1287
timestamp 1649977179
transform 1 0 119508 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1289
timestamp 1649977179
transform 1 0 119692 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1301
timestamp 1649977179
transform 1 0 120796 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1313
timestamp 1649977179
transform 1 0 121900 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1325
timestamp 1649977179
transform 1 0 123004 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1337
timestamp 1649977179
transform 1 0 124108 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1343
timestamp 1649977179
transform 1 0 124660 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1345
timestamp 1649977179
transform 1 0 124844 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1357
timestamp 1649977179
transform 1 0 125948 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1369
timestamp 1649977179
transform 1 0 127052 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1381
timestamp 1649977179
transform 1 0 128156 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1393
timestamp 1649977179
transform 1 0 129260 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1399
timestamp 1649977179
transform 1 0 129812 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1401
timestamp 1649977179
transform 1 0 129996 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1413
timestamp 1649977179
transform 1 0 131100 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1425
timestamp 1649977179
transform 1 0 132204 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1437
timestamp 1649977179
transform 1 0 133308 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1449
timestamp 1649977179
transform 1 0 134412 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1455
timestamp 1649977179
transform 1 0 134964 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1457
timestamp 1649977179
transform 1 0 135148 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1469
timestamp 1649977179
transform 1 0 136252 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1481
timestamp 1649977179
transform 1 0 137356 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1493
timestamp 1649977179
transform 1 0 138460 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1505
timestamp 1649977179
transform 1 0 139564 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1511
timestamp 1649977179
transform 1 0 140116 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1513
timestamp 1649977179
transform 1 0 140300 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1537
timestamp 1649977179
transform 1 0 142508 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1549
timestamp 1649977179
transform 1 0 143612 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1561
timestamp 1649977179
transform 1 0 144716 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1567
timestamp 1649977179
transform 1 0 145268 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1569
timestamp 1649977179
transform 1 0 145452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1581
timestamp 1649977179
transform 1 0 146556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1593
timestamp 1649977179
transform 1 0 147660 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1605
timestamp 1649977179
transform 1 0 148764 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1617
timestamp 1649977179
transform 1 0 149868 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1623
timestamp 1649977179
transform 1 0 150420 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1625
timestamp 1649977179
transform 1 0 150604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1637
timestamp 1649977179
transform 1 0 151708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1649
timestamp 1649977179
transform 1 0 152812 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1661
timestamp 1649977179
transform 1 0 153916 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1673
timestamp 1649977179
transform 1 0 155020 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1679
timestamp 1649977179
transform 1 0 155572 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1681
timestamp 1649977179
transform 1 0 155756 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1705
timestamp 1649977179
transform 1 0 157964 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1717
timestamp 1649977179
transform 1 0 159068 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1729
timestamp 1649977179
transform 1 0 160172 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1735
timestamp 1649977179
transform 1 0 160724 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1737
timestamp 1649977179
transform 1 0 160908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1749
timestamp 1649977179
transform 1 0 162012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1761
timestamp 1649977179
transform 1 0 163116 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1773
timestamp 1649977179
transform 1 0 164220 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1785
timestamp 1649977179
transform 1 0 165324 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1791
timestamp 1649977179
transform 1 0 165876 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1793
timestamp 1649977179
transform 1 0 166060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1805
timestamp 1649977179
transform 1 0 167164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1817
timestamp 1649977179
transform 1 0 168268 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1829
timestamp 1649977179
transform 1 0 169372 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1841
timestamp 1649977179
transform 1 0 170476 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1847
timestamp 1649977179
transform 1 0 171028 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1849
timestamp 1649977179
transform 1 0 171212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1861
timestamp 1649977179
transform 1 0 172316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1873
timestamp 1649977179
transform 1 0 173420 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1885
timestamp 1649977179
transform 1 0 174524 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1897
timestamp 1649977179
transform 1 0 175628 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1903
timestamp 1649977179
transform 1 0 176180 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1905
timestamp 1649977179
transform 1 0 176364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1917
timestamp 1649977179
transform 1 0 177468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1929
timestamp 1649977179
transform 1 0 178572 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1941
timestamp 1649977179
transform 1 0 179676 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1953
timestamp 1649977179
transform 1 0 180780 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1959
timestamp 1649977179
transform 1 0 181332 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1961
timestamp 1649977179
transform 1 0 181516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1973
timestamp 1649977179
transform 1 0 182620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1985
timestamp 1649977179
transform 1 0 183724 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1997
timestamp 1649977179
transform 1 0 184828 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2009
timestamp 1649977179
transform 1 0 185932 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2015
timestamp 1649977179
transform 1 0 186484 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2017
timestamp 1649977179
transform 1 0 186668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2029
timestamp 1649977179
transform 1 0 187772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2041
timestamp 1649977179
transform 1 0 188876 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2053
timestamp 1649977179
transform 1 0 189980 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2065
timestamp 1649977179
transform 1 0 191084 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2071
timestamp 1649977179
transform 1 0 191636 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_2073
timestamp 1649977179
transform 1 0 191820 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2077
timestamp 1649977179
transform 1 0 192188 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_2081
timestamp 1649977179
transform 1 0 192556 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2088
timestamp 1649977179
transform 1 0 193200 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2100
timestamp 1649977179
transform 1 0 194304 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2112
timestamp 1649977179
transform 1 0 195408 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_2124
timestamp 1649977179
transform 1 0 196512 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2129
timestamp 1649977179
transform 1 0 196972 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2141
timestamp 1649977179
transform 1 0 198076 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2153
timestamp 1649977179
transform 1 0 199180 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2165
timestamp 1649977179
transform 1 0 200284 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2177
timestamp 1649977179
transform 1 0 201388 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2183
timestamp 1649977179
transform 1 0 201940 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2185
timestamp 1649977179
transform 1 0 202124 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2197
timestamp 1649977179
transform 1 0 203228 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2209
timestamp 1649977179
transform 1 0 204332 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2221
timestamp 1649977179
transform 1 0 205436 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2233
timestamp 1649977179
transform 1 0 206540 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2239
timestamp 1649977179
transform 1 0 207092 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2241
timestamp 1649977179
transform 1 0 207276 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2253
timestamp 1649977179
transform 1 0 208380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2265
timestamp 1649977179
transform 1 0 209484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2277
timestamp 1649977179
transform 1 0 210588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2289
timestamp 1649977179
transform 1 0 211692 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2295
timestamp 1649977179
transform 1 0 212244 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2297
timestamp 1649977179
transform 1 0 212428 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2309
timestamp 1649977179
transform 1 0 213532 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2321
timestamp 1649977179
transform 1 0 214636 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2333
timestamp 1649977179
transform 1 0 215740 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2345
timestamp 1649977179
transform 1 0 216844 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2351
timestamp 1649977179
transform 1 0 217396 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2353
timestamp 1649977179
transform 1 0 217580 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2365
timestamp 1649977179
transform 1 0 218684 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2377
timestamp 1649977179
transform 1 0 219788 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2389
timestamp 1649977179
transform 1 0 220892 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2401
timestamp 1649977179
transform 1 0 221996 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2407
timestamp 1649977179
transform 1 0 222548 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2409
timestamp 1649977179
transform 1 0 222732 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2421
timestamp 1649977179
transform 1 0 223836 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2433
timestamp 1649977179
transform 1 0 224940 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2445
timestamp 1649977179
transform 1 0 226044 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2457
timestamp 1649977179
transform 1 0 227148 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2463
timestamp 1649977179
transform 1 0 227700 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2465
timestamp 1649977179
transform 1 0 227884 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2477
timestamp 1649977179
transform 1 0 228988 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2489
timestamp 1649977179
transform 1 0 230092 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2501
timestamp 1649977179
transform 1 0 231196 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2513
timestamp 1649977179
transform 1 0 232300 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2519
timestamp 1649977179
transform 1 0 232852 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2521
timestamp 1649977179
transform 1 0 233036 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2533
timestamp 1649977179
transform 1 0 234140 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2545
timestamp 1649977179
transform 1 0 235244 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2557
timestamp 1649977179
transform 1 0 236348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2569
timestamp 1649977179
transform 1 0 237452 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2575
timestamp 1649977179
transform 1 0 238004 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2577
timestamp 1649977179
transform 1 0 238188 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2589
timestamp 1649977179
transform 1 0 239292 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2601
timestamp 1649977179
transform 1 0 240396 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2613
timestamp 1649977179
transform 1 0 241500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2625
timestamp 1649977179
transform 1 0 242604 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2631
timestamp 1649977179
transform 1 0 243156 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2633
timestamp 1649977179
transform 1 0 243340 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2645
timestamp 1649977179
transform 1 0 244444 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2657
timestamp 1649977179
transform 1 0 245548 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2669
timestamp 1649977179
transform 1 0 246652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2681
timestamp 1649977179
transform 1 0 247756 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2687
timestamp 1649977179
transform 1 0 248308 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2689
timestamp 1649977179
transform 1 0 248492 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2701
timestamp 1649977179
transform 1 0 249596 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2713
timestamp 1649977179
transform 1 0 250700 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2725
timestamp 1649977179
transform 1 0 251804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2737
timestamp 1649977179
transform 1 0 252908 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2743
timestamp 1649977179
transform 1 0 253460 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2745
timestamp 1649977179
transform 1 0 253644 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2757
timestamp 1649977179
transform 1 0 254748 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2769
timestamp 1649977179
transform 1 0 255852 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2781
timestamp 1649977179
transform 1 0 256956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2793
timestamp 1649977179
transform 1 0 258060 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2799
timestamp 1649977179
transform 1 0 258612 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2801
timestamp 1649977179
transform 1 0 258796 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2813
timestamp 1649977179
transform 1 0 259900 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2825
timestamp 1649977179
transform 1 0 261004 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2837
timestamp 1649977179
transform 1 0 262108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2849
timestamp 1649977179
transform 1 0 263212 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2855
timestamp 1649977179
transform 1 0 263764 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2857
timestamp 1649977179
transform 1 0 263948 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2869
timestamp 1649977179
transform 1 0 265052 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2881
timestamp 1649977179
transform 1 0 266156 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2893
timestamp 1649977179
transform 1 0 267260 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_2902
timestamp 1649977179
transform 1 0 268088 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_2910
timestamp 1649977179
transform 1 0 268824 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2913
timestamp 1649977179
transform 1 0 269100 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2925
timestamp 1649977179
transform 1 0 270204 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2937
timestamp 1649977179
transform 1 0 271308 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2949
timestamp 1649977179
transform 1 0 272412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2961
timestamp 1649977179
transform 1 0 273516 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2967
timestamp 1649977179
transform 1 0 274068 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2969
timestamp 1649977179
transform 1 0 274252 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2981
timestamp 1649977179
transform 1 0 275356 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2993
timestamp 1649977179
transform 1 0 276460 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3005
timestamp 1649977179
transform 1 0 277564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3017
timestamp 1649977179
transform 1 0 278668 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3023
timestamp 1649977179
transform 1 0 279220 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3025
timestamp 1649977179
transform 1 0 279404 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3037
timestamp 1649977179
transform 1 0 280508 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3049
timestamp 1649977179
transform 1 0 281612 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3061
timestamp 1649977179
transform 1 0 282716 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3073
timestamp 1649977179
transform 1 0 283820 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3079
timestamp 1649977179
transform 1 0 284372 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3081
timestamp 1649977179
transform 1 0 284556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3093
timestamp 1649977179
transform 1 0 285660 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3105
timestamp 1649977179
transform 1 0 286764 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3117
timestamp 1649977179
transform 1 0 287868 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3129
timestamp 1649977179
transform 1 0 288972 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3135
timestamp 1649977179
transform 1 0 289524 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3137
timestamp 1649977179
transform 1 0 289708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3149
timestamp 1649977179
transform 1 0 290812 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3161
timestamp 1649977179
transform 1 0 291916 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3173
timestamp 1649977179
transform 1 0 293020 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3185
timestamp 1649977179
transform 1 0 294124 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3191
timestamp 1649977179
transform 1 0 294676 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3193
timestamp 1649977179
transform 1 0 294860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3205
timestamp 1649977179
transform 1 0 295964 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3217
timestamp 1649977179
transform 1 0 297068 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3229
timestamp 1649977179
transform 1 0 298172 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3241
timestamp 1649977179
transform 1 0 299276 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3247
timestamp 1649977179
transform 1 0 299828 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3249
timestamp 1649977179
transform 1 0 300012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3261
timestamp 1649977179
transform 1 0 301116 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3273
timestamp 1649977179
transform 1 0 302220 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3285
timestamp 1649977179
transform 1 0 303324 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3297
timestamp 1649977179
transform 1 0 304428 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3303
timestamp 1649977179
transform 1 0 304980 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3305
timestamp 1649977179
transform 1 0 305164 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1649977179
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1649977179
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1649977179
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1649977179
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1649977179
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1649977179
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1649977179
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1649977179
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1649977179
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1649977179
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1649977179
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1649977179
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_309
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_320
timestamp 1649977179
transform 1 0 30544 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_327
timestamp 1649977179
transform 1 0 31188 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_334
timestamp 1649977179
transform 1 0 31832 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_341
timestamp 1649977179
transform 1 0 32476 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_348
timestamp 1649977179
transform 1 0 33120 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_355
timestamp 1649977179
transform 1 0 33764 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1649977179
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1649977179
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1649977179
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1649977179
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1649977179
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1649977179
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1649977179
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1649977179
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1649977179
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1649977179
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1649977179
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1649977179
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1649977179
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1649977179
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1649977179
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1649977179
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1649977179
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1649977179
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1649977179
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1649977179
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1649977179
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1649977179
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1649977179
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1649977179
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1649977179
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_601
timestamp 1649977179
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_613
timestamp 1649977179
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_625
timestamp 1649977179
transform 1 0 58604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_637
timestamp 1649977179
transform 1 0 59708 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_643
timestamp 1649977179
transform 1 0 60260 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_645
timestamp 1649977179
transform 1 0 60444 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_657
timestamp 1649977179
transform 1 0 61548 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_669
timestamp 1649977179
transform 1 0 62652 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_681
timestamp 1649977179
transform 1 0 63756 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_693
timestamp 1649977179
transform 1 0 64860 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_699
timestamp 1649977179
transform 1 0 65412 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_701
timestamp 1649977179
transform 1 0 65596 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_713
timestamp 1649977179
transform 1 0 66700 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_725
timestamp 1649977179
transform 1 0 67804 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_737
timestamp 1649977179
transform 1 0 68908 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_749
timestamp 1649977179
transform 1 0 70012 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_755
timestamp 1649977179
transform 1 0 70564 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_757
timestamp 1649977179
transform 1 0 70748 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_769
timestamp 1649977179
transform 1 0 71852 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_781
timestamp 1649977179
transform 1 0 72956 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_793
timestamp 1649977179
transform 1 0 74060 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_805
timestamp 1649977179
transform 1 0 75164 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_811
timestamp 1649977179
transform 1 0 75716 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_813
timestamp 1649977179
transform 1 0 75900 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_825
timestamp 1649977179
transform 1 0 77004 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_837
timestamp 1649977179
transform 1 0 78108 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_849
timestamp 1649977179
transform 1 0 79212 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_861
timestamp 1649977179
transform 1 0 80316 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_867
timestamp 1649977179
transform 1 0 80868 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_869
timestamp 1649977179
transform 1 0 81052 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_881
timestamp 1649977179
transform 1 0 82156 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_893
timestamp 1649977179
transform 1 0 83260 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_905
timestamp 1649977179
transform 1 0 84364 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_917
timestamp 1649977179
transform 1 0 85468 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_923
timestamp 1649977179
transform 1 0 86020 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_925
timestamp 1649977179
transform 1 0 86204 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_937
timestamp 1649977179
transform 1 0 87308 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_949
timestamp 1649977179
transform 1 0 88412 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_961
timestamp 1649977179
transform 1 0 89516 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_973
timestamp 1649977179
transform 1 0 90620 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_979
timestamp 1649977179
transform 1 0 91172 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_981
timestamp 1649977179
transform 1 0 91356 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_993
timestamp 1649977179
transform 1 0 92460 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1005
timestamp 1649977179
transform 1 0 93564 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1017
timestamp 1649977179
transform 1 0 94668 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1029
timestamp 1649977179
transform 1 0 95772 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1035
timestamp 1649977179
transform 1 0 96324 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1037
timestamp 1649977179
transform 1 0 96508 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1049
timestamp 1649977179
transform 1 0 97612 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1061
timestamp 1649977179
transform 1 0 98716 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1073
timestamp 1649977179
transform 1 0 99820 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1085
timestamp 1649977179
transform 1 0 100924 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1091
timestamp 1649977179
transform 1 0 101476 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1093
timestamp 1649977179
transform 1 0 101660 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1105
timestamp 1649977179
transform 1 0 102764 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1117
timestamp 1649977179
transform 1 0 103868 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1129
timestamp 1649977179
transform 1 0 104972 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1141
timestamp 1649977179
transform 1 0 106076 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1147
timestamp 1649977179
transform 1 0 106628 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1149
timestamp 1649977179
transform 1 0 106812 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1161
timestamp 1649977179
transform 1 0 107916 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1173
timestamp 1649977179
transform 1 0 109020 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1185
timestamp 1649977179
transform 1 0 110124 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1197
timestamp 1649977179
transform 1 0 111228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1203
timestamp 1649977179
transform 1 0 111780 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1205
timestamp 1649977179
transform 1 0 111964 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1217
timestamp 1649977179
transform 1 0 113068 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1229
timestamp 1649977179
transform 1 0 114172 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1241
timestamp 1649977179
transform 1 0 115276 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1253
timestamp 1649977179
transform 1 0 116380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1259
timestamp 1649977179
transform 1 0 116932 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1261
timestamp 1649977179
transform 1 0 117116 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1273
timestamp 1649977179
transform 1 0 118220 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1285
timestamp 1649977179
transform 1 0 119324 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1297
timestamp 1649977179
transform 1 0 120428 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1309
timestamp 1649977179
transform 1 0 121532 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1315
timestamp 1649977179
transform 1 0 122084 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1317
timestamp 1649977179
transform 1 0 122268 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1329
timestamp 1649977179
transform 1 0 123372 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1341
timestamp 1649977179
transform 1 0 124476 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1353
timestamp 1649977179
transform 1 0 125580 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1365
timestamp 1649977179
transform 1 0 126684 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1371
timestamp 1649977179
transform 1 0 127236 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1373
timestamp 1649977179
transform 1 0 127420 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1385
timestamp 1649977179
transform 1 0 128524 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1397
timestamp 1649977179
transform 1 0 129628 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1409
timestamp 1649977179
transform 1 0 130732 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1421
timestamp 1649977179
transform 1 0 131836 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1427
timestamp 1649977179
transform 1 0 132388 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1429
timestamp 1649977179
transform 1 0 132572 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1441
timestamp 1649977179
transform 1 0 133676 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1453
timestamp 1649977179
transform 1 0 134780 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1465
timestamp 1649977179
transform 1 0 135884 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1477
timestamp 1649977179
transform 1 0 136988 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1483
timestamp 1649977179
transform 1 0 137540 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1485
timestamp 1649977179
transform 1 0 137724 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1497
timestamp 1649977179
transform 1 0 138828 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1509
timestamp 1649977179
transform 1 0 139932 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1513
timestamp 1649977179
transform 1 0 140300 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1534
timestamp 1649977179
transform 1 0 142232 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1541
timestamp 1649977179
transform 1 0 142876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1553
timestamp 1649977179
transform 1 0 143980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1565
timestamp 1649977179
transform 1 0 145084 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1577
timestamp 1649977179
transform 1 0 146188 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1589
timestamp 1649977179
transform 1 0 147292 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1595
timestamp 1649977179
transform 1 0 147844 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1597
timestamp 1649977179
transform 1 0 148028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1609
timestamp 1649977179
transform 1 0 149132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1621
timestamp 1649977179
transform 1 0 150236 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1633
timestamp 1649977179
transform 1 0 151340 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1645
timestamp 1649977179
transform 1 0 152444 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1651
timestamp 1649977179
transform 1 0 152996 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1653
timestamp 1649977179
transform 1 0 153180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1665
timestamp 1649977179
transform 1 0 154284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1677
timestamp 1649977179
transform 1 0 155388 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1683
timestamp 1649977179
transform 1 0 155940 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1704
timestamp 1649977179
transform 1 0 157872 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1709
timestamp 1649977179
transform 1 0 158332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1721
timestamp 1649977179
transform 1 0 159436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1733
timestamp 1649977179
transform 1 0 160540 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1745
timestamp 1649977179
transform 1 0 161644 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1757
timestamp 1649977179
transform 1 0 162748 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1763
timestamp 1649977179
transform 1 0 163300 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1765
timestamp 1649977179
transform 1 0 163484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1777
timestamp 1649977179
transform 1 0 164588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1789
timestamp 1649977179
transform 1 0 165692 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1801
timestamp 1649977179
transform 1 0 166796 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1813
timestamp 1649977179
transform 1 0 167900 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1819
timestamp 1649977179
transform 1 0 168452 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1821
timestamp 1649977179
transform 1 0 168636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1833
timestamp 1649977179
transform 1 0 169740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1845
timestamp 1649977179
transform 1 0 170844 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1857
timestamp 1649977179
transform 1 0 171948 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1869
timestamp 1649977179
transform 1 0 173052 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1875
timestamp 1649977179
transform 1 0 173604 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1877
timestamp 1649977179
transform 1 0 173788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1889
timestamp 1649977179
transform 1 0 174892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1901
timestamp 1649977179
transform 1 0 175996 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1913
timestamp 1649977179
transform 1 0 177100 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1925
timestamp 1649977179
transform 1 0 178204 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1931
timestamp 1649977179
transform 1 0 178756 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1933
timestamp 1649977179
transform 1 0 178940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1945
timestamp 1649977179
transform 1 0 180044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1957
timestamp 1649977179
transform 1 0 181148 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1969
timestamp 1649977179
transform 1 0 182252 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1981
timestamp 1649977179
transform 1 0 183356 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1987
timestamp 1649977179
transform 1 0 183908 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1989
timestamp 1649977179
transform 1 0 184092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2001
timestamp 1649977179
transform 1 0 185196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2013
timestamp 1649977179
transform 1 0 186300 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2025
timestamp 1649977179
transform 1 0 187404 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2037
timestamp 1649977179
transform 1 0 188508 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2043
timestamp 1649977179
transform 1 0 189060 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2045
timestamp 1649977179
transform 1 0 189244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2057
timestamp 1649977179
transform 1 0 190348 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_2069
timestamp 1649977179
transform 1 0 191452 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_2076
timestamp 1649977179
transform 1 0 192096 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_2083
timestamp 1649977179
transform 1 0 192740 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_2090
timestamp 1649977179
transform 1 0 193384 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_2098
timestamp 1649977179
transform 1 0 194120 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2101
timestamp 1649977179
transform 1 0 194396 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2113
timestamp 1649977179
transform 1 0 195500 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2125
timestamp 1649977179
transform 1 0 196604 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2137
timestamp 1649977179
transform 1 0 197708 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2149
timestamp 1649977179
transform 1 0 198812 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2155
timestamp 1649977179
transform 1 0 199364 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2157
timestamp 1649977179
transform 1 0 199548 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2169
timestamp 1649977179
transform 1 0 200652 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2181
timestamp 1649977179
transform 1 0 201756 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2193
timestamp 1649977179
transform 1 0 202860 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2205
timestamp 1649977179
transform 1 0 203964 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2211
timestamp 1649977179
transform 1 0 204516 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2213
timestamp 1649977179
transform 1 0 204700 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2225
timestamp 1649977179
transform 1 0 205804 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2237
timestamp 1649977179
transform 1 0 206908 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2249
timestamp 1649977179
transform 1 0 208012 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2261
timestamp 1649977179
transform 1 0 209116 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2267
timestamp 1649977179
transform 1 0 209668 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2269
timestamp 1649977179
transform 1 0 209852 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2281
timestamp 1649977179
transform 1 0 210956 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2293
timestamp 1649977179
transform 1 0 212060 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2305
timestamp 1649977179
transform 1 0 213164 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2317
timestamp 1649977179
transform 1 0 214268 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2323
timestamp 1649977179
transform 1 0 214820 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2325
timestamp 1649977179
transform 1 0 215004 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2337
timestamp 1649977179
transform 1 0 216108 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2349
timestamp 1649977179
transform 1 0 217212 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2361
timestamp 1649977179
transform 1 0 218316 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2373
timestamp 1649977179
transform 1 0 219420 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2379
timestamp 1649977179
transform 1 0 219972 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2381
timestamp 1649977179
transform 1 0 220156 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2393
timestamp 1649977179
transform 1 0 221260 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2405
timestamp 1649977179
transform 1 0 222364 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2417
timestamp 1649977179
transform 1 0 223468 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2429
timestamp 1649977179
transform 1 0 224572 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2435
timestamp 1649977179
transform 1 0 225124 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2437
timestamp 1649977179
transform 1 0 225308 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2449
timestamp 1649977179
transform 1 0 226412 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2461
timestamp 1649977179
transform 1 0 227516 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2473
timestamp 1649977179
transform 1 0 228620 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2485
timestamp 1649977179
transform 1 0 229724 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2491
timestamp 1649977179
transform 1 0 230276 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2493
timestamp 1649977179
transform 1 0 230460 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2505
timestamp 1649977179
transform 1 0 231564 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2517
timestamp 1649977179
transform 1 0 232668 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2529
timestamp 1649977179
transform 1 0 233772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2541
timestamp 1649977179
transform 1 0 234876 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2547
timestamp 1649977179
transform 1 0 235428 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2549
timestamp 1649977179
transform 1 0 235612 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2561
timestamp 1649977179
transform 1 0 236716 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2573
timestamp 1649977179
transform 1 0 237820 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2585
timestamp 1649977179
transform 1 0 238924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2597
timestamp 1649977179
transform 1 0 240028 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2603
timestamp 1649977179
transform 1 0 240580 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2605
timestamp 1649977179
transform 1 0 240764 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2617
timestamp 1649977179
transform 1 0 241868 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2629
timestamp 1649977179
transform 1 0 242972 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2641
timestamp 1649977179
transform 1 0 244076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2653
timestamp 1649977179
transform 1 0 245180 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2659
timestamp 1649977179
transform 1 0 245732 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2661
timestamp 1649977179
transform 1 0 245916 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2673
timestamp 1649977179
transform 1 0 247020 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2685
timestamp 1649977179
transform 1 0 248124 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2697
timestamp 1649977179
transform 1 0 249228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2709
timestamp 1649977179
transform 1 0 250332 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2715
timestamp 1649977179
transform 1 0 250884 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2717
timestamp 1649977179
transform 1 0 251068 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2729
timestamp 1649977179
transform 1 0 252172 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2741
timestamp 1649977179
transform 1 0 253276 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2753
timestamp 1649977179
transform 1 0 254380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2765
timestamp 1649977179
transform 1 0 255484 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2771
timestamp 1649977179
transform 1 0 256036 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2773
timestamp 1649977179
transform 1 0 256220 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2785
timestamp 1649977179
transform 1 0 257324 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2797
timestamp 1649977179
transform 1 0 258428 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2809
timestamp 1649977179
transform 1 0 259532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2821
timestamp 1649977179
transform 1 0 260636 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2827
timestamp 1649977179
transform 1 0 261188 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2829
timestamp 1649977179
transform 1 0 261372 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2841
timestamp 1649977179
transform 1 0 262476 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2853
timestamp 1649977179
transform 1 0 263580 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2865
timestamp 1649977179
transform 1 0 264684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2877
timestamp 1649977179
transform 1 0 265788 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2883
timestamp 1649977179
transform 1 0 266340 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2885
timestamp 1649977179
transform 1 0 266524 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_2894
timestamp 1649977179
transform 1 0 267352 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_2901
timestamp 1649977179
transform 1 0 267996 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_2908
timestamp 1649977179
transform 1 0 268640 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2915
timestamp 1649977179
transform 1 0 269284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2927
timestamp 1649977179
transform 1 0 270388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2939
timestamp 1649977179
transform 1 0 271492 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2941
timestamp 1649977179
transform 1 0 271676 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2953
timestamp 1649977179
transform 1 0 272780 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2965
timestamp 1649977179
transform 1 0 273884 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2977
timestamp 1649977179
transform 1 0 274988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2989
timestamp 1649977179
transform 1 0 276092 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2995
timestamp 1649977179
transform 1 0 276644 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_2997
timestamp 1649977179
transform 1 0 276828 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3009
timestamp 1649977179
transform 1 0 277932 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3021
timestamp 1649977179
transform 1 0 279036 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3033
timestamp 1649977179
transform 1 0 280140 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3045
timestamp 1649977179
transform 1 0 281244 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3051
timestamp 1649977179
transform 1 0 281796 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3053
timestamp 1649977179
transform 1 0 281980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3065
timestamp 1649977179
transform 1 0 283084 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3077
timestamp 1649977179
transform 1 0 284188 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3089
timestamp 1649977179
transform 1 0 285292 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3101
timestamp 1649977179
transform 1 0 286396 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3107
timestamp 1649977179
transform 1 0 286948 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3109
timestamp 1649977179
transform 1 0 287132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3121
timestamp 1649977179
transform 1 0 288236 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3133
timestamp 1649977179
transform 1 0 289340 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3145
timestamp 1649977179
transform 1 0 290444 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3157
timestamp 1649977179
transform 1 0 291548 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3163
timestamp 1649977179
transform 1 0 292100 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3165
timestamp 1649977179
transform 1 0 292284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3177
timestamp 1649977179
transform 1 0 293388 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3189
timestamp 1649977179
transform 1 0 294492 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3201
timestamp 1649977179
transform 1 0 295596 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3213
timestamp 1649977179
transform 1 0 296700 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3219
timestamp 1649977179
transform 1 0 297252 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3221
timestamp 1649977179
transform 1 0 297436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3233
timestamp 1649977179
transform 1 0 298540 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3245
timestamp 1649977179
transform 1 0 299644 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3257
timestamp 1649977179
transform 1 0 300748 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3269
timestamp 1649977179
transform 1 0 301852 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3275
timestamp 1649977179
transform 1 0 302404 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3277
timestamp 1649977179
transform 1 0 302588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3289
timestamp 1649977179
transform 1 0 303692 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3295
timestamp 1649977179
transform 1 0 304244 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3305
timestamp 1649977179
transform 1 0 305164 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1649977179
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1649977179
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1649977179
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1649977179
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1649977179
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1649977179
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1649977179
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1649977179
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1649977179
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1649977179
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1649977179
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1649977179
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1649977179
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1649977179
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_305
timestamp 1649977179
transform 1 0 29164 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_309
timestamp 1649977179
transform 1 0 29532 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_313
timestamp 1649977179
transform 1 0 29900 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_326
timestamp 1649977179
transform 1 0 31096 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_334
timestamp 1649977179
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_340
timestamp 1649977179
transform 1 0 32384 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_347
timestamp 1649977179
transform 1 0 33028 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_354
timestamp 1649977179
transform 1 0 33672 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_366
timestamp 1649977179
transform 1 0 34776 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_378
timestamp 1649977179
transform 1 0 35880 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_390
timestamp 1649977179
transform 1 0 36984 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1649977179
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1649977179
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1649977179
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1649977179
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1649977179
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1649977179
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1649977179
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1649977179
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1649977179
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1649977179
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1649977179
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1649977179
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1649977179
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1649977179
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1649977179
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1649977179
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1649977179
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1649977179
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1649977179
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1649977179
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_597
timestamp 1649977179
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1649977179
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1649977179
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_617
timestamp 1649977179
transform 1 0 57868 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_629
timestamp 1649977179
transform 1 0 58972 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_641
timestamp 1649977179
transform 1 0 60076 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_653
timestamp 1649977179
transform 1 0 61180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_665
timestamp 1649977179
transform 1 0 62284 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_671
timestamp 1649977179
transform 1 0 62836 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_673
timestamp 1649977179
transform 1 0 63020 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_685
timestamp 1649977179
transform 1 0 64124 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_697
timestamp 1649977179
transform 1 0 65228 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_709
timestamp 1649977179
transform 1 0 66332 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_721
timestamp 1649977179
transform 1 0 67436 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_727
timestamp 1649977179
transform 1 0 67988 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_729
timestamp 1649977179
transform 1 0 68172 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_741
timestamp 1649977179
transform 1 0 69276 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_753
timestamp 1649977179
transform 1 0 70380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_765
timestamp 1649977179
transform 1 0 71484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_777
timestamp 1649977179
transform 1 0 72588 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_783
timestamp 1649977179
transform 1 0 73140 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_785
timestamp 1649977179
transform 1 0 73324 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_797
timestamp 1649977179
transform 1 0 74428 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_809
timestamp 1649977179
transform 1 0 75532 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_821
timestamp 1649977179
transform 1 0 76636 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_833
timestamp 1649977179
transform 1 0 77740 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_839
timestamp 1649977179
transform 1 0 78292 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_841
timestamp 1649977179
transform 1 0 78476 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_853
timestamp 1649977179
transform 1 0 79580 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_865
timestamp 1649977179
transform 1 0 80684 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_877
timestamp 1649977179
transform 1 0 81788 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_889
timestamp 1649977179
transform 1 0 82892 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_895
timestamp 1649977179
transform 1 0 83444 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_897
timestamp 1649977179
transform 1 0 83628 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_909
timestamp 1649977179
transform 1 0 84732 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_921
timestamp 1649977179
transform 1 0 85836 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_933
timestamp 1649977179
transform 1 0 86940 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_945
timestamp 1649977179
transform 1 0 88044 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_951
timestamp 1649977179
transform 1 0 88596 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_953
timestamp 1649977179
transform 1 0 88780 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_965
timestamp 1649977179
transform 1 0 89884 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_977
timestamp 1649977179
transform 1 0 90988 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_989
timestamp 1649977179
transform 1 0 92092 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1001
timestamp 1649977179
transform 1 0 93196 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1007
timestamp 1649977179
transform 1 0 93748 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1009
timestamp 1649977179
transform 1 0 93932 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1021
timestamp 1649977179
transform 1 0 95036 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1033
timestamp 1649977179
transform 1 0 96140 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1045
timestamp 1649977179
transform 1 0 97244 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1057
timestamp 1649977179
transform 1 0 98348 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1063
timestamp 1649977179
transform 1 0 98900 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1065
timestamp 1649977179
transform 1 0 99084 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1077
timestamp 1649977179
transform 1 0 100188 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1089
timestamp 1649977179
transform 1 0 101292 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1096
timestamp 1649977179
transform 1 0 101936 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1108
timestamp 1649977179
transform 1 0 103040 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1121
timestamp 1649977179
transform 1 0 104236 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1133
timestamp 1649977179
transform 1 0 105340 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1145
timestamp 1649977179
transform 1 0 106444 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1157
timestamp 1649977179
transform 1 0 107548 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1169
timestamp 1649977179
transform 1 0 108652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1175
timestamp 1649977179
transform 1 0 109204 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1177
timestamp 1649977179
transform 1 0 109388 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1189
timestamp 1649977179
transform 1 0 110492 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1201
timestamp 1649977179
transform 1 0 111596 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1213
timestamp 1649977179
transform 1 0 112700 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1225
timestamp 1649977179
transform 1 0 113804 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1231
timestamp 1649977179
transform 1 0 114356 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1233
timestamp 1649977179
transform 1 0 114540 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1245
timestamp 1649977179
transform 1 0 115644 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1257
timestamp 1649977179
transform 1 0 116748 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1269
timestamp 1649977179
transform 1 0 117852 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1281
timestamp 1649977179
transform 1 0 118956 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1287
timestamp 1649977179
transform 1 0 119508 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1289
timestamp 1649977179
transform 1 0 119692 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1301
timestamp 1649977179
transform 1 0 120796 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1313
timestamp 1649977179
transform 1 0 121900 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1325
timestamp 1649977179
transform 1 0 123004 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1337
timestamp 1649977179
transform 1 0 124108 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1343
timestamp 1649977179
transform 1 0 124660 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1345
timestamp 1649977179
transform 1 0 124844 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1357
timestamp 1649977179
transform 1 0 125948 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1369
timestamp 1649977179
transform 1 0 127052 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1381
timestamp 1649977179
transform 1 0 128156 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1393
timestamp 1649977179
transform 1 0 129260 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1399
timestamp 1649977179
transform 1 0 129812 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1401
timestamp 1649977179
transform 1 0 129996 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1408
timestamp 1649977179
transform 1 0 130640 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1420
timestamp 1649977179
transform 1 0 131744 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1432
timestamp 1649977179
transform 1 0 132848 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1444
timestamp 1649977179
transform 1 0 133952 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1457
timestamp 1649977179
transform 1 0 135148 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1469
timestamp 1649977179
transform 1 0 136252 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1481
timestamp 1649977179
transform 1 0 137356 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1493
timestamp 1649977179
transform 1 0 138460 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1505
timestamp 1649977179
transform 1 0 139564 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1511
timestamp 1649977179
transform 1 0 140116 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1513
timestamp 1649977179
transform 1 0 140300 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1537
timestamp 1649977179
transform 1 0 142508 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1549
timestamp 1649977179
transform 1 0 143612 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1561
timestamp 1649977179
transform 1 0 144716 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1567
timestamp 1649977179
transform 1 0 145268 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1569
timestamp 1649977179
transform 1 0 145452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1581
timestamp 1649977179
transform 1 0 146556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1593
timestamp 1649977179
transform 1 0 147660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1605
timestamp 1649977179
transform 1 0 148764 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1609
timestamp 1649977179
transform 1 0 149132 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_1621
timestamp 1649977179
transform 1 0 150236 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1628
timestamp 1649977179
transform 1 0 150880 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1640
timestamp 1649977179
transform 1 0 151984 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1652
timestamp 1649977179
transform 1 0 153088 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1664
timestamp 1649977179
transform 1 0 154192 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1676
timestamp 1649977179
transform 1 0 155296 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1681
timestamp 1649977179
transform 1 0 155756 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1705
timestamp 1649977179
transform 1 0 157964 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1717
timestamp 1649977179
transform 1 0 159068 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1729
timestamp 1649977179
transform 1 0 160172 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1735
timestamp 1649977179
transform 1 0 160724 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1737
timestamp 1649977179
transform 1 0 160908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1749
timestamp 1649977179
transform 1 0 162012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1761
timestamp 1649977179
transform 1 0 163116 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1773
timestamp 1649977179
transform 1 0 164220 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1785
timestamp 1649977179
transform 1 0 165324 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1791
timestamp 1649977179
transform 1 0 165876 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1793
timestamp 1649977179
transform 1 0 166060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1805
timestamp 1649977179
transform 1 0 167164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1817
timestamp 1649977179
transform 1 0 168268 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1829
timestamp 1649977179
transform 1 0 169372 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1841
timestamp 1649977179
transform 1 0 170476 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1847
timestamp 1649977179
transform 1 0 171028 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1849
timestamp 1649977179
transform 1 0 171212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1861
timestamp 1649977179
transform 1 0 172316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1873
timestamp 1649977179
transform 1 0 173420 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1885
timestamp 1649977179
transform 1 0 174524 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1897
timestamp 1649977179
transform 1 0 175628 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1903
timestamp 1649977179
transform 1 0 176180 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1905
timestamp 1649977179
transform 1 0 176364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1917
timestamp 1649977179
transform 1 0 177468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1929
timestamp 1649977179
transform 1 0 178572 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1941
timestamp 1649977179
transform 1 0 179676 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1953
timestamp 1649977179
transform 1 0 180780 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1959
timestamp 1649977179
transform 1 0 181332 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1961
timestamp 1649977179
transform 1 0 181516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1973
timestamp 1649977179
transform 1 0 182620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1985
timestamp 1649977179
transform 1 0 183724 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1997
timestamp 1649977179
transform 1 0 184828 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_2009
timestamp 1649977179
transform 1 0 185932 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_2015
timestamp 1649977179
transform 1 0 186484 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_2017
timestamp 1649977179
transform 1 0 186668 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_2021
timestamp 1649977179
transform 1 0 187036 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2031
timestamp 1649977179
transform 1 0 187956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2043
timestamp 1649977179
transform 1 0 189060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_2055
timestamp 1649977179
transform 1 0 190164 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_2063
timestamp 1649977179
transform 1 0 190900 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_2068
timestamp 1649977179
transform 1 0 191360 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_2076
timestamp 1649977179
transform 1 0 192096 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_2086
timestamp 1649977179
transform 1 0 193016 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_2094
timestamp 1649977179
transform 1 0 193752 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2101
timestamp 1649977179
transform 1 0 194396 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2113
timestamp 1649977179
transform 1 0 195500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_2125
timestamp 1649977179
transform 1 0 196604 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2129
timestamp 1649977179
transform 1 0 196972 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2141
timestamp 1649977179
transform 1 0 198076 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2153
timestamp 1649977179
transform 1 0 199180 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2165
timestamp 1649977179
transform 1 0 200284 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_2177
timestamp 1649977179
transform 1 0 201388 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_2183
timestamp 1649977179
transform 1 0 201940 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_2185
timestamp 1649977179
transform 1 0 202124 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2196
timestamp 1649977179
transform 1 0 203136 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2208
timestamp 1649977179
transform 1 0 204240 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2220
timestamp 1649977179
transform 1 0 205344 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_2232
timestamp 1649977179
transform 1 0 206448 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2241
timestamp 1649977179
transform 1 0 207276 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2253
timestamp 1649977179
transform 1 0 208380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2265
timestamp 1649977179
transform 1 0 209484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2277
timestamp 1649977179
transform 1 0 210588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_2289
timestamp 1649977179
transform 1 0 211692 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_2295
timestamp 1649977179
transform 1 0 212244 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2297
timestamp 1649977179
transform 1 0 212428 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2309
timestamp 1649977179
transform 1 0 213532 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2321
timestamp 1649977179
transform 1 0 214636 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2333
timestamp 1649977179
transform 1 0 215740 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_2345
timestamp 1649977179
transform 1 0 216844 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_2351
timestamp 1649977179
transform 1 0 217396 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2353
timestamp 1649977179
transform 1 0 217580 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2365
timestamp 1649977179
transform 1 0 218684 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2377
timestamp 1649977179
transform 1 0 219788 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2389
timestamp 1649977179
transform 1 0 220892 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_2401
timestamp 1649977179
transform 1 0 221996 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_2407
timestamp 1649977179
transform 1 0 222548 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2409
timestamp 1649977179
transform 1 0 222732 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2421
timestamp 1649977179
transform 1 0 223836 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2433
timestamp 1649977179
transform 1 0 224940 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2445
timestamp 1649977179
transform 1 0 226044 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_2457
timestamp 1649977179
transform 1 0 227148 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_2463
timestamp 1649977179
transform 1 0 227700 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2465
timestamp 1649977179
transform 1 0 227884 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2477
timestamp 1649977179
transform 1 0 228988 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2489
timestamp 1649977179
transform 1 0 230092 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2501
timestamp 1649977179
transform 1 0 231196 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_2513
timestamp 1649977179
transform 1 0 232300 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_2519
timestamp 1649977179
transform 1 0 232852 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2521
timestamp 1649977179
transform 1 0 233036 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2533
timestamp 1649977179
transform 1 0 234140 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2545
timestamp 1649977179
transform 1 0 235244 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2557
timestamp 1649977179
transform 1 0 236348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_2569
timestamp 1649977179
transform 1 0 237452 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_2575
timestamp 1649977179
transform 1 0 238004 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2577
timestamp 1649977179
transform 1 0 238188 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2589
timestamp 1649977179
transform 1 0 239292 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2601
timestamp 1649977179
transform 1 0 240396 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2613
timestamp 1649977179
transform 1 0 241500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_2625
timestamp 1649977179
transform 1 0 242604 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_2631
timestamp 1649977179
transform 1 0 243156 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2633
timestamp 1649977179
transform 1 0 243340 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2645
timestamp 1649977179
transform 1 0 244444 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2657
timestamp 1649977179
transform 1 0 245548 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2669
timestamp 1649977179
transform 1 0 246652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_2681
timestamp 1649977179
transform 1 0 247756 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_2687
timestamp 1649977179
transform 1 0 248308 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2689
timestamp 1649977179
transform 1 0 248492 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2701
timestamp 1649977179
transform 1 0 249596 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2713
timestamp 1649977179
transform 1 0 250700 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2725
timestamp 1649977179
transform 1 0 251804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_2737
timestamp 1649977179
transform 1 0 252908 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_2743
timestamp 1649977179
transform 1 0 253460 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2748
timestamp 1649977179
transform 1 0 253920 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2760
timestamp 1649977179
transform 1 0 255024 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2772
timestamp 1649977179
transform 1 0 256128 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2784
timestamp 1649977179
transform 1 0 257232 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_2796
timestamp 1649977179
transform 1 0 258336 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2801
timestamp 1649977179
transform 1 0 258796 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2813
timestamp 1649977179
transform 1 0 259900 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2825
timestamp 1649977179
transform 1 0 261004 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2837
timestamp 1649977179
transform 1 0 262108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_2849
timestamp 1649977179
transform 1 0 263212 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_2855
timestamp 1649977179
transform 1 0 263764 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2857
timestamp 1649977179
transform 1 0 263948 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_2869
timestamp 1649977179
transform 1 0 265052 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_2880
timestamp 1649977179
transform 1 0 266064 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_2887
timestamp 1649977179
transform 1 0 266708 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_2894
timestamp 1649977179
transform 1 0 267352 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_2901
timestamp 1649977179
transform 1 0 267996 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_2908
timestamp 1649977179
transform 1 0 268640 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2916
timestamp 1649977179
transform 1 0 269376 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2928
timestamp 1649977179
transform 1 0 270480 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2940
timestamp 1649977179
transform 1 0 271584 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2952
timestamp 1649977179
transform 1 0 272688 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_2964
timestamp 1649977179
transform 1 0 273792 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2969
timestamp 1649977179
transform 1 0 274252 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2981
timestamp 1649977179
transform 1 0 275356 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_2993
timestamp 1649977179
transform 1 0 276460 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3005
timestamp 1649977179
transform 1 0 277564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3017
timestamp 1649977179
transform 1 0 278668 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3023
timestamp 1649977179
transform 1 0 279220 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3025
timestamp 1649977179
transform 1 0 279404 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3037
timestamp 1649977179
transform 1 0 280508 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3049
timestamp 1649977179
transform 1 0 281612 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3061
timestamp 1649977179
transform 1 0 282716 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3073
timestamp 1649977179
transform 1 0 283820 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3079
timestamp 1649977179
transform 1 0 284372 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3081
timestamp 1649977179
transform 1 0 284556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3093
timestamp 1649977179
transform 1 0 285660 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3105
timestamp 1649977179
transform 1 0 286764 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3117
timestamp 1649977179
transform 1 0 287868 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3129
timestamp 1649977179
transform 1 0 288972 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3135
timestamp 1649977179
transform 1 0 289524 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3137
timestamp 1649977179
transform 1 0 289708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3149
timestamp 1649977179
transform 1 0 290812 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3161
timestamp 1649977179
transform 1 0 291916 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3173
timestamp 1649977179
transform 1 0 293020 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3185
timestamp 1649977179
transform 1 0 294124 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3191
timestamp 1649977179
transform 1 0 294676 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3193
timestamp 1649977179
transform 1 0 294860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3205
timestamp 1649977179
transform 1 0 295964 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3217
timestamp 1649977179
transform 1 0 297068 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3229
timestamp 1649977179
transform 1 0 298172 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3241
timestamp 1649977179
transform 1 0 299276 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3247
timestamp 1649977179
transform 1 0 299828 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3249
timestamp 1649977179
transform 1 0 300012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3261
timestamp 1649977179
transform 1 0 301116 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3273
timestamp 1649977179
transform 1 0 302220 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3285
timestamp 1649977179
transform 1 0 303324 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3297
timestamp 1649977179
transform 1 0 304428 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3303
timestamp 1649977179
transform 1 0 304980 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3305
timestamp 1649977179
transform 1 0 305164 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1649977179
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1649977179
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1649977179
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1649977179
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1649977179
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1649977179
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1649977179
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1649977179
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1649977179
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1649977179
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1649977179
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1649977179
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_304
timestamp 1649977179
transform 1 0 29072 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_309
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_330
timestamp 1649977179
transform 1 0 31464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_343
timestamp 1649977179
transform 1 0 32660 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_351
timestamp 1649977179
transform 1 0 33396 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_355
timestamp 1649977179
transform 1 0 33764 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1649977179
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1649977179
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1649977179
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1649977179
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1649977179
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1649977179
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1649977179
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_421
timestamp 1649977179
transform 1 0 39836 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_425
timestamp 1649977179
transform 1 0 40204 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_429
timestamp 1649977179
transform 1 0 40572 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_436
timestamp 1649977179
transform 1 0 41216 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_443
timestamp 1649977179
transform 1 0 41860 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_450
timestamp 1649977179
transform 1 0 42504 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_462
timestamp 1649977179
transform 1 0 43608 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_474
timestamp 1649977179
transform 1 0 44712 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1649977179
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1649977179
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1649977179
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1649977179
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1649977179
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1649977179
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1649977179
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1649977179
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1649977179
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1649977179
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1649977179
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1649977179
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_592
timestamp 1649977179
transform 1 0 55568 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_598
timestamp 1649977179
transform 1 0 56120 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_602
timestamp 1649977179
transform 1 0 56488 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_614
timestamp 1649977179
transform 1 0 57592 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_626
timestamp 1649977179
transform 1 0 58696 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_638
timestamp 1649977179
transform 1 0 59800 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_645
timestamp 1649977179
transform 1 0 60444 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_657
timestamp 1649977179
transform 1 0 61548 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_669
timestamp 1649977179
transform 1 0 62652 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_681
timestamp 1649977179
transform 1 0 63756 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_693
timestamp 1649977179
transform 1 0 64860 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_699
timestamp 1649977179
transform 1 0 65412 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_701
timestamp 1649977179
transform 1 0 65596 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_713
timestamp 1649977179
transform 1 0 66700 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_725
timestamp 1649977179
transform 1 0 67804 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_737
timestamp 1649977179
transform 1 0 68908 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_749
timestamp 1649977179
transform 1 0 70012 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_755
timestamp 1649977179
transform 1 0 70564 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_757
timestamp 1649977179
transform 1 0 70748 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_769
timestamp 1649977179
transform 1 0 71852 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_781
timestamp 1649977179
transform 1 0 72956 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_793
timestamp 1649977179
transform 1 0 74060 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_805
timestamp 1649977179
transform 1 0 75164 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_811
timestamp 1649977179
transform 1 0 75716 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_813
timestamp 1649977179
transform 1 0 75900 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_822
timestamp 1649977179
transform 1 0 76728 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_834
timestamp 1649977179
transform 1 0 77832 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_841
timestamp 1649977179
transform 1 0 78476 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_853
timestamp 1649977179
transform 1 0 79580 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_865
timestamp 1649977179
transform 1 0 80684 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_869
timestamp 1649977179
transform 1 0 81052 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_881
timestamp 1649977179
transform 1 0 82156 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_893
timestamp 1649977179
transform 1 0 83260 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_905
timestamp 1649977179
transform 1 0 84364 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_917
timestamp 1649977179
transform 1 0 85468 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_923
timestamp 1649977179
transform 1 0 86020 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_928
timestamp 1649977179
transform 1 0 86480 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_935
timestamp 1649977179
transform 1 0 87124 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_939
timestamp 1649977179
transform 1 0 87492 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_943
timestamp 1649977179
transform 1 0 87860 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_950
timestamp 1649977179
transform 1 0 88504 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_962
timestamp 1649977179
transform 1 0 89608 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_974
timestamp 1649977179
transform 1 0 90712 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_981
timestamp 1649977179
transform 1 0 91356 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_993
timestamp 1649977179
transform 1 0 92460 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1005
timestamp 1649977179
transform 1 0 93564 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1017
timestamp 1649977179
transform 1 0 94668 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1029
timestamp 1649977179
transform 1 0 95772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1035
timestamp 1649977179
transform 1 0 96324 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1037
timestamp 1649977179
transform 1 0 96508 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1049
timestamp 1649977179
transform 1 0 97612 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1061
timestamp 1649977179
transform 1 0 98716 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1073
timestamp 1649977179
transform 1 0 99820 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1085
timestamp 1649977179
transform 1 0 100924 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1091
timestamp 1649977179
transform 1 0 101476 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1093
timestamp 1649977179
transform 1 0 101660 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1101
timestamp 1649977179
transform 1 0 102396 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1105
timestamp 1649977179
transform 1 0 102764 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1109
timestamp 1649977179
transform 1 0 103132 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1116
timestamp 1649977179
transform 1 0 103776 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1128
timestamp 1649977179
transform 1 0 104880 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1140
timestamp 1649977179
transform 1 0 105984 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1149
timestamp 1649977179
transform 1 0 106812 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1161
timestamp 1649977179
transform 1 0 107916 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1173
timestamp 1649977179
transform 1 0 109020 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1185
timestamp 1649977179
transform 1 0 110124 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1197
timestamp 1649977179
transform 1 0 111228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1203
timestamp 1649977179
transform 1 0 111780 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1205
timestamp 1649977179
transform 1 0 111964 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1217
timestamp 1649977179
transform 1 0 113068 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1229
timestamp 1649977179
transform 1 0 114172 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1244
timestamp 1649977179
transform 1 0 115552 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1248
timestamp 1649977179
transform 1 0 115920 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1252
timestamp 1649977179
transform 1 0 116288 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1264
timestamp 1649977179
transform 1 0 117392 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1276
timestamp 1649977179
transform 1 0 118496 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1288
timestamp 1649977179
transform 1 0 119600 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1300
timestamp 1649977179
transform 1 0 120704 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1312
timestamp 1649977179
transform 1 0 121808 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1317
timestamp 1649977179
transform 1 0 122268 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1329
timestamp 1649977179
transform 1 0 123372 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1341
timestamp 1649977179
transform 1 0 124476 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1353
timestamp 1649977179
transform 1 0 125580 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1365
timestamp 1649977179
transform 1 0 126684 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1371
timestamp 1649977179
transform 1 0 127236 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1373
timestamp 1649977179
transform 1 0 127420 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1385
timestamp 1649977179
transform 1 0 128524 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1397
timestamp 1649977179
transform 1 0 129628 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1405
timestamp 1649977179
transform 1 0 130364 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1409
timestamp 1649977179
transform 1 0 130732 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1416
timestamp 1649977179
transform 1 0 131376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1423
timestamp 1649977179
transform 1 0 132020 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1427
timestamp 1649977179
transform 1 0 132388 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1429
timestamp 1649977179
transform 1 0 132572 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1441
timestamp 1649977179
transform 1 0 133676 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1453
timestamp 1649977179
transform 1 0 134780 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1465
timestamp 1649977179
transform 1 0 135884 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1477
timestamp 1649977179
transform 1 0 136988 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1483
timestamp 1649977179
transform 1 0 137540 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1485
timestamp 1649977179
transform 1 0 137724 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1497
timestamp 1649977179
transform 1 0 138828 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1509
timestamp 1649977179
transform 1 0 139932 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1513
timestamp 1649977179
transform 1 0 140300 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1534
timestamp 1649977179
transform 1 0 142232 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1541
timestamp 1649977179
transform 1 0 142876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1553
timestamp 1649977179
transform 1 0 143980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1565
timestamp 1649977179
transform 1 0 145084 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1577
timestamp 1649977179
transform 1 0 146188 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1589
timestamp 1649977179
transform 1 0 147292 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1595
timestamp 1649977179
transform 1 0 147844 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1606
timestamp 1649977179
transform 1 0 148856 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1612
timestamp 1649977179
transform 1 0 149408 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1619
timestamp 1649977179
transform 1 0 150052 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1630
timestamp 1649977179
transform 1 0 151064 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1642
timestamp 1649977179
transform 1 0 152168 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1650
timestamp 1649977179
transform 1 0 152904 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1653
timestamp 1649977179
transform 1 0 153180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1665
timestamp 1649977179
transform 1 0 154284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1677
timestamp 1649977179
transform 1 0 155388 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1683
timestamp 1649977179
transform 1 0 155940 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1704
timestamp 1649977179
transform 1 0 157872 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1709
timestamp 1649977179
transform 1 0 158332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1721
timestamp 1649977179
transform 1 0 159436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1733
timestamp 1649977179
transform 1 0 160540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1745
timestamp 1649977179
transform 1 0 161644 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1752
timestamp 1649977179
transform 1 0 162288 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1759
timestamp 1649977179
transform 1 0 162932 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1763
timestamp 1649977179
transform 1 0 163300 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1768
timestamp 1649977179
transform 1 0 163760 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1780
timestamp 1649977179
transform 1 0 164864 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1792
timestamp 1649977179
transform 1 0 165968 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1804
timestamp 1649977179
transform 1 0 167072 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1816
timestamp 1649977179
transform 1 0 168176 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1821
timestamp 1649977179
transform 1 0 168636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1833
timestamp 1649977179
transform 1 0 169740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1845
timestamp 1649977179
transform 1 0 170844 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1857
timestamp 1649977179
transform 1 0 171948 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1869
timestamp 1649977179
transform 1 0 173052 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1875
timestamp 1649977179
transform 1 0 173604 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1877
timestamp 1649977179
transform 1 0 173788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1889
timestamp 1649977179
transform 1 0 174892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1901
timestamp 1649977179
transform 1 0 175996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1913
timestamp 1649977179
transform 1 0 177100 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1920
timestamp 1649977179
transform 1 0 177744 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1927
timestamp 1649977179
transform 1 0 178388 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1931
timestamp 1649977179
transform 1 0 178756 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1936
timestamp 1649977179
transform 1 0 179216 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1948
timestamp 1649977179
transform 1 0 180320 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1960
timestamp 1649977179
transform 1 0 181424 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1972
timestamp 1649977179
transform 1 0 182528 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1984
timestamp 1649977179
transform 1 0 183632 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1989
timestamp 1649977179
transform 1 0 184092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2001
timestamp 1649977179
transform 1 0 185196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2013
timestamp 1649977179
transform 1 0 186300 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2025
timestamp 1649977179
transform 1 0 187404 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_2037
timestamp 1649977179
transform 1 0 188508 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_2043
timestamp 1649977179
transform 1 0 189060 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_2045
timestamp 1649977179
transform 1 0 189244 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_2053
timestamp 1649977179
transform 1 0 189980 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2058
timestamp 1649977179
transform 1 0 190440 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_2065
timestamp 1649977179
transform 1 0 191084 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_2073
timestamp 1649977179
transform 1 0 191820 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2095
timestamp 1649977179
transform 1 0 193844 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_2099
timestamp 1649977179
transform 1 0 194212 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2110
timestamp 1649977179
transform 1 0 195224 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2117
timestamp 1649977179
transform 1 0 195868 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2129
timestamp 1649977179
transform 1 0 196972 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2141
timestamp 1649977179
transform 1 0 198076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_2153
timestamp 1649977179
transform 1 0 199180 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2157
timestamp 1649977179
transform 1 0 199548 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2169
timestamp 1649977179
transform 1 0 200652 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2181
timestamp 1649977179
transform 1 0 201756 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2188
timestamp 1649977179
transform 1 0 202400 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2195
timestamp 1649977179
transform 1 0 203044 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_2202
timestamp 1649977179
transform 1 0 203688 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_2210
timestamp 1649977179
transform 1 0 204424 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2216
timestamp 1649977179
transform 1 0 204976 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2228
timestamp 1649977179
transform 1 0 206080 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2240
timestamp 1649977179
transform 1 0 207184 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2252
timestamp 1649977179
transform 1 0 208288 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2264
timestamp 1649977179
transform 1 0 209392 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2269
timestamp 1649977179
transform 1 0 209852 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2281
timestamp 1649977179
transform 1 0 210956 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2293
timestamp 1649977179
transform 1 0 212060 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2305
timestamp 1649977179
transform 1 0 213164 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_2317
timestamp 1649977179
transform 1 0 214268 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_2323
timestamp 1649977179
transform 1 0 214820 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2325
timestamp 1649977179
transform 1 0 215004 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2337
timestamp 1649977179
transform 1 0 216108 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2349
timestamp 1649977179
transform 1 0 217212 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2361
timestamp 1649977179
transform 1 0 218316 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_2373
timestamp 1649977179
transform 1 0 219420 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_2379
timestamp 1649977179
transform 1 0 219972 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2381
timestamp 1649977179
transform 1 0 220156 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2393
timestamp 1649977179
transform 1 0 221260 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2405
timestamp 1649977179
transform 1 0 222364 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2417
timestamp 1649977179
transform 1 0 223468 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_2429
timestamp 1649977179
transform 1 0 224572 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_2435
timestamp 1649977179
transform 1 0 225124 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2437
timestamp 1649977179
transform 1 0 225308 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2449
timestamp 1649977179
transform 1 0 226412 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2461
timestamp 1649977179
transform 1 0 227516 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_2473
timestamp 1649977179
transform 1 0 228620 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_2482
timestamp 1649977179
transform 1 0 229448 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_2490
timestamp 1649977179
transform 1 0 230184 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2493
timestamp 1649977179
transform 1 0 230460 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2505
timestamp 1649977179
transform 1 0 231564 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2517
timestamp 1649977179
transform 1 0 232668 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2529
timestamp 1649977179
transform 1 0 233772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_2541
timestamp 1649977179
transform 1 0 234876 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_2547
timestamp 1649977179
transform 1 0 235428 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2549
timestamp 1649977179
transform 1 0 235612 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2561
timestamp 1649977179
transform 1 0 236716 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2573
timestamp 1649977179
transform 1 0 237820 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_2585
timestamp 1649977179
transform 1 0 238924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_2593
timestamp 1649977179
transform 1 0 239660 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_2598
timestamp 1649977179
transform 1 0 240120 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2608
timestamp 1649977179
transform 1 0 241040 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2615
timestamp 1649977179
transform 1 0 241684 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2622
timestamp 1649977179
transform 1 0 242328 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2634
timestamp 1649977179
transform 1 0 243432 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2646
timestamp 1649977179
transform 1 0 244536 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_2658
timestamp 1649977179
transform 1 0 245640 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2661
timestamp 1649977179
transform 1 0 245916 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2673
timestamp 1649977179
transform 1 0 247020 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2685
timestamp 1649977179
transform 1 0 248124 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2697
timestamp 1649977179
transform 1 0 249228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_2709
timestamp 1649977179
transform 1 0 250332 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_2715
timestamp 1649977179
transform 1 0 250884 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2717
timestamp 1649977179
transform 1 0 251068 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_2729
timestamp 1649977179
transform 1 0 252172 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2735
timestamp 1649977179
transform 1 0 252724 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2742
timestamp 1649977179
transform 1 0 253368 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2749
timestamp 1649977179
transform 1 0 254012 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2756
timestamp 1649977179
transform 1 0 254656 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2768
timestamp 1649977179
transform 1 0 255760 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2773
timestamp 1649977179
transform 1 0 256220 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2785
timestamp 1649977179
transform 1 0 257324 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2797
timestamp 1649977179
transform 1 0 258428 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2809
timestamp 1649977179
transform 1 0 259532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_2821
timestamp 1649977179
transform 1 0 260636 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_2827
timestamp 1649977179
transform 1 0 261188 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2829
timestamp 1649977179
transform 1 0 261372 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2841
timestamp 1649977179
transform 1 0 262476 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2853
timestamp 1649977179
transform 1 0 263580 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_2865
timestamp 1649977179
transform 1 0 264684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2870
timestamp 1649977179
transform 1 0 265144 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_2877
timestamp 1649977179
transform 1 0 265788 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_2883
timestamp 1649977179
transform 1 0 266340 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_2885
timestamp 1649977179
transform 1 0 266524 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2897
timestamp 1649977179
transform 1 0 267628 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_2904
timestamp 1649977179
transform 1 0 268272 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_2908
timestamp 1649977179
transform 1 0 268640 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_2919
timestamp 1649977179
transform 1 0 269652 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_2932
timestamp 1649977179
transform 1 0 270848 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2941
timestamp 1649977179
transform 1 0 271676 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2953
timestamp 1649977179
transform 1 0 272780 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2965
timestamp 1649977179
transform 1 0 273884 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2977
timestamp 1649977179
transform 1 0 274988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_2989
timestamp 1649977179
transform 1 0 276092 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_2995
timestamp 1649977179
transform 1 0 276644 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_2997
timestamp 1649977179
transform 1 0 276828 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3009
timestamp 1649977179
transform 1 0 277932 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3021
timestamp 1649977179
transform 1 0 279036 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3033
timestamp 1649977179
transform 1 0 280140 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3045
timestamp 1649977179
transform 1 0 281244 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3051
timestamp 1649977179
transform 1 0 281796 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3053
timestamp 1649977179
transform 1 0 281980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3065
timestamp 1649977179
transform 1 0 283084 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3077
timestamp 1649977179
transform 1 0 284188 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3089
timestamp 1649977179
transform 1 0 285292 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3101
timestamp 1649977179
transform 1 0 286396 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3107
timestamp 1649977179
transform 1 0 286948 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3109
timestamp 1649977179
transform 1 0 287132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3121
timestamp 1649977179
transform 1 0 288236 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3133
timestamp 1649977179
transform 1 0 289340 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3145
timestamp 1649977179
transform 1 0 290444 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3157
timestamp 1649977179
transform 1 0 291548 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3163
timestamp 1649977179
transform 1 0 292100 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3165
timestamp 1649977179
transform 1 0 292284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3177
timestamp 1649977179
transform 1 0 293388 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3189
timestamp 1649977179
transform 1 0 294492 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3201
timestamp 1649977179
transform 1 0 295596 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3213
timestamp 1649977179
transform 1 0 296700 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3219
timestamp 1649977179
transform 1 0 297252 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3221
timestamp 1649977179
transform 1 0 297436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3233
timestamp 1649977179
transform 1 0 298540 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3245
timestamp 1649977179
transform 1 0 299644 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3257
timestamp 1649977179
transform 1 0 300748 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3269
timestamp 1649977179
transform 1 0 301852 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3275
timestamp 1649977179
transform 1 0 302404 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3277
timestamp 1649977179
transform 1 0 302588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3289
timestamp 1649977179
transform 1 0 303692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_3301
timestamp 1649977179
transform 1 0 304796 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1649977179
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1649977179
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1649977179
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1649977179
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1649977179
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1649977179
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1649977179
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1649977179
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1649977179
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1649977179
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1649977179
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1649977179
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1649977179
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1649977179
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1649977179
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_289
timestamp 1649977179
transform 1 0 27692 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_293
timestamp 1649977179
transform 1 0 28060 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_306
timestamp 1649977179
transform 1 0 29256 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_330
timestamp 1649977179
transform 1 0 31464 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_346
timestamp 1649977179
transform 1 0 32936 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_357
timestamp 1649977179
transform 1 0 33948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_364
timestamp 1649977179
transform 1 0 34592 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_371
timestamp 1649977179
transform 1 0 35236 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_383
timestamp 1649977179
transform 1 0 36340 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1649977179
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1649977179
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_408
timestamp 1649977179
transform 1 0 38640 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_415
timestamp 1649977179
transform 1 0 39284 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_428
timestamp 1649977179
transform 1 0 40480 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_437
timestamp 1649977179
transform 1 0 41308 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_444
timestamp 1649977179
transform 1 0 41952 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_449
timestamp 1649977179
transform 1 0 42412 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_457
timestamp 1649977179
transform 1 0 43148 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1649977179
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1649977179
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1649977179
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1649977179
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1649977179
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1649977179
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1649977179
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1649977179
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1649977179
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1649977179
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1649977179
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_561
timestamp 1649977179
transform 1 0 52716 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_565
timestamp 1649977179
transform 1 0 53084 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_574
timestamp 1649977179
transform 1 0 53912 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_581
timestamp 1649977179
transform 1 0 54556 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_594
timestamp 1649977179
transform 1 0 55752 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_600
timestamp 1649977179
transform 1 0 56304 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_604
timestamp 1649977179
transform 1 0 56672 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_611
timestamp 1649977179
transform 1 0 57316 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1649977179
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_617
timestamp 1649977179
transform 1 0 57868 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_629
timestamp 1649977179
transform 1 0 58972 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_641
timestamp 1649977179
transform 1 0 60076 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_653
timestamp 1649977179
transform 1 0 61180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_665
timestamp 1649977179
transform 1 0 62284 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_671
timestamp 1649977179
transform 1 0 62836 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_673
timestamp 1649977179
transform 1 0 63020 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_685
timestamp 1649977179
transform 1 0 64124 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_697
timestamp 1649977179
transform 1 0 65228 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_709
timestamp 1649977179
transform 1 0 66332 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_721
timestamp 1649977179
transform 1 0 67436 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_727
timestamp 1649977179
transform 1 0 67988 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_729
timestamp 1649977179
transform 1 0 68172 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_741
timestamp 1649977179
transform 1 0 69276 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_753
timestamp 1649977179
transform 1 0 70380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_765
timestamp 1649977179
transform 1 0 71484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_777
timestamp 1649977179
transform 1 0 72588 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_783
timestamp 1649977179
transform 1 0 73140 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_785
timestamp 1649977179
transform 1 0 73324 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_797
timestamp 1649977179
transform 1 0 74428 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_818
timestamp 1649977179
transform 1 0 76360 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_17_827
timestamp 1649977179
transform 1 0 77188 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_836
timestamp 1649977179
transform 1 0 78016 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_844
timestamp 1649977179
transform 1 0 78752 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_856
timestamp 1649977179
transform 1 0 79856 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_868
timestamp 1649977179
transform 1 0 80960 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_880
timestamp 1649977179
transform 1 0 82064 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_892
timestamp 1649977179
transform 1 0 83168 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_897
timestamp 1649977179
transform 1 0 83628 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_908
timestamp 1649977179
transform 1 0 84640 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_915
timestamp 1649977179
transform 1 0 85284 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_928
timestamp 1649977179
transform 1 0 86480 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_932
timestamp 1649977179
transform 1 0 86848 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_937
timestamp 1649977179
transform 1 0 87308 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_945
timestamp 1649977179
transform 1 0 88044 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_951
timestamp 1649977179
transform 1 0 88596 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_956
timestamp 1649977179
transform 1 0 89056 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_968
timestamp 1649977179
transform 1 0 90160 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_980
timestamp 1649977179
transform 1 0 91264 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_992
timestamp 1649977179
transform 1 0 92368 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1004
timestamp 1649977179
transform 1 0 93472 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1009
timestamp 1649977179
transform 1 0 93932 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1021
timestamp 1649977179
transform 1 0 95036 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1033
timestamp 1649977179
transform 1 0 96140 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1045
timestamp 1649977179
transform 1 0 97244 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1057
timestamp 1649977179
transform 1 0 98348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1063
timestamp 1649977179
transform 1 0 98900 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1065
timestamp 1649977179
transform 1 0 99084 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1080
timestamp 1649977179
transform 1 0 100464 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1087
timestamp 1649977179
transform 1 0 101108 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1100
timestamp 1649977179
transform 1 0 102304 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1106
timestamp 1649977179
transform 1 0 102856 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1110
timestamp 1649977179
transform 1 0 103224 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1118
timestamp 1649977179
transform 1 0 103960 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1121
timestamp 1649977179
transform 1 0 104236 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1133
timestamp 1649977179
transform 1 0 105340 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1145
timestamp 1649977179
transform 1 0 106444 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1157
timestamp 1649977179
transform 1 0 107548 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1169
timestamp 1649977179
transform 1 0 108652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1175
timestamp 1649977179
transform 1 0 109204 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1177
timestamp 1649977179
transform 1 0 109388 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1189
timestamp 1649977179
transform 1 0 110492 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1201
timestamp 1649977179
transform 1 0 111596 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1213
timestamp 1649977179
transform 1 0 112700 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1228
timestamp 1649977179
transform 1 0 114080 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1233
timestamp 1649977179
transform 1 0 114540 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1243
timestamp 1649977179
transform 1 0 115460 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1254
timestamp 1649977179
transform 1 0 116472 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1261
timestamp 1649977179
transform 1 0 117116 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1268
timestamp 1649977179
transform 1 0 117760 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1280
timestamp 1649977179
transform 1 0 118864 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1289
timestamp 1649977179
transform 1 0 119692 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1301
timestamp 1649977179
transform 1 0 120796 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1313
timestamp 1649977179
transform 1 0 121900 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1325
timestamp 1649977179
transform 1 0 123004 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1337
timestamp 1649977179
transform 1 0 124108 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1343
timestamp 1649977179
transform 1 0 124660 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1345
timestamp 1649977179
transform 1 0 124844 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1357
timestamp 1649977179
transform 1 0 125948 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1369
timestamp 1649977179
transform 1 0 127052 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1381
timestamp 1649977179
transform 1 0 128156 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1396
timestamp 1649977179
transform 1 0 129536 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1401
timestamp 1649977179
transform 1 0 129996 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1405
timestamp 1649977179
transform 1 0 130364 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1415
timestamp 1649977179
transform 1 0 131284 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1423
timestamp 1649977179
transform 1 0 132020 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1430
timestamp 1649977179
transform 1 0 132664 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1442
timestamp 1649977179
transform 1 0 133768 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1454
timestamp 1649977179
transform 1 0 134872 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1457
timestamp 1649977179
transform 1 0 135148 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1469
timestamp 1649977179
transform 1 0 136252 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1481
timestamp 1649977179
transform 1 0 137356 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1493
timestamp 1649977179
transform 1 0 138460 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1505
timestamp 1649977179
transform 1 0 139564 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1511
timestamp 1649977179
transform 1 0 140116 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1513
timestamp 1649977179
transform 1 0 140300 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1525
timestamp 1649977179
transform 1 0 141404 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1537
timestamp 1649977179
transform 1 0 142508 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1549
timestamp 1649977179
transform 1 0 143612 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1561
timestamp 1649977179
transform 1 0 144716 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1567
timestamp 1649977179
transform 1 0 145268 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1569
timestamp 1649977179
transform 1 0 145452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1581
timestamp 1649977179
transform 1 0 146556 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_1589
timestamp 1649977179
transform 1 0 147292 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1595
timestamp 1649977179
transform 1 0 147844 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1599
timestamp 1649977179
transform 1 0 148212 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1620
timestamp 1649977179
transform 1 0 150144 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1625
timestamp 1649977179
transform 1 0 150604 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1629
timestamp 1649977179
transform 1 0 150972 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1633
timestamp 1649977179
transform 1 0 151340 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1639
timestamp 1649977179
transform 1 0 151892 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1643
timestamp 1649977179
transform 1 0 152260 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1650
timestamp 1649977179
transform 1 0 152904 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1662
timestamp 1649977179
transform 1 0 154008 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1674
timestamp 1649977179
transform 1 0 155112 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1681
timestamp 1649977179
transform 1 0 155756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1693
timestamp 1649977179
transform 1 0 156860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1705
timestamp 1649977179
transform 1 0 157964 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1717
timestamp 1649977179
transform 1 0 159068 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1729
timestamp 1649977179
transform 1 0 160172 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1735
timestamp 1649977179
transform 1 0 160724 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1740
timestamp 1649977179
transform 1 0 161184 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1747
timestamp 1649977179
transform 1 0 161828 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1754
timestamp 1649977179
transform 1 0 162472 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1761
timestamp 1649977179
transform 1 0 163116 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1768
timestamp 1649977179
transform 1 0 163760 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1775
timestamp 1649977179
transform 1 0 164404 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1782
timestamp 1649977179
transform 1 0 165048 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1790
timestamp 1649977179
transform 1 0 165784 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1793
timestamp 1649977179
transform 1 0 166060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1805
timestamp 1649977179
transform 1 0 167164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1817
timestamp 1649977179
transform 1 0 168268 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1829
timestamp 1649977179
transform 1 0 169372 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1841
timestamp 1649977179
transform 1 0 170476 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1847
timestamp 1649977179
transform 1 0 171028 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1849
timestamp 1649977179
transform 1 0 171212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1861
timestamp 1649977179
transform 1 0 172316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1873
timestamp 1649977179
transform 1 0 173420 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1885
timestamp 1649977179
transform 1 0 174524 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1897
timestamp 1649977179
transform 1 0 175628 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1903
timestamp 1649977179
transform 1 0 176180 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1905
timestamp 1649977179
transform 1 0 176364 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1909
timestamp 1649977179
transform 1 0 176732 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1917
timestamp 1649977179
transform 1 0 177468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1927
timestamp 1649977179
transform 1 0 178388 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1940
timestamp 1649977179
transform 1 0 179584 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1947
timestamp 1649977179
transform 1 0 180228 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1959
timestamp 1649977179
transform 1 0 181332 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1961
timestamp 1649977179
transform 1 0 181516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1973
timestamp 1649977179
transform 1 0 182620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1985
timestamp 1649977179
transform 1 0 183724 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1997
timestamp 1649977179
transform 1 0 184828 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_2009
timestamp 1649977179
transform 1 0 185932 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_2015
timestamp 1649977179
transform 1 0 186484 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2017
timestamp 1649977179
transform 1 0 186668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2029
timestamp 1649977179
transform 1 0 187772 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_2041
timestamp 1649977179
transform 1 0 188876 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2050
timestamp 1649977179
transform 1 0 189704 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2057
timestamp 1649977179
transform 1 0 190348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_2064
timestamp 1649977179
transform 1 0 190992 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2093
timestamp 1649977179
transform 1 0 193660 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2117
timestamp 1649977179
transform 1 0 195868 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2124
timestamp 1649977179
transform 1 0 196512 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2129
timestamp 1649977179
transform 1 0 196972 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2141
timestamp 1649977179
transform 1 0 198076 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2153
timestamp 1649977179
transform 1 0 199180 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2165
timestamp 1649977179
transform 1 0 200284 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_2177
timestamp 1649977179
transform 1 0 201388 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_2183
timestamp 1649977179
transform 1 0 201940 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_2185
timestamp 1649977179
transform 1 0 202124 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2189
timestamp 1649977179
transform 1 0 202492 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2196
timestamp 1649977179
transform 1 0 203136 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_2200
timestamp 1649977179
transform 1 0 203504 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2210
timestamp 1649977179
transform 1 0 204424 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2223
timestamp 1649977179
transform 1 0 205620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2235
timestamp 1649977179
transform 1 0 206724 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_2239
timestamp 1649977179
transform 1 0 207092 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2241
timestamp 1649977179
transform 1 0 207276 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2253
timestamp 1649977179
transform 1 0 208380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2265
timestamp 1649977179
transform 1 0 209484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2277
timestamp 1649977179
transform 1 0 210588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_2289
timestamp 1649977179
transform 1 0 211692 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_2295
timestamp 1649977179
transform 1 0 212244 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2297
timestamp 1649977179
transform 1 0 212428 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2309
timestamp 1649977179
transform 1 0 213532 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2321
timestamp 1649977179
transform 1 0 214636 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2333
timestamp 1649977179
transform 1 0 215740 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_2345
timestamp 1649977179
transform 1 0 216844 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_2351
timestamp 1649977179
transform 1 0 217396 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2353
timestamp 1649977179
transform 1 0 217580 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2365
timestamp 1649977179
transform 1 0 218684 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2377
timestamp 1649977179
transform 1 0 219788 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2389
timestamp 1649977179
transform 1 0 220892 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_2401
timestamp 1649977179
transform 1 0 221996 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_2407
timestamp 1649977179
transform 1 0 222548 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2409
timestamp 1649977179
transform 1 0 222732 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2421
timestamp 1649977179
transform 1 0 223836 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2433
timestamp 1649977179
transform 1 0 224940 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2445
timestamp 1649977179
transform 1 0 226044 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_2457
timestamp 1649977179
transform 1 0 227148 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_2463
timestamp 1649977179
transform 1 0 227700 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2474
timestamp 1649977179
transform 1 0 228712 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2487
timestamp 1649977179
transform 1 0 229908 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2494
timestamp 1649977179
transform 1 0 230552 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2501
timestamp 1649977179
transform 1 0 231196 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2508
timestamp 1649977179
transform 1 0 231840 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2521
timestamp 1649977179
transform 1 0 233036 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2533
timestamp 1649977179
transform 1 0 234140 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2545
timestamp 1649977179
transform 1 0 235244 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2557
timestamp 1649977179
transform 1 0 236348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_2569
timestamp 1649977179
transform 1 0 237452 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_2575
timestamp 1649977179
transform 1 0 238004 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2577
timestamp 1649977179
transform 1 0 238188 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_2585
timestamp 1649977179
transform 1 0 238924 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_2593
timestamp 1649977179
transform 1 0 239660 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2604
timestamp 1649977179
transform 1 0 240672 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2611
timestamp 1649977179
transform 1 0 241316 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2618
timestamp 1649977179
transform 1 0 241960 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_2625
timestamp 1649977179
transform 1 0 242604 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_2631
timestamp 1649977179
transform 1 0 243156 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2633
timestamp 1649977179
transform 1 0 243340 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2645
timestamp 1649977179
transform 1 0 244444 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2657
timestamp 1649977179
transform 1 0 245548 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2669
timestamp 1649977179
transform 1 0 246652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_2681
timestamp 1649977179
transform 1 0 247756 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_2687
timestamp 1649977179
transform 1 0 248308 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2689
timestamp 1649977179
transform 1 0 248492 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2701
timestamp 1649977179
transform 1 0 249596 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2713
timestamp 1649977179
transform 1 0 250700 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_2728
timestamp 1649977179
transform 1 0 252080 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_2732
timestamp 1649977179
transform 1 0 252448 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_2738
timestamp 1649977179
transform 1 0 253000 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2754
timestamp 1649977179
transform 1 0 254472 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2761
timestamp 1649977179
transform 1 0 255116 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2768
timestamp 1649977179
transform 1 0 255760 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2780
timestamp 1649977179
transform 1 0 256864 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_2792
timestamp 1649977179
transform 1 0 257968 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2801
timestamp 1649977179
transform 1 0 258796 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2813
timestamp 1649977179
transform 1 0 259900 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2825
timestamp 1649977179
transform 1 0 261004 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2837
timestamp 1649977179
transform 1 0 262108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_2849
timestamp 1649977179
transform 1 0 263212 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_2855
timestamp 1649977179
transform 1 0 263764 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2857
timestamp 1649977179
transform 1 0 263948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2864
timestamp 1649977179
transform 1 0 264592 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2871
timestamp 1649977179
transform 1 0 265236 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2895
timestamp 1649977179
transform 1 0 267444 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2908
timestamp 1649977179
transform 1 0 268640 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2933
timestamp 1649977179
transform 1 0 270940 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2940
timestamp 1649977179
transform 1 0 271584 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2952
timestamp 1649977179
transform 1 0 272688 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_2964
timestamp 1649977179
transform 1 0 273792 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2969
timestamp 1649977179
transform 1 0 274252 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2981
timestamp 1649977179
transform 1 0 275356 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_2993
timestamp 1649977179
transform 1 0 276460 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3005
timestamp 1649977179
transform 1 0 277564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3017
timestamp 1649977179
transform 1 0 278668 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3023
timestamp 1649977179
transform 1 0 279220 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3025
timestamp 1649977179
transform 1 0 279404 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3037
timestamp 1649977179
transform 1 0 280508 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3049
timestamp 1649977179
transform 1 0 281612 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3061
timestamp 1649977179
transform 1 0 282716 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3073
timestamp 1649977179
transform 1 0 283820 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3079
timestamp 1649977179
transform 1 0 284372 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3081
timestamp 1649977179
transform 1 0 284556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3093
timestamp 1649977179
transform 1 0 285660 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3105
timestamp 1649977179
transform 1 0 286764 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3117
timestamp 1649977179
transform 1 0 287868 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3129
timestamp 1649977179
transform 1 0 288972 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3135
timestamp 1649977179
transform 1 0 289524 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3137
timestamp 1649977179
transform 1 0 289708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3149
timestamp 1649977179
transform 1 0 290812 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3161
timestamp 1649977179
transform 1 0 291916 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3173
timestamp 1649977179
transform 1 0 293020 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3185
timestamp 1649977179
transform 1 0 294124 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3191
timestamp 1649977179
transform 1 0 294676 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3193
timestamp 1649977179
transform 1 0 294860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3205
timestamp 1649977179
transform 1 0 295964 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3217
timestamp 1649977179
transform 1 0 297068 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3229
timestamp 1649977179
transform 1 0 298172 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3241
timestamp 1649977179
transform 1 0 299276 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3247
timestamp 1649977179
transform 1 0 299828 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3249
timestamp 1649977179
transform 1 0 300012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3261
timestamp 1649977179
transform 1 0 301116 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3273
timestamp 1649977179
transform 1 0 302220 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3285
timestamp 1649977179
transform 1 0 303324 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3297
timestamp 1649977179
transform 1 0 304428 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3303
timestamp 1649977179
transform 1 0 304980 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3305
timestamp 1649977179
transform 1 0 305164 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1649977179
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1649977179
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1649977179
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1649977179
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1649977179
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1649977179
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1649977179
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1649977179
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1649977179
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_277
timestamp 1649977179
transform 1 0 26588 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_281
timestamp 1649977179
transform 1 0 26956 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_291
timestamp 1649977179
transform 1 0 27876 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_304
timestamp 1649977179
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_329
timestamp 1649977179
transform 1 0 31372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_353
timestamp 1649977179
transform 1 0 33580 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_360
timestamp 1649977179
transform 1 0 34224 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_368
timestamp 1649977179
transform 1 0 34960 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_375
timestamp 1649977179
transform 1 0 35604 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_381
timestamp 1649977179
transform 1 0 36156 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_386
timestamp 1649977179
transform 1 0 36616 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_394
timestamp 1649977179
transform 1 0 37352 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_409
timestamp 1649977179
transform 1 0 38732 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_416
timestamp 1649977179
transform 1 0 39376 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_421
timestamp 1649977179
transform 1 0 39836 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_434
timestamp 1649977179
transform 1 0 41032 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_458
timestamp 1649977179
transform 1 0 43240 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_466
timestamp 1649977179
transform 1 0 43976 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_474
timestamp 1649977179
transform 1 0 44712 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1649977179
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1649977179
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1649977179
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1649977179
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1649977179
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1649977179
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1649977179
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1649977179
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_577
timestamp 1649977179
transform 1 0 54188 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_584
timestamp 1649977179
transform 1 0 54832 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_589
timestamp 1649977179
transform 1 0 55292 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_594
timestamp 1649977179
transform 1 0 55752 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_607
timestamp 1649977179
transform 1 0 56948 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_614
timestamp 1649977179
transform 1 0 57592 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_621
timestamp 1649977179
transform 1 0 58236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_633
timestamp 1649977179
transform 1 0 59340 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_641
timestamp 1649977179
transform 1 0 60076 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_645
timestamp 1649977179
transform 1 0 60444 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_657
timestamp 1649977179
transform 1 0 61548 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_669
timestamp 1649977179
transform 1 0 62652 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_681
timestamp 1649977179
transform 1 0 63756 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_693
timestamp 1649977179
transform 1 0 64860 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_699
timestamp 1649977179
transform 1 0 65412 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_701
timestamp 1649977179
transform 1 0 65596 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_713
timestamp 1649977179
transform 1 0 66700 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_725
timestamp 1649977179
transform 1 0 67804 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_737
timestamp 1649977179
transform 1 0 68908 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_749
timestamp 1649977179
transform 1 0 70012 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_755
timestamp 1649977179
transform 1 0 70564 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_757
timestamp 1649977179
transform 1 0 70748 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_769
timestamp 1649977179
transform 1 0 71852 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_781
timestamp 1649977179
transform 1 0 72956 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_793
timestamp 1649977179
transform 1 0 74060 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_808
timestamp 1649977179
transform 1 0 75440 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_813
timestamp 1649977179
transform 1 0 75900 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_826
timestamp 1649977179
transform 1 0 77096 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_839
timestamp 1649977179
transform 1 0 78292 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_847
timestamp 1649977179
transform 1 0 79028 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_852
timestamp 1649977179
transform 1 0 79488 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_858
timestamp 1649977179
transform 1 0 80040 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_862
timestamp 1649977179
transform 1 0 80408 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_869
timestamp 1649977179
transform 1 0 81052 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_881
timestamp 1649977179
transform 1 0 82156 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_893
timestamp 1649977179
transform 1 0 83260 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_910
timestamp 1649977179
transform 1 0 84824 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_916
timestamp 1649977179
transform 1 0 85376 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_920
timestamp 1649977179
transform 1 0 85744 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_925
timestamp 1649977179
transform 1 0 86204 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_936
timestamp 1649977179
transform 1 0 87216 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_949
timestamp 1649977179
transform 1 0 88412 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_956
timestamp 1649977179
transform 1 0 89056 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_963
timestamp 1649977179
transform 1 0 89700 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_970
timestamp 1649977179
transform 1 0 90344 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_978
timestamp 1649977179
transform 1 0 91080 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_981
timestamp 1649977179
transform 1 0 91356 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_993
timestamp 1649977179
transform 1 0 92460 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1005
timestamp 1649977179
transform 1 0 93564 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1017
timestamp 1649977179
transform 1 0 94668 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1029
timestamp 1649977179
transform 1 0 95772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1035
timestamp 1649977179
transform 1 0 96324 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1037
timestamp 1649977179
transform 1 0 96508 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1049
timestamp 1649977179
transform 1 0 97612 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1061
timestamp 1649977179
transform 1 0 98716 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1068
timestamp 1649977179
transform 1 0 99360 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1075
timestamp 1649977179
transform 1 0 100004 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1088
timestamp 1649977179
transform 1 0 101200 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1093
timestamp 1649977179
transform 1 0 101660 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1099
timestamp 1649977179
transform 1 0 102212 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1112
timestamp 1649977179
transform 1 0 103408 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1119
timestamp 1649977179
transform 1 0 104052 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1126
timestamp 1649977179
transform 1 0 104696 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1133
timestamp 1649977179
transform 1 0 105340 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_1145
timestamp 1649977179
transform 1 0 106444 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1149
timestamp 1649977179
transform 1 0 106812 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1161
timestamp 1649977179
transform 1 0 107916 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1173
timestamp 1649977179
transform 1 0 109020 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1185
timestamp 1649977179
transform 1 0 110124 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1197
timestamp 1649977179
transform 1 0 111228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1203
timestamp 1649977179
transform 1 0 111780 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1205
timestamp 1649977179
transform 1 0 111964 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1220
timestamp 1649977179
transform 1 0 113344 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1227
timestamp 1649977179
transform 1 0 113988 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1251
timestamp 1649977179
transform 1 0 116196 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1259
timestamp 1649977179
transform 1 0 116932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1270
timestamp 1649977179
transform 1 0 117944 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1277
timestamp 1649977179
transform 1 0 118588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1289
timestamp 1649977179
transform 1 0 119692 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1301
timestamp 1649977179
transform 1 0 120796 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_1313
timestamp 1649977179
transform 1 0 121900 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1317
timestamp 1649977179
transform 1 0 122268 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1329
timestamp 1649977179
transform 1 0 123372 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1341
timestamp 1649977179
transform 1 0 124476 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1353
timestamp 1649977179
transform 1 0 125580 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1365
timestamp 1649977179
transform 1 0 126684 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1371
timestamp 1649977179
transform 1 0 127236 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_1373
timestamp 1649977179
transform 1 0 127420 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1379
timestamp 1649977179
transform 1 0 127972 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1383
timestamp 1649977179
transform 1 0 128340 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1387
timestamp 1649977179
transform 1 0 128708 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1411
timestamp 1649977179
transform 1 0 130916 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1424
timestamp 1649977179
transform 1 0 132112 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1432
timestamp 1649977179
transform 1 0 132848 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1444
timestamp 1649977179
transform 1 0 133952 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1456
timestamp 1649977179
transform 1 0 135056 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1468
timestamp 1649977179
transform 1 0 136160 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1480
timestamp 1649977179
transform 1 0 137264 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1491
timestamp 1649977179
transform 1 0 138276 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1503
timestamp 1649977179
transform 1 0 139380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1515
timestamp 1649977179
transform 1 0 140484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1527
timestamp 1649977179
transform 1 0 141588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1539
timestamp 1649977179
transform 1 0 142692 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1541
timestamp 1649977179
transform 1 0 142876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1553
timestamp 1649977179
transform 1 0 143980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1565
timestamp 1649977179
transform 1 0 145084 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1571
timestamp 1649977179
transform 1 0 145636 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1578
timestamp 1649977179
transform 1 0 146280 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_1586
timestamp 1649977179
transform 1 0 147016 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1592
timestamp 1649977179
transform 1 0 147568 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_1597
timestamp 1649977179
transform 1 0 148028 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1603
timestamp 1649977179
transform 1 0 148580 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1611
timestamp 1649977179
transform 1 0 149316 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1632
timestamp 1649977179
transform 1 0 151248 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1648
timestamp 1649977179
transform 1 0 152720 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1653
timestamp 1649977179
transform 1 0 153180 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1666
timestamp 1649977179
transform 1 0 154376 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1678
timestamp 1649977179
transform 1 0 155480 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1690
timestamp 1649977179
transform 1 0 156584 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1702
timestamp 1649977179
transform 1 0 157688 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1709
timestamp 1649977179
transform 1 0 158332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1721
timestamp 1649977179
transform 1 0 159436 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1730
timestamp 1649977179
transform 1 0 160264 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1745
timestamp 1649977179
transform 1 0 161644 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1758
timestamp 1649977179
transform 1 0 162840 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1765
timestamp 1649977179
transform 1 0 163484 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1786
timestamp 1649977179
transform 1 0 165416 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1794
timestamp 1649977179
transform 1 0 166152 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1806
timestamp 1649977179
transform 1 0 167256 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1818
timestamp 1649977179
transform 1 0 168360 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1821
timestamp 1649977179
transform 1 0 168636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1833
timestamp 1649977179
transform 1 0 169740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1845
timestamp 1649977179
transform 1 0 170844 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1857
timestamp 1649977179
transform 1 0 171948 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1869
timestamp 1649977179
transform 1 0 173052 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1875
timestamp 1649977179
transform 1 0 173604 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1877
timestamp 1649977179
transform 1 0 173788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1889
timestamp 1649977179
transform 1 0 174892 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_1897
timestamp 1649977179
transform 1 0 175628 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1903
timestamp 1649977179
transform 1 0 176180 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1916
timestamp 1649977179
transform 1 0 177376 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1920
timestamp 1649977179
transform 1 0 177744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1925
timestamp 1649977179
transform 1 0 178204 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1931
timestamp 1649977179
transform 1 0 178756 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1933
timestamp 1649977179
transform 1 0 178940 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1955
timestamp 1649977179
transform 1 0 180964 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1962
timestamp 1649977179
transform 1 0 181608 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1974
timestamp 1649977179
transform 1 0 182712 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1986
timestamp 1649977179
transform 1 0 183816 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1989
timestamp 1649977179
transform 1 0 184092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2001
timestamp 1649977179
transform 1 0 185196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2013
timestamp 1649977179
transform 1 0 186300 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2025
timestamp 1649977179
transform 1 0 187404 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2040
timestamp 1649977179
transform 1 0 188784 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_2045
timestamp 1649977179
transform 1 0 189244 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2051
timestamp 1649977179
transform 1 0 189796 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2058
timestamp 1649977179
transform 1 0 190440 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2082
timestamp 1649977179
transform 1 0 192648 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2095
timestamp 1649977179
transform 1 0 193844 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_2099
timestamp 1649977179
transform 1 0 194212 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_2124
timestamp 1649977179
transform 1 0 196512 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2138
timestamp 1649977179
transform 1 0 197800 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_2150
timestamp 1649977179
transform 1 0 198904 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2157
timestamp 1649977179
transform 1 0 199548 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2169
timestamp 1649977179
transform 1 0 200652 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2176
timestamp 1649977179
transform 1 0 201296 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_2183
timestamp 1649977179
transform 1 0 201940 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_2191
timestamp 1649977179
transform 1 0 202676 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_2202
timestamp 1649977179
transform 1 0 203688 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_2210
timestamp 1649977179
transform 1 0 204424 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2233
timestamp 1649977179
transform 1 0 206540 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2245
timestamp 1649977179
transform 1 0 207644 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_2257
timestamp 1649977179
transform 1 0 208748 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_2265
timestamp 1649977179
transform 1 0 209484 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2269
timestamp 1649977179
transform 1 0 209852 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2281
timestamp 1649977179
transform 1 0 210956 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2293
timestamp 1649977179
transform 1 0 212060 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2305
timestamp 1649977179
transform 1 0 213164 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_2317
timestamp 1649977179
transform 1 0 214268 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_2323
timestamp 1649977179
transform 1 0 214820 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2325
timestamp 1649977179
transform 1 0 215004 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2337
timestamp 1649977179
transform 1 0 216108 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2349
timestamp 1649977179
transform 1 0 217212 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2361
timestamp 1649977179
transform 1 0 218316 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_2373
timestamp 1649977179
transform 1 0 219420 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_2379
timestamp 1649977179
transform 1 0 219972 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2381
timestamp 1649977179
transform 1 0 220156 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2393
timestamp 1649977179
transform 1 0 221260 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2405
timestamp 1649977179
transform 1 0 222364 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2417
timestamp 1649977179
transform 1 0 223468 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_2429
timestamp 1649977179
transform 1 0 224572 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_2435
timestamp 1649977179
transform 1 0 225124 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2437
timestamp 1649977179
transform 1 0 225308 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2449
timestamp 1649977179
transform 1 0 226412 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2481
timestamp 1649977179
transform 1 0 229356 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2488
timestamp 1649977179
transform 1 0 230000 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2493
timestamp 1649977179
transform 1 0 230460 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_2497
timestamp 1649977179
transform 1 0 230828 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2507
timestamp 1649977179
transform 1 0 231748 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2514
timestamp 1649977179
transform 1 0 232392 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2526
timestamp 1649977179
transform 1 0 233496 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_2538
timestamp 1649977179
transform 1 0 234600 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_2546
timestamp 1649977179
transform 1 0 235336 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2549
timestamp 1649977179
transform 1 0 235612 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2561
timestamp 1649977179
transform 1 0 236716 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_2573
timestamp 1649977179
transform 1 0 237820 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2579
timestamp 1649977179
transform 1 0 238372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2592
timestamp 1649977179
transform 1 0 239568 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2599
timestamp 1649977179
transform 1 0 240212 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_2603
timestamp 1649977179
transform 1 0 240580 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_2605
timestamp 1649977179
transform 1 0 240764 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_2615
timestamp 1649977179
transform 1 0 241684 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_2621
timestamp 1649977179
transform 1 0 242236 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2631
timestamp 1649977179
transform 1 0 243156 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2638
timestamp 1649977179
transform 1 0 243800 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2645
timestamp 1649977179
transform 1 0 244444 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_2657
timestamp 1649977179
transform 1 0 245548 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2661
timestamp 1649977179
transform 1 0 245916 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2673
timestamp 1649977179
transform 1 0 247020 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_2685
timestamp 1649977179
transform 1 0 248124 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_2693
timestamp 1649977179
transform 1 0 248860 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2698
timestamp 1649977179
transform 1 0 249320 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_2710
timestamp 1649977179
transform 1 0 250424 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2720
timestamp 1649977179
transform 1 0 251344 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_2724
timestamp 1649977179
transform 1 0 251712 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2729
timestamp 1649977179
transform 1 0 252172 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2753
timestamp 1649977179
transform 1 0 254380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_2766
timestamp 1649977179
transform 1 0 255576 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2776
timestamp 1649977179
transform 1 0 256496 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2783
timestamp 1649977179
transform 1 0 257140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2795
timestamp 1649977179
transform 1 0 258244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2807
timestamp 1649977179
transform 1 0 259348 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_2819
timestamp 1649977179
transform 1 0 260452 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_2827
timestamp 1649977179
transform 1 0 261188 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2829
timestamp 1649977179
transform 1 0 261372 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2844
timestamp 1649977179
transform 1 0 262752 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_2856
timestamp 1649977179
transform 1 0 263856 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2860
timestamp 1649977179
transform 1 0 264224 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2867
timestamp 1649977179
transform 1 0 264868 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2880
timestamp 1649977179
transform 1 0 266064 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2905
timestamp 1649977179
transform 1 0 268364 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2929
timestamp 1649977179
transform 1 0 270572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_2936
timestamp 1649977179
transform 1 0 271216 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2950
timestamp 1649977179
transform 1 0 272504 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2962
timestamp 1649977179
transform 1 0 273608 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2974
timestamp 1649977179
transform 1 0 274712 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_2986
timestamp 1649977179
transform 1 0 275816 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_2994
timestamp 1649977179
transform 1 0 276552 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_2997
timestamp 1649977179
transform 1 0 276828 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3009
timestamp 1649977179
transform 1 0 277932 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3021
timestamp 1649977179
transform 1 0 279036 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3033
timestamp 1649977179
transform 1 0 280140 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3045
timestamp 1649977179
transform 1 0 281244 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3051
timestamp 1649977179
transform 1 0 281796 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3053
timestamp 1649977179
transform 1 0 281980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3065
timestamp 1649977179
transform 1 0 283084 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3077
timestamp 1649977179
transform 1 0 284188 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3089
timestamp 1649977179
transform 1 0 285292 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3101
timestamp 1649977179
transform 1 0 286396 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3107
timestamp 1649977179
transform 1 0 286948 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3109
timestamp 1649977179
transform 1 0 287132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3121
timestamp 1649977179
transform 1 0 288236 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3133
timestamp 1649977179
transform 1 0 289340 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3145
timestamp 1649977179
transform 1 0 290444 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3157
timestamp 1649977179
transform 1 0 291548 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3163
timestamp 1649977179
transform 1 0 292100 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3165
timestamp 1649977179
transform 1 0 292284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3177
timestamp 1649977179
transform 1 0 293388 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3189
timestamp 1649977179
transform 1 0 294492 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3201
timestamp 1649977179
transform 1 0 295596 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3213
timestamp 1649977179
transform 1 0 296700 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3219
timestamp 1649977179
transform 1 0 297252 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3221
timestamp 1649977179
transform 1 0 297436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3233
timestamp 1649977179
transform 1 0 298540 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3245
timestamp 1649977179
transform 1 0 299644 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3257
timestamp 1649977179
transform 1 0 300748 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3269
timestamp 1649977179
transform 1 0 301852 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3275
timestamp 1649977179
transform 1 0 302404 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3277
timestamp 1649977179
transform 1 0 302588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3289
timestamp 1649977179
transform 1 0 303692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3301
timestamp 1649977179
transform 1 0 304796 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1649977179
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1649977179
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1649977179
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1649977179
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1649977179
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1649977179
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1649977179
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1649977179
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_261
timestamp 1649977179
transform 1 0 25116 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_269
timestamp 1649977179
transform 1 0 25852 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_274
timestamp 1649977179
transform 1 0 26312 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_281
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_285
timestamp 1649977179
transform 1 0 27324 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_295
timestamp 1649977179
transform 1 0 28244 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_308
timestamp 1649977179
transform 1 0 29440 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_332
timestamp 1649977179
transform 1 0 31648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_357
timestamp 1649977179
transform 1 0 33948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_370
timestamp 1649977179
transform 1 0 35144 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_377
timestamp 1649977179
transform 1 0 35788 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_383
timestamp 1649977179
transform 1 0 36340 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_388
timestamp 1649977179
transform 1 0 36800 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_397
timestamp 1649977179
transform 1 0 37628 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_410
timestamp 1649977179
transform 1 0 38824 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_416
timestamp 1649977179
transform 1 0 39376 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_437
timestamp 1649977179
transform 1 0 41308 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_444
timestamp 1649977179
transform 1 0 41952 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_452
timestamp 1649977179
transform 1 0 42688 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_465
timestamp 1649977179
transform 1 0 43884 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_471
timestamp 1649977179
transform 1 0 44436 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_475
timestamp 1649977179
transform 1 0 44804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_487
timestamp 1649977179
transform 1 0 45908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_499
timestamp 1649977179
transform 1 0 47012 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1649977179
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1649977179
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1649977179
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1649977179
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1649977179
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_556
timestamp 1649977179
transform 1 0 52256 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_561
timestamp 1649977179
transform 1 0 52716 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_566
timestamp 1649977179
transform 1 0 53176 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_579
timestamp 1649977179
transform 1 0 54372 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_603
timestamp 1649977179
transform 1 0 56580 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_611
timestamp 1649977179
transform 1 0 57316 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1649977179
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_617
timestamp 1649977179
transform 1 0 57868 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_629
timestamp 1649977179
transform 1 0 58972 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_641
timestamp 1649977179
transform 1 0 60076 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_653
timestamp 1649977179
transform 1 0 61180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_665
timestamp 1649977179
transform 1 0 62284 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_671
timestamp 1649977179
transform 1 0 62836 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_673
timestamp 1649977179
transform 1 0 63020 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_685
timestamp 1649977179
transform 1 0 64124 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_697
timestamp 1649977179
transform 1 0 65228 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_709
timestamp 1649977179
transform 1 0 66332 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_721
timestamp 1649977179
transform 1 0 67436 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_727
timestamp 1649977179
transform 1 0 67988 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_729
timestamp 1649977179
transform 1 0 68172 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_741
timestamp 1649977179
transform 1 0 69276 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_753
timestamp 1649977179
transform 1 0 70380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_765
timestamp 1649977179
transform 1 0 71484 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_771
timestamp 1649977179
transform 1 0 72036 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_775
timestamp 1649977179
transform 1 0 72404 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_783
timestamp 1649977179
transform 1 0 73140 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_785
timestamp 1649977179
transform 1 0 73324 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_797
timestamp 1649977179
transform 1 0 74428 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_801
timestamp 1649977179
transform 1 0 74796 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_805
timestamp 1649977179
transform 1 0 75164 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_829
timestamp 1649977179
transform 1 0 77372 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_836
timestamp 1649977179
transform 1 0 78016 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_844
timestamp 1649977179
transform 1 0 78752 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_851
timestamp 1649977179
transform 1 0 79396 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_875
timestamp 1649977179
transform 1 0 81604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_887
timestamp 1649977179
transform 1 0 82708 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_895
timestamp 1649977179
transform 1 0 83444 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_897
timestamp 1649977179
transform 1 0 83628 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_921
timestamp 1649977179
transform 1 0 85836 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_945
timestamp 1649977179
transform 1 0 88044 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_951
timestamp 1649977179
transform 1 0 88596 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_953
timestamp 1649977179
transform 1 0 88780 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_966
timestamp 1649977179
transform 1 0 89976 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_974
timestamp 1649977179
transform 1 0 90712 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_981
timestamp 1649977179
transform 1 0 91356 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_993
timestamp 1649977179
transform 1 0 92460 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_1005
timestamp 1649977179
transform 1 0 93564 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1009
timestamp 1649977179
transform 1 0 93932 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1021
timestamp 1649977179
transform 1 0 95036 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1033
timestamp 1649977179
transform 1 0 96140 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1045
timestamp 1649977179
transform 1 0 97244 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1060
timestamp 1649977179
transform 1 0 98624 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1065
timestamp 1649977179
transform 1 0 99084 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1086
timestamp 1649977179
transform 1 0 101016 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1110
timestamp 1649977179
transform 1 0 103224 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1118
timestamp 1649977179
transform 1 0 103960 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1130
timestamp 1649977179
transform 1 0 105064 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1138
timestamp 1649977179
transform 1 0 105800 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1142
timestamp 1649977179
transform 1 0 106168 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1154
timestamp 1649977179
transform 1 0 107272 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1166
timestamp 1649977179
transform 1 0 108376 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1174
timestamp 1649977179
transform 1 0 109112 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1177
timestamp 1649977179
transform 1 0 109388 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1189
timestamp 1649977179
transform 1 0 110492 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_1201
timestamp 1649977179
transform 1 0 111596 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1213
timestamp 1649977179
transform 1 0 112700 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1220
timestamp 1649977179
transform 1 0 113344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1228
timestamp 1649977179
transform 1 0 114080 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1237
timestamp 1649977179
transform 1 0 114908 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1250
timestamp 1649977179
transform 1 0 116104 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1274
timestamp 1649977179
transform 1 0 118312 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1281
timestamp 1649977179
transform 1 0 118956 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1287
timestamp 1649977179
transform 1 0 119508 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1289
timestamp 1649977179
transform 1 0 119692 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1301
timestamp 1649977179
transform 1 0 120796 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1313
timestamp 1649977179
transform 1 0 121900 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1325
timestamp 1649977179
transform 1 0 123004 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1337
timestamp 1649977179
transform 1 0 124108 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1343
timestamp 1649977179
transform 1 0 124660 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1345
timestamp 1649977179
transform 1 0 124844 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1357
timestamp 1649977179
transform 1 0 125948 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1368
timestamp 1649977179
transform 1 0 126960 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1376
timestamp 1649977179
transform 1 0 127696 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1383
timestamp 1649977179
transform 1 0 128340 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1396
timestamp 1649977179
transform 1 0 129536 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1401
timestamp 1649977179
transform 1 0 129996 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1406
timestamp 1649977179
transform 1 0 130456 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1430
timestamp 1649977179
transform 1 0 132664 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1434
timestamp 1649977179
transform 1 0 133032 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1444
timestamp 1649977179
transform 1 0 133952 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1451
timestamp 1649977179
transform 1 0 134596 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1455
timestamp 1649977179
transform 1 0 134964 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1457
timestamp 1649977179
transform 1 0 135148 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1463
timestamp 1649977179
transform 1 0 135700 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1475
timestamp 1649977179
transform 1 0 136804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1487
timestamp 1649977179
transform 1 0 137908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1499
timestamp 1649977179
transform 1 0 139012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1511
timestamp 1649977179
transform 1 0 140116 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1513
timestamp 1649977179
transform 1 0 140300 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1525
timestamp 1649977179
transform 1 0 141404 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1537
timestamp 1649977179
transform 1 0 142508 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1541
timestamp 1649977179
transform 1 0 142876 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1548
timestamp 1649977179
transform 1 0 143520 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1560
timestamp 1649977179
transform 1 0 144624 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1578
timestamp 1649977179
transform 1 0 146280 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1587
timestamp 1649977179
transform 1 0 147108 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1611
timestamp 1649977179
transform 1 0 149316 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1620
timestamp 1649977179
transform 1 0 150144 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1625
timestamp 1649977179
transform 1 0 150604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1629
timestamp 1649977179
transform 1 0 150972 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1639
timestamp 1649977179
transform 1 0 151892 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1645
timestamp 1649977179
transform 1 0 152444 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1649
timestamp 1649977179
transform 1 0 152812 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1653
timestamp 1649977179
transform 1 0 153180 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1657
timestamp 1649977179
transform 1 0 153548 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1661
timestamp 1649977179
transform 1 0 153916 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1665
timestamp 1649977179
transform 1 0 154284 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1676
timestamp 1649977179
transform 1 0 155296 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1681
timestamp 1649977179
transform 1 0 155756 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1685
timestamp 1649977179
transform 1 0 156124 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1689
timestamp 1649977179
transform 1 0 156492 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1693
timestamp 1649977179
transform 1 0 156860 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1697
timestamp 1649977179
transform 1 0 157228 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1709
timestamp 1649977179
transform 1 0 158332 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1713
timestamp 1649977179
transform 1 0 158700 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1723
timestamp 1649977179
transform 1 0 159620 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1731
timestamp 1649977179
transform 1 0 160356 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1735
timestamp 1649977179
transform 1 0 160724 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1737
timestamp 1649977179
transform 1 0 160908 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1743
timestamp 1649977179
transform 1 0 161460 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1767
timestamp 1649977179
transform 1 0 163668 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1780
timestamp 1649977179
transform 1 0 164864 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1788
timestamp 1649977179
transform 1 0 165600 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1793
timestamp 1649977179
transform 1 0 166060 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1801
timestamp 1649977179
transform 1 0 166796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1808
timestamp 1649977179
transform 1 0 167440 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1815
timestamp 1649977179
transform 1 0 168084 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1827
timestamp 1649977179
transform 1 0 169188 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1839
timestamp 1649977179
transform 1 0 170292 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1847
timestamp 1649977179
transform 1 0 171028 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1849
timestamp 1649977179
transform 1 0 171212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1861
timestamp 1649977179
transform 1 0 172316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1873
timestamp 1649977179
transform 1 0 173420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1885
timestamp 1649977179
transform 1 0 174524 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1889
timestamp 1649977179
transform 1 0 174892 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1893
timestamp 1649977179
transform 1 0 175260 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1900
timestamp 1649977179
transform 1 0 175904 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1925
timestamp 1649977179
transform 1 0 178204 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1949
timestamp 1649977179
transform 1 0 180412 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1956
timestamp 1649977179
transform 1 0 181056 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1964
timestamp 1649977179
transform 1 0 181792 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1971
timestamp 1649977179
transform 1 0 182436 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1983
timestamp 1649977179
transform 1 0 183540 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1995
timestamp 1649977179
transform 1 0 184644 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_2007
timestamp 1649977179
transform 1 0 185748 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_2015
timestamp 1649977179
transform 1 0 186484 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2017
timestamp 1649977179
transform 1 0 186668 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_2029
timestamp 1649977179
transform 1 0 187772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2033
timestamp 1649977179
transform 1 0 188140 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2041
timestamp 1649977179
transform 1 0 188876 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_2049
timestamp 1649977179
transform 1 0 189612 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_2057
timestamp 1649977179
transform 1 0 190348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2068
timestamp 1649977179
transform 1 0 191360 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2082
timestamp 1649977179
transform 1 0 192648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2109
timestamp 1649977179
transform 1 0 195132 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_2122
timestamp 1649977179
transform 1 0 196328 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_2138
timestamp 1649977179
transform 1 0 197800 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2145
timestamp 1649977179
transform 1 0 198444 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_2157
timestamp 1649977179
transform 1 0 199548 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_2165
timestamp 1649977179
transform 1 0 200284 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2170
timestamp 1649977179
transform 1 0 200744 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_2177
timestamp 1649977179
transform 1 0 201388 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_2183
timestamp 1649977179
transform 1 0 201940 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2185
timestamp 1649977179
transform 1 0 202124 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_2189
timestamp 1649977179
transform 1 0 202492 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2210
timestamp 1649977179
transform 1 0 204424 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_2234
timestamp 1649977179
transform 1 0 206632 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2244
timestamp 1649977179
transform 1 0 207552 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2256
timestamp 1649977179
transform 1 0 208656 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2268
timestamp 1649977179
transform 1 0 209760 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2280
timestamp 1649977179
transform 1 0 210864 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2292
timestamp 1649977179
transform 1 0 211968 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2297
timestamp 1649977179
transform 1 0 212428 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2309
timestamp 1649977179
transform 1 0 213532 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2321
timestamp 1649977179
transform 1 0 214636 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2333
timestamp 1649977179
transform 1 0 215740 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_2345
timestamp 1649977179
transform 1 0 216844 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_2351
timestamp 1649977179
transform 1 0 217396 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2353
timestamp 1649977179
transform 1 0 217580 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2365
timestamp 1649977179
transform 1 0 218684 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2377
timestamp 1649977179
transform 1 0 219788 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2389
timestamp 1649977179
transform 1 0 220892 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_2401
timestamp 1649977179
transform 1 0 221996 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_2407
timestamp 1649977179
transform 1 0 222548 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2409
timestamp 1649977179
transform 1 0 222732 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2421
timestamp 1649977179
transform 1 0 223836 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2433
timestamp 1649977179
transform 1 0 224940 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2445
timestamp 1649977179
transform 1 0 226044 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_2449
timestamp 1649977179
transform 1 0 226412 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2453
timestamp 1649977179
transform 1 0 226780 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2460
timestamp 1649977179
transform 1 0 227424 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2485
timestamp 1649977179
transform 1 0 229724 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2492
timestamp 1649977179
transform 1 0 230368 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2516
timestamp 1649977179
transform 1 0 232576 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2524
timestamp 1649977179
transform 1 0 233312 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2536
timestamp 1649977179
transform 1 0 234416 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2548
timestamp 1649977179
transform 1 0 235520 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_2560
timestamp 1649977179
transform 1 0 236624 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2565
timestamp 1649977179
transform 1 0 237084 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2572
timestamp 1649977179
transform 1 0 237728 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_2577
timestamp 1649977179
transform 1 0 238188 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2600
timestamp 1649977179
transform 1 0 240304 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_2624
timestamp 1649977179
transform 1 0 242512 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2633
timestamp 1649977179
transform 1 0 243340 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2641
timestamp 1649977179
transform 1 0 244076 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2649
timestamp 1649977179
transform 1 0 244812 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2656
timestamp 1649977179
transform 1 0 245456 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2668
timestamp 1649977179
transform 1 0 246560 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_2680
timestamp 1649977179
transform 1 0 247664 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2689
timestamp 1649977179
transform 1 0 248492 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_2701
timestamp 1649977179
transform 1 0 249596 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_2710
timestamp 1649977179
transform 1 0 250424 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_2718
timestamp 1649977179
transform 1 0 251160 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2723
timestamp 1649977179
transform 1 0 251620 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_2736
timestamp 1649977179
transform 1 0 252816 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2765
timestamp 1649977179
transform 1 0 255484 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2778
timestamp 1649977179
transform 1 0 256680 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2785
timestamp 1649977179
transform 1 0 257324 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_2797
timestamp 1649977179
transform 1 0 258428 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2801
timestamp 1649977179
transform 1 0 258796 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2813
timestamp 1649977179
transform 1 0 259900 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_2825
timestamp 1649977179
transform 1 0 261004 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_2831
timestamp 1649977179
transform 1 0 261556 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2836
timestamp 1649977179
transform 1 0 262016 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2844
timestamp 1649977179
transform 1 0 262752 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2852
timestamp 1649977179
transform 1 0 263488 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2860
timestamp 1649977179
transform 1 0 264224 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2867
timestamp 1649977179
transform 1 0 264868 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2891
timestamp 1649977179
transform 1 0 267076 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_2904
timestamp 1649977179
transform 1 0 268272 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2933
timestamp 1649977179
transform 1 0 270940 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_2946
timestamp 1649977179
transform 1 0 272136 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_2959
timestamp 1649977179
transform 1 0 273332 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_2967
timestamp 1649977179
transform 1 0 274068 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2969
timestamp 1649977179
transform 1 0 274252 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2981
timestamp 1649977179
transform 1 0 275356 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_2993
timestamp 1649977179
transform 1 0 276460 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3005
timestamp 1649977179
transform 1 0 277564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3017
timestamp 1649977179
transform 1 0 278668 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3023
timestamp 1649977179
transform 1 0 279220 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3025
timestamp 1649977179
transform 1 0 279404 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3037
timestamp 1649977179
transform 1 0 280508 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3049
timestamp 1649977179
transform 1 0 281612 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3061
timestamp 1649977179
transform 1 0 282716 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3073
timestamp 1649977179
transform 1 0 283820 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3079
timestamp 1649977179
transform 1 0 284372 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3081
timestamp 1649977179
transform 1 0 284556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3093
timestamp 1649977179
transform 1 0 285660 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3105
timestamp 1649977179
transform 1 0 286764 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3117
timestamp 1649977179
transform 1 0 287868 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3129
timestamp 1649977179
transform 1 0 288972 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3135
timestamp 1649977179
transform 1 0 289524 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3137
timestamp 1649977179
transform 1 0 289708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3149
timestamp 1649977179
transform 1 0 290812 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3161
timestamp 1649977179
transform 1 0 291916 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3173
timestamp 1649977179
transform 1 0 293020 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3185
timestamp 1649977179
transform 1 0 294124 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3191
timestamp 1649977179
transform 1 0 294676 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3193
timestamp 1649977179
transform 1 0 294860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3205
timestamp 1649977179
transform 1 0 295964 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3217
timestamp 1649977179
transform 1 0 297068 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3229
timestamp 1649977179
transform 1 0 298172 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3241
timestamp 1649977179
transform 1 0 299276 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3247
timestamp 1649977179
transform 1 0 299828 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3249
timestamp 1649977179
transform 1 0 300012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3261
timestamp 1649977179
transform 1 0 301116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3273
timestamp 1649977179
transform 1 0 302220 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3280
timestamp 1649977179
transform 1 0 302864 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3292
timestamp 1649977179
transform 1 0 303968 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3296
timestamp 1649977179
transform 1 0 304336 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3300
timestamp 1649977179
transform 1 0 304704 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3305
timestamp 1649977179
transform 1 0 305164 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_8
timestamp 1649977179
transform 1 0 1840 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp 1649977179
transform 1 0 2944 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_37
timestamp 1649977179
transform 1 0 4508 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_57
timestamp 1649977179
transform 1 0 6348 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_69
timestamp 1649977179
transform 1 0 7452 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_74
timestamp 1649977179
transform 1 0 7912 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1649977179
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_108
timestamp 1649977179
transform 1 0 11040 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_113
timestamp 1649977179
transform 1 0 11500 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_125
timestamp 1649977179
transform 1 0 12604 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_137
timestamp 1649977179
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_144
timestamp 1649977179
transform 1 0 14352 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_156
timestamp 1649977179
transform 1 0 15456 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_169
timestamp 1649977179
transform 1 0 16652 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_174
timestamp 1649977179
transform 1 0 17112 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_186
timestamp 1649977179
transform 1 0 18216 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1649977179
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_208
timestamp 1649977179
transform 1 0 20240 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_220
timestamp 1649977179
transform 1 0 21344 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_225
timestamp 1649977179
transform 1 0 21804 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_237
timestamp 1649977179
transform 1 0 22908 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_241
timestamp 1649977179
transform 1 0 23276 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_249
timestamp 1649977179
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_265
timestamp 1649977179
transform 1 0 25484 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_276
timestamp 1649977179
transform 1 0 26496 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_281
timestamp 1649977179
transform 1 0 26956 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_304
timestamp 1649977179
transform 1 0 29072 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_309
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_332
timestamp 1649977179
transform 1 0 31648 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_337
timestamp 1649977179
transform 1 0 32108 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_360
timestamp 1649977179
transform 1 0 34224 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_385
timestamp 1649977179
transform 1 0 36524 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_391
timestamp 1649977179
transform 1 0 37076 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_393
timestamp 1649977179
transform 1 0 37260 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_416
timestamp 1649977179
transform 1 0 39376 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_421
timestamp 1649977179
transform 1 0 39836 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_444
timestamp 1649977179
transform 1 0 41952 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_449
timestamp 1649977179
transform 1 0 42412 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_470
timestamp 1649977179
transform 1 0 44344 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_486
timestamp 1649977179
transform 1 0 45816 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_498
timestamp 1649977179
transform 1 0 46920 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_508
timestamp 1649977179
transform 1 0 47840 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_520
timestamp 1649977179
transform 1 0 48944 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_533
timestamp 1649977179
transform 1 0 50140 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_538
timestamp 1649977179
transform 1 0 50600 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_551
timestamp 1649977179
transform 1 0 51796 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_559
timestamp 1649977179
transform 1 0 52532 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_561
timestamp 1649977179
transform 1 0 52716 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_584
timestamp 1649977179
transform 1 0 54832 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_589
timestamp 1649977179
transform 1 0 55292 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_612
timestamp 1649977179
transform 1 0 57408 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_637
timestamp 1649977179
transform 1 0 59708 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_643
timestamp 1649977179
transform 1 0 60260 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_648
timestamp 1649977179
transform 1 0 60720 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_660
timestamp 1649977179
transform 1 0 61824 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_676
timestamp 1649977179
transform 1 0 63296 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_688
timestamp 1649977179
transform 1 0 64400 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_701
timestamp 1649977179
transform 1 0 65596 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_708
timestamp 1649977179
transform 1 0 66240 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_720
timestamp 1649977179
transform 1 0 67344 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_729
timestamp 1649977179
transform 1 0 68172 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_737
timestamp 1649977179
transform 1 0 68908 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_742
timestamp 1649977179
transform 1 0 69368 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_754
timestamp 1649977179
transform 1 0 70472 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_757
timestamp 1649977179
transform 1 0 70748 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_769
timestamp 1649977179
transform 1 0 71852 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_780
timestamp 1649977179
transform 1 0 72864 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_785
timestamp 1649977179
transform 1 0 73324 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_808
timestamp 1649977179
transform 1 0 75440 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_813
timestamp 1649977179
transform 1 0 75900 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_836
timestamp 1649977179
transform 1 0 78016 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_861
timestamp 1649977179
transform 1 0 80316 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_867
timestamp 1649977179
transform 1 0 80868 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_878
timestamp 1649977179
transform 1 0 81880 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_885
timestamp 1649977179
transform 1 0 82524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_892
timestamp 1649977179
transform 1 0 83168 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_897
timestamp 1649977179
transform 1 0 83628 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_920
timestamp 1649977179
transform 1 0 85744 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_925
timestamp 1649977179
transform 1 0 86204 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_948
timestamp 1649977179
transform 1 0 88320 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_973
timestamp 1649977179
transform 1 0 90620 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_979
timestamp 1649977179
transform 1 0 91172 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_981
timestamp 1649977179
transform 1 0 91356 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_989
timestamp 1649977179
transform 1 0 92092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1001
timestamp 1649977179
transform 1 0 93196 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1007
timestamp 1649977179
transform 1 0 93748 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1012
timestamp 1649977179
transform 1 0 94208 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1024
timestamp 1649977179
transform 1 0 95312 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1037
timestamp 1649977179
transform 1 0 96508 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1042
timestamp 1649977179
transform 1 0 96968 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1057
timestamp 1649977179
transform 1 0 98348 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1063
timestamp 1649977179
transform 1 0 98900 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1065
timestamp 1649977179
transform 1 0 99084 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1088
timestamp 1649977179
transform 1 0 101200 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1093
timestamp 1649977179
transform 1 0 101660 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1116
timestamp 1649977179
transform 1 0 103776 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1141
timestamp 1649977179
transform 1 0 106076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1147
timestamp 1649977179
transform 1 0 106628 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1149
timestamp 1649977179
transform 1 0 106812 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1161
timestamp 1649977179
transform 1 0 107916 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1173
timestamp 1649977179
transform 1 0 109020 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1180
timestamp 1649977179
transform 1 0 109664 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1192
timestamp 1649977179
transform 1 0 110768 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1196
timestamp 1649977179
transform 1 0 111136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1200
timestamp 1649977179
transform 1 0 111504 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1205
timestamp 1649977179
transform 1 0 111964 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1228
timestamp 1649977179
transform 1 0 114080 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1233
timestamp 1649977179
transform 1 0 114540 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1256
timestamp 1649977179
transform 1 0 116656 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1261
timestamp 1649977179
transform 1 0 117116 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1284
timestamp 1649977179
transform 1 0 119232 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1298
timestamp 1649977179
transform 1 0 120520 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1309
timestamp 1649977179
transform 1 0 121532 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1315
timestamp 1649977179
transform 1 0 122084 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1317
timestamp 1649977179
transform 1 0 122268 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1329
timestamp 1649977179
transform 1 0 123372 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1340
timestamp 1649977179
transform 1 0 124384 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1345
timestamp 1649977179
transform 1 0 124844 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1355
timestamp 1649977179
transform 1 0 125764 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1368
timestamp 1649977179
transform 1 0 126960 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1373
timestamp 1649977179
transform 1 0 127420 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1394
timestamp 1649977179
transform 1 0 129352 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1401
timestamp 1649977179
transform 1 0 129996 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1424
timestamp 1649977179
transform 1 0 132112 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1449
timestamp 1649977179
transform 1 0 134412 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1455
timestamp 1649977179
transform 1 0 134964 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1457
timestamp 1649977179
transform 1 0 135148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1469
timestamp 1649977179
transform 1 0 136252 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1476
timestamp 1649977179
transform 1 0 136896 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1485
timestamp 1649977179
transform 1 0 137724 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1497
timestamp 1649977179
transform 1 0 138828 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1509
timestamp 1649977179
transform 1 0 139932 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1516
timestamp 1649977179
transform 1 0 140576 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1528
timestamp 1649977179
transform 1 0 141680 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1544
timestamp 1649977179
transform 1 0 143152 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1556
timestamp 1649977179
transform 1 0 144256 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1560
timestamp 1649977179
transform 1 0 144624 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1564
timestamp 1649977179
transform 1 0 144992 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1569
timestamp 1649977179
transform 1 0 145452 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1592
timestamp 1649977179
transform 1 0 147568 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1620
timestamp 1649977179
transform 1 0 150144 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1625
timestamp 1649977179
transform 1 0 150604 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1648
timestamp 1649977179
transform 1 0 152720 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1653
timestamp 1649977179
transform 1 0 153180 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1676
timestamp 1649977179
transform 1 0 155296 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1684
timestamp 1649977179
transform 1 0 156032 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1691
timestamp 1649977179
transform 1 0 156676 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1699
timestamp 1649977179
transform 1 0 157412 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1704
timestamp 1649977179
transform 1 0 157872 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1709
timestamp 1649977179
transform 1 0 158332 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1732
timestamp 1649977179
transform 1 0 160448 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1757
timestamp 1649977179
transform 1 0 162748 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1763
timestamp 1649977179
transform 1 0 163300 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1785
timestamp 1649977179
transform 1 0 165324 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1791
timestamp 1649977179
transform 1 0 165876 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1802
timestamp 1649977179
transform 1 0 166888 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1810
timestamp 1649977179
transform 1 0 167624 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1818
timestamp 1649977179
transform 1 0 168360 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1821
timestamp 1649977179
transform 1 0 168636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1833
timestamp 1649977179
transform 1 0 169740 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1839
timestamp 1649977179
transform 1 0 170292 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1843
timestamp 1649977179
transform 1 0 170660 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1847
timestamp 1649977179
transform 1 0 171028 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1849
timestamp 1649977179
transform 1 0 171212 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1861
timestamp 1649977179
transform 1 0 172316 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1872
timestamp 1649977179
transform 1 0 173328 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1886
timestamp 1649977179
transform 1 0 174616 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1894
timestamp 1649977179
transform 1 0 175352 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1900
timestamp 1649977179
transform 1 0 175904 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1925
timestamp 1649977179
transform 1 0 178204 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1931
timestamp 1649977179
transform 1 0 178756 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1953
timestamp 1649977179
transform 1 0 180780 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1959
timestamp 1649977179
transform 1 0 181332 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1970
timestamp 1649977179
transform 1 0 182344 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1977
timestamp 1649977179
transform 1 0 182988 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1985
timestamp 1649977179
transform 1 0 183724 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1989
timestamp 1649977179
transform 1 0 184092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2001
timestamp 1649977179
transform 1 0 185196 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2010
timestamp 1649977179
transform 1 0 186024 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2017
timestamp 1649977179
transform 1 0 186668 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2023
timestamp 1649977179
transform 1 0 187220 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2027
timestamp 1649977179
transform 1 0 187588 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2040
timestamp 1649977179
transform 1 0 188784 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_2045
timestamp 1649977179
transform 1 0 189244 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2068
timestamp 1649977179
transform 1 0 191360 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2096
timestamp 1649977179
transform 1 0 193936 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2124
timestamp 1649977179
transform 1 0 196512 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_2129
timestamp 1649977179
transform 1 0 196972 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2137
timestamp 1649977179
transform 1 0 197708 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_2140
timestamp 1649977179
transform 1 0 197984 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2151
timestamp 1649977179
transform 1 0 198996 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2155
timestamp 1649977179
transform 1 0 199364 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_2157
timestamp 1649977179
transform 1 0 199548 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2163
timestamp 1649977179
transform 1 0 200100 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_2176
timestamp 1649977179
transform 1 0 201296 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2205
timestamp 1649977179
transform 1 0 203964 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2211
timestamp 1649977179
transform 1 0 204516 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2233
timestamp 1649977179
transform 1 0 206540 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2239
timestamp 1649977179
transform 1 0 207092 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_2250
timestamp 1649977179
transform 1 0 208104 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2262
timestamp 1649977179
transform 1 0 209208 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2269
timestamp 1649977179
transform 1 0 209852 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2273
timestamp 1649977179
transform 1 0 210220 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_2277
timestamp 1649977179
transform 1 0 210588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2289
timestamp 1649977179
transform 1 0 211692 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2295
timestamp 1649977179
transform 1 0 212244 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_2297
timestamp 1649977179
transform 1 0 212428 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_2305
timestamp 1649977179
transform 1 0 213164 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_2310
timestamp 1649977179
transform 1 0 213624 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_2322
timestamp 1649977179
transform 1 0 214728 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_2325
timestamp 1649977179
transform 1 0 215004 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_2337
timestamp 1649977179
transform 1 0 216108 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_2343
timestamp 1649977179
transform 1 0 216660 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2351
timestamp 1649977179
transform 1 0 217396 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_2353
timestamp 1649977179
transform 1 0 217580 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_2365
timestamp 1649977179
transform 1 0 218684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_2377
timestamp 1649977179
transform 1 0 219788 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_2384
timestamp 1649977179
transform 1 0 220432 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_2396
timestamp 1649977179
transform 1 0 221536 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2412
timestamp 1649977179
transform 1 0 223008 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2418
timestamp 1649977179
transform 1 0 223560 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_2428
timestamp 1649977179
transform 1 0 224480 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2437
timestamp 1649977179
transform 1 0 225308 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2444
timestamp 1649977179
transform 1 0 225952 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2450
timestamp 1649977179
transform 1 0 226504 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2460
timestamp 1649977179
transform 1 0 227424 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2485
timestamp 1649977179
transform 1 0 229724 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2491
timestamp 1649977179
transform 1 0 230276 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2513
timestamp 1649977179
transform 1 0 232300 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2519
timestamp 1649977179
transform 1 0 232852 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2524
timestamp 1649977179
transform 1 0 233312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_2531
timestamp 1649977179
transform 1 0 233956 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_2539
timestamp 1649977179
transform 1 0 234692 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2544
timestamp 1649977179
transform 1 0 235152 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_2549
timestamp 1649977179
transform 1 0 235612 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2570
timestamp 1649977179
transform 1 0 237544 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2597
timestamp 1649977179
transform 1 0 240028 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2603
timestamp 1649977179
transform 1 0 240580 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2625
timestamp 1649977179
transform 1 0 242604 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2631
timestamp 1649977179
transform 1 0 243156 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2653
timestamp 1649977179
transform 1 0 245180 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2659
timestamp 1649977179
transform 1 0 245732 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_2661
timestamp 1649977179
transform 1 0 245916 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2673
timestamp 1649977179
transform 1 0 247020 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_2677
timestamp 1649977179
transform 1 0 247388 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_2685
timestamp 1649977179
transform 1 0 248124 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_2689
timestamp 1649977179
transform 1 0 248492 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_2697
timestamp 1649977179
transform 1 0 249228 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2709
timestamp 1649977179
transform 1 0 250332 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2715
timestamp 1649977179
transform 1 0 250884 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2737
timestamp 1649977179
transform 1 0 252908 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2743
timestamp 1649977179
transform 1 0 253460 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2765
timestamp 1649977179
transform 1 0 255484 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2771
timestamp 1649977179
transform 1 0 256036 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2793
timestamp 1649977179
transform 1 0 258060 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2799
timestamp 1649977179
transform 1 0 258612 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2801
timestamp 1649977179
transform 1 0 258796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2807
timestamp 1649977179
transform 1 0 259348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_2811
timestamp 1649977179
transform 1 0 259716 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2823
timestamp 1649977179
transform 1 0 260820 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2827
timestamp 1649977179
transform 1 0 261188 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2829
timestamp 1649977179
transform 1 0 261372 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2837
timestamp 1649977179
transform 1 0 262108 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2852
timestamp 1649977179
transform 1 0 263488 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_2857
timestamp 1649977179
transform 1 0 263948 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2880
timestamp 1649977179
transform 1 0 266064 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2908
timestamp 1649977179
transform 1 0 268640 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2933
timestamp 1649977179
transform 1 0 270940 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2939
timestamp 1649977179
transform 1 0 271492 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_2961
timestamp 1649977179
transform 1 0 273516 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2967
timestamp 1649977179
transform 1 0 274068 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2972
timestamp 1649977179
transform 1 0 274528 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_2979
timestamp 1649977179
transform 1 0 275172 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_2991
timestamp 1649977179
transform 1 0 276276 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_2995
timestamp 1649977179
transform 1 0 276644 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_2997
timestamp 1649977179
transform 1 0 276828 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3005
timestamp 1649977179
transform 1 0 277564 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3011
timestamp 1649977179
transform 1 0 278116 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3023
timestamp 1649977179
transform 1 0 279220 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3025
timestamp 1649977179
transform 1 0 279404 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3037
timestamp 1649977179
transform 1 0 280508 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3044
timestamp 1649977179
transform 1 0 281152 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3053
timestamp 1649977179
transform 1 0 281980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3065
timestamp 1649977179
transform 1 0 283084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3077
timestamp 1649977179
transform 1 0 284188 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3084
timestamp 1649977179
transform 1 0 284832 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3096
timestamp 1649977179
transform 1 0 285936 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3112
timestamp 1649977179
transform 1 0 287408 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3124
timestamp 1649977179
transform 1 0 288512 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3137
timestamp 1649977179
transform 1 0 289708 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3144
timestamp 1649977179
transform 1 0 290352 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3156
timestamp 1649977179
transform 1 0 291456 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3165
timestamp 1649977179
transform 1 0 292284 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3173
timestamp 1649977179
transform 1 0 293020 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3178
timestamp 1649977179
transform 1 0 293480 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3190
timestamp 1649977179
transform 1 0 294584 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3193
timestamp 1649977179
transform 1 0 294860 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3201
timestamp 1649977179
transform 1 0 295596 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3206
timestamp 1649977179
transform 1 0 296056 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3211
timestamp 1649977179
transform 1 0 296516 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3219
timestamp 1649977179
transform 1 0 297252 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3221
timestamp 1649977179
transform 1 0 297436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3233
timestamp 1649977179
transform 1 0 298540 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3244
timestamp 1649977179
transform 1 0 299552 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3249
timestamp 1649977179
transform 1 0 300012 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3261
timestamp 1649977179
transform 1 0 301116 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3266
timestamp 1649977179
transform 1 0 301576 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3270
timestamp 1649977179
transform 1 0 301944 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3274
timestamp 1649977179
transform 1 0 302312 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3277
timestamp 1649977179
transform 1 0 302588 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3283
timestamp 1649977179
transform 1 0 303140 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3287
timestamp 1649977179
transform 1 0 303508 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3300
timestamp 1649977179
transform 1 0 304704 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3305
timestamp 1649977179
transform 1 0 305164 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 305808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 305808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 305808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 305808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 305808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 305808 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 305808 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 305808 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 305808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 305808 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 305808 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 305808 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 305808 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 305808 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 305808 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 305808 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 305808 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 305808 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 305808 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 305808 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 305808 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1649977179
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1649977179
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1649977179
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1649977179
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1649977179
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1649977179
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1649977179
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1649977179
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1649977179
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1649977179
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1649977179
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1649977179
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1649977179
transform 1 0 70656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 73232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 75808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 78384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 80960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 83536 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 86112 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 88688 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 91264 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 93840 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 96416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 98992 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 101568 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 104144 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 106720 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 109296 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 111872 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 114448 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 117024 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 119600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 122176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 124752 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 127328 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 129904 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 132480 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 135056 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 137632 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 140208 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 142784 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 145360 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 147936 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 150512 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 153088 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 155664 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 158240 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 160816 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 163392 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 165968 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 168544 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 171120 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 173696 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 176272 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 178848 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 181424 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 184000 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 186576 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 189152 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 191728 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 194304 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 196880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 199456 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 202032 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 204608 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 207184 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 209760 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 212336 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 214912 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 217488 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 220064 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 222640 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 225216 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 227792 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 230368 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 232944 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 235520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 238096 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 240672 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 243248 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 245824 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 248400 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 250976 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 253552 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 256128 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 258704 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 261280 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 263856 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 266432 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 269008 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 271584 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 274160 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 276736 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 279312 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 281888 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 284464 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 287040 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 289616 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 292192 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 294768 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 297344 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 299920 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 302496 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 305072 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 73232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 78384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 83536 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 88688 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 93840 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 98992 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 104144 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 109296 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 114448 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 119600 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 124752 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 129904 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 135056 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 140208 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 145360 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 150512 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 155664 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 160816 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 165968 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 171120 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 176272 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1649977179
transform 1 0 181424 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1649977179
transform 1 0 186576 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1649977179
transform 1 0 191728 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1649977179
transform 1 0 196880 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1649977179
transform 1 0 202032 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1649977179
transform 1 0 207184 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1649977179
transform 1 0 212336 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1649977179
transform 1 0 217488 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1649977179
transform 1 0 222640 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1649977179
transform 1 0 227792 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1649977179
transform 1 0 232944 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 238096 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 243248 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 248400 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 253552 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 258704 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 263856 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 269008 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 274160 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 279312 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 284464 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 289616 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 294768 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 299920 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 305072 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 70656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 75808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 80960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 86112 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 91264 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 96416 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 101568 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 106720 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 111872 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 117024 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 122176 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 127328 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 132480 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 137632 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 142784 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 147936 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 153088 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 158240 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 163392 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 168544 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 173696 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 178848 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 184000 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 189152 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 194304 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 199456 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 204608 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 209760 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 214912 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 220064 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 225216 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 230368 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 235520 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 240672 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 245824 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 250976 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 256128 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 261280 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 266432 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 271584 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 276736 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 281888 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 287040 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 292192 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 297344 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 302496 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 73232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 78384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 83536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 88688 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 93840 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 98992 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 104144 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 109296 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 114448 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 119600 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 124752 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 129904 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 135056 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 140208 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 145360 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 150512 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 155664 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 160816 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 165968 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 171120 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 176272 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 181424 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 186576 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 191728 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 196880 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 202032 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 207184 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 212336 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 217488 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 222640 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 227792 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 232944 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 238096 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 243248 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 248400 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 253552 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 258704 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 263856 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 269008 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 274160 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 279312 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 284464 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 289616 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 294768 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 299920 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 305072 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 70656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 75808 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 80960 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 86112 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 91264 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 96416 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 101568 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 106720 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 111872 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 117024 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 122176 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 127328 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 132480 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 137632 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 142784 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 147936 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 153088 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 158240 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 163392 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 168544 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 173696 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 178848 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 184000 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 189152 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 194304 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 199456 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 204608 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 209760 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 214912 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 220064 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 225216 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 230368 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 235520 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 240672 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 245824 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 250976 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 256128 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 261280 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 266432 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 271584 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 276736 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 281888 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 287040 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 292192 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 297344 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 302496 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 73232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 78384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 83536 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 88688 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 93840 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 98992 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 104144 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 109296 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 114448 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 119600 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 124752 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 129904 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 135056 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 140208 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 145360 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 150512 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 155664 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 160816 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 165968 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 171120 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 176272 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 181424 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 186576 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 191728 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 196880 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 202032 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 207184 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 212336 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 217488 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 222640 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 227792 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 232944 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 238096 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 243248 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 248400 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 253552 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 258704 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 263856 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 269008 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 274160 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 279312 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 284464 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 289616 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 294768 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 299920 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 305072 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 70656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 75808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 80960 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 86112 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 91264 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 96416 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 101568 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 106720 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 111872 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 117024 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 122176 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 127328 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 132480 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 137632 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 142784 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 147936 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 153088 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 158240 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 163392 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 168544 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 173696 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 178848 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 184000 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 189152 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 194304 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 199456 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 204608 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 209760 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 214912 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 220064 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 225216 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 230368 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 235520 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 240672 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 245824 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 250976 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 256128 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 261280 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 266432 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 271584 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 276736 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 281888 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 287040 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 292192 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 297344 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 302496 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 73232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 78384 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 83536 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 88688 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 93840 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 98992 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 104144 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 109296 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 114448 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1649977179
transform 1 0 119600 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1649977179
transform 1 0 124752 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1649977179
transform 1 0 129904 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1649977179
transform 1 0 135056 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1649977179
transform 1 0 140208 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1649977179
transform 1 0 145360 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1649977179
transform 1 0 150512 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1649977179
transform 1 0 155664 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1649977179
transform 1 0 160816 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1649977179
transform 1 0 165968 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1649977179
transform 1 0 171120 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1649977179
transform 1 0 176272 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1649977179
transform 1 0 181424 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1649977179
transform 1 0 186576 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1649977179
transform 1 0 191728 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1649977179
transform 1 0 196880 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1649977179
transform 1 0 202032 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1649977179
transform 1 0 207184 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1649977179
transform 1 0 212336 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1649977179
transform 1 0 217488 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1649977179
transform 1 0 222640 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1649977179
transform 1 0 227792 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1649977179
transform 1 0 232944 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1649977179
transform 1 0 238096 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1649977179
transform 1 0 243248 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1649977179
transform 1 0 248400 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1649977179
transform 1 0 253552 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1649977179
transform 1 0 258704 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1649977179
transform 1 0 263856 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1649977179
transform 1 0 269008 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1649977179
transform 1 0 274160 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1649977179
transform 1 0 279312 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1649977179
transform 1 0 284464 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1649977179
transform 1 0 289616 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1649977179
transform 1 0 294768 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1649977179
transform 1 0 299920 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1649977179
transform 1 0 305072 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1649977179
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1649977179
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1649977179
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1649977179
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1649977179
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1649977179
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1649977179
transform 1 0 70656 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1649977179
transform 1 0 75808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1649977179
transform 1 0 80960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1649977179
transform 1 0 86112 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1649977179
transform 1 0 91264 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1649977179
transform 1 0 96416 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1649977179
transform 1 0 101568 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1649977179
transform 1 0 106720 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1649977179
transform 1 0 111872 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1649977179
transform 1 0 117024 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1649977179
transform 1 0 122176 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1649977179
transform 1 0 127328 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1649977179
transform 1 0 132480 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1649977179
transform 1 0 137632 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1649977179
transform 1 0 142784 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1649977179
transform 1 0 147936 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1649977179
transform 1 0 153088 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1649977179
transform 1 0 158240 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1649977179
transform 1 0 163392 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1649977179
transform 1 0 168544 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1649977179
transform 1 0 173696 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1649977179
transform 1 0 178848 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1649977179
transform 1 0 184000 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1649977179
transform 1 0 189152 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1649977179
transform 1 0 194304 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1649977179
transform 1 0 199456 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1649977179
transform 1 0 204608 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1649977179
transform 1 0 209760 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1649977179
transform 1 0 214912 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1649977179
transform 1 0 220064 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1649977179
transform 1 0 225216 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1649977179
transform 1 0 230368 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1649977179
transform 1 0 235520 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1649977179
transform 1 0 240672 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1649977179
transform 1 0 245824 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1649977179
transform 1 0 250976 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1649977179
transform 1 0 256128 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1649977179
transform 1 0 261280 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1649977179
transform 1 0 266432 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1649977179
transform 1 0 271584 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1649977179
transform 1 0 276736 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1649977179
transform 1 0 281888 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1649977179
transform 1 0 287040 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1649977179
transform 1 0 292192 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1649977179
transform 1 0 297344 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1649977179
transform 1 0 302496 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1649977179
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1649977179
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1649977179
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1649977179
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1649977179
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1649977179
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1649977179
transform 1 0 73232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1649977179
transform 1 0 78384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1649977179
transform 1 0 83536 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1649977179
transform 1 0 88688 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1649977179
transform 1 0 93840 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1649977179
transform 1 0 98992 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1649977179
transform 1 0 104144 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1649977179
transform 1 0 109296 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1649977179
transform 1 0 114448 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1649977179
transform 1 0 119600 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1649977179
transform 1 0 124752 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1649977179
transform 1 0 129904 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1649977179
transform 1 0 135056 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1649977179
transform 1 0 140208 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1649977179
transform 1 0 145360 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1649977179
transform 1 0 150512 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1649977179
transform 1 0 155664 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1649977179
transform 1 0 160816 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1649977179
transform 1 0 165968 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1649977179
transform 1 0 171120 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1649977179
transform 1 0 176272 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1649977179
transform 1 0 181424 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1649977179
transform 1 0 186576 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1649977179
transform 1 0 191728 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1649977179
transform 1 0 196880 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1649977179
transform 1 0 202032 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1649977179
transform 1 0 207184 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1649977179
transform 1 0 212336 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1649977179
transform 1 0 217488 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1649977179
transform 1 0 222640 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1649977179
transform 1 0 227792 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1649977179
transform 1 0 232944 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1649977179
transform 1 0 238096 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1649977179
transform 1 0 243248 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1649977179
transform 1 0 248400 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1649977179
transform 1 0 253552 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1649977179
transform 1 0 258704 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1649977179
transform 1 0 263856 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1649977179
transform 1 0 269008 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1649977179
transform 1 0 274160 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1649977179
transform 1 0 279312 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1649977179
transform 1 0 284464 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1649977179
transform 1 0 289616 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1649977179
transform 1 0 294768 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1649977179
transform 1 0 299920 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1649977179
transform 1 0 305072 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1649977179
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1649977179
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1649977179
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1649977179
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1649977179
transform 1 0 60352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1649977179
transform 1 0 65504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1649977179
transform 1 0 70656 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1649977179
transform 1 0 75808 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1649977179
transform 1 0 80960 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1649977179
transform 1 0 86112 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1649977179
transform 1 0 91264 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1649977179
transform 1 0 96416 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1649977179
transform 1 0 101568 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1649977179
transform 1 0 106720 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1649977179
transform 1 0 111872 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1649977179
transform 1 0 117024 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1649977179
transform 1 0 122176 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1649977179
transform 1 0 127328 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1649977179
transform 1 0 132480 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1649977179
transform 1 0 137632 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1649977179
transform 1 0 142784 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1649977179
transform 1 0 147936 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1649977179
transform 1 0 153088 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1649977179
transform 1 0 158240 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1649977179
transform 1 0 163392 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1649977179
transform 1 0 168544 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1649977179
transform 1 0 173696 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1649977179
transform 1 0 178848 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1649977179
transform 1 0 184000 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1649977179
transform 1 0 189152 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1649977179
transform 1 0 194304 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1649977179
transform 1 0 199456 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1649977179
transform 1 0 204608 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1649977179
transform 1 0 209760 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1649977179
transform 1 0 214912 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1649977179
transform 1 0 220064 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1649977179
transform 1 0 225216 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1649977179
transform 1 0 230368 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1649977179
transform 1 0 235520 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1649977179
transform 1 0 240672 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1649977179
transform 1 0 245824 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1649977179
transform 1 0 250976 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1649977179
transform 1 0 256128 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1649977179
transform 1 0 261280 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1649977179
transform 1 0 266432 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1649977179
transform 1 0 271584 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1649977179
transform 1 0 276736 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1649977179
transform 1 0 281888 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1649977179
transform 1 0 287040 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1649977179
transform 1 0 292192 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1649977179
transform 1 0 297344 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1649977179
transform 1 0 302496 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1649977179
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1649977179
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1649977179
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1649977179
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1649977179
transform 1 0 62928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1649977179
transform 1 0 68080 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1649977179
transform 1 0 73232 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1649977179
transform 1 0 78384 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1649977179
transform 1 0 83536 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1649977179
transform 1 0 88688 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1649977179
transform 1 0 93840 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1649977179
transform 1 0 98992 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1649977179
transform 1 0 104144 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1649977179
transform 1 0 109296 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1649977179
transform 1 0 114448 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1649977179
transform 1 0 119600 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1649977179
transform 1 0 124752 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1649977179
transform 1 0 129904 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1649977179
transform 1 0 135056 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1649977179
transform 1 0 140208 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1649977179
transform 1 0 145360 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1649977179
transform 1 0 150512 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1649977179
transform 1 0 155664 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1649977179
transform 1 0 160816 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1649977179
transform 1 0 165968 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1649977179
transform 1 0 171120 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1649977179
transform 1 0 176272 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1649977179
transform 1 0 181424 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1649977179
transform 1 0 186576 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1649977179
transform 1 0 191728 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1649977179
transform 1 0 196880 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1649977179
transform 1 0 202032 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1649977179
transform 1 0 207184 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1649977179
transform 1 0 212336 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1649977179
transform 1 0 217488 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1649977179
transform 1 0 222640 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1649977179
transform 1 0 227792 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1649977179
transform 1 0 232944 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1649977179
transform 1 0 238096 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1649977179
transform 1 0 243248 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1649977179
transform 1 0 248400 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1649977179
transform 1 0 253552 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1649977179
transform 1 0 258704 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1649977179
transform 1 0 263856 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1649977179
transform 1 0 269008 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1649977179
transform 1 0 274160 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1649977179
transform 1 0 279312 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1649977179
transform 1 0 284464 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1649977179
transform 1 0 289616 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1649977179
transform 1 0 294768 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1649977179
transform 1 0 299920 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1649977179
transform 1 0 305072 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1649977179
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1649977179
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1649977179
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1649977179
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1649977179
transform 1 0 60352 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1649977179
transform 1 0 65504 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1649977179
transform 1 0 70656 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1649977179
transform 1 0 75808 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1649977179
transform 1 0 80960 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1649977179
transform 1 0 86112 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1649977179
transform 1 0 91264 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1649977179
transform 1 0 96416 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1649977179
transform 1 0 101568 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1649977179
transform 1 0 106720 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1649977179
transform 1 0 111872 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1649977179
transform 1 0 117024 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1649977179
transform 1 0 122176 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1649977179
transform 1 0 127328 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1649977179
transform 1 0 132480 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1649977179
transform 1 0 137632 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1649977179
transform 1 0 142784 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1649977179
transform 1 0 147936 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1649977179
transform 1 0 153088 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1649977179
transform 1 0 158240 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1649977179
transform 1 0 163392 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1649977179
transform 1 0 168544 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1649977179
transform 1 0 173696 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1649977179
transform 1 0 178848 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1649977179
transform 1 0 184000 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1649977179
transform 1 0 189152 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1649977179
transform 1 0 194304 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1649977179
transform 1 0 199456 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1649977179
transform 1 0 204608 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1649977179
transform 1 0 209760 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1649977179
transform 1 0 214912 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1649977179
transform 1 0 220064 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1649977179
transform 1 0 225216 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1649977179
transform 1 0 230368 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1649977179
transform 1 0 235520 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1649977179
transform 1 0 240672 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1649977179
transform 1 0 245824 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1649977179
transform 1 0 250976 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1649977179
transform 1 0 256128 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1649977179
transform 1 0 261280 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1649977179
transform 1 0 266432 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1649977179
transform 1 0 271584 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1649977179
transform 1 0 276736 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1649977179
transform 1 0 281888 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1649977179
transform 1 0 287040 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1649977179
transform 1 0 292192 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1649977179
transform 1 0 297344 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1649977179
transform 1 0 302496 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1649977179
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1649977179
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1649977179
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1649977179
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1649977179
transform 1 0 62928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1649977179
transform 1 0 68080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1649977179
transform 1 0 73232 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1649977179
transform 1 0 78384 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1649977179
transform 1 0 83536 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1649977179
transform 1 0 88688 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1649977179
transform 1 0 93840 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1649977179
transform 1 0 98992 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1649977179
transform 1 0 104144 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1649977179
transform 1 0 109296 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1649977179
transform 1 0 114448 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1649977179
transform 1 0 119600 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1649977179
transform 1 0 124752 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1649977179
transform 1 0 129904 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1649977179
transform 1 0 135056 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1649977179
transform 1 0 140208 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1649977179
transform 1 0 145360 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1649977179
transform 1 0 150512 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1649977179
transform 1 0 155664 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1649977179
transform 1 0 160816 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1649977179
transform 1 0 165968 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1649977179
transform 1 0 171120 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1649977179
transform 1 0 176272 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1649977179
transform 1 0 181424 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1649977179
transform 1 0 186576 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1649977179
transform 1 0 191728 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1649977179
transform 1 0 196880 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1649977179
transform 1 0 202032 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1649977179
transform 1 0 207184 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1649977179
transform 1 0 212336 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1649977179
transform 1 0 217488 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1649977179
transform 1 0 222640 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1649977179
transform 1 0 227792 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1649977179
transform 1 0 232944 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1649977179
transform 1 0 238096 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1649977179
transform 1 0 243248 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1649977179
transform 1 0 248400 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1649977179
transform 1 0 253552 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1649977179
transform 1 0 258704 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1649977179
transform 1 0 263856 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1649977179
transform 1 0 269008 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1649977179
transform 1 0 274160 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1649977179
transform 1 0 279312 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1649977179
transform 1 0 284464 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1649977179
transform 1 0 289616 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1649977179
transform 1 0 294768 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1649977179
transform 1 0 299920 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1649977179
transform 1 0 305072 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1649977179
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1649977179
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1649977179
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1649977179
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1649977179
transform 1 0 60352 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1649977179
transform 1 0 65504 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1649977179
transform 1 0 70656 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1649977179
transform 1 0 75808 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1649977179
transform 1 0 80960 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1649977179
transform 1 0 86112 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1649977179
transform 1 0 91264 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1649977179
transform 1 0 96416 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1649977179
transform 1 0 101568 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1649977179
transform 1 0 106720 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1649977179
transform 1 0 111872 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1649977179
transform 1 0 117024 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1649977179
transform 1 0 122176 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1649977179
transform 1 0 127328 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1649977179
transform 1 0 132480 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1649977179
transform 1 0 137632 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1649977179
transform 1 0 142784 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1649977179
transform 1 0 147936 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1649977179
transform 1 0 153088 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1649977179
transform 1 0 158240 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1649977179
transform 1 0 163392 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1649977179
transform 1 0 168544 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1649977179
transform 1 0 173696 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1649977179
transform 1 0 178848 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1649977179
transform 1 0 184000 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1649977179
transform 1 0 189152 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1649977179
transform 1 0 194304 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1649977179
transform 1 0 199456 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1649977179
transform 1 0 204608 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1649977179
transform 1 0 209760 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1649977179
transform 1 0 214912 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1649977179
transform 1 0 220064 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1649977179
transform 1 0 225216 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1649977179
transform 1 0 230368 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1649977179
transform 1 0 235520 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1649977179
transform 1 0 240672 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1649977179
transform 1 0 245824 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1649977179
transform 1 0 250976 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1649977179
transform 1 0 256128 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1649977179
transform 1 0 261280 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1649977179
transform 1 0 266432 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1649977179
transform 1 0 271584 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1649977179
transform 1 0 276736 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1649977179
transform 1 0 281888 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1649977179
transform 1 0 287040 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1649977179
transform 1 0 292192 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1649977179
transform 1 0 297344 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1649977179
transform 1 0 302496 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1649977179
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1649977179
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1649977179
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1649977179
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1649977179
transform 1 0 62928 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1649977179
transform 1 0 68080 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1649977179
transform 1 0 73232 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1649977179
transform 1 0 78384 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1649977179
transform 1 0 83536 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1649977179
transform 1 0 88688 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1649977179
transform 1 0 93840 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1649977179
transform 1 0 98992 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1649977179
transform 1 0 104144 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1649977179
transform 1 0 109296 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1649977179
transform 1 0 114448 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1649977179
transform 1 0 119600 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1649977179
transform 1 0 124752 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1649977179
transform 1 0 129904 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1649977179
transform 1 0 135056 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1649977179
transform 1 0 140208 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1649977179
transform 1 0 145360 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1649977179
transform 1 0 150512 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1649977179
transform 1 0 155664 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1649977179
transform 1 0 160816 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1649977179
transform 1 0 165968 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1649977179
transform 1 0 171120 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1649977179
transform 1 0 176272 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1649977179
transform 1 0 181424 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1649977179
transform 1 0 186576 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1649977179
transform 1 0 191728 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1649977179
transform 1 0 196880 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1649977179
transform 1 0 202032 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1649977179
transform 1 0 207184 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1649977179
transform 1 0 212336 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1649977179
transform 1 0 217488 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1649977179
transform 1 0 222640 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1649977179
transform 1 0 227792 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1649977179
transform 1 0 232944 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1649977179
transform 1 0 238096 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1649977179
transform 1 0 243248 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1649977179
transform 1 0 248400 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1649977179
transform 1 0 253552 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1649977179
transform 1 0 258704 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1649977179
transform 1 0 263856 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1649977179
transform 1 0 269008 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1649977179
transform 1 0 274160 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1649977179
transform 1 0 279312 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1649977179
transform 1 0 284464 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1649977179
transform 1 0 289616 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1649977179
transform 1 0 294768 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1649977179
transform 1 0 299920 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1649977179
transform 1 0 305072 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1649977179
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1649977179
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1649977179
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1649977179
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1649977179
transform 1 0 60352 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1649977179
transform 1 0 65504 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1649977179
transform 1 0 70656 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1649977179
transform 1 0 75808 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1649977179
transform 1 0 80960 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1649977179
transform 1 0 86112 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1649977179
transform 1 0 91264 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1649977179
transform 1 0 96416 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1649977179
transform 1 0 101568 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1649977179
transform 1 0 106720 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1649977179
transform 1 0 111872 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1649977179
transform 1 0 117024 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1649977179
transform 1 0 122176 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1649977179
transform 1 0 127328 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1649977179
transform 1 0 132480 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1649977179
transform 1 0 137632 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1649977179
transform 1 0 142784 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1649977179
transform 1 0 147936 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1649977179
transform 1 0 153088 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1649977179
transform 1 0 158240 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1649977179
transform 1 0 163392 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1649977179
transform 1 0 168544 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1649977179
transform 1 0 173696 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1649977179
transform 1 0 178848 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1649977179
transform 1 0 184000 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1649977179
transform 1 0 189152 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1649977179
transform 1 0 194304 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1649977179
transform 1 0 199456 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1649977179
transform 1 0 204608 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1649977179
transform 1 0 209760 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1649977179
transform 1 0 214912 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1649977179
transform 1 0 220064 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1649977179
transform 1 0 225216 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1649977179
transform 1 0 230368 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1649977179
transform 1 0 235520 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1649977179
transform 1 0 240672 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1649977179
transform 1 0 245824 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1649977179
transform 1 0 250976 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1649977179
transform 1 0 256128 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1649977179
transform 1 0 261280 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1649977179
transform 1 0 266432 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1649977179
transform 1 0 271584 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1649977179
transform 1 0 276736 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1649977179
transform 1 0 281888 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1649977179
transform 1 0 287040 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1649977179
transform 1 0 292192 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1649977179
transform 1 0 297344 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1649977179
transform 1 0 302496 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1649977179
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1649977179
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1649977179
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1649977179
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1649977179
transform 1 0 62928 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1649977179
transform 1 0 68080 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1649977179
transform 1 0 73232 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1649977179
transform 1 0 78384 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1649977179
transform 1 0 83536 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1649977179
transform 1 0 88688 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1649977179
transform 1 0 93840 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1649977179
transform 1 0 98992 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1649977179
transform 1 0 104144 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1649977179
transform 1 0 109296 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1649977179
transform 1 0 114448 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1649977179
transform 1 0 119600 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1649977179
transform 1 0 124752 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1649977179
transform 1 0 129904 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1649977179
transform 1 0 135056 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1649977179
transform 1 0 140208 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1649977179
transform 1 0 145360 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1649977179
transform 1 0 150512 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1649977179
transform 1 0 155664 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1649977179
transform 1 0 160816 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1649977179
transform 1 0 165968 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1649977179
transform 1 0 171120 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1649977179
transform 1 0 176272 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1649977179
transform 1 0 181424 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1649977179
transform 1 0 186576 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1649977179
transform 1 0 191728 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1649977179
transform 1 0 196880 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1649977179
transform 1 0 202032 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1649977179
transform 1 0 207184 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1649977179
transform 1 0 212336 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1649977179
transform 1 0 217488 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1649977179
transform 1 0 222640 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1649977179
transform 1 0 227792 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1649977179
transform 1 0 232944 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1649977179
transform 1 0 238096 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1649977179
transform 1 0 243248 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1649977179
transform 1 0 248400 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1649977179
transform 1 0 253552 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1649977179
transform 1 0 258704 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1649977179
transform 1 0 263856 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1649977179
transform 1 0 269008 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1649977179
transform 1 0 274160 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1649977179
transform 1 0 279312 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1649977179
transform 1 0 284464 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1649977179
transform 1 0 289616 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1649977179
transform 1 0 294768 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1649977179
transform 1 0 299920 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1649977179
transform 1 0 305072 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1649977179
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1649977179
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1649977179
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1649977179
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1649977179
transform 1 0 60352 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1649977179
transform 1 0 65504 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1649977179
transform 1 0 70656 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1649977179
transform 1 0 75808 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1649977179
transform 1 0 80960 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1649977179
transform 1 0 86112 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1649977179
transform 1 0 91264 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1649977179
transform 1 0 96416 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1649977179
transform 1 0 101568 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1649977179
transform 1 0 106720 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1649977179
transform 1 0 111872 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1649977179
transform 1 0 117024 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1649977179
transform 1 0 122176 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1649977179
transform 1 0 127328 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1649977179
transform 1 0 132480 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1649977179
transform 1 0 137632 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1649977179
transform 1 0 142784 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1649977179
transform 1 0 147936 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1649977179
transform 1 0 153088 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1649977179
transform 1 0 158240 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1649977179
transform 1 0 163392 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1649977179
transform 1 0 168544 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1649977179
transform 1 0 173696 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1649977179
transform 1 0 178848 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1649977179
transform 1 0 184000 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1649977179
transform 1 0 189152 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1649977179
transform 1 0 194304 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1649977179
transform 1 0 199456 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1649977179
transform 1 0 204608 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1649977179
transform 1 0 209760 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1649977179
transform 1 0 214912 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1649977179
transform 1 0 220064 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1649977179
transform 1 0 225216 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1649977179
transform 1 0 230368 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1649977179
transform 1 0 235520 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1649977179
transform 1 0 240672 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1649977179
transform 1 0 245824 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1649977179
transform 1 0 250976 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1649977179
transform 1 0 256128 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1649977179
transform 1 0 261280 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1649977179
transform 1 0 266432 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1649977179
transform 1 0 271584 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1649977179
transform 1 0 276736 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1649977179
transform 1 0 281888 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1649977179
transform 1 0 287040 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1649977179
transform 1 0 292192 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1649977179
transform 1 0 297344 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1649977179
transform 1 0 302496 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1649977179
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1649977179
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1649977179
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1649977179
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1649977179
transform 1 0 62928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1649977179
transform 1 0 68080 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1649977179
transform 1 0 73232 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1649977179
transform 1 0 78384 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1649977179
transform 1 0 83536 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1649977179
transform 1 0 88688 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1649977179
transform 1 0 93840 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1649977179
transform 1 0 98992 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1649977179
transform 1 0 104144 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1649977179
transform 1 0 109296 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1649977179
transform 1 0 114448 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1649977179
transform 1 0 119600 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1649977179
transform 1 0 124752 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1649977179
transform 1 0 129904 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1649977179
transform 1 0 135056 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1649977179
transform 1 0 140208 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1649977179
transform 1 0 145360 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1649977179
transform 1 0 150512 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1649977179
transform 1 0 155664 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1649977179
transform 1 0 160816 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1649977179
transform 1 0 165968 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1649977179
transform 1 0 171120 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1649977179
transform 1 0 176272 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1649977179
transform 1 0 181424 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1649977179
transform 1 0 186576 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1649977179
transform 1 0 191728 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1649977179
transform 1 0 196880 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1649977179
transform 1 0 202032 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1649977179
transform 1 0 207184 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1649977179
transform 1 0 212336 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1649977179
transform 1 0 217488 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1649977179
transform 1 0 222640 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1649977179
transform 1 0 227792 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1649977179
transform 1 0 232944 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1649977179
transform 1 0 238096 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1649977179
transform 1 0 243248 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1649977179
transform 1 0 248400 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1649977179
transform 1 0 253552 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1649977179
transform 1 0 258704 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1649977179
transform 1 0 263856 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1649977179
transform 1 0 269008 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1649977179
transform 1 0 274160 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1649977179
transform 1 0 279312 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1649977179
transform 1 0 284464 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1649977179
transform 1 0 289616 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1649977179
transform 1 0 294768 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1649977179
transform 1 0 299920 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1649977179
transform 1 0 305072 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1649977179
transform 1 0 6256 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1649977179
transform 1 0 11408 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1649977179
transform 1 0 16560 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1649977179
transform 1 0 21712 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1649977179
transform 1 0 26864 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1649977179
transform 1 0 32016 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1649977179
transform 1 0 37168 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1649977179
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1649977179
transform 1 0 42320 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1649977179
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1649977179
transform 1 0 47472 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1649977179
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1649977179
transform 1 0 52624 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1649977179
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1649977179
transform 1 0 57776 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1649977179
transform 1 0 60352 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1649977179
transform 1 0 62928 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1649977179
transform 1 0 65504 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1649977179
transform 1 0 68080 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1649977179
transform 1 0 70656 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1649977179
transform 1 0 73232 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1649977179
transform 1 0 75808 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1649977179
transform 1 0 78384 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1649977179
transform 1 0 80960 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1649977179
transform 1 0 83536 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1649977179
transform 1 0 86112 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1649977179
transform 1 0 88688 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1649977179
transform 1 0 91264 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1649977179
transform 1 0 93840 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1649977179
transform 1 0 96416 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1649977179
transform 1 0 98992 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1649977179
transform 1 0 101568 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1649977179
transform 1 0 104144 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1649977179
transform 1 0 106720 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1649977179
transform 1 0 109296 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1649977179
transform 1 0 111872 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1649977179
transform 1 0 114448 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1649977179
transform 1 0 117024 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1649977179
transform 1 0 119600 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1649977179
transform 1 0 122176 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1649977179
transform 1 0 124752 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1649977179
transform 1 0 127328 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1649977179
transform 1 0 129904 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1649977179
transform 1 0 132480 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1649977179
transform 1 0 135056 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1649977179
transform 1 0 137632 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1649977179
transform 1 0 140208 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1649977179
transform 1 0 142784 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1649977179
transform 1 0 145360 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1649977179
transform 1 0 147936 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1649977179
transform 1 0 150512 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1649977179
transform 1 0 153088 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1649977179
transform 1 0 155664 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1649977179
transform 1 0 158240 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1649977179
transform 1 0 160816 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1649977179
transform 1 0 163392 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1649977179
transform 1 0 165968 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1649977179
transform 1 0 168544 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1649977179
transform 1 0 171120 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1649977179
transform 1 0 173696 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1649977179
transform 1 0 176272 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1649977179
transform 1 0 178848 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1649977179
transform 1 0 181424 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1649977179
transform 1 0 184000 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1649977179
transform 1 0 186576 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1649977179
transform 1 0 189152 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1649977179
transform 1 0 191728 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1649977179
transform 1 0 194304 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1649977179
transform 1 0 196880 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1649977179
transform 1 0 199456 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1649977179
transform 1 0 202032 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1649977179
transform 1 0 204608 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1649977179
transform 1 0 207184 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1649977179
transform 1 0 209760 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1649977179
transform 1 0 212336 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1649977179
transform 1 0 214912 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1649977179
transform 1 0 217488 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1649977179
transform 1 0 220064 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1649977179
transform 1 0 222640 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1649977179
transform 1 0 225216 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1649977179
transform 1 0 227792 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1649977179
transform 1 0 230368 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1649977179
transform 1 0 232944 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1649977179
transform 1 0 235520 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1649977179
transform 1 0 238096 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1649977179
transform 1 0 240672 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1649977179
transform 1 0 243248 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1649977179
transform 1 0 245824 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1649977179
transform 1 0 248400 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1649977179
transform 1 0 250976 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1649977179
transform 1 0 253552 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1649977179
transform 1 0 256128 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1649977179
transform 1 0 258704 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1649977179
transform 1 0 261280 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1649977179
transform 1 0 263856 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1649977179
transform 1 0 266432 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1649977179
transform 1 0 269008 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1649977179
transform 1 0 271584 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1649977179
transform 1 0 274160 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1649977179
transform 1 0 276736 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1649977179
transform 1 0 279312 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1649977179
transform 1 0 281888 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1649977179
transform 1 0 284464 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1649977179
transform 1 0 287040 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1649977179
transform 1 0 289616 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1649977179
transform 1 0 292192 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1649977179
transform 1 0 294768 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1649977179
transform 1 0 297344 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1649977179
transform 1 0 299920 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1649977179
transform 1 0 302496 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1649977179
transform 1 0 305072 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  _348_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 137724 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _349_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 56948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _350_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 58144 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _351_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 56212 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _352_
timestamp 1649977179
transform 1 0 56120 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _353_
timestamp 1649977179
transform 1 0 57960 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _354_
timestamp 1649977179
transform 1 0 54924 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _355_
timestamp 1649977179
transform 1 0 55292 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _356_
timestamp 1649977179
transform 1 0 53544 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _357_
timestamp 1649977179
transform 1 0 51980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _358_
timestamp 1649977179
transform 1 0 50968 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _359_
timestamp 1649977179
transform 1 0 52808 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _360_
timestamp 1649977179
transform 1 0 43608 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _361_
timestamp 1649977179
transform 1 0 43056 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _362_
timestamp 1649977179
transform 1 0 41676 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _363_
timestamp 1649977179
transform 1 0 44988 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _364_
timestamp 1649977179
transform 1 0 41584 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _365_
timestamp 1649977179
transform 1 0 40204 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _366_
timestamp 1649977179
transform 1 0 40296 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _367_
timestamp 1649977179
transform 1 0 39652 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _368_
timestamp 1649977179
transform 1 0 39008 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _369_
timestamp 1649977179
transform 1 0 37996 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _370_
timestamp 1649977179
transform 1 0 38456 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _371_
timestamp 1649977179
transform 1 0 36984 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _372_
timestamp 1649977179
transform 1 0 34316 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _373_
timestamp 1649977179
transform 1 0 33948 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _374_
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _375_
timestamp 1649977179
transform 1 0 32752 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _376_
timestamp 1649977179
transform 1 0 31832 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _377_
timestamp 1649977179
transform 1 0 33396 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _378_
timestamp 1649977179
transform 1 0 28612 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _379_
timestamp 1649977179
transform 1 0 34960 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _380_
timestamp 1649977179
transform 1 0 30268 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _381_
timestamp 1649977179
transform 1 0 32108 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _382_
timestamp 1649977179
transform 1 0 36248 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _383_
timestamp 1649977179
transform 1 0 28244 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _384_
timestamp 1649977179
transform 1 0 30912 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _385_
timestamp 1649977179
transform 1 0 28428 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _386_
timestamp 1649977179
transform 1 0 29624 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _387_
timestamp 1649977179
transform 1 0 25668 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _388_
timestamp 1649977179
transform 1 0 28796 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _389_
timestamp 1649977179
transform 1 0 27048 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _390_
timestamp 1649977179
transform 1 0 30268 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _391_
timestamp 1649977179
transform 1 0 27416 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _392_
timestamp 1649977179
transform 1 0 31096 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _393_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 145728 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _394_
timestamp 1649977179
transform 1 0 154468 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _395_
timestamp 1649977179
transform 1 0 150788 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _396_
timestamp 1649977179
transform 1 0 195500 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _397_
timestamp 1649977179
transform 1 0 188508 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _398_
timestamp 1649977179
transform 1 0 194396 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _399_
timestamp 1649977179
transform 1 0 193108 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _400_
timestamp 1649977179
transform 1 0 196972 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _401_
timestamp 1649977179
transform 1 0 192280 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _402_
timestamp 1649977179
transform 1 0 198168 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _403_
timestamp 1649977179
transform 1 0 196236 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _404_
timestamp 1649977179
transform 1 0 248952 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _405_
timestamp 1649977179
transform 1 0 262384 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _406_
timestamp 1649977179
transform 1 0 268824 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _407_
timestamp 1649977179
transform 1 0 267720 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _408_
timestamp 1649977179
transform 1 0 272504 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _409_
timestamp 1649977179
transform 1 0 268364 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _410_
timestamp 1649977179
transform 1 0 271676 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _411_
timestamp 1649977179
transform 1 0 267076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _412_
timestamp 1649977179
transform 1 0 270020 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _413_
timestamp 1649977179
transform 1 0 267720 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _414_
timestamp 1649977179
transform 1 0 271308 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _415_
timestamp 1649977179
transform 1 0 267996 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _416_
timestamp 1649977179
transform 1 0 261740 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _417_
timestamp 1649977179
transform 1 0 267812 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _418_
timestamp 1649977179
transform 1 0 265788 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _419_
timestamp 1649977179
transform 1 0 266800 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _420_
timestamp 1649977179
transform 1 0 264960 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _421_
timestamp 1649977179
transform 1 0 267444 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _422_
timestamp 1649977179
transform 1 0 263948 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _423_
timestamp 1649977179
transform 1 0 265236 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _424_
timestamp 1649977179
transform 1 0 264592 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _425_
timestamp 1649977179
transform 1 0 262660 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _426_
timestamp 1649977179
transform 1 0 264592 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _427_
timestamp 1649977179
transform 1 0 251804 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _428_
timestamp 1649977179
transform 1 0 255852 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _429_
timestamp 1649977179
transform 1 0 253644 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _430_
timestamp 1649977179
transform 1 0 254748 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _431_
timestamp 1649977179
transform 1 0 253736 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _432_
timestamp 1649977179
transform 1 0 253644 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _433_
timestamp 1649977179
transform 1 0 253092 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _434_
timestamp 1649977179
transform 1 0 251988 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _435_
timestamp 1649977179
transform 1 0 251804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _436_
timestamp 1649977179
transform 1 0 249504 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _437_
timestamp 1649977179
transform 1 0 251068 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _438_
timestamp 1649977179
transform 1 0 243708 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _439_
timestamp 1649977179
transform 1 0 242328 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _440_
timestamp 1649977179
transform 1 0 243524 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _441_
timestamp 1649977179
transform 1 0 240856 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _442_
timestamp 1649977179
transform 1 0 241408 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _443_
timestamp 1649977179
transform 1 0 239844 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _444_
timestamp 1649977179
transform 1 0 241040 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _445_
timestamp 1649977179
transform 1 0 238740 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _446_
timestamp 1649977179
transform 1 0 239936 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _447_
timestamp 1649977179
transform 1 0 236716 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _448_
timestamp 1649977179
transform 1 0 236808 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _449_
timestamp 1649977179
transform 1 0 238556 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _450_
timestamp 1649977179
transform 1 0 230920 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _451_
timestamp 1649977179
transform 1 0 231564 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _452_
timestamp 1649977179
transform 1 0 229080 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _453_
timestamp 1649977179
transform 1 0 229172 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _454_
timestamp 1649977179
transform 1 0 227884 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _455_
timestamp 1649977179
transform 1 0 230092 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _456_
timestamp 1649977179
transform 1 0 226596 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _457_
timestamp 1649977179
transform 1 0 227148 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _458_
timestamp 1649977179
transform 1 0 223652 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _459_
timestamp 1649977179
transform 1 0 226504 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _460_
timestamp 1649977179
transform 1 0 165784 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _461_
timestamp 1649977179
transform 1 0 193384 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _462_
timestamp 1649977179
transform 1 0 207276 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _463_
timestamp 1649977179
transform 1 0 202124 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _464_
timestamp 1649977179
transform 1 0 204792 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _465_
timestamp 1649977179
transform 1 0 202860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _466_
timestamp 1649977179
transform 1 0 203596 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _467_
timestamp 1649977179
transform 1 0 199824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _468_
timestamp 1649977179
transform 1 0 202860 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _469_
timestamp 1649977179
transform 1 0 202860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _470_
timestamp 1649977179
transform 1 0 200468 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _471_
timestamp 1649977179
transform 1 0 201664 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _472_
timestamp 1649977179
transform 1 0 189244 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _473_
timestamp 1649977179
transform 1 0 196972 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _474_
timestamp 1649977179
transform 1 0 192464 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _475_
timestamp 1649977179
transform 1 0 193016 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _476_
timestamp 1649977179
transform 1 0 189428 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _477_
timestamp 1649977179
transform 1 0 190532 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _478_
timestamp 1649977179
transform 1 0 191084 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _479_
timestamp 1649977179
transform 1 0 191820 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _480_
timestamp 1649977179
transform 1 0 191820 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _481_
timestamp 1649977179
transform 1 0 187956 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _482_
timestamp 1649977179
transform 1 0 190164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _483_
timestamp 1649977179
transform 1 0 175536 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _484_
timestamp 1649977179
transform 1 0 181516 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _485_
timestamp 1649977179
transform 1 0 178940 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _486_
timestamp 1649977179
transform 1 0 178756 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _487_
timestamp 1649977179
transform 1 0 180780 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _488_
timestamp 1649977179
transform 1 0 177560 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _489_
timestamp 1649977179
transform 1 0 174984 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _490_
timestamp 1649977179
transform 1 0 176548 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _491_
timestamp 1649977179
transform 1 0 176456 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _492_
timestamp 1649977179
transform 1 0 173788 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _493_
timestamp 1649977179
transform 1 0 175628 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _494_
timestamp 1649977179
transform 1 0 167256 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _495_
timestamp 1649977179
transform 1 0 166060 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _496_
timestamp 1649977179
transform 1 0 162656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _497_
timestamp 1649977179
transform 1 0 164036 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _498_
timestamp 1649977179
transform 1 0 163484 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _499_
timestamp 1649977179
transform 1 0 162012 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _500_
timestamp 1649977179
transform 1 0 162012 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _501_
timestamp 1649977179
transform 1 0 160816 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _502_
timestamp 1649977179
transform 1 0 160908 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _503_
timestamp 1649977179
transform 1 0 158792 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _504_
timestamp 1649977179
transform 1 0 159988 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _505_
timestamp 1649977179
transform 1 0 161092 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _506_
timestamp 1649977179
transform 1 0 153272 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _507_
timestamp 1649977179
transform 1 0 154100 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _508_
timestamp 1649977179
transform 1 0 151064 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _509_
timestamp 1649977179
transform 1 0 151064 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _510_
timestamp 1649977179
transform 1 0 151616 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _511_
timestamp 1649977179
transform 1 0 148856 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _512_
timestamp 1649977179
transform 1 0 148028 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _513_
timestamp 1649977179
transform 1 0 147292 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _514_
timestamp 1649977179
transform 1 0 145452 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _515_
timestamp 1649977179
transform 1 0 147568 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _516_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 131652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _517_
timestamp 1649977179
transform 1 0 125396 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _518_
timestamp 1649977179
transform 1 0 133124 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _519_
timestamp 1649977179
transform 1 0 131744 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _520_
timestamp 1649977179
transform 1 0 131284 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _521_
timestamp 1649977179
transform 1 0 132388 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _522_
timestamp 1649977179
transform 1 0 130456 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _523_
timestamp 1649977179
transform 1 0 128064 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _524_
timestamp 1649977179
transform 1 0 128708 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _525_
timestamp 1649977179
transform 1 0 128432 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _526_
timestamp 1649977179
transform 1 0 126132 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _527_
timestamp 1649977179
transform 1 0 127696 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _528_
timestamp 1649977179
transform 1 0 113712 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _529_
timestamp 1649977179
transform 1 0 119692 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _530_
timestamp 1649977179
transform 1 0 117116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _531_
timestamp 1649977179
transform 1 0 117116 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _532_
timestamp 1649977179
transform 1 0 116196 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _533_
timestamp 1649977179
transform 1 0 115276 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _534_
timestamp 1649977179
transform 1 0 116012 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _535_
timestamp 1649977179
transform 1 0 114632 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _536_
timestamp 1649977179
transform 1 0 113804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _537_
timestamp 1649977179
transform 1 0 111872 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _538_
timestamp 1649977179
transform 1 0 113068 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _539_
timestamp 1649977179
transform 1 0 102028 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _540_
timestamp 1649977179
transform 1 0 104236 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _541_
timestamp 1649977179
transform 1 0 102948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _542_
timestamp 1649977179
transform 1 0 102580 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _543_
timestamp 1649977179
transform 1 0 103500 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _544_
timestamp 1649977179
transform 1 0 101476 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _545_
timestamp 1649977179
transform 1 0 101660 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _546_
timestamp 1649977179
transform 1 0 100372 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _547_
timestamp 1649977179
transform 1 0 100188 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _548_
timestamp 1649977179
transform 1 0 97520 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _549_
timestamp 1649977179
transform 1 0 99084 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _550_
timestamp 1649977179
transform 1 0 90344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _551_
timestamp 1649977179
transform 1 0 89148 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _552_
timestamp 1649977179
transform 1 0 88228 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _553_
timestamp 1649977179
transform 1 0 87584 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _554_
timestamp 1649977179
transform 1 0 87584 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _555_
timestamp 1649977179
transform 1 0 86388 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _556_
timestamp 1649977179
transform 1 0 82892 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _557_
timestamp 1649977179
transform 1 0 85652 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _558_
timestamp 1649977179
transform 1 0 86204 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _559_
timestamp 1649977179
transform 1 0 83996 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _560_
timestamp 1649977179
transform 1 0 85008 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _561_
timestamp 1649977179
transform 1 0 87676 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _562_
timestamp 1649977179
transform 1 0 81052 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _563_
timestamp 1649977179
transform 1 0 79120 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _564_
timestamp 1649977179
transform 1 0 77464 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _565_
timestamp 1649977179
transform 1 0 78200 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _566_
timestamp 1649977179
transform 1 0 76268 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _567_
timestamp 1649977179
transform 1 0 76912 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _568_
timestamp 1649977179
transform 1 0 75532 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _569_
timestamp 1649977179
transform 1 0 74888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _570_
timestamp 1649977179
transform 1 0 72036 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _571_
timestamp 1649977179
transform 1 0 76452 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _572_
timestamp 1649977179
transform 1 0 135332 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _573_
timestamp 1649977179
transform 1 0 86940 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _574_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 77740 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _575_
timestamp 1649977179
transform 1 0 77740 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _576_
timestamp 1649977179
transform 1 0 78476 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _577_
timestamp 1649977179
transform 1 0 79212 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _578_
timestamp 1649977179
transform 1 0 80132 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _579_
timestamp 1649977179
transform 1 0 91724 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _580_
timestamp 1649977179
transform 1 0 86848 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _581_
timestamp 1649977179
transform 1 0 85468 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _582_
timestamp 1649977179
transform 1 0 90068 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _583_
timestamp 1649977179
transform 1 0 88780 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _584_
timestamp 1649977179
transform 1 0 88780 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _585_
timestamp 1649977179
transform 1 0 101844 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _586_
timestamp 1649977179
transform 1 0 99728 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _587_
timestamp 1649977179
transform 1 0 100832 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _588_
timestamp 1649977179
transform 1 0 105064 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _589_
timestamp 1649977179
transform 1 0 104420 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _590_
timestamp 1649977179
transform 1 0 103776 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _591_
timestamp 1649977179
transform 1 0 114540 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _592_
timestamp 1649977179
transform 1 0 115276 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _593_
timestamp 1649977179
transform 1 0 113068 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _594_
timestamp 1649977179
transform 1 0 118312 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _595_
timestamp 1649977179
transform 1 0 116840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _596_
timestamp 1649977179
transform 1 0 117484 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _597_
timestamp 1649977179
transform 1 0 127328 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _598_
timestamp 1649977179
transform 1 0 129260 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _599_
timestamp 1649977179
transform 1 0 130364 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _600_
timestamp 1649977179
transform 1 0 131100 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _601_
timestamp 1649977179
transform 1 0 132572 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _602_
timestamp 1649977179
transform 1 0 130180 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _603_
timestamp 1649977179
transform 1 0 165232 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _604_
timestamp 1649977179
transform 1 0 159988 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _605_
timestamp 1649977179
transform 1 0 148304 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _606_
timestamp 1649977179
transform 1 0 150604 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _607_
timestamp 1649977179
transform 1 0 149868 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _608_
timestamp 1649977179
transform 1 0 152444 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _609_
timestamp 1649977179
transform 1 0 152628 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _610_
timestamp 1649977179
transform 1 0 166428 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _611_
timestamp 1649977179
transform 1 0 162196 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _612_
timestamp 1649977179
transform 1 0 162840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _613_
timestamp 1649977179
transform 1 0 163484 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _614_
timestamp 1649977179
transform 1 0 164772 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _615_
timestamp 1649977179
transform 1 0 164128 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _616_
timestamp 1649977179
transform 1 0 177836 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _617_
timestamp 1649977179
transform 1 0 177468 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _618_
timestamp 1649977179
transform 1 0 178112 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _619_
timestamp 1649977179
transform 1 0 179952 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _620_
timestamp 1649977179
transform 1 0 181516 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _621_
timestamp 1649977179
transform 1 0 182160 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _622_
timestamp 1649977179
transform 1 0 188508 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _623_
timestamp 1649977179
transform 1 0 187312 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _624_
timestamp 1649977179
transform 1 0 190164 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _625_
timestamp 1649977179
transform 1 0 194120 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _626_
timestamp 1649977179
transform 1 0 192924 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _627_
timestamp 1649977179
transform 1 0 196696 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _628_
timestamp 1649977179
transform 1 0 192648 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _629_
timestamp 1649977179
transform 1 0 202216 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _630_
timestamp 1649977179
transform 1 0 202768 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _631_
timestamp 1649977179
transform 1 0 203412 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _632_
timestamp 1649977179
transform 1 0 201020 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _633_
timestamp 1649977179
transform 1 0 200468 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _634_
timestamp 1649977179
transform 1 0 252632 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _635_
timestamp 1649977179
transform 1 0 238004 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _636_
timestamp 1649977179
transform 1 0 233036 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _637_
timestamp 1649977179
transform 1 0 230276 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _638_
timestamp 1649977179
transform 1 0 230920 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _639_
timestamp 1649977179
transform 1 0 232116 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _640_
timestamp 1649977179
transform 1 0 233036 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _641_
timestamp 1649977179
transform 1 0 244444 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _642_
timestamp 1649977179
transform 1 0 239844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _643_
timestamp 1649977179
transform 1 0 240764 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _644_
timestamp 1649977179
transform 1 0 241684 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _645_
timestamp 1649977179
transform 1 0 242052 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _646_
timestamp 1649977179
transform 1 0 245180 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _647_
timestamp 1649977179
transform 1 0 251252 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _648_
timestamp 1649977179
transform 1 0 252448 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _649_
timestamp 1649977179
transform 1 0 254840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _650_
timestamp 1649977179
transform 1 0 255484 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _651_
timestamp 1649977179
transform 1 0 257048 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _652_
timestamp 1649977179
transform 1 0 256220 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _653_
timestamp 1649977179
transform 1 0 261648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _654_
timestamp 1649977179
transform 1 0 263948 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _655_
timestamp 1649977179
transform 1 0 266432 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _656_
timestamp 1649977179
transform 1 0 264316 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _657_
timestamp 1649977179
transform 1 0 264868 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _658_
timestamp 1649977179
transform 1 0 267076 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _659_
timestamp 1649977179
transform 1 0 263120 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _660_
timestamp 1649977179
transform 1 0 270940 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _661_
timestamp 1649977179
transform 1 0 268364 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _662_
timestamp 1649977179
transform 1 0 269100 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _663_
timestamp 1649977179
transform 1 0 267812 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _664_
timestamp 1649977179
transform 1 0 271308 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _665_
timestamp 1649977179
transform 1 0 142968 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _666_
timestamp 1649977179
transform 1 0 149500 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _667_
timestamp 1649977179
transform 1 0 189520 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _668_
timestamp 1649977179
transform 1 0 190808 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _669_
timestamp 1649977179
transform 1 0 190072 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _670_
timestamp 1649977179
transform 1 0 190716 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _671_
timestamp 1649977179
transform 1 0 156400 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _672_
timestamp 1649977179
transform 1 0 36432 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _673_
timestamp 1649977179
transform 1 0 31556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _674_
timestamp 1649977179
transform 1 0 32108 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _675_
timestamp 1649977179
transform 1 0 33488 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _676_
timestamp 1649977179
transform 1 0 32752 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _677_
timestamp 1649977179
transform 1 0 32200 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _678_
timestamp 1649977179
transform 1 0 37260 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _679_
timestamp 1649977179
transform 1 0 33488 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _680_
timestamp 1649977179
transform 1 0 35328 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _681_
timestamp 1649977179
transform 1 0 34316 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _682_
timestamp 1649977179
transform 1 0 33672 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _683_
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _684_
timestamp 1649977179
transform 1 0 42780 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _685_
timestamp 1649977179
transform 1 0 39100 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _686_
timestamp 1649977179
transform 1 0 40940 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _687_
timestamp 1649977179
transform 1 0 41032 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _688_
timestamp 1649977179
transform 1 0 41676 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _689_
timestamp 1649977179
transform 1 0 42412 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _690_
timestamp 1649977179
transform 1 0 55384 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _691_
timestamp 1649977179
transform 1 0 52900 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _692_
timestamp 1649977179
transform 1 0 54280 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _693_
timestamp 1649977179
transform 1 0 54556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _694_
timestamp 1649977179
transform 1 0 56396 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _695_
timestamp 1649977179
transform 1 0 57040 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _696_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 73600 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _697_
timestamp 1649977179
transform 1 0 75532 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _698_
timestamp 1649977179
transform 1 0 76176 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _699_
timestamp 1649977179
transform 1 0 78476 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _700_
timestamp 1649977179
transform 1 0 79764 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _701_
timestamp 1649977179
transform 1 0 83996 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _702_
timestamp 1649977179
transform 1 0 83904 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _703_
timestamp 1649977179
transform 1 0 86204 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _704_
timestamp 1649977179
transform 1 0 86480 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _705_
timestamp 1649977179
transform 1 0 88780 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _706_
timestamp 1649977179
transform 1 0 99176 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _707_
timestamp 1649977179
transform 1 0 99360 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _708_
timestamp 1649977179
transform 1 0 101384 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _709_
timestamp 1649977179
transform 1 0 101936 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _710_
timestamp 1649977179
transform 1 0 104236 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _711_
timestamp 1649977179
transform 1 0 112240 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _712_
timestamp 1649977179
transform 1 0 114356 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _713_
timestamp 1649977179
transform 1 0 114816 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _714_
timestamp 1649977179
transform 1 0 116472 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _715_
timestamp 1649977179
transform 1 0 117392 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _716_
timestamp 1649977179
transform 1 0 127512 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _717_
timestamp 1649977179
transform 1 0 129076 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _718_
timestamp 1649977179
transform 1 0 130272 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _719_
timestamp 1649977179
transform 1 0 130824 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _720_
timestamp 1649977179
transform 1 0 132572 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _721_
timestamp 1649977179
transform 1 0 145728 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _722_
timestamp 1649977179
transform 1 0 147476 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _723_
timestamp 1649977179
transform 1 0 148304 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _724_
timestamp 1649977179
transform 1 0 150880 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _725_
timestamp 1649977179
transform 1 0 153456 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _726_
timestamp 1649977179
transform 1 0 158608 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _727_
timestamp 1649977179
transform 1 0 160908 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _728_
timestamp 1649977179
transform 1 0 161828 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _729_
timestamp 1649977179
transform 1 0 163484 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _730_
timestamp 1649977179
transform 1 0 163576 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _731_
timestamp 1649977179
transform 1 0 176364 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _732_
timestamp 1649977179
transform 1 0 176364 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _733_
timestamp 1649977179
transform 1 0 178940 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _734_
timestamp 1649977179
transform 1 0 178572 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _735_
timestamp 1649977179
transform 1 0 179124 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _736_
timestamp 1649977179
transform 1 0 189520 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _737_
timestamp 1649977179
transform 1 0 190808 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _738_
timestamp 1649977179
transform 1 0 191820 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _739_
timestamp 1649977179
transform 1 0 192004 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _740_
timestamp 1649977179
transform 1 0 194028 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _741_
timestamp 1649977179
transform 1 0 202124 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _742_
timestamp 1649977179
transform 1 0 202584 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _743_
timestamp 1649977179
transform 1 0 204700 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _744_
timestamp 1649977179
transform 1 0 204792 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _745_
timestamp 1649977179
transform 1 0 204700 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _746_
timestamp 1649977179
transform 1 0 227884 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _747_
timestamp 1649977179
transform 1 0 227884 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _748_
timestamp 1649977179
transform 1 0 227516 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _749_
timestamp 1649977179
transform 1 0 230460 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _750_
timestamp 1649977179
transform 1 0 230736 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _751_
timestamp 1649977179
transform 1 0 238188 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _752_
timestamp 1649977179
transform 1 0 238464 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _753_
timestamp 1649977179
transform 1 0 240764 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _754_
timestamp 1649977179
transform 1 0 240672 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _755_
timestamp 1649977179
transform 1 0 243340 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _756_
timestamp 1649977179
transform 1 0 251068 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _757_
timestamp 1649977179
transform 1 0 253644 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _758_
timestamp 1649977179
transform 1 0 252540 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _759_
timestamp 1649977179
transform 1 0 253644 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _760_
timestamp 1649977179
transform 1 0 256220 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _761_
timestamp 1649977179
transform 1 0 264224 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _762_
timestamp 1649977179
transform 1 0 265236 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _763_
timestamp 1649977179
transform 1 0 265604 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _764_
timestamp 1649977179
transform 1 0 266524 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _765_
timestamp 1649977179
transform 1 0 269100 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _766_
timestamp 1649977179
transform 1 0 269100 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _767_
timestamp 1649977179
transform 1 0 268732 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _768_
timestamp 1649977179
transform 1 0 271676 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _769_
timestamp 1649977179
transform 1 0 269100 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _770_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 266524 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _771_
timestamp 1649977179
transform 1 0 194396 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _772_
timestamp 1649977179
transform 1 0 194396 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _773_
timestamp 1649977179
transform 1 0 191820 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _774_
timestamp 1649977179
transform 1 0 193016 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _775_
timestamp 1649977179
transform 1 0 148028 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _776_
timestamp 1649977179
transform 1 0 29624 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _777_
timestamp 1649977179
transform 1 0 27232 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _778_
timestamp 1649977179
transform 1 0 29624 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _779_
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _780_
timestamp 1649977179
transform 1 0 29808 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _781_
timestamp 1649977179
transform 1 0 29808 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _782_
timestamp 1649977179
transform 1 0 31740 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _783_
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _784_
timestamp 1649977179
transform 1 0 32384 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _785_
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _786_
timestamp 1649977179
transform 1 0 37536 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _787_
timestamp 1649977179
transform 1 0 39468 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _788_
timestamp 1649977179
transform 1 0 40112 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _789_
timestamp 1649977179
transform 1 0 41400 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _790_
timestamp 1649977179
transform 1 0 42504 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _791_
timestamp 1649977179
transform 1 0 52348 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _792_
timestamp 1649977179
transform 1 0 52992 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _793_
timestamp 1649977179
transform 1 0 54740 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _794_
timestamp 1649977179
transform 1 0 55568 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _795_
timestamp 1649977179
transform 1 0 57868 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_6  _796_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 187128 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 149408 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1649977179
transform 1 0 140668 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1649977179
transform 1 0 140392 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1649977179
transform 1 0 140392 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1649977179
transform 1 0 140668 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1649977179
transform 1 0 156124 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1649977179
transform 1 0 156032 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1649977179
transform 1 0 156032 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1649977179
transform 1 0 156124 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 303692 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  input2
timestamp 1649977179
transform 1 0 303876 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  input3
timestamp 1649977179
transform 1 0 304336 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  output4
timestamp 1649977179
transform 1 0 1564 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output5
timestamp 1649977179
transform 1 0 32844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output6
timestamp 1649977179
transform 1 0 35512 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output7
timestamp 1649977179
transform 1 0 38364 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output8
timestamp 1649977179
transform 1 0 42228 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output9
timestamp 1649977179
transform 1 0 44528 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output10
timestamp 1649977179
transform 1 0 47564 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output11
timestamp 1649977179
transform 1 0 50324 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output12
timestamp 1649977179
transform 1 0 53636 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output13
timestamp 1649977179
transform 1 0 57316 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output14
timestamp 1649977179
transform 1 0 60444 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output15
timestamp 1649977179
transform 1 0 4600 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output16
timestamp 1649977179
transform 1 0 63020 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output17
timestamp 1649977179
transform 1 0 65964 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output18
timestamp 1649977179
transform 1 0 69092 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output19
timestamp 1649977179
transform 1 0 72128 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output20
timestamp 1649977179
transform 1 0 75164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output21
timestamp 1649977179
transform 1 0 78476 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output22
timestamp 1649977179
transform 1 0 82248 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output23
timestamp 1649977179
transform 1 0 84364 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output24
timestamp 1649977179
transform 1 0 89424 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output25
timestamp 1649977179
transform 1 0 91080 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output26
timestamp 1649977179
transform 1 0 7636 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output27
timestamp 1649977179
transform 1 0 93932 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output28
timestamp 1649977179
transform 1 0 96692 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output29
timestamp 1649977179
transform 1 0 98348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output30
timestamp 1649977179
transform 1 0 102856 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output31
timestamp 1649977179
transform 1 0 105892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output32
timestamp 1649977179
transform 1 0 109388 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output33
timestamp 1649977179
transform 1 0 111228 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output34
timestamp 1649977179
transform 1 0 113712 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output35
timestamp 1649977179
transform 1 0 118680 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output36
timestamp 1649977179
transform 1 0 121256 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output37
timestamp 1649977179
transform 1 0 10764 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output38
timestamp 1649977179
transform 1 0 124108 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output39
timestamp 1649977179
transform 1 0 126684 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output40
timestamp 1649977179
transform 1 0 130456 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output41
timestamp 1649977179
transform 1 0 134320 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output42
timestamp 1649977179
transform 1 0 136620 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output43
timestamp 1649977179
transform 1 0 140300 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output44
timestamp 1649977179
transform 1 0 142876 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output45
timestamp 1649977179
transform 1 0 144716 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output46
timestamp 1649977179
transform 1 0 146832 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output47
timestamp 1649977179
transform 1 0 151984 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output48
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output49
timestamp 1649977179
transform 1 0 155756 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output50
timestamp 1649977179
transform 1 0 157596 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output51
timestamp 1649977179
transform 1 0 161552 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output52
timestamp 1649977179
transform 1 0 167164 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output53
timestamp 1649977179
transform 1 0 167808 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output54
timestamp 1649977179
transform 1 0 170384 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output55
timestamp 1649977179
transform 1 0 173052 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output56
timestamp 1649977179
transform 1 0 175904 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output57
timestamp 1649977179
transform 1 0 181332 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output58
timestamp 1649977179
transform 1 0 182712 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output59
timestamp 1649977179
transform 1 0 16836 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output60
timestamp 1649977179
transform 1 0 185748 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output61
timestamp 1649977179
transform 1 0 187864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output62
timestamp 1649977179
transform 1 0 191820 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output63
timestamp 1649977179
transform 1 0 195592 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output64
timestamp 1649977179
transform 1 0 198168 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output65
timestamp 1649977179
transform 1 0 201112 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output66
timestamp 1649977179
transform 1 0 204700 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output67
timestamp 1649977179
transform 1 0 207276 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output68
timestamp 1649977179
transform 1 0 210312 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output69
timestamp 1649977179
transform 1 0 213348 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output70
timestamp 1649977179
transform 1 0 19964 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output71
timestamp 1649977179
transform 1 0 216384 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output72
timestamp 1649977179
transform 1 0 220156 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output73
timestamp 1649977179
transform 1 0 222732 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output74
timestamp 1649977179
transform 1 0 225676 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output75
timestamp 1649977179
transform 1 0 229724 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output76
timestamp 1649977179
transform 1 0 233680 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output77
timestamp 1649977179
transform 1 0 234876 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output78
timestamp 1649977179
transform 1 0 237452 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output79
timestamp 1649977179
transform 1 0 242328 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output80
timestamp 1649977179
transform 1 0 244168 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output81
timestamp 1649977179
transform 1 0 23000 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output82
timestamp 1649977179
transform 1 0 247112 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output83
timestamp 1649977179
transform 1 0 250148 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output84
timestamp 1649977179
transform 1 0 254380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output85
timestamp 1649977179
transform 1 0 256864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output86
timestamp 1649977179
transform 1 0 259440 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output87
timestamp 1649977179
transform 1 0 262476 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output88
timestamp 1649977179
transform 1 0 265512 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output89
timestamp 1649977179
transform 1 0 269008 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output90
timestamp 1649977179
transform 1 0 274252 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output91
timestamp 1649977179
transform 1 0 274896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output92
timestamp 1649977179
transform 1 0 26036 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output93
timestamp 1649977179
transform 1 0 277840 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output94
timestamp 1649977179
transform 1 0 280876 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output95
timestamp 1649977179
transform 1 0 284556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output96
timestamp 1649977179
transform 1 0 287132 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output97
timestamp 1649977179
transform 1 0 290076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output98
timestamp 1649977179
transform 1 0 293204 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output99
timestamp 1649977179
transform 1 0 296240 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output100
timestamp 1649977179
transform 1 0 299276 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output101
timestamp 1649977179
transform 1 0 302588 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output102
timestamp 1649977179
transform 1 0 304428 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output103
timestamp 1649977179
transform 1 0 27784 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output104
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
<< labels >>
rlabel metal4 s -1076 -4 -756 15780 4 GND
port 0 nsew ground bidirectional
rlabel metal5 s -1076 -4 307988 316 6 GND
port 0 nsew ground bidirectional
rlabel metal5 s -1076 15460 307988 15780 6 GND
port 0 nsew ground bidirectional
rlabel metal4 s 307668 -4 307988 15780 6 GND
port 0 nsew ground bidirectional
rlabel metal4 s 77142 -4 77462 15780 6 GND
port 0 nsew ground bidirectional
rlabel metal4 s 153340 -4 153660 15780 6 GND
port 0 nsew ground bidirectional
rlabel metal4 s 229538 -4 229858 15780 6 GND
port 0 nsew ground bidirectional
rlabel metal5 s -1076 4928 307988 5248 6 GND
port 0 nsew ground bidirectional
rlabel metal5 s -1076 7840 307988 8160 6 GND
port 0 nsew ground bidirectional
rlabel metal5 s -1076 10752 307988 11072 6 GND
port 0 nsew ground bidirectional
rlabel metal2 s 1490 15200 1546 16000 6 ROW_SEL[0]
port 1 nsew signal tristate
rlabel metal2 s 32126 15200 32182 16000 6 ROW_SEL[10]
port 2 nsew signal tristate
rlabel metal2 s 35254 15200 35310 16000 6 ROW_SEL[11]
port 3 nsew signal tristate
rlabel metal2 s 38290 15200 38346 16000 6 ROW_SEL[12]
port 4 nsew signal tristate
rlabel metal2 s 41326 15200 41382 16000 6 ROW_SEL[13]
port 5 nsew signal tristate
rlabel metal2 s 44454 15200 44510 16000 6 ROW_SEL[14]
port 6 nsew signal tristate
rlabel metal2 s 47490 15200 47546 16000 6 ROW_SEL[15]
port 7 nsew signal tristate
rlabel metal2 s 50526 15200 50582 16000 6 ROW_SEL[16]
port 8 nsew signal tristate
rlabel metal2 s 53654 15200 53710 16000 6 ROW_SEL[17]
port 9 nsew signal tristate
rlabel metal2 s 56690 15200 56746 16000 6 ROW_SEL[18]
port 10 nsew signal tristate
rlabel metal2 s 59818 15200 59874 16000 6 ROW_SEL[19]
port 11 nsew signal tristate
rlabel metal2 s 4526 15200 4582 16000 6 ROW_SEL[1]
port 12 nsew signal tristate
rlabel metal2 s 62854 15200 62910 16000 6 ROW_SEL[20]
port 13 nsew signal tristate
rlabel metal2 s 65890 15200 65946 16000 6 ROW_SEL[21]
port 14 nsew signal tristate
rlabel metal2 s 69018 15200 69074 16000 6 ROW_SEL[22]
port 15 nsew signal tristate
rlabel metal2 s 72054 15200 72110 16000 6 ROW_SEL[23]
port 16 nsew signal tristate
rlabel metal2 s 75090 15200 75146 16000 6 ROW_SEL[24]
port 17 nsew signal tristate
rlabel metal2 s 78218 15200 78274 16000 6 ROW_SEL[25]
port 18 nsew signal tristate
rlabel metal2 s 81254 15200 81310 16000 6 ROW_SEL[26]
port 19 nsew signal tristate
rlabel metal2 s 84290 15200 84346 16000 6 ROW_SEL[27]
port 20 nsew signal tristate
rlabel metal2 s 87418 15200 87474 16000 6 ROW_SEL[28]
port 21 nsew signal tristate
rlabel metal2 s 90454 15200 90510 16000 6 ROW_SEL[29]
port 22 nsew signal tristate
rlabel metal2 s 7562 15200 7618 16000 6 ROW_SEL[2]
port 23 nsew signal tristate
rlabel metal2 s 93582 15200 93638 16000 6 ROW_SEL[30]
port 24 nsew signal tristate
rlabel metal2 s 96618 15200 96674 16000 6 ROW_SEL[31]
port 25 nsew signal tristate
rlabel metal2 s 99654 15200 99710 16000 6 ROW_SEL[32]
port 26 nsew signal tristate
rlabel metal2 s 102782 15200 102838 16000 6 ROW_SEL[33]
port 27 nsew signal tristate
rlabel metal2 s 105818 15200 105874 16000 6 ROW_SEL[34]
port 28 nsew signal tristate
rlabel metal2 s 108854 15200 108910 16000 6 ROW_SEL[35]
port 29 nsew signal tristate
rlabel metal2 s 111982 15200 112038 16000 6 ROW_SEL[36]
port 30 nsew signal tristate
rlabel metal2 s 115018 15200 115074 16000 6 ROW_SEL[37]
port 31 nsew signal tristate
rlabel metal2 s 118146 15200 118202 16000 6 ROW_SEL[38]
port 32 nsew signal tristate
rlabel metal2 s 121182 15200 121238 16000 6 ROW_SEL[39]
port 33 nsew signal tristate
rlabel metal2 s 10690 15200 10746 16000 6 ROW_SEL[3]
port 34 nsew signal tristate
rlabel metal2 s 124218 15200 124274 16000 6 ROW_SEL[40]
port 35 nsew signal tristate
rlabel metal2 s 127346 15200 127402 16000 6 ROW_SEL[41]
port 36 nsew signal tristate
rlabel metal2 s 130382 15200 130438 16000 6 ROW_SEL[42]
port 37 nsew signal tristate
rlabel metal2 s 133418 15200 133474 16000 6 ROW_SEL[43]
port 38 nsew signal tristate
rlabel metal2 s 136546 15200 136602 16000 6 ROW_SEL[44]
port 39 nsew signal tristate
rlabel metal2 s 139582 15200 139638 16000 6 ROW_SEL[45]
port 40 nsew signal tristate
rlabel metal2 s 142710 15200 142766 16000 6 ROW_SEL[46]
port 41 nsew signal tristate
rlabel metal2 s 145746 15200 145802 16000 6 ROW_SEL[47]
port 42 nsew signal tristate
rlabel metal2 s 148782 15200 148838 16000 6 ROW_SEL[48]
port 43 nsew signal tristate
rlabel metal2 s 151910 15200 151966 16000 6 ROW_SEL[49]
port 44 nsew signal tristate
rlabel metal2 s 13726 15200 13782 16000 6 ROW_SEL[4]
port 45 nsew signal tristate
rlabel metal2 s 154946 15200 155002 16000 6 ROW_SEL[50]
port 46 nsew signal tristate
rlabel metal2 s 157982 15200 158038 16000 6 ROW_SEL[51]
port 47 nsew signal tristate
rlabel metal2 s 161110 15200 161166 16000 6 ROW_SEL[52]
port 48 nsew signal tristate
rlabel metal2 s 164146 15200 164202 16000 6 ROW_SEL[53]
port 49 nsew signal tristate
rlabel metal2 s 167182 15200 167238 16000 6 ROW_SEL[54]
port 50 nsew signal tristate
rlabel metal2 s 170310 15200 170366 16000 6 ROW_SEL[55]
port 51 nsew signal tristate
rlabel metal2 s 173346 15200 173402 16000 6 ROW_SEL[56]
port 52 nsew signal tristate
rlabel metal2 s 176474 15200 176530 16000 6 ROW_SEL[57]
port 53 nsew signal tristate
rlabel metal2 s 179510 15200 179566 16000 6 ROW_SEL[58]
port 54 nsew signal tristate
rlabel metal2 s 182546 15200 182602 16000 6 ROW_SEL[59]
port 55 nsew signal tristate
rlabel metal2 s 16762 15200 16818 16000 6 ROW_SEL[5]
port 56 nsew signal tristate
rlabel metal2 s 185674 15200 185730 16000 6 ROW_SEL[60]
port 57 nsew signal tristate
rlabel metal2 s 188710 15200 188766 16000 6 ROW_SEL[61]
port 58 nsew signal tristate
rlabel metal2 s 191746 15200 191802 16000 6 ROW_SEL[62]
port 59 nsew signal tristate
rlabel metal2 s 194874 15200 194930 16000 6 ROW_SEL[63]
port 60 nsew signal tristate
rlabel metal2 s 197910 15200 197966 16000 6 ROW_SEL[64]
port 61 nsew signal tristate
rlabel metal2 s 201038 15200 201094 16000 6 ROW_SEL[65]
port 62 nsew signal tristate
rlabel metal2 s 204074 15200 204130 16000 6 ROW_SEL[66]
port 63 nsew signal tristate
rlabel metal2 s 207110 15200 207166 16000 6 ROW_SEL[67]
port 64 nsew signal tristate
rlabel metal2 s 210238 15200 210294 16000 6 ROW_SEL[68]
port 65 nsew signal tristate
rlabel metal2 s 213274 15200 213330 16000 6 ROW_SEL[69]
port 66 nsew signal tristate
rlabel metal2 s 19890 15200 19946 16000 6 ROW_SEL[6]
port 67 nsew signal tristate
rlabel metal2 s 216310 15200 216366 16000 6 ROW_SEL[70]
port 68 nsew signal tristate
rlabel metal2 s 219438 15200 219494 16000 6 ROW_SEL[71]
port 69 nsew signal tristate
rlabel metal2 s 222474 15200 222530 16000 6 ROW_SEL[72]
port 70 nsew signal tristate
rlabel metal2 s 225602 15200 225658 16000 6 ROW_SEL[73]
port 71 nsew signal tristate
rlabel metal2 s 228638 15200 228694 16000 6 ROW_SEL[74]
port 72 nsew signal tristate
rlabel metal2 s 231674 15200 231730 16000 6 ROW_SEL[75]
port 73 nsew signal tristate
rlabel metal2 s 234802 15200 234858 16000 6 ROW_SEL[76]
port 74 nsew signal tristate
rlabel metal2 s 237838 15200 237894 16000 6 ROW_SEL[77]
port 75 nsew signal tristate
rlabel metal2 s 240874 15200 240930 16000 6 ROW_SEL[78]
port 76 nsew signal tristate
rlabel metal2 s 244002 15200 244058 16000 6 ROW_SEL[79]
port 77 nsew signal tristate
rlabel metal2 s 22926 15200 22982 16000 6 ROW_SEL[7]
port 78 nsew signal tristate
rlabel metal2 s 247038 15200 247094 16000 6 ROW_SEL[80]
port 79 nsew signal tristate
rlabel metal2 s 250074 15200 250130 16000 6 ROW_SEL[81]
port 80 nsew signal tristate
rlabel metal2 s 253202 15200 253258 16000 6 ROW_SEL[82]
port 81 nsew signal tristate
rlabel metal2 s 256238 15200 256294 16000 6 ROW_SEL[83]
port 82 nsew signal tristate
rlabel metal2 s 259366 15200 259422 16000 6 ROW_SEL[84]
port 83 nsew signal tristate
rlabel metal2 s 262402 15200 262458 16000 6 ROW_SEL[85]
port 84 nsew signal tristate
rlabel metal2 s 265438 15200 265494 16000 6 ROW_SEL[86]
port 85 nsew signal tristate
rlabel metal2 s 268566 15200 268622 16000 6 ROW_SEL[87]
port 86 nsew signal tristate
rlabel metal2 s 271602 15200 271658 16000 6 ROW_SEL[88]
port 87 nsew signal tristate
rlabel metal2 s 274638 15200 274694 16000 6 ROW_SEL[89]
port 88 nsew signal tristate
rlabel metal2 s 25962 15200 26018 16000 6 ROW_SEL[8]
port 89 nsew signal tristate
rlabel metal2 s 277766 15200 277822 16000 6 ROW_SEL[90]
port 90 nsew signal tristate
rlabel metal2 s 280802 15200 280858 16000 6 ROW_SEL[91]
port 91 nsew signal tristate
rlabel metal2 s 283930 15200 283986 16000 6 ROW_SEL[92]
port 92 nsew signal tristate
rlabel metal2 s 286966 15200 287022 16000 6 ROW_SEL[93]
port 93 nsew signal tristate
rlabel metal2 s 290002 15200 290058 16000 6 ROW_SEL[94]
port 94 nsew signal tristate
rlabel metal2 s 293130 15200 293186 16000 6 ROW_SEL[95]
port 95 nsew signal tristate
rlabel metal2 s 296166 15200 296222 16000 6 ROW_SEL[96]
port 96 nsew signal tristate
rlabel metal2 s 299202 15200 299258 16000 6 ROW_SEL[97]
port 97 nsew signal tristate
rlabel metal2 s 302330 15200 302386 16000 6 ROW_SEL[98]
port 98 nsew signal tristate
rlabel metal2 s 305366 15200 305422 16000 6 ROW_SEL[99]
port 99 nsew signal tristate
rlabel metal2 s 29090 15200 29146 16000 6 ROW_SEL[9]
port 100 nsew signal tristate
rlabel metal4 s -416 656 -96 15120 4 VDD
port 101 nsew power bidirectional
rlabel metal5 s -416 656 307328 976 6 VDD
port 101 nsew power bidirectional
rlabel metal5 s -416 14800 307328 15120 6 VDD
port 101 nsew power bidirectional
rlabel metal4 s 307008 656 307328 15120 6 VDD
port 101 nsew power bidirectional
rlabel metal4 s 39043 -4 39363 15780 6 VDD
port 101 nsew power bidirectional
rlabel metal4 s 115241 -4 115561 15780 6 VDD
port 101 nsew power bidirectional
rlabel metal4 s 191439 -4 191759 15780 6 VDD
port 101 nsew power bidirectional
rlabel metal4 s 267637 -4 267957 15780 6 VDD
port 101 nsew power bidirectional
rlabel metal5 s -1076 3472 307988 3792 6 VDD
port 101 nsew power bidirectional
rlabel metal5 s -1076 6384 307988 6704 6 VDD
port 101 nsew power bidirectional
rlabel metal5 s -1076 9296 307988 9616 6 VDD
port 101 nsew power bidirectional
rlabel metal5 s -1076 12208 307988 12528 6 VDD
port 101 nsew power bidirectional
rlabel metal3 s 306200 1912 307000 2032 6 clk
port 102 nsew signal input
rlabel metal3 s 306200 13880 307000 14000 6 data_in
port 103 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 data_out
port 104 nsew signal tristate
rlabel metal3 s 306200 5856 307000 5976 6 ena
port 105 nsew signal input
rlabel metal3 s 306200 9936 307000 10056 6 rst
port 106 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 307000 16000
<< end >>
