magic
tech sky130A
magscale 1 2
timestamp 1654740282
<< checkpaint >>
rect 20160 -181440 300705 3783
rect 40320 -297711 300705 -181440
<< nmoslvt >>
rect 540 -297800 2140 -297400
rect 3540 -297800 5140 -297400
rect 6540 -297800 8140 -297400
rect 9540 -297800 11140 -297400
rect 12540 -297800 14140 -297400
rect 15540 -297800 17140 -297400
rect 18540 -297800 20140 -297400
rect 21540 -297800 23140 -297400
rect 24540 -297800 26140 -297400
rect 27540 -297800 29140 -297400
rect 30540 -297800 32140 -297400
rect 33540 -297800 35140 -297400
rect 36540 -297800 38140 -297400
rect 39540 -297800 41140 -297400
rect 42540 -297800 44140 -297400
rect 45540 -297800 47140 -297400
rect 48540 -297800 50140 -297400
rect 51540 -297800 53140 -297400
rect 54540 -297800 56140 -297400
rect 57540 -297800 59140 -297400
rect 60540 -297800 62140 -297400
rect 63540 -297800 65140 -297400
rect 66540 -297800 68140 -297400
rect 69540 -297800 71140 -297400
rect 72540 -297800 74140 -297400
rect 75540 -297800 77140 -297400
rect 78540 -297800 80140 -297400
rect 81540 -297800 83140 -297400
rect 84540 -297800 86140 -297400
rect 87540 -297800 89140 -297400
rect 90540 -297800 92140 -297400
rect 93540 -297800 95140 -297400
rect 96540 -297800 98140 -297400
rect 99540 -297800 101140 -297400
rect 102540 -297800 104140 -297400
rect 105540 -297800 107140 -297400
rect 108540 -297800 110140 -297400
rect 111540 -297800 113140 -297400
rect 114540 -297800 116140 -297400
rect 117540 -297800 119140 -297400
rect 120540 -297800 122140 -297400
rect 123540 -297800 125140 -297400
rect 126540 -297800 128140 -297400
rect 129540 -297800 131140 -297400
rect 132540 -297800 134140 -297400
rect 135540 -297800 137140 -297400
rect 138540 -297800 140140 -297400
rect 141540 -297800 143140 -297400
rect 144540 -297800 146140 -297400
rect 147540 -297800 149140 -297400
rect 150540 -297800 152140 -297400
rect 153540 -297800 155140 -297400
rect 156540 -297800 158140 -297400
rect 159540 -297800 161140 -297400
rect 162540 -297800 164140 -297400
rect 165540 -297800 167140 -297400
rect 168540 -297800 170140 -297400
rect 171540 -297800 173140 -297400
rect 174540 -297800 176140 -297400
rect 177540 -297800 179140 -297400
rect 180540 -297800 182140 -297400
rect 183540 -297800 185140 -297400
rect 186540 -297800 188140 -297400
rect 189540 -297800 191140 -297400
rect 192540 -297800 194140 -297400
rect 195540 -297800 197140 -297400
rect 198540 -297800 200140 -297400
rect 201540 -297800 203140 -297400
rect 204540 -297800 206140 -297400
rect 207540 -297800 209140 -297400
rect 210540 -297800 212140 -297400
rect 213540 -297800 215140 -297400
rect 216540 -297800 218140 -297400
rect 219540 -297800 221140 -297400
rect 222540 -297800 224140 -297400
rect 225540 -297800 227140 -297400
rect 228540 -297800 230140 -297400
rect 231540 -297800 233140 -297400
rect 234540 -297800 236140 -297400
rect 237540 -297800 239140 -297400
rect 240540 -297800 242140 -297400
rect 243540 -297800 245140 -297400
rect 246540 -297800 248140 -297400
rect 249540 -297800 251140 -297400
rect 252540 -297800 254140 -297400
rect 255540 -297800 257140 -297400
rect 258540 -297800 260140 -297400
rect 261540 -297800 263140 -297400
rect 264540 -297800 266140 -297400
rect 267540 -297800 269140 -297400
rect 270540 -297800 272140 -297400
rect 273540 -297800 275140 -297400
rect 276540 -297800 278140 -297400
rect 279540 -297800 281140 -297400
rect 282540 -297800 284140 -297400
rect 285540 -297800 287140 -297400
rect 288540 -297800 290140 -297400
rect 291540 -297800 293140 -297400
rect 294540 -297800 296140 -297400
rect 297540 -297800 299140 -297400
<< ndiff >>
rect 540 -297320 2140 -297300
rect 540 -297380 560 -297320
rect 2120 -297380 2140 -297320
rect 540 -297400 2140 -297380
rect 3540 -297320 5140 -297300
rect 3540 -297380 3560 -297320
rect 5120 -297380 5140 -297320
rect 3540 -297400 5140 -297380
rect 6540 -297320 8140 -297300
rect 6540 -297380 6560 -297320
rect 8120 -297380 8140 -297320
rect 6540 -297400 8140 -297380
rect 9540 -297320 11140 -297300
rect 9540 -297380 9560 -297320
rect 11120 -297380 11140 -297320
rect 9540 -297400 11140 -297380
rect 12540 -297320 14140 -297300
rect 12540 -297380 12560 -297320
rect 14120 -297380 14140 -297320
rect 12540 -297400 14140 -297380
rect 15540 -297320 17140 -297300
rect 15540 -297380 15560 -297320
rect 17120 -297380 17140 -297320
rect 15540 -297400 17140 -297380
rect 18540 -297320 20140 -297300
rect 18540 -297380 18560 -297320
rect 20120 -297380 20140 -297320
rect 18540 -297400 20140 -297380
rect 21540 -297320 23140 -297300
rect 21540 -297380 21560 -297320
rect 23120 -297380 23140 -297320
rect 21540 -297400 23140 -297380
rect 24540 -297320 26140 -297300
rect 24540 -297380 24560 -297320
rect 26120 -297380 26140 -297320
rect 24540 -297400 26140 -297380
rect 27540 -297320 29140 -297300
rect 27540 -297380 27560 -297320
rect 29120 -297380 29140 -297320
rect 27540 -297400 29140 -297380
rect 30540 -297320 32140 -297300
rect 30540 -297380 30560 -297320
rect 32120 -297380 32140 -297320
rect 30540 -297400 32140 -297380
rect 33540 -297320 35140 -297300
rect 33540 -297380 33560 -297320
rect 35120 -297380 35140 -297320
rect 33540 -297400 35140 -297380
rect 36540 -297320 38140 -297300
rect 36540 -297380 36560 -297320
rect 38120 -297380 38140 -297320
rect 36540 -297400 38140 -297380
rect 39540 -297320 41140 -297300
rect 39540 -297380 39560 -297320
rect 41120 -297380 41140 -297320
rect 39540 -297400 41140 -297380
rect 42540 -297320 44140 -297300
rect 42540 -297380 42560 -297320
rect 44120 -297380 44140 -297320
rect 42540 -297400 44140 -297380
rect 45540 -297320 47140 -297300
rect 45540 -297380 45560 -297320
rect 47120 -297380 47140 -297320
rect 45540 -297400 47140 -297380
rect 48540 -297320 50140 -297300
rect 48540 -297380 48560 -297320
rect 50120 -297380 50140 -297320
rect 48540 -297400 50140 -297380
rect 51540 -297320 53140 -297300
rect 51540 -297380 51560 -297320
rect 53120 -297380 53140 -297320
rect 51540 -297400 53140 -297380
rect 54540 -297320 56140 -297300
rect 54540 -297380 54560 -297320
rect 56120 -297380 56140 -297320
rect 54540 -297400 56140 -297380
rect 57540 -297320 59140 -297300
rect 57540 -297380 57560 -297320
rect 59120 -297380 59140 -297320
rect 57540 -297400 59140 -297380
rect 60540 -297320 62140 -297300
rect 60540 -297380 60560 -297320
rect 62120 -297380 62140 -297320
rect 60540 -297400 62140 -297380
rect 63540 -297320 65140 -297300
rect 63540 -297380 63560 -297320
rect 65120 -297380 65140 -297320
rect 63540 -297400 65140 -297380
rect 66540 -297320 68140 -297300
rect 66540 -297380 66560 -297320
rect 68120 -297380 68140 -297320
rect 66540 -297400 68140 -297380
rect 69540 -297320 71140 -297300
rect 69540 -297380 69560 -297320
rect 71120 -297380 71140 -297320
rect 69540 -297400 71140 -297380
rect 72540 -297320 74140 -297300
rect 72540 -297380 72560 -297320
rect 74120 -297380 74140 -297320
rect 72540 -297400 74140 -297380
rect 75540 -297320 77140 -297300
rect 75540 -297380 75560 -297320
rect 77120 -297380 77140 -297320
rect 75540 -297400 77140 -297380
rect 78540 -297320 80140 -297300
rect 78540 -297380 78560 -297320
rect 80120 -297380 80140 -297320
rect 78540 -297400 80140 -297380
rect 81540 -297320 83140 -297300
rect 81540 -297380 81560 -297320
rect 83120 -297380 83140 -297320
rect 81540 -297400 83140 -297380
rect 84540 -297320 86140 -297300
rect 84540 -297380 84560 -297320
rect 86120 -297380 86140 -297320
rect 84540 -297400 86140 -297380
rect 87540 -297320 89140 -297300
rect 87540 -297380 87560 -297320
rect 89120 -297380 89140 -297320
rect 87540 -297400 89140 -297380
rect 90540 -297320 92140 -297300
rect 90540 -297380 90560 -297320
rect 92120 -297380 92140 -297320
rect 90540 -297400 92140 -297380
rect 93540 -297320 95140 -297300
rect 93540 -297380 93560 -297320
rect 95120 -297380 95140 -297320
rect 93540 -297400 95140 -297380
rect 96540 -297320 98140 -297300
rect 96540 -297380 96560 -297320
rect 98120 -297380 98140 -297320
rect 96540 -297400 98140 -297380
rect 99540 -297320 101140 -297300
rect 99540 -297380 99560 -297320
rect 101120 -297380 101140 -297320
rect 99540 -297400 101140 -297380
rect 102540 -297320 104140 -297300
rect 102540 -297380 102560 -297320
rect 104120 -297380 104140 -297320
rect 102540 -297400 104140 -297380
rect 105540 -297320 107140 -297300
rect 105540 -297380 105560 -297320
rect 107120 -297380 107140 -297320
rect 105540 -297400 107140 -297380
rect 108540 -297320 110140 -297300
rect 108540 -297380 108560 -297320
rect 110120 -297380 110140 -297320
rect 108540 -297400 110140 -297380
rect 111540 -297320 113140 -297300
rect 111540 -297380 111560 -297320
rect 113120 -297380 113140 -297320
rect 111540 -297400 113140 -297380
rect 114540 -297320 116140 -297300
rect 114540 -297380 114560 -297320
rect 116120 -297380 116140 -297320
rect 114540 -297400 116140 -297380
rect 117540 -297320 119140 -297300
rect 117540 -297380 117560 -297320
rect 119120 -297380 119140 -297320
rect 117540 -297400 119140 -297380
rect 120540 -297320 122140 -297300
rect 120540 -297380 120560 -297320
rect 122120 -297380 122140 -297320
rect 120540 -297400 122140 -297380
rect 123540 -297320 125140 -297300
rect 123540 -297380 123560 -297320
rect 125120 -297380 125140 -297320
rect 123540 -297400 125140 -297380
rect 126540 -297320 128140 -297300
rect 126540 -297380 126560 -297320
rect 128120 -297380 128140 -297320
rect 126540 -297400 128140 -297380
rect 129540 -297320 131140 -297300
rect 129540 -297380 129560 -297320
rect 131120 -297380 131140 -297320
rect 129540 -297400 131140 -297380
rect 132540 -297320 134140 -297300
rect 132540 -297380 132560 -297320
rect 134120 -297380 134140 -297320
rect 132540 -297400 134140 -297380
rect 135540 -297320 137140 -297300
rect 135540 -297380 135560 -297320
rect 137120 -297380 137140 -297320
rect 135540 -297400 137140 -297380
rect 138540 -297320 140140 -297300
rect 138540 -297380 138560 -297320
rect 140120 -297380 140140 -297320
rect 138540 -297400 140140 -297380
rect 141540 -297320 143140 -297300
rect 141540 -297380 141560 -297320
rect 143120 -297380 143140 -297320
rect 141540 -297400 143140 -297380
rect 144540 -297320 146140 -297300
rect 144540 -297380 144560 -297320
rect 146120 -297380 146140 -297320
rect 144540 -297400 146140 -297380
rect 147540 -297320 149140 -297300
rect 147540 -297380 147560 -297320
rect 149120 -297380 149140 -297320
rect 147540 -297400 149140 -297380
rect 150540 -297320 152140 -297300
rect 150540 -297380 150560 -297320
rect 152120 -297380 152140 -297320
rect 150540 -297400 152140 -297380
rect 153540 -297320 155140 -297300
rect 153540 -297380 153560 -297320
rect 155120 -297380 155140 -297320
rect 153540 -297400 155140 -297380
rect 156540 -297320 158140 -297300
rect 156540 -297380 156560 -297320
rect 158120 -297380 158140 -297320
rect 156540 -297400 158140 -297380
rect 159540 -297320 161140 -297300
rect 159540 -297380 159560 -297320
rect 161120 -297380 161140 -297320
rect 159540 -297400 161140 -297380
rect 162540 -297320 164140 -297300
rect 162540 -297380 162560 -297320
rect 164120 -297380 164140 -297320
rect 162540 -297400 164140 -297380
rect 165540 -297320 167140 -297300
rect 165540 -297380 165560 -297320
rect 167120 -297380 167140 -297320
rect 165540 -297400 167140 -297380
rect 168540 -297320 170140 -297300
rect 168540 -297380 168560 -297320
rect 170120 -297380 170140 -297320
rect 168540 -297400 170140 -297380
rect 171540 -297320 173140 -297300
rect 171540 -297380 171560 -297320
rect 173120 -297380 173140 -297320
rect 171540 -297400 173140 -297380
rect 174540 -297320 176140 -297300
rect 174540 -297380 174560 -297320
rect 176120 -297380 176140 -297320
rect 174540 -297400 176140 -297380
rect 177540 -297320 179140 -297300
rect 177540 -297380 177560 -297320
rect 179120 -297380 179140 -297320
rect 177540 -297400 179140 -297380
rect 180540 -297320 182140 -297300
rect 180540 -297380 180560 -297320
rect 182120 -297380 182140 -297320
rect 180540 -297400 182140 -297380
rect 183540 -297320 185140 -297300
rect 183540 -297380 183560 -297320
rect 185120 -297380 185140 -297320
rect 183540 -297400 185140 -297380
rect 186540 -297320 188140 -297300
rect 186540 -297380 186560 -297320
rect 188120 -297380 188140 -297320
rect 186540 -297400 188140 -297380
rect 189540 -297320 191140 -297300
rect 189540 -297380 189560 -297320
rect 191120 -297380 191140 -297320
rect 189540 -297400 191140 -297380
rect 192540 -297320 194140 -297300
rect 192540 -297380 192560 -297320
rect 194120 -297380 194140 -297320
rect 192540 -297400 194140 -297380
rect 195540 -297320 197140 -297300
rect 195540 -297380 195560 -297320
rect 197120 -297380 197140 -297320
rect 195540 -297400 197140 -297380
rect 198540 -297320 200140 -297300
rect 198540 -297380 198560 -297320
rect 200120 -297380 200140 -297320
rect 198540 -297400 200140 -297380
rect 201540 -297320 203140 -297300
rect 201540 -297380 201560 -297320
rect 203120 -297380 203140 -297320
rect 201540 -297400 203140 -297380
rect 204540 -297320 206140 -297300
rect 204540 -297380 204560 -297320
rect 206120 -297380 206140 -297320
rect 204540 -297400 206140 -297380
rect 207540 -297320 209140 -297300
rect 207540 -297380 207560 -297320
rect 209120 -297380 209140 -297320
rect 207540 -297400 209140 -297380
rect 210540 -297320 212140 -297300
rect 210540 -297380 210560 -297320
rect 212120 -297380 212140 -297320
rect 210540 -297400 212140 -297380
rect 213540 -297320 215140 -297300
rect 213540 -297380 213560 -297320
rect 215120 -297380 215140 -297320
rect 213540 -297400 215140 -297380
rect 216540 -297320 218140 -297300
rect 216540 -297380 216560 -297320
rect 218120 -297380 218140 -297320
rect 216540 -297400 218140 -297380
rect 219540 -297320 221140 -297300
rect 219540 -297380 219560 -297320
rect 221120 -297380 221140 -297320
rect 219540 -297400 221140 -297380
rect 222540 -297320 224140 -297300
rect 222540 -297380 222560 -297320
rect 224120 -297380 224140 -297320
rect 222540 -297400 224140 -297380
rect 225540 -297320 227140 -297300
rect 225540 -297380 225560 -297320
rect 227120 -297380 227140 -297320
rect 225540 -297400 227140 -297380
rect 228540 -297320 230140 -297300
rect 228540 -297380 228560 -297320
rect 230120 -297380 230140 -297320
rect 228540 -297400 230140 -297380
rect 231540 -297320 233140 -297300
rect 231540 -297380 231560 -297320
rect 233120 -297380 233140 -297320
rect 231540 -297400 233140 -297380
rect 234540 -297320 236140 -297300
rect 234540 -297380 234560 -297320
rect 236120 -297380 236140 -297320
rect 234540 -297400 236140 -297380
rect 237540 -297320 239140 -297300
rect 237540 -297380 237560 -297320
rect 239120 -297380 239140 -297320
rect 237540 -297400 239140 -297380
rect 240540 -297320 242140 -297300
rect 240540 -297380 240560 -297320
rect 242120 -297380 242140 -297320
rect 240540 -297400 242140 -297380
rect 243540 -297320 245140 -297300
rect 243540 -297380 243560 -297320
rect 245120 -297380 245140 -297320
rect 243540 -297400 245140 -297380
rect 246540 -297320 248140 -297300
rect 246540 -297380 246560 -297320
rect 248120 -297380 248140 -297320
rect 246540 -297400 248140 -297380
rect 249540 -297320 251140 -297300
rect 249540 -297380 249560 -297320
rect 251120 -297380 251140 -297320
rect 249540 -297400 251140 -297380
rect 252540 -297320 254140 -297300
rect 252540 -297380 252560 -297320
rect 254120 -297380 254140 -297320
rect 252540 -297400 254140 -297380
rect 255540 -297320 257140 -297300
rect 255540 -297380 255560 -297320
rect 257120 -297380 257140 -297320
rect 255540 -297400 257140 -297380
rect 258540 -297320 260140 -297300
rect 258540 -297380 258560 -297320
rect 260120 -297380 260140 -297320
rect 258540 -297400 260140 -297380
rect 261540 -297320 263140 -297300
rect 261540 -297380 261560 -297320
rect 263120 -297380 263140 -297320
rect 261540 -297400 263140 -297380
rect 264540 -297320 266140 -297300
rect 264540 -297380 264560 -297320
rect 266120 -297380 266140 -297320
rect 264540 -297400 266140 -297380
rect 267540 -297320 269140 -297300
rect 267540 -297380 267560 -297320
rect 269120 -297380 269140 -297320
rect 267540 -297400 269140 -297380
rect 270540 -297320 272140 -297300
rect 270540 -297380 270560 -297320
rect 272120 -297380 272140 -297320
rect 270540 -297400 272140 -297380
rect 273540 -297320 275140 -297300
rect 273540 -297380 273560 -297320
rect 275120 -297380 275140 -297320
rect 273540 -297400 275140 -297380
rect 276540 -297320 278140 -297300
rect 276540 -297380 276560 -297320
rect 278120 -297380 278140 -297320
rect 276540 -297400 278140 -297380
rect 279540 -297320 281140 -297300
rect 279540 -297380 279560 -297320
rect 281120 -297380 281140 -297320
rect 279540 -297400 281140 -297380
rect 282540 -297320 284140 -297300
rect 282540 -297380 282560 -297320
rect 284120 -297380 284140 -297320
rect 282540 -297400 284140 -297380
rect 285540 -297320 287140 -297300
rect 285540 -297380 285560 -297320
rect 287120 -297380 287140 -297320
rect 285540 -297400 287140 -297380
rect 288540 -297320 290140 -297300
rect 288540 -297380 288560 -297320
rect 290120 -297380 290140 -297320
rect 288540 -297400 290140 -297380
rect 291540 -297320 293140 -297300
rect 291540 -297380 291560 -297320
rect 293120 -297380 293140 -297320
rect 291540 -297400 293140 -297380
rect 294540 -297320 296140 -297300
rect 294540 -297380 294560 -297320
rect 296120 -297380 296140 -297320
rect 294540 -297400 296140 -297380
rect 297540 -297320 299140 -297300
rect 297540 -297380 297560 -297320
rect 299120 -297380 299140 -297320
rect 297540 -297400 299140 -297380
rect 540 -297830 2140 -297800
rect 540 -297870 560 -297830
rect 2120 -297870 2140 -297830
rect 540 -297880 2140 -297870
rect 3540 -297830 5140 -297800
rect 3540 -297870 3560 -297830
rect 5120 -297870 5140 -297830
rect 3540 -297880 5140 -297870
rect 6540 -297830 8140 -297800
rect 6540 -297870 6560 -297830
rect 8120 -297870 8140 -297830
rect 6540 -297880 8140 -297870
rect 9540 -297830 11140 -297800
rect 9540 -297870 9560 -297830
rect 11120 -297870 11140 -297830
rect 9540 -297880 11140 -297870
rect 12540 -297830 14140 -297800
rect 12540 -297870 12560 -297830
rect 14120 -297870 14140 -297830
rect 12540 -297880 14140 -297870
rect 15540 -297830 17140 -297800
rect 15540 -297870 15560 -297830
rect 17120 -297870 17140 -297830
rect 15540 -297880 17140 -297870
rect 18540 -297830 20140 -297800
rect 18540 -297870 18560 -297830
rect 20120 -297870 20140 -297830
rect 18540 -297880 20140 -297870
rect 21540 -297830 23140 -297800
rect 21540 -297870 21560 -297830
rect 23120 -297870 23140 -297830
rect 21540 -297880 23140 -297870
rect 24540 -297830 26140 -297800
rect 24540 -297870 24560 -297830
rect 26120 -297870 26140 -297830
rect 24540 -297880 26140 -297870
rect 27540 -297830 29140 -297800
rect 27540 -297870 27560 -297830
rect 29120 -297870 29140 -297830
rect 27540 -297880 29140 -297870
rect 30540 -297830 32140 -297800
rect 30540 -297870 30560 -297830
rect 32120 -297870 32140 -297830
rect 30540 -297880 32140 -297870
rect 33540 -297830 35140 -297800
rect 33540 -297870 33560 -297830
rect 35120 -297870 35140 -297830
rect 33540 -297880 35140 -297870
rect 36540 -297830 38140 -297800
rect 36540 -297870 36560 -297830
rect 38120 -297870 38140 -297830
rect 36540 -297880 38140 -297870
rect 39540 -297830 41140 -297800
rect 39540 -297870 39560 -297830
rect 41120 -297870 41140 -297830
rect 39540 -297880 41140 -297870
rect 42540 -297830 44140 -297800
rect 42540 -297870 42560 -297830
rect 44120 -297870 44140 -297830
rect 42540 -297880 44140 -297870
rect 45540 -297830 47140 -297800
rect 45540 -297870 45560 -297830
rect 47120 -297870 47140 -297830
rect 45540 -297880 47140 -297870
rect 48540 -297830 50140 -297800
rect 48540 -297870 48560 -297830
rect 50120 -297870 50140 -297830
rect 48540 -297880 50140 -297870
rect 51540 -297830 53140 -297800
rect 51540 -297870 51560 -297830
rect 53120 -297870 53140 -297830
rect 51540 -297880 53140 -297870
rect 54540 -297830 56140 -297800
rect 54540 -297870 54560 -297830
rect 56120 -297870 56140 -297830
rect 54540 -297880 56140 -297870
rect 57540 -297830 59140 -297800
rect 57540 -297870 57560 -297830
rect 59120 -297870 59140 -297830
rect 57540 -297880 59140 -297870
rect 60540 -297830 62140 -297800
rect 60540 -297870 60560 -297830
rect 62120 -297870 62140 -297830
rect 60540 -297880 62140 -297870
rect 63540 -297830 65140 -297800
rect 63540 -297870 63560 -297830
rect 65120 -297870 65140 -297830
rect 63540 -297880 65140 -297870
rect 66540 -297830 68140 -297800
rect 66540 -297870 66560 -297830
rect 68120 -297870 68140 -297830
rect 66540 -297880 68140 -297870
rect 69540 -297830 71140 -297800
rect 69540 -297870 69560 -297830
rect 71120 -297870 71140 -297830
rect 69540 -297880 71140 -297870
rect 72540 -297830 74140 -297800
rect 72540 -297870 72560 -297830
rect 74120 -297870 74140 -297830
rect 72540 -297880 74140 -297870
rect 75540 -297830 77140 -297800
rect 75540 -297870 75560 -297830
rect 77120 -297870 77140 -297830
rect 75540 -297880 77140 -297870
rect 78540 -297830 80140 -297800
rect 78540 -297870 78560 -297830
rect 80120 -297870 80140 -297830
rect 78540 -297880 80140 -297870
rect 81540 -297830 83140 -297800
rect 81540 -297870 81560 -297830
rect 83120 -297870 83140 -297830
rect 81540 -297880 83140 -297870
rect 84540 -297830 86140 -297800
rect 84540 -297870 84560 -297830
rect 86120 -297870 86140 -297830
rect 84540 -297880 86140 -297870
rect 87540 -297830 89140 -297800
rect 87540 -297870 87560 -297830
rect 89120 -297870 89140 -297830
rect 87540 -297880 89140 -297870
rect 90540 -297830 92140 -297800
rect 90540 -297870 90560 -297830
rect 92120 -297870 92140 -297830
rect 90540 -297880 92140 -297870
rect 93540 -297830 95140 -297800
rect 93540 -297870 93560 -297830
rect 95120 -297870 95140 -297830
rect 93540 -297880 95140 -297870
rect 96540 -297830 98140 -297800
rect 96540 -297870 96560 -297830
rect 98120 -297870 98140 -297830
rect 96540 -297880 98140 -297870
rect 99540 -297830 101140 -297800
rect 99540 -297870 99560 -297830
rect 101120 -297870 101140 -297830
rect 99540 -297880 101140 -297870
rect 102540 -297830 104140 -297800
rect 102540 -297870 102560 -297830
rect 104120 -297870 104140 -297830
rect 102540 -297880 104140 -297870
rect 105540 -297830 107140 -297800
rect 105540 -297870 105560 -297830
rect 107120 -297870 107140 -297830
rect 105540 -297880 107140 -297870
rect 108540 -297830 110140 -297800
rect 108540 -297870 108560 -297830
rect 110120 -297870 110140 -297830
rect 108540 -297880 110140 -297870
rect 111540 -297830 113140 -297800
rect 111540 -297870 111560 -297830
rect 113120 -297870 113140 -297830
rect 111540 -297880 113140 -297870
rect 114540 -297830 116140 -297800
rect 114540 -297870 114560 -297830
rect 116120 -297870 116140 -297830
rect 114540 -297880 116140 -297870
rect 117540 -297830 119140 -297800
rect 117540 -297870 117560 -297830
rect 119120 -297870 119140 -297830
rect 117540 -297880 119140 -297870
rect 120540 -297830 122140 -297800
rect 120540 -297870 120560 -297830
rect 122120 -297870 122140 -297830
rect 120540 -297880 122140 -297870
rect 123540 -297830 125140 -297800
rect 123540 -297870 123560 -297830
rect 125120 -297870 125140 -297830
rect 123540 -297880 125140 -297870
rect 126540 -297830 128140 -297800
rect 126540 -297870 126560 -297830
rect 128120 -297870 128140 -297830
rect 126540 -297880 128140 -297870
rect 129540 -297830 131140 -297800
rect 129540 -297870 129560 -297830
rect 131120 -297870 131140 -297830
rect 129540 -297880 131140 -297870
rect 132540 -297830 134140 -297800
rect 132540 -297870 132560 -297830
rect 134120 -297870 134140 -297830
rect 132540 -297880 134140 -297870
rect 135540 -297830 137140 -297800
rect 135540 -297870 135560 -297830
rect 137120 -297870 137140 -297830
rect 135540 -297880 137140 -297870
rect 138540 -297830 140140 -297800
rect 138540 -297870 138560 -297830
rect 140120 -297870 140140 -297830
rect 138540 -297880 140140 -297870
rect 141540 -297830 143140 -297800
rect 141540 -297870 141560 -297830
rect 143120 -297870 143140 -297830
rect 141540 -297880 143140 -297870
rect 144540 -297830 146140 -297800
rect 144540 -297870 144560 -297830
rect 146120 -297870 146140 -297830
rect 144540 -297880 146140 -297870
rect 147540 -297830 149140 -297800
rect 147540 -297870 147560 -297830
rect 149120 -297870 149140 -297830
rect 147540 -297880 149140 -297870
rect 150540 -297830 152140 -297800
rect 150540 -297870 150560 -297830
rect 152120 -297870 152140 -297830
rect 150540 -297880 152140 -297870
rect 153540 -297830 155140 -297800
rect 153540 -297870 153560 -297830
rect 155120 -297870 155140 -297830
rect 153540 -297880 155140 -297870
rect 156540 -297830 158140 -297800
rect 156540 -297870 156560 -297830
rect 158120 -297870 158140 -297830
rect 156540 -297880 158140 -297870
rect 159540 -297830 161140 -297800
rect 159540 -297870 159560 -297830
rect 161120 -297870 161140 -297830
rect 159540 -297880 161140 -297870
rect 162540 -297830 164140 -297800
rect 162540 -297870 162560 -297830
rect 164120 -297870 164140 -297830
rect 162540 -297880 164140 -297870
rect 165540 -297830 167140 -297800
rect 165540 -297870 165560 -297830
rect 167120 -297870 167140 -297830
rect 165540 -297880 167140 -297870
rect 168540 -297830 170140 -297800
rect 168540 -297870 168560 -297830
rect 170120 -297870 170140 -297830
rect 168540 -297880 170140 -297870
rect 171540 -297830 173140 -297800
rect 171540 -297870 171560 -297830
rect 173120 -297870 173140 -297830
rect 171540 -297880 173140 -297870
rect 174540 -297830 176140 -297800
rect 174540 -297870 174560 -297830
rect 176120 -297870 176140 -297830
rect 174540 -297880 176140 -297870
rect 177540 -297830 179140 -297800
rect 177540 -297870 177560 -297830
rect 179120 -297870 179140 -297830
rect 177540 -297880 179140 -297870
rect 180540 -297830 182140 -297800
rect 180540 -297870 180560 -297830
rect 182120 -297870 182140 -297830
rect 180540 -297880 182140 -297870
rect 183540 -297830 185140 -297800
rect 183540 -297870 183560 -297830
rect 185120 -297870 185140 -297830
rect 183540 -297880 185140 -297870
rect 186540 -297830 188140 -297800
rect 186540 -297870 186560 -297830
rect 188120 -297870 188140 -297830
rect 186540 -297880 188140 -297870
rect 189540 -297830 191140 -297800
rect 189540 -297870 189560 -297830
rect 191120 -297870 191140 -297830
rect 189540 -297880 191140 -297870
rect 192540 -297830 194140 -297800
rect 192540 -297870 192560 -297830
rect 194120 -297870 194140 -297830
rect 192540 -297880 194140 -297870
rect 195540 -297830 197140 -297800
rect 195540 -297870 195560 -297830
rect 197120 -297870 197140 -297830
rect 195540 -297880 197140 -297870
rect 198540 -297830 200140 -297800
rect 198540 -297870 198560 -297830
rect 200120 -297870 200140 -297830
rect 198540 -297880 200140 -297870
rect 201540 -297830 203140 -297800
rect 201540 -297870 201560 -297830
rect 203120 -297870 203140 -297830
rect 201540 -297880 203140 -297870
rect 204540 -297830 206140 -297800
rect 204540 -297870 204560 -297830
rect 206120 -297870 206140 -297830
rect 204540 -297880 206140 -297870
rect 207540 -297830 209140 -297800
rect 207540 -297870 207560 -297830
rect 209120 -297870 209140 -297830
rect 207540 -297880 209140 -297870
rect 210540 -297830 212140 -297800
rect 210540 -297870 210560 -297830
rect 212120 -297870 212140 -297830
rect 210540 -297880 212140 -297870
rect 213540 -297830 215140 -297800
rect 213540 -297870 213560 -297830
rect 215120 -297870 215140 -297830
rect 213540 -297880 215140 -297870
rect 216540 -297830 218140 -297800
rect 216540 -297870 216560 -297830
rect 218120 -297870 218140 -297830
rect 216540 -297880 218140 -297870
rect 219540 -297830 221140 -297800
rect 219540 -297870 219560 -297830
rect 221120 -297870 221140 -297830
rect 219540 -297880 221140 -297870
rect 222540 -297830 224140 -297800
rect 222540 -297870 222560 -297830
rect 224120 -297870 224140 -297830
rect 222540 -297880 224140 -297870
rect 225540 -297830 227140 -297800
rect 225540 -297870 225560 -297830
rect 227120 -297870 227140 -297830
rect 225540 -297880 227140 -297870
rect 228540 -297830 230140 -297800
rect 228540 -297870 228560 -297830
rect 230120 -297870 230140 -297830
rect 228540 -297880 230140 -297870
rect 231540 -297830 233140 -297800
rect 231540 -297870 231560 -297830
rect 233120 -297870 233140 -297830
rect 231540 -297880 233140 -297870
rect 234540 -297830 236140 -297800
rect 234540 -297870 234560 -297830
rect 236120 -297870 236140 -297830
rect 234540 -297880 236140 -297870
rect 237540 -297830 239140 -297800
rect 237540 -297870 237560 -297830
rect 239120 -297870 239140 -297830
rect 237540 -297880 239140 -297870
rect 240540 -297830 242140 -297800
rect 240540 -297870 240560 -297830
rect 242120 -297870 242140 -297830
rect 240540 -297880 242140 -297870
rect 243540 -297830 245140 -297800
rect 243540 -297870 243560 -297830
rect 245120 -297870 245140 -297830
rect 243540 -297880 245140 -297870
rect 246540 -297830 248140 -297800
rect 246540 -297870 246560 -297830
rect 248120 -297870 248140 -297830
rect 246540 -297880 248140 -297870
rect 249540 -297830 251140 -297800
rect 249540 -297870 249560 -297830
rect 251120 -297870 251140 -297830
rect 249540 -297880 251140 -297870
rect 252540 -297830 254140 -297800
rect 252540 -297870 252560 -297830
rect 254120 -297870 254140 -297830
rect 252540 -297880 254140 -297870
rect 255540 -297830 257140 -297800
rect 255540 -297870 255560 -297830
rect 257120 -297870 257140 -297830
rect 255540 -297880 257140 -297870
rect 258540 -297830 260140 -297800
rect 258540 -297870 258560 -297830
rect 260120 -297870 260140 -297830
rect 258540 -297880 260140 -297870
rect 261540 -297830 263140 -297800
rect 261540 -297870 261560 -297830
rect 263120 -297870 263140 -297830
rect 261540 -297880 263140 -297870
rect 264540 -297830 266140 -297800
rect 264540 -297870 264560 -297830
rect 266120 -297870 266140 -297830
rect 264540 -297880 266140 -297870
rect 267540 -297830 269140 -297800
rect 267540 -297870 267560 -297830
rect 269120 -297870 269140 -297830
rect 267540 -297880 269140 -297870
rect 270540 -297830 272140 -297800
rect 270540 -297870 270560 -297830
rect 272120 -297870 272140 -297830
rect 270540 -297880 272140 -297870
rect 273540 -297830 275140 -297800
rect 273540 -297870 273560 -297830
rect 275120 -297870 275140 -297830
rect 273540 -297880 275140 -297870
rect 276540 -297830 278140 -297800
rect 276540 -297870 276560 -297830
rect 278120 -297870 278140 -297830
rect 276540 -297880 278140 -297870
rect 279540 -297830 281140 -297800
rect 279540 -297870 279560 -297830
rect 281120 -297870 281140 -297830
rect 279540 -297880 281140 -297870
rect 282540 -297830 284140 -297800
rect 282540 -297870 282560 -297830
rect 284120 -297870 284140 -297830
rect 282540 -297880 284140 -297870
rect 285540 -297830 287140 -297800
rect 285540 -297870 285560 -297830
rect 287120 -297870 287140 -297830
rect 285540 -297880 287140 -297870
rect 288540 -297830 290140 -297800
rect 288540 -297870 288560 -297830
rect 290120 -297870 290140 -297830
rect 288540 -297880 290140 -297870
rect 291540 -297830 293140 -297800
rect 291540 -297870 291560 -297830
rect 293120 -297870 293140 -297830
rect 291540 -297880 293140 -297870
rect 294540 -297830 296140 -297800
rect 294540 -297870 294560 -297830
rect 296120 -297870 296140 -297830
rect 294540 -297880 296140 -297870
rect 297540 -297830 299140 -297800
rect 297540 -297870 297560 -297830
rect 299120 -297870 299140 -297830
rect 297540 -297880 299140 -297870
<< ndiffc >>
rect 560 -297380 2120 -297320
rect 3560 -297380 5120 -297320
rect 6560 -297380 8120 -297320
rect 9560 -297380 11120 -297320
rect 12560 -297380 14120 -297320
rect 15560 -297380 17120 -297320
rect 18560 -297380 20120 -297320
rect 21560 -297380 23120 -297320
rect 24560 -297380 26120 -297320
rect 27560 -297380 29120 -297320
rect 30560 -297380 32120 -297320
rect 33560 -297380 35120 -297320
rect 36560 -297380 38120 -297320
rect 39560 -297380 41120 -297320
rect 42560 -297380 44120 -297320
rect 45560 -297380 47120 -297320
rect 48560 -297380 50120 -297320
rect 51560 -297380 53120 -297320
rect 54560 -297380 56120 -297320
rect 57560 -297380 59120 -297320
rect 60560 -297380 62120 -297320
rect 63560 -297380 65120 -297320
rect 66560 -297380 68120 -297320
rect 69560 -297380 71120 -297320
rect 72560 -297380 74120 -297320
rect 75560 -297380 77120 -297320
rect 78560 -297380 80120 -297320
rect 81560 -297380 83120 -297320
rect 84560 -297380 86120 -297320
rect 87560 -297380 89120 -297320
rect 90560 -297380 92120 -297320
rect 93560 -297380 95120 -297320
rect 96560 -297380 98120 -297320
rect 99560 -297380 101120 -297320
rect 102560 -297380 104120 -297320
rect 105560 -297380 107120 -297320
rect 108560 -297380 110120 -297320
rect 111560 -297380 113120 -297320
rect 114560 -297380 116120 -297320
rect 117560 -297380 119120 -297320
rect 120560 -297380 122120 -297320
rect 123560 -297380 125120 -297320
rect 126560 -297380 128120 -297320
rect 129560 -297380 131120 -297320
rect 132560 -297380 134120 -297320
rect 135560 -297380 137120 -297320
rect 138560 -297380 140120 -297320
rect 141560 -297380 143120 -297320
rect 144560 -297380 146120 -297320
rect 147560 -297380 149120 -297320
rect 150560 -297380 152120 -297320
rect 153560 -297380 155120 -297320
rect 156560 -297380 158120 -297320
rect 159560 -297380 161120 -297320
rect 162560 -297380 164120 -297320
rect 165560 -297380 167120 -297320
rect 168560 -297380 170120 -297320
rect 171560 -297380 173120 -297320
rect 174560 -297380 176120 -297320
rect 177560 -297380 179120 -297320
rect 180560 -297380 182120 -297320
rect 183560 -297380 185120 -297320
rect 186560 -297380 188120 -297320
rect 189560 -297380 191120 -297320
rect 192560 -297380 194120 -297320
rect 195560 -297380 197120 -297320
rect 198560 -297380 200120 -297320
rect 201560 -297380 203120 -297320
rect 204560 -297380 206120 -297320
rect 207560 -297380 209120 -297320
rect 210560 -297380 212120 -297320
rect 213560 -297380 215120 -297320
rect 216560 -297380 218120 -297320
rect 219560 -297380 221120 -297320
rect 222560 -297380 224120 -297320
rect 225560 -297380 227120 -297320
rect 228560 -297380 230120 -297320
rect 231560 -297380 233120 -297320
rect 234560 -297380 236120 -297320
rect 237560 -297380 239120 -297320
rect 240560 -297380 242120 -297320
rect 243560 -297380 245120 -297320
rect 246560 -297380 248120 -297320
rect 249560 -297380 251120 -297320
rect 252560 -297380 254120 -297320
rect 255560 -297380 257120 -297320
rect 258560 -297380 260120 -297320
rect 261560 -297380 263120 -297320
rect 264560 -297380 266120 -297320
rect 267560 -297380 269120 -297320
rect 270560 -297380 272120 -297320
rect 273560 -297380 275120 -297320
rect 276560 -297380 278120 -297320
rect 279560 -297380 281120 -297320
rect 282560 -297380 284120 -297320
rect 285560 -297380 287120 -297320
rect 288560 -297380 290120 -297320
rect 291560 -297380 293120 -297320
rect 294560 -297380 296120 -297320
rect 297560 -297380 299120 -297320
rect 560 -297870 2120 -297830
rect 3560 -297870 5120 -297830
rect 6560 -297870 8120 -297830
rect 9560 -297870 11120 -297830
rect 12560 -297870 14120 -297830
rect 15560 -297870 17120 -297830
rect 18560 -297870 20120 -297830
rect 21560 -297870 23120 -297830
rect 24560 -297870 26120 -297830
rect 27560 -297870 29120 -297830
rect 30560 -297870 32120 -297830
rect 33560 -297870 35120 -297830
rect 36560 -297870 38120 -297830
rect 39560 -297870 41120 -297830
rect 42560 -297870 44120 -297830
rect 45560 -297870 47120 -297830
rect 48560 -297870 50120 -297830
rect 51560 -297870 53120 -297830
rect 54560 -297870 56120 -297830
rect 57560 -297870 59120 -297830
rect 60560 -297870 62120 -297830
rect 63560 -297870 65120 -297830
rect 66560 -297870 68120 -297830
rect 69560 -297870 71120 -297830
rect 72560 -297870 74120 -297830
rect 75560 -297870 77120 -297830
rect 78560 -297870 80120 -297830
rect 81560 -297870 83120 -297830
rect 84560 -297870 86120 -297830
rect 87560 -297870 89120 -297830
rect 90560 -297870 92120 -297830
rect 93560 -297870 95120 -297830
rect 96560 -297870 98120 -297830
rect 99560 -297870 101120 -297830
rect 102560 -297870 104120 -297830
rect 105560 -297870 107120 -297830
rect 108560 -297870 110120 -297830
rect 111560 -297870 113120 -297830
rect 114560 -297870 116120 -297830
rect 117560 -297870 119120 -297830
rect 120560 -297870 122120 -297830
rect 123560 -297870 125120 -297830
rect 126560 -297870 128120 -297830
rect 129560 -297870 131120 -297830
rect 132560 -297870 134120 -297830
rect 135560 -297870 137120 -297830
rect 138560 -297870 140120 -297830
rect 141560 -297870 143120 -297830
rect 144560 -297870 146120 -297830
rect 147560 -297870 149120 -297830
rect 150560 -297870 152120 -297830
rect 153560 -297870 155120 -297830
rect 156560 -297870 158120 -297830
rect 159560 -297870 161120 -297830
rect 162560 -297870 164120 -297830
rect 165560 -297870 167120 -297830
rect 168560 -297870 170120 -297830
rect 171560 -297870 173120 -297830
rect 174560 -297870 176120 -297830
rect 177560 -297870 179120 -297830
rect 180560 -297870 182120 -297830
rect 183560 -297870 185120 -297830
rect 186560 -297870 188120 -297830
rect 189560 -297870 191120 -297830
rect 192560 -297870 194120 -297830
rect 195560 -297870 197120 -297830
rect 198560 -297870 200120 -297830
rect 201560 -297870 203120 -297830
rect 204560 -297870 206120 -297830
rect 207560 -297870 209120 -297830
rect 210560 -297870 212120 -297830
rect 213560 -297870 215120 -297830
rect 216560 -297870 218120 -297830
rect 219560 -297870 221120 -297830
rect 222560 -297870 224120 -297830
rect 225560 -297870 227120 -297830
rect 228560 -297870 230120 -297830
rect 231560 -297870 233120 -297830
rect 234560 -297870 236120 -297830
rect 237560 -297870 239120 -297830
rect 240560 -297870 242120 -297830
rect 243560 -297870 245120 -297830
rect 246560 -297870 248120 -297830
rect 249560 -297870 251120 -297830
rect 252560 -297870 254120 -297830
rect 255560 -297870 257120 -297830
rect 258560 -297870 260120 -297830
rect 261560 -297870 263120 -297830
rect 264560 -297870 266120 -297830
rect 267560 -297870 269120 -297830
rect 270560 -297870 272120 -297830
rect 273560 -297870 275120 -297830
rect 276560 -297870 278120 -297830
rect 279560 -297870 281120 -297830
rect 282560 -297870 284120 -297830
rect 285560 -297870 287120 -297830
rect 288560 -297870 290120 -297830
rect 291560 -297870 293120 -297830
rect 294560 -297870 296120 -297830
rect 297560 -297870 299120 -297830
<< poly >>
rect 510 -297490 540 -297400
rect 220 -297500 540 -297490
rect 220 -297700 240 -297500
rect 420 -297700 540 -297500
rect 220 -297710 540 -297700
rect 510 -297800 540 -297710
rect 2140 -297800 2170 -297400
rect 3510 -297490 3540 -297400
rect 3220 -297500 3540 -297490
rect 3220 -297700 3240 -297500
rect 3420 -297700 3540 -297500
rect 3220 -297710 3540 -297700
rect 3510 -297800 3540 -297710
rect 5140 -297800 5170 -297400
rect 6510 -297490 6540 -297400
rect 6220 -297500 6540 -297490
rect 6220 -297700 6240 -297500
rect 6420 -297700 6540 -297500
rect 6220 -297710 6540 -297700
rect 6510 -297800 6540 -297710
rect 8140 -297800 8170 -297400
rect 9510 -297490 9540 -297400
rect 9220 -297500 9540 -297490
rect 9220 -297700 9240 -297500
rect 9420 -297700 9540 -297500
rect 9220 -297710 9540 -297700
rect 9510 -297800 9540 -297710
rect 11140 -297800 11170 -297400
rect 12510 -297490 12540 -297400
rect 12220 -297500 12540 -297490
rect 12220 -297700 12240 -297500
rect 12420 -297700 12540 -297500
rect 12220 -297710 12540 -297700
rect 12510 -297800 12540 -297710
rect 14140 -297800 14170 -297400
rect 15510 -297490 15540 -297400
rect 15220 -297500 15540 -297490
rect 15220 -297700 15240 -297500
rect 15420 -297700 15540 -297500
rect 15220 -297710 15540 -297700
rect 15510 -297800 15540 -297710
rect 17140 -297800 17170 -297400
rect 18510 -297490 18540 -297400
rect 18220 -297500 18540 -297490
rect 18220 -297700 18240 -297500
rect 18420 -297700 18540 -297500
rect 18220 -297710 18540 -297700
rect 18510 -297800 18540 -297710
rect 20140 -297800 20170 -297400
rect 21510 -297490 21540 -297400
rect 21220 -297500 21540 -297490
rect 21220 -297700 21240 -297500
rect 21420 -297700 21540 -297500
rect 21220 -297710 21540 -297700
rect 21510 -297800 21540 -297710
rect 23140 -297800 23170 -297400
rect 24510 -297490 24540 -297400
rect 24220 -297500 24540 -297490
rect 24220 -297700 24240 -297500
rect 24420 -297700 24540 -297500
rect 24220 -297710 24540 -297700
rect 24510 -297800 24540 -297710
rect 26140 -297800 26170 -297400
rect 27510 -297490 27540 -297400
rect 27220 -297500 27540 -297490
rect 27220 -297700 27240 -297500
rect 27420 -297700 27540 -297500
rect 27220 -297710 27540 -297700
rect 27510 -297800 27540 -297710
rect 29140 -297800 29170 -297400
rect 30510 -297490 30540 -297400
rect 30220 -297500 30540 -297490
rect 30220 -297700 30240 -297500
rect 30420 -297700 30540 -297500
rect 30220 -297710 30540 -297700
rect 30510 -297800 30540 -297710
rect 32140 -297800 32170 -297400
rect 33510 -297490 33540 -297400
rect 33220 -297500 33540 -297490
rect 33220 -297700 33240 -297500
rect 33420 -297700 33540 -297500
rect 33220 -297710 33540 -297700
rect 33510 -297800 33540 -297710
rect 35140 -297800 35170 -297400
rect 36510 -297490 36540 -297400
rect 36220 -297500 36540 -297490
rect 36220 -297700 36240 -297500
rect 36420 -297700 36540 -297500
rect 36220 -297710 36540 -297700
rect 36510 -297800 36540 -297710
rect 38140 -297800 38170 -297400
rect 39510 -297490 39540 -297400
rect 39220 -297500 39540 -297490
rect 39220 -297700 39240 -297500
rect 39420 -297700 39540 -297500
rect 39220 -297710 39540 -297700
rect 39510 -297800 39540 -297710
rect 41140 -297800 41170 -297400
rect 42510 -297490 42540 -297400
rect 42220 -297500 42540 -297490
rect 42220 -297700 42240 -297500
rect 42420 -297700 42540 -297500
rect 42220 -297710 42540 -297700
rect 42510 -297800 42540 -297710
rect 44140 -297800 44170 -297400
rect 45510 -297490 45540 -297400
rect 45220 -297500 45540 -297490
rect 45220 -297700 45240 -297500
rect 45420 -297700 45540 -297500
rect 45220 -297710 45540 -297700
rect 45510 -297800 45540 -297710
rect 47140 -297800 47170 -297400
rect 48510 -297490 48540 -297400
rect 48220 -297500 48540 -297490
rect 48220 -297700 48240 -297500
rect 48420 -297700 48540 -297500
rect 48220 -297710 48540 -297700
rect 48510 -297800 48540 -297710
rect 50140 -297800 50170 -297400
rect 51510 -297490 51540 -297400
rect 51220 -297500 51540 -297490
rect 51220 -297700 51240 -297500
rect 51420 -297700 51540 -297500
rect 51220 -297710 51540 -297700
rect 51510 -297800 51540 -297710
rect 53140 -297800 53170 -297400
rect 54510 -297490 54540 -297400
rect 54220 -297500 54540 -297490
rect 54220 -297700 54240 -297500
rect 54420 -297700 54540 -297500
rect 54220 -297710 54540 -297700
rect 54510 -297800 54540 -297710
rect 56140 -297800 56170 -297400
rect 57510 -297490 57540 -297400
rect 57220 -297500 57540 -297490
rect 57220 -297700 57240 -297500
rect 57420 -297700 57540 -297500
rect 57220 -297710 57540 -297700
rect 57510 -297800 57540 -297710
rect 59140 -297800 59170 -297400
rect 60510 -297490 60540 -297400
rect 60220 -297500 60540 -297490
rect 60220 -297700 60240 -297500
rect 60420 -297700 60540 -297500
rect 60220 -297710 60540 -297700
rect 60510 -297800 60540 -297710
rect 62140 -297800 62170 -297400
rect 63510 -297490 63540 -297400
rect 63220 -297500 63540 -297490
rect 63220 -297700 63240 -297500
rect 63420 -297700 63540 -297500
rect 63220 -297710 63540 -297700
rect 63510 -297800 63540 -297710
rect 65140 -297800 65170 -297400
rect 66510 -297490 66540 -297400
rect 66220 -297500 66540 -297490
rect 66220 -297700 66240 -297500
rect 66420 -297700 66540 -297500
rect 66220 -297710 66540 -297700
rect 66510 -297800 66540 -297710
rect 68140 -297800 68170 -297400
rect 69510 -297490 69540 -297400
rect 69220 -297500 69540 -297490
rect 69220 -297700 69240 -297500
rect 69420 -297700 69540 -297500
rect 69220 -297710 69540 -297700
rect 69510 -297800 69540 -297710
rect 71140 -297800 71170 -297400
rect 72510 -297490 72540 -297400
rect 72220 -297500 72540 -297490
rect 72220 -297700 72240 -297500
rect 72420 -297700 72540 -297500
rect 72220 -297710 72540 -297700
rect 72510 -297800 72540 -297710
rect 74140 -297800 74170 -297400
rect 75510 -297490 75540 -297400
rect 75220 -297500 75540 -297490
rect 75220 -297700 75240 -297500
rect 75420 -297700 75540 -297500
rect 75220 -297710 75540 -297700
rect 75510 -297800 75540 -297710
rect 77140 -297800 77170 -297400
rect 78510 -297490 78540 -297400
rect 78220 -297500 78540 -297490
rect 78220 -297700 78240 -297500
rect 78420 -297700 78540 -297500
rect 78220 -297710 78540 -297700
rect 78510 -297800 78540 -297710
rect 80140 -297800 80170 -297400
rect 81510 -297490 81540 -297400
rect 81220 -297500 81540 -297490
rect 81220 -297700 81240 -297500
rect 81420 -297700 81540 -297500
rect 81220 -297710 81540 -297700
rect 81510 -297800 81540 -297710
rect 83140 -297800 83170 -297400
rect 84510 -297490 84540 -297400
rect 84220 -297500 84540 -297490
rect 84220 -297700 84240 -297500
rect 84420 -297700 84540 -297500
rect 84220 -297710 84540 -297700
rect 84510 -297800 84540 -297710
rect 86140 -297800 86170 -297400
rect 87510 -297490 87540 -297400
rect 87220 -297500 87540 -297490
rect 87220 -297700 87240 -297500
rect 87420 -297700 87540 -297500
rect 87220 -297710 87540 -297700
rect 87510 -297800 87540 -297710
rect 89140 -297800 89170 -297400
rect 90510 -297490 90540 -297400
rect 90220 -297500 90540 -297490
rect 90220 -297700 90240 -297500
rect 90420 -297700 90540 -297500
rect 90220 -297710 90540 -297700
rect 90510 -297800 90540 -297710
rect 92140 -297800 92170 -297400
rect 93510 -297490 93540 -297400
rect 93220 -297500 93540 -297490
rect 93220 -297700 93240 -297500
rect 93420 -297700 93540 -297500
rect 93220 -297710 93540 -297700
rect 93510 -297800 93540 -297710
rect 95140 -297800 95170 -297400
rect 96510 -297490 96540 -297400
rect 96220 -297500 96540 -297490
rect 96220 -297700 96240 -297500
rect 96420 -297700 96540 -297500
rect 96220 -297710 96540 -297700
rect 96510 -297800 96540 -297710
rect 98140 -297800 98170 -297400
rect 99510 -297490 99540 -297400
rect 99220 -297500 99540 -297490
rect 99220 -297700 99240 -297500
rect 99420 -297700 99540 -297500
rect 99220 -297710 99540 -297700
rect 99510 -297800 99540 -297710
rect 101140 -297800 101170 -297400
rect 102510 -297490 102540 -297400
rect 102220 -297500 102540 -297490
rect 102220 -297700 102240 -297500
rect 102420 -297700 102540 -297500
rect 102220 -297710 102540 -297700
rect 102510 -297800 102540 -297710
rect 104140 -297800 104170 -297400
rect 105510 -297490 105540 -297400
rect 105220 -297500 105540 -297490
rect 105220 -297700 105240 -297500
rect 105420 -297700 105540 -297500
rect 105220 -297710 105540 -297700
rect 105510 -297800 105540 -297710
rect 107140 -297800 107170 -297400
rect 108510 -297490 108540 -297400
rect 108220 -297500 108540 -297490
rect 108220 -297700 108240 -297500
rect 108420 -297700 108540 -297500
rect 108220 -297710 108540 -297700
rect 108510 -297800 108540 -297710
rect 110140 -297800 110170 -297400
rect 111510 -297490 111540 -297400
rect 111220 -297500 111540 -297490
rect 111220 -297700 111240 -297500
rect 111420 -297700 111540 -297500
rect 111220 -297710 111540 -297700
rect 111510 -297800 111540 -297710
rect 113140 -297800 113170 -297400
rect 114510 -297490 114540 -297400
rect 114220 -297500 114540 -297490
rect 114220 -297700 114240 -297500
rect 114420 -297700 114540 -297500
rect 114220 -297710 114540 -297700
rect 114510 -297800 114540 -297710
rect 116140 -297800 116170 -297400
rect 117510 -297490 117540 -297400
rect 117220 -297500 117540 -297490
rect 117220 -297700 117240 -297500
rect 117420 -297700 117540 -297500
rect 117220 -297710 117540 -297700
rect 117510 -297800 117540 -297710
rect 119140 -297800 119170 -297400
rect 120510 -297490 120540 -297400
rect 120220 -297500 120540 -297490
rect 120220 -297700 120240 -297500
rect 120420 -297700 120540 -297500
rect 120220 -297710 120540 -297700
rect 120510 -297800 120540 -297710
rect 122140 -297800 122170 -297400
rect 123510 -297490 123540 -297400
rect 123220 -297500 123540 -297490
rect 123220 -297700 123240 -297500
rect 123420 -297700 123540 -297500
rect 123220 -297710 123540 -297700
rect 123510 -297800 123540 -297710
rect 125140 -297800 125170 -297400
rect 126510 -297490 126540 -297400
rect 126220 -297500 126540 -297490
rect 126220 -297700 126240 -297500
rect 126420 -297700 126540 -297500
rect 126220 -297710 126540 -297700
rect 126510 -297800 126540 -297710
rect 128140 -297800 128170 -297400
rect 129510 -297490 129540 -297400
rect 129220 -297500 129540 -297490
rect 129220 -297700 129240 -297500
rect 129420 -297700 129540 -297500
rect 129220 -297710 129540 -297700
rect 129510 -297800 129540 -297710
rect 131140 -297800 131170 -297400
rect 132510 -297490 132540 -297400
rect 132220 -297500 132540 -297490
rect 132220 -297700 132240 -297500
rect 132420 -297700 132540 -297500
rect 132220 -297710 132540 -297700
rect 132510 -297800 132540 -297710
rect 134140 -297800 134170 -297400
rect 135510 -297490 135540 -297400
rect 135220 -297500 135540 -297490
rect 135220 -297700 135240 -297500
rect 135420 -297700 135540 -297500
rect 135220 -297710 135540 -297700
rect 135510 -297800 135540 -297710
rect 137140 -297800 137170 -297400
rect 138510 -297490 138540 -297400
rect 138220 -297500 138540 -297490
rect 138220 -297700 138240 -297500
rect 138420 -297700 138540 -297500
rect 138220 -297710 138540 -297700
rect 138510 -297800 138540 -297710
rect 140140 -297800 140170 -297400
rect 141510 -297490 141540 -297400
rect 141220 -297500 141540 -297490
rect 141220 -297700 141240 -297500
rect 141420 -297700 141540 -297500
rect 141220 -297710 141540 -297700
rect 141510 -297800 141540 -297710
rect 143140 -297800 143170 -297400
rect 144510 -297490 144540 -297400
rect 144220 -297500 144540 -297490
rect 144220 -297700 144240 -297500
rect 144420 -297700 144540 -297500
rect 144220 -297710 144540 -297700
rect 144510 -297800 144540 -297710
rect 146140 -297800 146170 -297400
rect 147510 -297490 147540 -297400
rect 147220 -297500 147540 -297490
rect 147220 -297700 147240 -297500
rect 147420 -297700 147540 -297500
rect 147220 -297710 147540 -297700
rect 147510 -297800 147540 -297710
rect 149140 -297800 149170 -297400
rect 150510 -297490 150540 -297400
rect 150220 -297500 150540 -297490
rect 150220 -297700 150240 -297500
rect 150420 -297700 150540 -297500
rect 150220 -297710 150540 -297700
rect 150510 -297800 150540 -297710
rect 152140 -297800 152170 -297400
rect 153510 -297490 153540 -297400
rect 153220 -297500 153540 -297490
rect 153220 -297700 153240 -297500
rect 153420 -297700 153540 -297500
rect 153220 -297710 153540 -297700
rect 153510 -297800 153540 -297710
rect 155140 -297800 155170 -297400
rect 156510 -297490 156540 -297400
rect 156220 -297500 156540 -297490
rect 156220 -297700 156240 -297500
rect 156420 -297700 156540 -297500
rect 156220 -297710 156540 -297700
rect 156510 -297800 156540 -297710
rect 158140 -297800 158170 -297400
rect 159510 -297490 159540 -297400
rect 159220 -297500 159540 -297490
rect 159220 -297700 159240 -297500
rect 159420 -297700 159540 -297500
rect 159220 -297710 159540 -297700
rect 159510 -297800 159540 -297710
rect 161140 -297800 161170 -297400
rect 162510 -297490 162540 -297400
rect 162220 -297500 162540 -297490
rect 162220 -297700 162240 -297500
rect 162420 -297700 162540 -297500
rect 162220 -297710 162540 -297700
rect 162510 -297800 162540 -297710
rect 164140 -297800 164170 -297400
rect 165510 -297490 165540 -297400
rect 165220 -297500 165540 -297490
rect 165220 -297700 165240 -297500
rect 165420 -297700 165540 -297500
rect 165220 -297710 165540 -297700
rect 165510 -297800 165540 -297710
rect 167140 -297800 167170 -297400
rect 168510 -297490 168540 -297400
rect 168220 -297500 168540 -297490
rect 168220 -297700 168240 -297500
rect 168420 -297700 168540 -297500
rect 168220 -297710 168540 -297700
rect 168510 -297800 168540 -297710
rect 170140 -297800 170170 -297400
rect 171510 -297490 171540 -297400
rect 171220 -297500 171540 -297490
rect 171220 -297700 171240 -297500
rect 171420 -297700 171540 -297500
rect 171220 -297710 171540 -297700
rect 171510 -297800 171540 -297710
rect 173140 -297800 173170 -297400
rect 174510 -297490 174540 -297400
rect 174220 -297500 174540 -297490
rect 174220 -297700 174240 -297500
rect 174420 -297700 174540 -297500
rect 174220 -297710 174540 -297700
rect 174510 -297800 174540 -297710
rect 176140 -297800 176170 -297400
rect 177510 -297490 177540 -297400
rect 177220 -297500 177540 -297490
rect 177220 -297700 177240 -297500
rect 177420 -297700 177540 -297500
rect 177220 -297710 177540 -297700
rect 177510 -297800 177540 -297710
rect 179140 -297800 179170 -297400
rect 180510 -297490 180540 -297400
rect 180220 -297500 180540 -297490
rect 180220 -297700 180240 -297500
rect 180420 -297700 180540 -297500
rect 180220 -297710 180540 -297700
rect 180510 -297800 180540 -297710
rect 182140 -297800 182170 -297400
rect 183510 -297490 183540 -297400
rect 183220 -297500 183540 -297490
rect 183220 -297700 183240 -297500
rect 183420 -297700 183540 -297500
rect 183220 -297710 183540 -297700
rect 183510 -297800 183540 -297710
rect 185140 -297800 185170 -297400
rect 186510 -297490 186540 -297400
rect 186220 -297500 186540 -297490
rect 186220 -297700 186240 -297500
rect 186420 -297700 186540 -297500
rect 186220 -297710 186540 -297700
rect 186510 -297800 186540 -297710
rect 188140 -297800 188170 -297400
rect 189510 -297490 189540 -297400
rect 189220 -297500 189540 -297490
rect 189220 -297700 189240 -297500
rect 189420 -297700 189540 -297500
rect 189220 -297710 189540 -297700
rect 189510 -297800 189540 -297710
rect 191140 -297800 191170 -297400
rect 192510 -297490 192540 -297400
rect 192220 -297500 192540 -297490
rect 192220 -297700 192240 -297500
rect 192420 -297700 192540 -297500
rect 192220 -297710 192540 -297700
rect 192510 -297800 192540 -297710
rect 194140 -297800 194170 -297400
rect 195510 -297490 195540 -297400
rect 195220 -297500 195540 -297490
rect 195220 -297700 195240 -297500
rect 195420 -297700 195540 -297500
rect 195220 -297710 195540 -297700
rect 195510 -297800 195540 -297710
rect 197140 -297800 197170 -297400
rect 198510 -297490 198540 -297400
rect 198220 -297500 198540 -297490
rect 198220 -297700 198240 -297500
rect 198420 -297700 198540 -297500
rect 198220 -297710 198540 -297700
rect 198510 -297800 198540 -297710
rect 200140 -297800 200170 -297400
rect 201510 -297490 201540 -297400
rect 201220 -297500 201540 -297490
rect 201220 -297700 201240 -297500
rect 201420 -297700 201540 -297500
rect 201220 -297710 201540 -297700
rect 201510 -297800 201540 -297710
rect 203140 -297800 203170 -297400
rect 204510 -297490 204540 -297400
rect 204220 -297500 204540 -297490
rect 204220 -297700 204240 -297500
rect 204420 -297700 204540 -297500
rect 204220 -297710 204540 -297700
rect 204510 -297800 204540 -297710
rect 206140 -297800 206170 -297400
rect 207510 -297490 207540 -297400
rect 207220 -297500 207540 -297490
rect 207220 -297700 207240 -297500
rect 207420 -297700 207540 -297500
rect 207220 -297710 207540 -297700
rect 207510 -297800 207540 -297710
rect 209140 -297800 209170 -297400
rect 210510 -297490 210540 -297400
rect 210220 -297500 210540 -297490
rect 210220 -297700 210240 -297500
rect 210420 -297700 210540 -297500
rect 210220 -297710 210540 -297700
rect 210510 -297800 210540 -297710
rect 212140 -297800 212170 -297400
rect 213510 -297490 213540 -297400
rect 213220 -297500 213540 -297490
rect 213220 -297700 213240 -297500
rect 213420 -297700 213540 -297500
rect 213220 -297710 213540 -297700
rect 213510 -297800 213540 -297710
rect 215140 -297800 215170 -297400
rect 216510 -297490 216540 -297400
rect 216220 -297500 216540 -297490
rect 216220 -297700 216240 -297500
rect 216420 -297700 216540 -297500
rect 216220 -297710 216540 -297700
rect 216510 -297800 216540 -297710
rect 218140 -297800 218170 -297400
rect 219510 -297490 219540 -297400
rect 219220 -297500 219540 -297490
rect 219220 -297700 219240 -297500
rect 219420 -297700 219540 -297500
rect 219220 -297710 219540 -297700
rect 219510 -297800 219540 -297710
rect 221140 -297800 221170 -297400
rect 222510 -297490 222540 -297400
rect 222220 -297500 222540 -297490
rect 222220 -297700 222240 -297500
rect 222420 -297700 222540 -297500
rect 222220 -297710 222540 -297700
rect 222510 -297800 222540 -297710
rect 224140 -297800 224170 -297400
rect 225510 -297490 225540 -297400
rect 225220 -297500 225540 -297490
rect 225220 -297700 225240 -297500
rect 225420 -297700 225540 -297500
rect 225220 -297710 225540 -297700
rect 225510 -297800 225540 -297710
rect 227140 -297800 227170 -297400
rect 228510 -297490 228540 -297400
rect 228220 -297500 228540 -297490
rect 228220 -297700 228240 -297500
rect 228420 -297700 228540 -297500
rect 228220 -297710 228540 -297700
rect 228510 -297800 228540 -297710
rect 230140 -297800 230170 -297400
rect 231510 -297490 231540 -297400
rect 231220 -297500 231540 -297490
rect 231220 -297700 231240 -297500
rect 231420 -297700 231540 -297500
rect 231220 -297710 231540 -297700
rect 231510 -297800 231540 -297710
rect 233140 -297800 233170 -297400
rect 234510 -297490 234540 -297400
rect 234220 -297500 234540 -297490
rect 234220 -297700 234240 -297500
rect 234420 -297700 234540 -297500
rect 234220 -297710 234540 -297700
rect 234510 -297800 234540 -297710
rect 236140 -297800 236170 -297400
rect 237510 -297490 237540 -297400
rect 237220 -297500 237540 -297490
rect 237220 -297700 237240 -297500
rect 237420 -297700 237540 -297500
rect 237220 -297710 237540 -297700
rect 237510 -297800 237540 -297710
rect 239140 -297800 239170 -297400
rect 240510 -297490 240540 -297400
rect 240220 -297500 240540 -297490
rect 240220 -297700 240240 -297500
rect 240420 -297700 240540 -297500
rect 240220 -297710 240540 -297700
rect 240510 -297800 240540 -297710
rect 242140 -297800 242170 -297400
rect 243510 -297490 243540 -297400
rect 243220 -297500 243540 -297490
rect 243220 -297700 243240 -297500
rect 243420 -297700 243540 -297500
rect 243220 -297710 243540 -297700
rect 243510 -297800 243540 -297710
rect 245140 -297800 245170 -297400
rect 246510 -297490 246540 -297400
rect 246220 -297500 246540 -297490
rect 246220 -297700 246240 -297500
rect 246420 -297700 246540 -297500
rect 246220 -297710 246540 -297700
rect 246510 -297800 246540 -297710
rect 248140 -297800 248170 -297400
rect 249510 -297490 249540 -297400
rect 249220 -297500 249540 -297490
rect 249220 -297700 249240 -297500
rect 249420 -297700 249540 -297500
rect 249220 -297710 249540 -297700
rect 249510 -297800 249540 -297710
rect 251140 -297800 251170 -297400
rect 252510 -297490 252540 -297400
rect 252220 -297500 252540 -297490
rect 252220 -297700 252240 -297500
rect 252420 -297700 252540 -297500
rect 252220 -297710 252540 -297700
rect 252510 -297800 252540 -297710
rect 254140 -297800 254170 -297400
rect 255510 -297490 255540 -297400
rect 255220 -297500 255540 -297490
rect 255220 -297700 255240 -297500
rect 255420 -297700 255540 -297500
rect 255220 -297710 255540 -297700
rect 255510 -297800 255540 -297710
rect 257140 -297800 257170 -297400
rect 258510 -297490 258540 -297400
rect 258220 -297500 258540 -297490
rect 258220 -297700 258240 -297500
rect 258420 -297700 258540 -297500
rect 258220 -297710 258540 -297700
rect 258510 -297800 258540 -297710
rect 260140 -297800 260170 -297400
rect 261510 -297490 261540 -297400
rect 261220 -297500 261540 -297490
rect 261220 -297700 261240 -297500
rect 261420 -297700 261540 -297500
rect 261220 -297710 261540 -297700
rect 261510 -297800 261540 -297710
rect 263140 -297800 263170 -297400
rect 264510 -297490 264540 -297400
rect 264220 -297500 264540 -297490
rect 264220 -297700 264240 -297500
rect 264420 -297700 264540 -297500
rect 264220 -297710 264540 -297700
rect 264510 -297800 264540 -297710
rect 266140 -297800 266170 -297400
rect 267510 -297490 267540 -297400
rect 267220 -297500 267540 -297490
rect 267220 -297700 267240 -297500
rect 267420 -297700 267540 -297500
rect 267220 -297710 267540 -297700
rect 267510 -297800 267540 -297710
rect 269140 -297800 269170 -297400
rect 270510 -297490 270540 -297400
rect 270220 -297500 270540 -297490
rect 270220 -297700 270240 -297500
rect 270420 -297700 270540 -297500
rect 270220 -297710 270540 -297700
rect 270510 -297800 270540 -297710
rect 272140 -297800 272170 -297400
rect 273510 -297490 273540 -297400
rect 273220 -297500 273540 -297490
rect 273220 -297700 273240 -297500
rect 273420 -297700 273540 -297500
rect 273220 -297710 273540 -297700
rect 273510 -297800 273540 -297710
rect 275140 -297800 275170 -297400
rect 276510 -297490 276540 -297400
rect 276220 -297500 276540 -297490
rect 276220 -297700 276240 -297500
rect 276420 -297700 276540 -297500
rect 276220 -297710 276540 -297700
rect 276510 -297800 276540 -297710
rect 278140 -297800 278170 -297400
rect 279510 -297490 279540 -297400
rect 279220 -297500 279540 -297490
rect 279220 -297700 279240 -297500
rect 279420 -297700 279540 -297500
rect 279220 -297710 279540 -297700
rect 279510 -297800 279540 -297710
rect 281140 -297800 281170 -297400
rect 282510 -297490 282540 -297400
rect 282220 -297500 282540 -297490
rect 282220 -297700 282240 -297500
rect 282420 -297700 282540 -297500
rect 282220 -297710 282540 -297700
rect 282510 -297800 282540 -297710
rect 284140 -297800 284170 -297400
rect 285510 -297490 285540 -297400
rect 285220 -297500 285540 -297490
rect 285220 -297700 285240 -297500
rect 285420 -297700 285540 -297500
rect 285220 -297710 285540 -297700
rect 285510 -297800 285540 -297710
rect 287140 -297800 287170 -297400
rect 288510 -297490 288540 -297400
rect 288220 -297500 288540 -297490
rect 288220 -297700 288240 -297500
rect 288420 -297700 288540 -297500
rect 288220 -297710 288540 -297700
rect 288510 -297800 288540 -297710
rect 290140 -297800 290170 -297400
rect 291510 -297490 291540 -297400
rect 291220 -297500 291540 -297490
rect 291220 -297700 291240 -297500
rect 291420 -297700 291540 -297500
rect 291220 -297710 291540 -297700
rect 291510 -297800 291540 -297710
rect 293140 -297800 293170 -297400
rect 294510 -297490 294540 -297400
rect 294220 -297500 294540 -297490
rect 294220 -297700 294240 -297500
rect 294420 -297700 294540 -297500
rect 294220 -297710 294540 -297700
rect 294510 -297800 294540 -297710
rect 296140 -297800 296170 -297400
rect 297510 -297490 297540 -297400
rect 297220 -297500 297540 -297490
rect 297220 -297700 297240 -297500
rect 297420 -297700 297540 -297500
rect 297220 -297710 297540 -297700
rect 297510 -297800 297540 -297710
rect 299140 -297800 299170 -297400
<< polycont >>
rect 240 -297700 420 -297500
rect 3240 -297700 3420 -297500
rect 6240 -297700 6420 -297500
rect 9240 -297700 9420 -297500
rect 12240 -297700 12420 -297500
rect 15240 -297700 15420 -297500
rect 18240 -297700 18420 -297500
rect 21240 -297700 21420 -297500
rect 24240 -297700 24420 -297500
rect 27240 -297700 27420 -297500
rect 30240 -297700 30420 -297500
rect 33240 -297700 33420 -297500
rect 36240 -297700 36420 -297500
rect 39240 -297700 39420 -297500
rect 42240 -297700 42420 -297500
rect 45240 -297700 45420 -297500
rect 48240 -297700 48420 -297500
rect 51240 -297700 51420 -297500
rect 54240 -297700 54420 -297500
rect 57240 -297700 57420 -297500
rect 60240 -297700 60420 -297500
rect 63240 -297700 63420 -297500
rect 66240 -297700 66420 -297500
rect 69240 -297700 69420 -297500
rect 72240 -297700 72420 -297500
rect 75240 -297700 75420 -297500
rect 78240 -297700 78420 -297500
rect 81240 -297700 81420 -297500
rect 84240 -297700 84420 -297500
rect 87240 -297700 87420 -297500
rect 90240 -297700 90420 -297500
rect 93240 -297700 93420 -297500
rect 96240 -297700 96420 -297500
rect 99240 -297700 99420 -297500
rect 102240 -297700 102420 -297500
rect 105240 -297700 105420 -297500
rect 108240 -297700 108420 -297500
rect 111240 -297700 111420 -297500
rect 114240 -297700 114420 -297500
rect 117240 -297700 117420 -297500
rect 120240 -297700 120420 -297500
rect 123240 -297700 123420 -297500
rect 126240 -297700 126420 -297500
rect 129240 -297700 129420 -297500
rect 132240 -297700 132420 -297500
rect 135240 -297700 135420 -297500
rect 138240 -297700 138420 -297500
rect 141240 -297700 141420 -297500
rect 144240 -297700 144420 -297500
rect 147240 -297700 147420 -297500
rect 150240 -297700 150420 -297500
rect 153240 -297700 153420 -297500
rect 156240 -297700 156420 -297500
rect 159240 -297700 159420 -297500
rect 162240 -297700 162420 -297500
rect 165240 -297700 165420 -297500
rect 168240 -297700 168420 -297500
rect 171240 -297700 171420 -297500
rect 174240 -297700 174420 -297500
rect 177240 -297700 177420 -297500
rect 180240 -297700 180420 -297500
rect 183240 -297700 183420 -297500
rect 186240 -297700 186420 -297500
rect 189240 -297700 189420 -297500
rect 192240 -297700 192420 -297500
rect 195240 -297700 195420 -297500
rect 198240 -297700 198420 -297500
rect 201240 -297700 201420 -297500
rect 204240 -297700 204420 -297500
rect 207240 -297700 207420 -297500
rect 210240 -297700 210420 -297500
rect 213240 -297700 213420 -297500
rect 216240 -297700 216420 -297500
rect 219240 -297700 219420 -297500
rect 222240 -297700 222420 -297500
rect 225240 -297700 225420 -297500
rect 228240 -297700 228420 -297500
rect 231240 -297700 231420 -297500
rect 234240 -297700 234420 -297500
rect 237240 -297700 237420 -297500
rect 240240 -297700 240420 -297500
rect 243240 -297700 243420 -297500
rect 246240 -297700 246420 -297500
rect 249240 -297700 249420 -297500
rect 252240 -297700 252420 -297500
rect 255240 -297700 255420 -297500
rect 258240 -297700 258420 -297500
rect 261240 -297700 261420 -297500
rect 264240 -297700 264420 -297500
rect 267240 -297700 267420 -297500
rect 270240 -297700 270420 -297500
rect 273240 -297700 273420 -297500
rect 276240 -297700 276420 -297500
rect 279240 -297700 279420 -297500
rect 282240 -297700 282420 -297500
rect 285240 -297700 285420 -297500
rect 288240 -297700 288420 -297500
rect 291240 -297700 291420 -297500
rect 294240 -297700 294420 -297500
rect 297240 -297700 297420 -297500
<< locali >>
rect 540 -297290 560 -297230
rect 2120 -297290 2140 -297230
rect 540 -297320 2140 -297290
rect 540 -297380 560 -297320
rect 2120 -297380 2140 -297320
rect 3540 -297290 3560 -297230
rect 5120 -297290 5140 -297230
rect 3540 -297320 5140 -297290
rect 3540 -297380 3560 -297320
rect 5120 -297380 5140 -297320
rect 6540 -297290 6560 -297230
rect 8120 -297290 8140 -297230
rect 6540 -297320 8140 -297290
rect 6540 -297380 6560 -297320
rect 8120 -297380 8140 -297320
rect 9540 -297290 9560 -297230
rect 11120 -297290 11140 -297230
rect 9540 -297320 11140 -297290
rect 9540 -297380 9560 -297320
rect 11120 -297380 11140 -297320
rect 12540 -297290 12560 -297230
rect 14120 -297290 14140 -297230
rect 12540 -297320 14140 -297290
rect 12540 -297380 12560 -297320
rect 14120 -297380 14140 -297320
rect 15540 -297290 15560 -297230
rect 17120 -297290 17140 -297230
rect 15540 -297320 17140 -297290
rect 15540 -297380 15560 -297320
rect 17120 -297380 17140 -297320
rect 18540 -297290 18560 -297230
rect 20120 -297290 20140 -297230
rect 18540 -297320 20140 -297290
rect 18540 -297380 18560 -297320
rect 20120 -297380 20140 -297320
rect 21540 -297290 21560 -297230
rect 23120 -297290 23140 -297230
rect 21540 -297320 23140 -297290
rect 21540 -297380 21560 -297320
rect 23120 -297380 23140 -297320
rect 24540 -297290 24560 -297230
rect 26120 -297290 26140 -297230
rect 24540 -297320 26140 -297290
rect 24540 -297380 24560 -297320
rect 26120 -297380 26140 -297320
rect 27540 -297290 27560 -297230
rect 29120 -297290 29140 -297230
rect 27540 -297320 29140 -297290
rect 27540 -297380 27560 -297320
rect 29120 -297380 29140 -297320
rect 30540 -297290 30560 -297230
rect 32120 -297290 32140 -297230
rect 30540 -297320 32140 -297290
rect 30540 -297380 30560 -297320
rect 32120 -297380 32140 -297320
rect 33540 -297290 33560 -297230
rect 35120 -297290 35140 -297230
rect 33540 -297320 35140 -297290
rect 33540 -297380 33560 -297320
rect 35120 -297380 35140 -297320
rect 36540 -297290 36560 -297230
rect 38120 -297290 38140 -297230
rect 36540 -297320 38140 -297290
rect 36540 -297380 36560 -297320
rect 38120 -297380 38140 -297320
rect 39540 -297290 39560 -297230
rect 41120 -297290 41140 -297230
rect 39540 -297320 41140 -297290
rect 39540 -297380 39560 -297320
rect 41120 -297380 41140 -297320
rect 42540 -297290 42560 -297230
rect 44120 -297290 44140 -297230
rect 42540 -297320 44140 -297290
rect 42540 -297380 42560 -297320
rect 44120 -297380 44140 -297320
rect 45540 -297290 45560 -297230
rect 47120 -297290 47140 -297230
rect 45540 -297320 47140 -297290
rect 45540 -297380 45560 -297320
rect 47120 -297380 47140 -297320
rect 48540 -297290 48560 -297230
rect 50120 -297290 50140 -297230
rect 48540 -297320 50140 -297290
rect 48540 -297380 48560 -297320
rect 50120 -297380 50140 -297320
rect 51540 -297290 51560 -297230
rect 53120 -297290 53140 -297230
rect 51540 -297320 53140 -297290
rect 51540 -297380 51560 -297320
rect 53120 -297380 53140 -297320
rect 54540 -297290 54560 -297230
rect 56120 -297290 56140 -297230
rect 54540 -297320 56140 -297290
rect 54540 -297380 54560 -297320
rect 56120 -297380 56140 -297320
rect 57540 -297290 57560 -297230
rect 59120 -297290 59140 -297230
rect 57540 -297320 59140 -297290
rect 57540 -297380 57560 -297320
rect 59120 -297380 59140 -297320
rect 60540 -297290 60560 -297230
rect 62120 -297290 62140 -297230
rect 60540 -297320 62140 -297290
rect 60540 -297380 60560 -297320
rect 62120 -297380 62140 -297320
rect 63540 -297290 63560 -297230
rect 65120 -297290 65140 -297230
rect 63540 -297320 65140 -297290
rect 63540 -297380 63560 -297320
rect 65120 -297380 65140 -297320
rect 66540 -297290 66560 -297230
rect 68120 -297290 68140 -297230
rect 66540 -297320 68140 -297290
rect 66540 -297380 66560 -297320
rect 68120 -297380 68140 -297320
rect 69540 -297290 69560 -297230
rect 71120 -297290 71140 -297230
rect 69540 -297320 71140 -297290
rect 69540 -297380 69560 -297320
rect 71120 -297380 71140 -297320
rect 72540 -297290 72560 -297230
rect 74120 -297290 74140 -297230
rect 72540 -297320 74140 -297290
rect 72540 -297380 72560 -297320
rect 74120 -297380 74140 -297320
rect 75540 -297290 75560 -297230
rect 77120 -297290 77140 -297230
rect 75540 -297320 77140 -297290
rect 75540 -297380 75560 -297320
rect 77120 -297380 77140 -297320
rect 78540 -297290 78560 -297230
rect 80120 -297290 80140 -297230
rect 78540 -297320 80140 -297290
rect 78540 -297380 78560 -297320
rect 80120 -297380 80140 -297320
rect 81540 -297290 81560 -297230
rect 83120 -297290 83140 -297230
rect 81540 -297320 83140 -297290
rect 81540 -297380 81560 -297320
rect 83120 -297380 83140 -297320
rect 84540 -297290 84560 -297230
rect 86120 -297290 86140 -297230
rect 84540 -297320 86140 -297290
rect 84540 -297380 84560 -297320
rect 86120 -297380 86140 -297320
rect 87540 -297290 87560 -297230
rect 89120 -297290 89140 -297230
rect 87540 -297320 89140 -297290
rect 87540 -297380 87560 -297320
rect 89120 -297380 89140 -297320
rect 90540 -297290 90560 -297230
rect 92120 -297290 92140 -297230
rect 90540 -297320 92140 -297290
rect 90540 -297380 90560 -297320
rect 92120 -297380 92140 -297320
rect 93540 -297290 93560 -297230
rect 95120 -297290 95140 -297230
rect 93540 -297320 95140 -297290
rect 93540 -297380 93560 -297320
rect 95120 -297380 95140 -297320
rect 96540 -297290 96560 -297230
rect 98120 -297290 98140 -297230
rect 96540 -297320 98140 -297290
rect 96540 -297380 96560 -297320
rect 98120 -297380 98140 -297320
rect 99540 -297290 99560 -297230
rect 101120 -297290 101140 -297230
rect 99540 -297320 101140 -297290
rect 99540 -297380 99560 -297320
rect 101120 -297380 101140 -297320
rect 102540 -297290 102560 -297230
rect 104120 -297290 104140 -297230
rect 102540 -297320 104140 -297290
rect 102540 -297380 102560 -297320
rect 104120 -297380 104140 -297320
rect 105540 -297290 105560 -297230
rect 107120 -297290 107140 -297230
rect 105540 -297320 107140 -297290
rect 105540 -297380 105560 -297320
rect 107120 -297380 107140 -297320
rect 108540 -297290 108560 -297230
rect 110120 -297290 110140 -297230
rect 108540 -297320 110140 -297290
rect 108540 -297380 108560 -297320
rect 110120 -297380 110140 -297320
rect 111540 -297290 111560 -297230
rect 113120 -297290 113140 -297230
rect 111540 -297320 113140 -297290
rect 111540 -297380 111560 -297320
rect 113120 -297380 113140 -297320
rect 114540 -297290 114560 -297230
rect 116120 -297290 116140 -297230
rect 114540 -297320 116140 -297290
rect 114540 -297380 114560 -297320
rect 116120 -297380 116140 -297320
rect 117540 -297290 117560 -297230
rect 119120 -297290 119140 -297230
rect 117540 -297320 119140 -297290
rect 117540 -297380 117560 -297320
rect 119120 -297380 119140 -297320
rect 120540 -297290 120560 -297230
rect 122120 -297290 122140 -297230
rect 120540 -297320 122140 -297290
rect 120540 -297380 120560 -297320
rect 122120 -297380 122140 -297320
rect 123540 -297290 123560 -297230
rect 125120 -297290 125140 -297230
rect 123540 -297320 125140 -297290
rect 123540 -297380 123560 -297320
rect 125120 -297380 125140 -297320
rect 126540 -297290 126560 -297230
rect 128120 -297290 128140 -297230
rect 126540 -297320 128140 -297290
rect 126540 -297380 126560 -297320
rect 128120 -297380 128140 -297320
rect 129540 -297290 129560 -297230
rect 131120 -297290 131140 -297230
rect 129540 -297320 131140 -297290
rect 129540 -297380 129560 -297320
rect 131120 -297380 131140 -297320
rect 132540 -297290 132560 -297230
rect 134120 -297290 134140 -297230
rect 132540 -297320 134140 -297290
rect 132540 -297380 132560 -297320
rect 134120 -297380 134140 -297320
rect 135540 -297290 135560 -297230
rect 137120 -297290 137140 -297230
rect 135540 -297320 137140 -297290
rect 135540 -297380 135560 -297320
rect 137120 -297380 137140 -297320
rect 138540 -297290 138560 -297230
rect 140120 -297290 140140 -297230
rect 138540 -297320 140140 -297290
rect 138540 -297380 138560 -297320
rect 140120 -297380 140140 -297320
rect 141540 -297290 141560 -297230
rect 143120 -297290 143140 -297230
rect 141540 -297320 143140 -297290
rect 141540 -297380 141560 -297320
rect 143120 -297380 143140 -297320
rect 144540 -297290 144560 -297230
rect 146120 -297290 146140 -297230
rect 144540 -297320 146140 -297290
rect 144540 -297380 144560 -297320
rect 146120 -297380 146140 -297320
rect 147540 -297290 147560 -297230
rect 149120 -297290 149140 -297230
rect 147540 -297320 149140 -297290
rect 147540 -297380 147560 -297320
rect 149120 -297380 149140 -297320
rect 150540 -297290 150560 -297230
rect 152120 -297290 152140 -297230
rect 150540 -297320 152140 -297290
rect 150540 -297380 150560 -297320
rect 152120 -297380 152140 -297320
rect 153540 -297290 153560 -297230
rect 155120 -297290 155140 -297230
rect 153540 -297320 155140 -297290
rect 153540 -297380 153560 -297320
rect 155120 -297380 155140 -297320
rect 156540 -297290 156560 -297230
rect 158120 -297290 158140 -297230
rect 156540 -297320 158140 -297290
rect 156540 -297380 156560 -297320
rect 158120 -297380 158140 -297320
rect 159540 -297290 159560 -297230
rect 161120 -297290 161140 -297230
rect 159540 -297320 161140 -297290
rect 159540 -297380 159560 -297320
rect 161120 -297380 161140 -297320
rect 162540 -297290 162560 -297230
rect 164120 -297290 164140 -297230
rect 162540 -297320 164140 -297290
rect 162540 -297380 162560 -297320
rect 164120 -297380 164140 -297320
rect 165540 -297290 165560 -297230
rect 167120 -297290 167140 -297230
rect 165540 -297320 167140 -297290
rect 165540 -297380 165560 -297320
rect 167120 -297380 167140 -297320
rect 168540 -297290 168560 -297230
rect 170120 -297290 170140 -297230
rect 168540 -297320 170140 -297290
rect 168540 -297380 168560 -297320
rect 170120 -297380 170140 -297320
rect 171540 -297290 171560 -297230
rect 173120 -297290 173140 -297230
rect 171540 -297320 173140 -297290
rect 171540 -297380 171560 -297320
rect 173120 -297380 173140 -297320
rect 174540 -297290 174560 -297230
rect 176120 -297290 176140 -297230
rect 174540 -297320 176140 -297290
rect 174540 -297380 174560 -297320
rect 176120 -297380 176140 -297320
rect 177540 -297290 177560 -297230
rect 179120 -297290 179140 -297230
rect 177540 -297320 179140 -297290
rect 177540 -297380 177560 -297320
rect 179120 -297380 179140 -297320
rect 180540 -297290 180560 -297230
rect 182120 -297290 182140 -297230
rect 180540 -297320 182140 -297290
rect 180540 -297380 180560 -297320
rect 182120 -297380 182140 -297320
rect 183540 -297290 183560 -297230
rect 185120 -297290 185140 -297230
rect 183540 -297320 185140 -297290
rect 183540 -297380 183560 -297320
rect 185120 -297380 185140 -297320
rect 186540 -297290 186560 -297230
rect 188120 -297290 188140 -297230
rect 186540 -297320 188140 -297290
rect 186540 -297380 186560 -297320
rect 188120 -297380 188140 -297320
rect 189540 -297290 189560 -297230
rect 191120 -297290 191140 -297230
rect 189540 -297320 191140 -297290
rect 189540 -297380 189560 -297320
rect 191120 -297380 191140 -297320
rect 192540 -297290 192560 -297230
rect 194120 -297290 194140 -297230
rect 192540 -297320 194140 -297290
rect 192540 -297380 192560 -297320
rect 194120 -297380 194140 -297320
rect 195540 -297290 195560 -297230
rect 197120 -297290 197140 -297230
rect 195540 -297320 197140 -297290
rect 195540 -297380 195560 -297320
rect 197120 -297380 197140 -297320
rect 198540 -297290 198560 -297230
rect 200120 -297290 200140 -297230
rect 198540 -297320 200140 -297290
rect 198540 -297380 198560 -297320
rect 200120 -297380 200140 -297320
rect 201540 -297290 201560 -297230
rect 203120 -297290 203140 -297230
rect 201540 -297320 203140 -297290
rect 201540 -297380 201560 -297320
rect 203120 -297380 203140 -297320
rect 204540 -297290 204560 -297230
rect 206120 -297290 206140 -297230
rect 204540 -297320 206140 -297290
rect 204540 -297380 204560 -297320
rect 206120 -297380 206140 -297320
rect 207540 -297290 207560 -297230
rect 209120 -297290 209140 -297230
rect 207540 -297320 209140 -297290
rect 207540 -297380 207560 -297320
rect 209120 -297380 209140 -297320
rect 210540 -297290 210560 -297230
rect 212120 -297290 212140 -297230
rect 210540 -297320 212140 -297290
rect 210540 -297380 210560 -297320
rect 212120 -297380 212140 -297320
rect 213540 -297290 213560 -297230
rect 215120 -297290 215140 -297230
rect 213540 -297320 215140 -297290
rect 213540 -297380 213560 -297320
rect 215120 -297380 215140 -297320
rect 216540 -297290 216560 -297230
rect 218120 -297290 218140 -297230
rect 216540 -297320 218140 -297290
rect 216540 -297380 216560 -297320
rect 218120 -297380 218140 -297320
rect 219540 -297290 219560 -297230
rect 221120 -297290 221140 -297230
rect 219540 -297320 221140 -297290
rect 219540 -297380 219560 -297320
rect 221120 -297380 221140 -297320
rect 222540 -297290 222560 -297230
rect 224120 -297290 224140 -297230
rect 222540 -297320 224140 -297290
rect 222540 -297380 222560 -297320
rect 224120 -297380 224140 -297320
rect 225540 -297290 225560 -297230
rect 227120 -297290 227140 -297230
rect 225540 -297320 227140 -297290
rect 225540 -297380 225560 -297320
rect 227120 -297380 227140 -297320
rect 228540 -297290 228560 -297230
rect 230120 -297290 230140 -297230
rect 228540 -297320 230140 -297290
rect 228540 -297380 228560 -297320
rect 230120 -297380 230140 -297320
rect 231540 -297290 231560 -297230
rect 233120 -297290 233140 -297230
rect 231540 -297320 233140 -297290
rect 231540 -297380 231560 -297320
rect 233120 -297380 233140 -297320
rect 234540 -297290 234560 -297230
rect 236120 -297290 236140 -297230
rect 234540 -297320 236140 -297290
rect 234540 -297380 234560 -297320
rect 236120 -297380 236140 -297320
rect 237540 -297290 237560 -297230
rect 239120 -297290 239140 -297230
rect 237540 -297320 239140 -297290
rect 237540 -297380 237560 -297320
rect 239120 -297380 239140 -297320
rect 240540 -297290 240560 -297230
rect 242120 -297290 242140 -297230
rect 240540 -297320 242140 -297290
rect 240540 -297380 240560 -297320
rect 242120 -297380 242140 -297320
rect 243540 -297290 243560 -297230
rect 245120 -297290 245140 -297230
rect 243540 -297320 245140 -297290
rect 243540 -297380 243560 -297320
rect 245120 -297380 245140 -297320
rect 246540 -297290 246560 -297230
rect 248120 -297290 248140 -297230
rect 246540 -297320 248140 -297290
rect 246540 -297380 246560 -297320
rect 248120 -297380 248140 -297320
rect 249540 -297290 249560 -297230
rect 251120 -297290 251140 -297230
rect 249540 -297320 251140 -297290
rect 249540 -297380 249560 -297320
rect 251120 -297380 251140 -297320
rect 252540 -297290 252560 -297230
rect 254120 -297290 254140 -297230
rect 252540 -297320 254140 -297290
rect 252540 -297380 252560 -297320
rect 254120 -297380 254140 -297320
rect 255540 -297290 255560 -297230
rect 257120 -297290 257140 -297230
rect 255540 -297320 257140 -297290
rect 255540 -297380 255560 -297320
rect 257120 -297380 257140 -297320
rect 258540 -297290 258560 -297230
rect 260120 -297290 260140 -297230
rect 258540 -297320 260140 -297290
rect 258540 -297380 258560 -297320
rect 260120 -297380 260140 -297320
rect 261540 -297290 261560 -297230
rect 263120 -297290 263140 -297230
rect 261540 -297320 263140 -297290
rect 261540 -297380 261560 -297320
rect 263120 -297380 263140 -297320
rect 264540 -297290 264560 -297230
rect 266120 -297290 266140 -297230
rect 264540 -297320 266140 -297290
rect 264540 -297380 264560 -297320
rect 266120 -297380 266140 -297320
rect 267540 -297290 267560 -297230
rect 269120 -297290 269140 -297230
rect 267540 -297320 269140 -297290
rect 267540 -297380 267560 -297320
rect 269120 -297380 269140 -297320
rect 270540 -297290 270560 -297230
rect 272120 -297290 272140 -297230
rect 270540 -297320 272140 -297290
rect 270540 -297380 270560 -297320
rect 272120 -297380 272140 -297320
rect 273540 -297290 273560 -297230
rect 275120 -297290 275140 -297230
rect 273540 -297320 275140 -297290
rect 273540 -297380 273560 -297320
rect 275120 -297380 275140 -297320
rect 276540 -297290 276560 -297230
rect 278120 -297290 278140 -297230
rect 276540 -297320 278140 -297290
rect 276540 -297380 276560 -297320
rect 278120 -297380 278140 -297320
rect 279540 -297290 279560 -297230
rect 281120 -297290 281140 -297230
rect 279540 -297320 281140 -297290
rect 279540 -297380 279560 -297320
rect 281120 -297380 281140 -297320
rect 282540 -297290 282560 -297230
rect 284120 -297290 284140 -297230
rect 282540 -297320 284140 -297290
rect 282540 -297380 282560 -297320
rect 284120 -297380 284140 -297320
rect 285540 -297290 285560 -297230
rect 287120 -297290 287140 -297230
rect 285540 -297320 287140 -297290
rect 285540 -297380 285560 -297320
rect 287120 -297380 287140 -297320
rect 288540 -297290 288560 -297230
rect 290120 -297290 290140 -297230
rect 288540 -297320 290140 -297290
rect 288540 -297380 288560 -297320
rect 290120 -297380 290140 -297320
rect 291540 -297290 291560 -297230
rect 293120 -297290 293140 -297230
rect 291540 -297320 293140 -297290
rect 291540 -297380 291560 -297320
rect 293120 -297380 293140 -297320
rect 294540 -297290 294560 -297230
rect 296120 -297290 296140 -297230
rect 294540 -297320 296140 -297290
rect 294540 -297380 294560 -297320
rect 296120 -297380 296140 -297320
rect 297540 -297290 297560 -297230
rect 299120 -297290 299140 -297230
rect 297540 -297320 299140 -297290
rect 297540 -297380 297560 -297320
rect 299120 -297380 299140 -297320
rect 220 -297500 440 -297490
rect 220 -297700 240 -297500
rect 420 -297700 440 -297500
rect 220 -297710 440 -297700
rect 3220 -297500 3440 -297490
rect 3220 -297700 3240 -297500
rect 3420 -297700 3440 -297500
rect 3220 -297710 3440 -297700
rect 6220 -297500 6440 -297490
rect 6220 -297700 6240 -297500
rect 6420 -297700 6440 -297500
rect 6220 -297710 6440 -297700
rect 9220 -297500 9440 -297490
rect 9220 -297700 9240 -297500
rect 9420 -297700 9440 -297500
rect 9220 -297710 9440 -297700
rect 12220 -297500 12440 -297490
rect 12220 -297700 12240 -297500
rect 12420 -297700 12440 -297500
rect 12220 -297710 12440 -297700
rect 15220 -297500 15440 -297490
rect 15220 -297700 15240 -297500
rect 15420 -297700 15440 -297500
rect 15220 -297710 15440 -297700
rect 18220 -297500 18440 -297490
rect 18220 -297700 18240 -297500
rect 18420 -297700 18440 -297500
rect 18220 -297710 18440 -297700
rect 21220 -297500 21440 -297490
rect 21220 -297700 21240 -297500
rect 21420 -297700 21440 -297500
rect 21220 -297710 21440 -297700
rect 24220 -297500 24440 -297490
rect 24220 -297700 24240 -297500
rect 24420 -297700 24440 -297500
rect 24220 -297710 24440 -297700
rect 27220 -297500 27440 -297490
rect 27220 -297700 27240 -297500
rect 27420 -297700 27440 -297500
rect 27220 -297710 27440 -297700
rect 30220 -297500 30440 -297490
rect 30220 -297700 30240 -297500
rect 30420 -297700 30440 -297500
rect 30220 -297710 30440 -297700
rect 33220 -297500 33440 -297490
rect 33220 -297700 33240 -297500
rect 33420 -297700 33440 -297500
rect 33220 -297710 33440 -297700
rect 36220 -297500 36440 -297490
rect 36220 -297700 36240 -297500
rect 36420 -297700 36440 -297500
rect 36220 -297710 36440 -297700
rect 39220 -297500 39440 -297490
rect 39220 -297700 39240 -297500
rect 39420 -297700 39440 -297500
rect 39220 -297710 39440 -297700
rect 42220 -297500 42440 -297490
rect 42220 -297700 42240 -297500
rect 42420 -297700 42440 -297500
rect 42220 -297710 42440 -297700
rect 45220 -297500 45440 -297490
rect 45220 -297700 45240 -297500
rect 45420 -297700 45440 -297500
rect 45220 -297710 45440 -297700
rect 48220 -297500 48440 -297490
rect 48220 -297700 48240 -297500
rect 48420 -297700 48440 -297500
rect 48220 -297710 48440 -297700
rect 51220 -297500 51440 -297490
rect 51220 -297700 51240 -297500
rect 51420 -297700 51440 -297500
rect 51220 -297710 51440 -297700
rect 54220 -297500 54440 -297490
rect 54220 -297700 54240 -297500
rect 54420 -297700 54440 -297500
rect 54220 -297710 54440 -297700
rect 57220 -297500 57440 -297490
rect 57220 -297700 57240 -297500
rect 57420 -297700 57440 -297500
rect 57220 -297710 57440 -297700
rect 60220 -297500 60440 -297490
rect 60220 -297700 60240 -297500
rect 60420 -297700 60440 -297500
rect 60220 -297710 60440 -297700
rect 63220 -297500 63440 -297490
rect 63220 -297700 63240 -297500
rect 63420 -297700 63440 -297500
rect 63220 -297710 63440 -297700
rect 66220 -297500 66440 -297490
rect 66220 -297700 66240 -297500
rect 66420 -297700 66440 -297500
rect 66220 -297710 66440 -297700
rect 69220 -297500 69440 -297490
rect 69220 -297700 69240 -297500
rect 69420 -297700 69440 -297500
rect 69220 -297710 69440 -297700
rect 72220 -297500 72440 -297490
rect 72220 -297700 72240 -297500
rect 72420 -297700 72440 -297500
rect 72220 -297710 72440 -297700
rect 75220 -297500 75440 -297490
rect 75220 -297700 75240 -297500
rect 75420 -297700 75440 -297500
rect 75220 -297710 75440 -297700
rect 78220 -297500 78440 -297490
rect 78220 -297700 78240 -297500
rect 78420 -297700 78440 -297500
rect 78220 -297710 78440 -297700
rect 81220 -297500 81440 -297490
rect 81220 -297700 81240 -297500
rect 81420 -297700 81440 -297500
rect 81220 -297710 81440 -297700
rect 84220 -297500 84440 -297490
rect 84220 -297700 84240 -297500
rect 84420 -297700 84440 -297500
rect 84220 -297710 84440 -297700
rect 87220 -297500 87440 -297490
rect 87220 -297700 87240 -297500
rect 87420 -297700 87440 -297500
rect 87220 -297710 87440 -297700
rect 90220 -297500 90440 -297490
rect 90220 -297700 90240 -297500
rect 90420 -297700 90440 -297500
rect 90220 -297710 90440 -297700
rect 93220 -297500 93440 -297490
rect 93220 -297700 93240 -297500
rect 93420 -297700 93440 -297500
rect 93220 -297710 93440 -297700
rect 96220 -297500 96440 -297490
rect 96220 -297700 96240 -297500
rect 96420 -297700 96440 -297500
rect 96220 -297710 96440 -297700
rect 99220 -297500 99440 -297490
rect 99220 -297700 99240 -297500
rect 99420 -297700 99440 -297500
rect 99220 -297710 99440 -297700
rect 102220 -297500 102440 -297490
rect 102220 -297700 102240 -297500
rect 102420 -297700 102440 -297500
rect 102220 -297710 102440 -297700
rect 105220 -297500 105440 -297490
rect 105220 -297700 105240 -297500
rect 105420 -297700 105440 -297500
rect 105220 -297710 105440 -297700
rect 108220 -297500 108440 -297490
rect 108220 -297700 108240 -297500
rect 108420 -297700 108440 -297500
rect 108220 -297710 108440 -297700
rect 111220 -297500 111440 -297490
rect 111220 -297700 111240 -297500
rect 111420 -297700 111440 -297500
rect 111220 -297710 111440 -297700
rect 114220 -297500 114440 -297490
rect 114220 -297700 114240 -297500
rect 114420 -297700 114440 -297500
rect 114220 -297710 114440 -297700
rect 117220 -297500 117440 -297490
rect 117220 -297700 117240 -297500
rect 117420 -297700 117440 -297500
rect 117220 -297710 117440 -297700
rect 120220 -297500 120440 -297490
rect 120220 -297700 120240 -297500
rect 120420 -297700 120440 -297500
rect 120220 -297710 120440 -297700
rect 123220 -297500 123440 -297490
rect 123220 -297700 123240 -297500
rect 123420 -297700 123440 -297500
rect 123220 -297710 123440 -297700
rect 126220 -297500 126440 -297490
rect 126220 -297700 126240 -297500
rect 126420 -297700 126440 -297500
rect 126220 -297710 126440 -297700
rect 129220 -297500 129440 -297490
rect 129220 -297700 129240 -297500
rect 129420 -297700 129440 -297500
rect 129220 -297710 129440 -297700
rect 132220 -297500 132440 -297490
rect 132220 -297700 132240 -297500
rect 132420 -297700 132440 -297500
rect 132220 -297710 132440 -297700
rect 135220 -297500 135440 -297490
rect 135220 -297700 135240 -297500
rect 135420 -297700 135440 -297500
rect 135220 -297710 135440 -297700
rect 138220 -297500 138440 -297490
rect 138220 -297700 138240 -297500
rect 138420 -297700 138440 -297500
rect 138220 -297710 138440 -297700
rect 141220 -297500 141440 -297490
rect 141220 -297700 141240 -297500
rect 141420 -297700 141440 -297500
rect 141220 -297710 141440 -297700
rect 144220 -297500 144440 -297490
rect 144220 -297700 144240 -297500
rect 144420 -297700 144440 -297500
rect 144220 -297710 144440 -297700
rect 147220 -297500 147440 -297490
rect 147220 -297700 147240 -297500
rect 147420 -297700 147440 -297500
rect 147220 -297710 147440 -297700
rect 150220 -297500 150440 -297490
rect 150220 -297700 150240 -297500
rect 150420 -297700 150440 -297500
rect 150220 -297710 150440 -297700
rect 153220 -297500 153440 -297490
rect 153220 -297700 153240 -297500
rect 153420 -297700 153440 -297500
rect 153220 -297710 153440 -297700
rect 156220 -297500 156440 -297490
rect 156220 -297700 156240 -297500
rect 156420 -297700 156440 -297500
rect 156220 -297710 156440 -297700
rect 159220 -297500 159440 -297490
rect 159220 -297700 159240 -297500
rect 159420 -297700 159440 -297500
rect 159220 -297710 159440 -297700
rect 162220 -297500 162440 -297490
rect 162220 -297700 162240 -297500
rect 162420 -297700 162440 -297500
rect 162220 -297710 162440 -297700
rect 165220 -297500 165440 -297490
rect 165220 -297700 165240 -297500
rect 165420 -297700 165440 -297500
rect 165220 -297710 165440 -297700
rect 168220 -297500 168440 -297490
rect 168220 -297700 168240 -297500
rect 168420 -297700 168440 -297500
rect 168220 -297710 168440 -297700
rect 171220 -297500 171440 -297490
rect 171220 -297700 171240 -297500
rect 171420 -297700 171440 -297500
rect 171220 -297710 171440 -297700
rect 174220 -297500 174440 -297490
rect 174220 -297700 174240 -297500
rect 174420 -297700 174440 -297500
rect 174220 -297710 174440 -297700
rect 177220 -297500 177440 -297490
rect 177220 -297700 177240 -297500
rect 177420 -297700 177440 -297500
rect 177220 -297710 177440 -297700
rect 180220 -297500 180440 -297490
rect 180220 -297700 180240 -297500
rect 180420 -297700 180440 -297500
rect 180220 -297710 180440 -297700
rect 183220 -297500 183440 -297490
rect 183220 -297700 183240 -297500
rect 183420 -297700 183440 -297500
rect 183220 -297710 183440 -297700
rect 186220 -297500 186440 -297490
rect 186220 -297700 186240 -297500
rect 186420 -297700 186440 -297500
rect 186220 -297710 186440 -297700
rect 189220 -297500 189440 -297490
rect 189220 -297700 189240 -297500
rect 189420 -297700 189440 -297500
rect 189220 -297710 189440 -297700
rect 192220 -297500 192440 -297490
rect 192220 -297700 192240 -297500
rect 192420 -297700 192440 -297500
rect 192220 -297710 192440 -297700
rect 195220 -297500 195440 -297490
rect 195220 -297700 195240 -297500
rect 195420 -297700 195440 -297500
rect 195220 -297710 195440 -297700
rect 198220 -297500 198440 -297490
rect 198220 -297700 198240 -297500
rect 198420 -297700 198440 -297500
rect 198220 -297710 198440 -297700
rect 201220 -297500 201440 -297490
rect 201220 -297700 201240 -297500
rect 201420 -297700 201440 -297500
rect 201220 -297710 201440 -297700
rect 204220 -297500 204440 -297490
rect 204220 -297700 204240 -297500
rect 204420 -297700 204440 -297500
rect 204220 -297710 204440 -297700
rect 207220 -297500 207440 -297490
rect 207220 -297700 207240 -297500
rect 207420 -297700 207440 -297500
rect 207220 -297710 207440 -297700
rect 210220 -297500 210440 -297490
rect 210220 -297700 210240 -297500
rect 210420 -297700 210440 -297500
rect 210220 -297710 210440 -297700
rect 213220 -297500 213440 -297490
rect 213220 -297700 213240 -297500
rect 213420 -297700 213440 -297500
rect 213220 -297710 213440 -297700
rect 216220 -297500 216440 -297490
rect 216220 -297700 216240 -297500
rect 216420 -297700 216440 -297500
rect 216220 -297710 216440 -297700
rect 219220 -297500 219440 -297490
rect 219220 -297700 219240 -297500
rect 219420 -297700 219440 -297500
rect 219220 -297710 219440 -297700
rect 222220 -297500 222440 -297490
rect 222220 -297700 222240 -297500
rect 222420 -297700 222440 -297500
rect 222220 -297710 222440 -297700
rect 225220 -297500 225440 -297490
rect 225220 -297700 225240 -297500
rect 225420 -297700 225440 -297500
rect 225220 -297710 225440 -297700
rect 228220 -297500 228440 -297490
rect 228220 -297700 228240 -297500
rect 228420 -297700 228440 -297500
rect 228220 -297710 228440 -297700
rect 231220 -297500 231440 -297490
rect 231220 -297700 231240 -297500
rect 231420 -297700 231440 -297500
rect 231220 -297710 231440 -297700
rect 234220 -297500 234440 -297490
rect 234220 -297700 234240 -297500
rect 234420 -297700 234440 -297500
rect 234220 -297710 234440 -297700
rect 237220 -297500 237440 -297490
rect 237220 -297700 237240 -297500
rect 237420 -297700 237440 -297500
rect 237220 -297710 237440 -297700
rect 240220 -297500 240440 -297490
rect 240220 -297700 240240 -297500
rect 240420 -297700 240440 -297500
rect 240220 -297710 240440 -297700
rect 243220 -297500 243440 -297490
rect 243220 -297700 243240 -297500
rect 243420 -297700 243440 -297500
rect 243220 -297710 243440 -297700
rect 246220 -297500 246440 -297490
rect 246220 -297700 246240 -297500
rect 246420 -297700 246440 -297500
rect 246220 -297710 246440 -297700
rect 249220 -297500 249440 -297490
rect 249220 -297700 249240 -297500
rect 249420 -297700 249440 -297500
rect 249220 -297710 249440 -297700
rect 252220 -297500 252440 -297490
rect 252220 -297700 252240 -297500
rect 252420 -297700 252440 -297500
rect 252220 -297710 252440 -297700
rect 255220 -297500 255440 -297490
rect 255220 -297700 255240 -297500
rect 255420 -297700 255440 -297500
rect 255220 -297710 255440 -297700
rect 258220 -297500 258440 -297490
rect 258220 -297700 258240 -297500
rect 258420 -297700 258440 -297500
rect 258220 -297710 258440 -297700
rect 261220 -297500 261440 -297490
rect 261220 -297700 261240 -297500
rect 261420 -297700 261440 -297500
rect 261220 -297710 261440 -297700
rect 264220 -297500 264440 -297490
rect 264220 -297700 264240 -297500
rect 264420 -297700 264440 -297500
rect 264220 -297710 264440 -297700
rect 267220 -297500 267440 -297490
rect 267220 -297700 267240 -297500
rect 267420 -297700 267440 -297500
rect 267220 -297710 267440 -297700
rect 270220 -297500 270440 -297490
rect 270220 -297700 270240 -297500
rect 270420 -297700 270440 -297500
rect 270220 -297710 270440 -297700
rect 273220 -297500 273440 -297490
rect 273220 -297700 273240 -297500
rect 273420 -297700 273440 -297500
rect 273220 -297710 273440 -297700
rect 276220 -297500 276440 -297490
rect 276220 -297700 276240 -297500
rect 276420 -297700 276440 -297500
rect 276220 -297710 276440 -297700
rect 279220 -297500 279440 -297490
rect 279220 -297700 279240 -297500
rect 279420 -297700 279440 -297500
rect 279220 -297710 279440 -297700
rect 282220 -297500 282440 -297490
rect 282220 -297700 282240 -297500
rect 282420 -297700 282440 -297500
rect 282220 -297710 282440 -297700
rect 285220 -297500 285440 -297490
rect 285220 -297700 285240 -297500
rect 285420 -297700 285440 -297500
rect 285220 -297710 285440 -297700
rect 288220 -297500 288440 -297490
rect 288220 -297700 288240 -297500
rect 288420 -297700 288440 -297500
rect 288220 -297710 288440 -297700
rect 291220 -297500 291440 -297490
rect 291220 -297700 291240 -297500
rect 291420 -297700 291440 -297500
rect 291220 -297710 291440 -297700
rect 294220 -297500 294440 -297490
rect 294220 -297700 294240 -297500
rect 294420 -297700 294440 -297500
rect 294220 -297710 294440 -297700
rect 297220 -297500 297440 -297490
rect 297220 -297700 297240 -297500
rect 297420 -297700 297440 -297500
rect 297220 -297710 297440 -297700
rect 540 -297830 2140 -297800
rect 540 -297870 560 -297830
rect 2120 -297870 2140 -297830
rect 540 -297920 2140 -297870
rect 540 -297980 560 -297920
rect 2120 -297980 2140 -297920
rect 540 -298000 2140 -297980
rect 3540 -297830 5140 -297800
rect 3540 -297870 3560 -297830
rect 5120 -297870 5140 -297830
rect 3540 -297920 5140 -297870
rect 3540 -297980 3560 -297920
rect 5120 -297980 5140 -297920
rect 3540 -298000 5140 -297980
rect 6540 -297830 8140 -297800
rect 6540 -297870 6560 -297830
rect 8120 -297870 8140 -297830
rect 6540 -297920 8140 -297870
rect 6540 -297980 6560 -297920
rect 8120 -297980 8140 -297920
rect 6540 -298000 8140 -297980
rect 9540 -297830 11140 -297800
rect 9540 -297870 9560 -297830
rect 11120 -297870 11140 -297830
rect 9540 -297920 11140 -297870
rect 9540 -297980 9560 -297920
rect 11120 -297980 11140 -297920
rect 9540 -298000 11140 -297980
rect 12540 -297830 14140 -297800
rect 12540 -297870 12560 -297830
rect 14120 -297870 14140 -297830
rect 12540 -297920 14140 -297870
rect 12540 -297980 12560 -297920
rect 14120 -297980 14140 -297920
rect 12540 -298000 14140 -297980
rect 15540 -297830 17140 -297800
rect 15540 -297870 15560 -297830
rect 17120 -297870 17140 -297830
rect 15540 -297920 17140 -297870
rect 15540 -297980 15560 -297920
rect 17120 -297980 17140 -297920
rect 15540 -298000 17140 -297980
rect 18540 -297830 20140 -297800
rect 18540 -297870 18560 -297830
rect 20120 -297870 20140 -297830
rect 18540 -297920 20140 -297870
rect 18540 -297980 18560 -297920
rect 20120 -297980 20140 -297920
rect 18540 -298000 20140 -297980
rect 21540 -297830 23140 -297800
rect 21540 -297870 21560 -297830
rect 23120 -297870 23140 -297830
rect 21540 -297920 23140 -297870
rect 21540 -297980 21560 -297920
rect 23120 -297980 23140 -297920
rect 21540 -298000 23140 -297980
rect 24540 -297830 26140 -297800
rect 24540 -297870 24560 -297830
rect 26120 -297870 26140 -297830
rect 24540 -297920 26140 -297870
rect 24540 -297980 24560 -297920
rect 26120 -297980 26140 -297920
rect 24540 -298000 26140 -297980
rect 27540 -297830 29140 -297800
rect 27540 -297870 27560 -297830
rect 29120 -297870 29140 -297830
rect 27540 -297920 29140 -297870
rect 27540 -297980 27560 -297920
rect 29120 -297980 29140 -297920
rect 27540 -298000 29140 -297980
rect 30540 -297830 32140 -297800
rect 30540 -297870 30560 -297830
rect 32120 -297870 32140 -297830
rect 30540 -297920 32140 -297870
rect 30540 -297980 30560 -297920
rect 32120 -297980 32140 -297920
rect 30540 -298000 32140 -297980
rect 33540 -297830 35140 -297800
rect 33540 -297870 33560 -297830
rect 35120 -297870 35140 -297830
rect 33540 -297920 35140 -297870
rect 33540 -297980 33560 -297920
rect 35120 -297980 35140 -297920
rect 33540 -298000 35140 -297980
rect 36540 -297830 38140 -297800
rect 36540 -297870 36560 -297830
rect 38120 -297870 38140 -297830
rect 36540 -297920 38140 -297870
rect 36540 -297980 36560 -297920
rect 38120 -297980 38140 -297920
rect 36540 -298000 38140 -297980
rect 39540 -297830 41140 -297800
rect 39540 -297870 39560 -297830
rect 41120 -297870 41140 -297830
rect 39540 -297920 41140 -297870
rect 39540 -297980 39560 -297920
rect 41120 -297980 41140 -297920
rect 39540 -298000 41140 -297980
rect 42540 -297830 44140 -297800
rect 42540 -297870 42560 -297830
rect 44120 -297870 44140 -297830
rect 42540 -297920 44140 -297870
rect 42540 -297980 42560 -297920
rect 44120 -297980 44140 -297920
rect 42540 -298000 44140 -297980
rect 45540 -297830 47140 -297800
rect 45540 -297870 45560 -297830
rect 47120 -297870 47140 -297830
rect 45540 -297920 47140 -297870
rect 45540 -297980 45560 -297920
rect 47120 -297980 47140 -297920
rect 45540 -298000 47140 -297980
rect 48540 -297830 50140 -297800
rect 48540 -297870 48560 -297830
rect 50120 -297870 50140 -297830
rect 48540 -297920 50140 -297870
rect 48540 -297980 48560 -297920
rect 50120 -297980 50140 -297920
rect 48540 -298000 50140 -297980
rect 51540 -297830 53140 -297800
rect 51540 -297870 51560 -297830
rect 53120 -297870 53140 -297830
rect 51540 -297920 53140 -297870
rect 51540 -297980 51560 -297920
rect 53120 -297980 53140 -297920
rect 51540 -298000 53140 -297980
rect 54540 -297830 56140 -297800
rect 54540 -297870 54560 -297830
rect 56120 -297870 56140 -297830
rect 54540 -297920 56140 -297870
rect 54540 -297980 54560 -297920
rect 56120 -297980 56140 -297920
rect 54540 -298000 56140 -297980
rect 57540 -297830 59140 -297800
rect 57540 -297870 57560 -297830
rect 59120 -297870 59140 -297830
rect 57540 -297920 59140 -297870
rect 57540 -297980 57560 -297920
rect 59120 -297980 59140 -297920
rect 57540 -298000 59140 -297980
rect 60540 -297830 62140 -297800
rect 60540 -297870 60560 -297830
rect 62120 -297870 62140 -297830
rect 60540 -297920 62140 -297870
rect 60540 -297980 60560 -297920
rect 62120 -297980 62140 -297920
rect 60540 -298000 62140 -297980
rect 63540 -297830 65140 -297800
rect 63540 -297870 63560 -297830
rect 65120 -297870 65140 -297830
rect 63540 -297920 65140 -297870
rect 63540 -297980 63560 -297920
rect 65120 -297980 65140 -297920
rect 63540 -298000 65140 -297980
rect 66540 -297830 68140 -297800
rect 66540 -297870 66560 -297830
rect 68120 -297870 68140 -297830
rect 66540 -297920 68140 -297870
rect 66540 -297980 66560 -297920
rect 68120 -297980 68140 -297920
rect 66540 -298000 68140 -297980
rect 69540 -297830 71140 -297800
rect 69540 -297870 69560 -297830
rect 71120 -297870 71140 -297830
rect 69540 -297920 71140 -297870
rect 69540 -297980 69560 -297920
rect 71120 -297980 71140 -297920
rect 69540 -298000 71140 -297980
rect 72540 -297830 74140 -297800
rect 72540 -297870 72560 -297830
rect 74120 -297870 74140 -297830
rect 72540 -297920 74140 -297870
rect 72540 -297980 72560 -297920
rect 74120 -297980 74140 -297920
rect 72540 -298000 74140 -297980
rect 75540 -297830 77140 -297800
rect 75540 -297870 75560 -297830
rect 77120 -297870 77140 -297830
rect 75540 -297920 77140 -297870
rect 75540 -297980 75560 -297920
rect 77120 -297980 77140 -297920
rect 75540 -298000 77140 -297980
rect 78540 -297830 80140 -297800
rect 78540 -297870 78560 -297830
rect 80120 -297870 80140 -297830
rect 78540 -297920 80140 -297870
rect 78540 -297980 78560 -297920
rect 80120 -297980 80140 -297920
rect 78540 -298000 80140 -297980
rect 81540 -297830 83140 -297800
rect 81540 -297870 81560 -297830
rect 83120 -297870 83140 -297830
rect 81540 -297920 83140 -297870
rect 81540 -297980 81560 -297920
rect 83120 -297980 83140 -297920
rect 81540 -298000 83140 -297980
rect 84540 -297830 86140 -297800
rect 84540 -297870 84560 -297830
rect 86120 -297870 86140 -297830
rect 84540 -297920 86140 -297870
rect 84540 -297980 84560 -297920
rect 86120 -297980 86140 -297920
rect 84540 -298000 86140 -297980
rect 87540 -297830 89140 -297800
rect 87540 -297870 87560 -297830
rect 89120 -297870 89140 -297830
rect 87540 -297920 89140 -297870
rect 87540 -297980 87560 -297920
rect 89120 -297980 89140 -297920
rect 87540 -298000 89140 -297980
rect 90540 -297830 92140 -297800
rect 90540 -297870 90560 -297830
rect 92120 -297870 92140 -297830
rect 90540 -297920 92140 -297870
rect 90540 -297980 90560 -297920
rect 92120 -297980 92140 -297920
rect 90540 -298000 92140 -297980
rect 93540 -297830 95140 -297800
rect 93540 -297870 93560 -297830
rect 95120 -297870 95140 -297830
rect 93540 -297920 95140 -297870
rect 93540 -297980 93560 -297920
rect 95120 -297980 95140 -297920
rect 93540 -298000 95140 -297980
rect 96540 -297830 98140 -297800
rect 96540 -297870 96560 -297830
rect 98120 -297870 98140 -297830
rect 96540 -297920 98140 -297870
rect 96540 -297980 96560 -297920
rect 98120 -297980 98140 -297920
rect 96540 -298000 98140 -297980
rect 99540 -297830 101140 -297800
rect 99540 -297870 99560 -297830
rect 101120 -297870 101140 -297830
rect 99540 -297920 101140 -297870
rect 99540 -297980 99560 -297920
rect 101120 -297980 101140 -297920
rect 99540 -298000 101140 -297980
rect 102540 -297830 104140 -297800
rect 102540 -297870 102560 -297830
rect 104120 -297870 104140 -297830
rect 102540 -297920 104140 -297870
rect 102540 -297980 102560 -297920
rect 104120 -297980 104140 -297920
rect 102540 -298000 104140 -297980
rect 105540 -297830 107140 -297800
rect 105540 -297870 105560 -297830
rect 107120 -297870 107140 -297830
rect 105540 -297920 107140 -297870
rect 105540 -297980 105560 -297920
rect 107120 -297980 107140 -297920
rect 105540 -298000 107140 -297980
rect 108540 -297830 110140 -297800
rect 108540 -297870 108560 -297830
rect 110120 -297870 110140 -297830
rect 108540 -297920 110140 -297870
rect 108540 -297980 108560 -297920
rect 110120 -297980 110140 -297920
rect 108540 -298000 110140 -297980
rect 111540 -297830 113140 -297800
rect 111540 -297870 111560 -297830
rect 113120 -297870 113140 -297830
rect 111540 -297920 113140 -297870
rect 111540 -297980 111560 -297920
rect 113120 -297980 113140 -297920
rect 111540 -298000 113140 -297980
rect 114540 -297830 116140 -297800
rect 114540 -297870 114560 -297830
rect 116120 -297870 116140 -297830
rect 114540 -297920 116140 -297870
rect 114540 -297980 114560 -297920
rect 116120 -297980 116140 -297920
rect 114540 -298000 116140 -297980
rect 117540 -297830 119140 -297800
rect 117540 -297870 117560 -297830
rect 119120 -297870 119140 -297830
rect 117540 -297920 119140 -297870
rect 117540 -297980 117560 -297920
rect 119120 -297980 119140 -297920
rect 117540 -298000 119140 -297980
rect 120540 -297830 122140 -297800
rect 120540 -297870 120560 -297830
rect 122120 -297870 122140 -297830
rect 120540 -297920 122140 -297870
rect 120540 -297980 120560 -297920
rect 122120 -297980 122140 -297920
rect 120540 -298000 122140 -297980
rect 123540 -297830 125140 -297800
rect 123540 -297870 123560 -297830
rect 125120 -297870 125140 -297830
rect 123540 -297920 125140 -297870
rect 123540 -297980 123560 -297920
rect 125120 -297980 125140 -297920
rect 123540 -298000 125140 -297980
rect 126540 -297830 128140 -297800
rect 126540 -297870 126560 -297830
rect 128120 -297870 128140 -297830
rect 126540 -297920 128140 -297870
rect 126540 -297980 126560 -297920
rect 128120 -297980 128140 -297920
rect 126540 -298000 128140 -297980
rect 129540 -297830 131140 -297800
rect 129540 -297870 129560 -297830
rect 131120 -297870 131140 -297830
rect 129540 -297920 131140 -297870
rect 129540 -297980 129560 -297920
rect 131120 -297980 131140 -297920
rect 129540 -298000 131140 -297980
rect 132540 -297830 134140 -297800
rect 132540 -297870 132560 -297830
rect 134120 -297870 134140 -297830
rect 132540 -297920 134140 -297870
rect 132540 -297980 132560 -297920
rect 134120 -297980 134140 -297920
rect 132540 -298000 134140 -297980
rect 135540 -297830 137140 -297800
rect 135540 -297870 135560 -297830
rect 137120 -297870 137140 -297830
rect 135540 -297920 137140 -297870
rect 135540 -297980 135560 -297920
rect 137120 -297980 137140 -297920
rect 135540 -298000 137140 -297980
rect 138540 -297830 140140 -297800
rect 138540 -297870 138560 -297830
rect 140120 -297870 140140 -297830
rect 138540 -297920 140140 -297870
rect 138540 -297980 138560 -297920
rect 140120 -297980 140140 -297920
rect 138540 -298000 140140 -297980
rect 141540 -297830 143140 -297800
rect 141540 -297870 141560 -297830
rect 143120 -297870 143140 -297830
rect 141540 -297920 143140 -297870
rect 141540 -297980 141560 -297920
rect 143120 -297980 143140 -297920
rect 141540 -298000 143140 -297980
rect 144540 -297830 146140 -297800
rect 144540 -297870 144560 -297830
rect 146120 -297870 146140 -297830
rect 144540 -297920 146140 -297870
rect 144540 -297980 144560 -297920
rect 146120 -297980 146140 -297920
rect 144540 -298000 146140 -297980
rect 147540 -297830 149140 -297800
rect 147540 -297870 147560 -297830
rect 149120 -297870 149140 -297830
rect 147540 -297920 149140 -297870
rect 147540 -297980 147560 -297920
rect 149120 -297980 149140 -297920
rect 147540 -298000 149140 -297980
rect 150540 -297830 152140 -297800
rect 150540 -297870 150560 -297830
rect 152120 -297870 152140 -297830
rect 150540 -297920 152140 -297870
rect 150540 -297980 150560 -297920
rect 152120 -297980 152140 -297920
rect 150540 -298000 152140 -297980
rect 153540 -297830 155140 -297800
rect 153540 -297870 153560 -297830
rect 155120 -297870 155140 -297830
rect 153540 -297920 155140 -297870
rect 153540 -297980 153560 -297920
rect 155120 -297980 155140 -297920
rect 153540 -298000 155140 -297980
rect 156540 -297830 158140 -297800
rect 156540 -297870 156560 -297830
rect 158120 -297870 158140 -297830
rect 156540 -297920 158140 -297870
rect 156540 -297980 156560 -297920
rect 158120 -297980 158140 -297920
rect 156540 -298000 158140 -297980
rect 159540 -297830 161140 -297800
rect 159540 -297870 159560 -297830
rect 161120 -297870 161140 -297830
rect 159540 -297920 161140 -297870
rect 159540 -297980 159560 -297920
rect 161120 -297980 161140 -297920
rect 159540 -298000 161140 -297980
rect 162540 -297830 164140 -297800
rect 162540 -297870 162560 -297830
rect 164120 -297870 164140 -297830
rect 162540 -297920 164140 -297870
rect 162540 -297980 162560 -297920
rect 164120 -297980 164140 -297920
rect 162540 -298000 164140 -297980
rect 165540 -297830 167140 -297800
rect 165540 -297870 165560 -297830
rect 167120 -297870 167140 -297830
rect 165540 -297920 167140 -297870
rect 165540 -297980 165560 -297920
rect 167120 -297980 167140 -297920
rect 165540 -298000 167140 -297980
rect 168540 -297830 170140 -297800
rect 168540 -297870 168560 -297830
rect 170120 -297870 170140 -297830
rect 168540 -297920 170140 -297870
rect 168540 -297980 168560 -297920
rect 170120 -297980 170140 -297920
rect 168540 -298000 170140 -297980
rect 171540 -297830 173140 -297800
rect 171540 -297870 171560 -297830
rect 173120 -297870 173140 -297830
rect 171540 -297920 173140 -297870
rect 171540 -297980 171560 -297920
rect 173120 -297980 173140 -297920
rect 171540 -298000 173140 -297980
rect 174540 -297830 176140 -297800
rect 174540 -297870 174560 -297830
rect 176120 -297870 176140 -297830
rect 174540 -297920 176140 -297870
rect 174540 -297980 174560 -297920
rect 176120 -297980 176140 -297920
rect 174540 -298000 176140 -297980
rect 177540 -297830 179140 -297800
rect 177540 -297870 177560 -297830
rect 179120 -297870 179140 -297830
rect 177540 -297920 179140 -297870
rect 177540 -297980 177560 -297920
rect 179120 -297980 179140 -297920
rect 177540 -298000 179140 -297980
rect 180540 -297830 182140 -297800
rect 180540 -297870 180560 -297830
rect 182120 -297870 182140 -297830
rect 180540 -297920 182140 -297870
rect 180540 -297980 180560 -297920
rect 182120 -297980 182140 -297920
rect 180540 -298000 182140 -297980
rect 183540 -297830 185140 -297800
rect 183540 -297870 183560 -297830
rect 185120 -297870 185140 -297830
rect 183540 -297920 185140 -297870
rect 183540 -297980 183560 -297920
rect 185120 -297980 185140 -297920
rect 183540 -298000 185140 -297980
rect 186540 -297830 188140 -297800
rect 186540 -297870 186560 -297830
rect 188120 -297870 188140 -297830
rect 186540 -297920 188140 -297870
rect 186540 -297980 186560 -297920
rect 188120 -297980 188140 -297920
rect 186540 -298000 188140 -297980
rect 189540 -297830 191140 -297800
rect 189540 -297870 189560 -297830
rect 191120 -297870 191140 -297830
rect 189540 -297920 191140 -297870
rect 189540 -297980 189560 -297920
rect 191120 -297980 191140 -297920
rect 189540 -298000 191140 -297980
rect 192540 -297830 194140 -297800
rect 192540 -297870 192560 -297830
rect 194120 -297870 194140 -297830
rect 192540 -297920 194140 -297870
rect 192540 -297980 192560 -297920
rect 194120 -297980 194140 -297920
rect 192540 -298000 194140 -297980
rect 195540 -297830 197140 -297800
rect 195540 -297870 195560 -297830
rect 197120 -297870 197140 -297830
rect 195540 -297920 197140 -297870
rect 195540 -297980 195560 -297920
rect 197120 -297980 197140 -297920
rect 195540 -298000 197140 -297980
rect 198540 -297830 200140 -297800
rect 198540 -297870 198560 -297830
rect 200120 -297870 200140 -297830
rect 198540 -297920 200140 -297870
rect 198540 -297980 198560 -297920
rect 200120 -297980 200140 -297920
rect 198540 -298000 200140 -297980
rect 201540 -297830 203140 -297800
rect 201540 -297870 201560 -297830
rect 203120 -297870 203140 -297830
rect 201540 -297920 203140 -297870
rect 201540 -297980 201560 -297920
rect 203120 -297980 203140 -297920
rect 201540 -298000 203140 -297980
rect 204540 -297830 206140 -297800
rect 204540 -297870 204560 -297830
rect 206120 -297870 206140 -297830
rect 204540 -297920 206140 -297870
rect 204540 -297980 204560 -297920
rect 206120 -297980 206140 -297920
rect 204540 -298000 206140 -297980
rect 207540 -297830 209140 -297800
rect 207540 -297870 207560 -297830
rect 209120 -297870 209140 -297830
rect 207540 -297920 209140 -297870
rect 207540 -297980 207560 -297920
rect 209120 -297980 209140 -297920
rect 207540 -298000 209140 -297980
rect 210540 -297830 212140 -297800
rect 210540 -297870 210560 -297830
rect 212120 -297870 212140 -297830
rect 210540 -297920 212140 -297870
rect 210540 -297980 210560 -297920
rect 212120 -297980 212140 -297920
rect 210540 -298000 212140 -297980
rect 213540 -297830 215140 -297800
rect 213540 -297870 213560 -297830
rect 215120 -297870 215140 -297830
rect 213540 -297920 215140 -297870
rect 213540 -297980 213560 -297920
rect 215120 -297980 215140 -297920
rect 213540 -298000 215140 -297980
rect 216540 -297830 218140 -297800
rect 216540 -297870 216560 -297830
rect 218120 -297870 218140 -297830
rect 216540 -297920 218140 -297870
rect 216540 -297980 216560 -297920
rect 218120 -297980 218140 -297920
rect 216540 -298000 218140 -297980
rect 219540 -297830 221140 -297800
rect 219540 -297870 219560 -297830
rect 221120 -297870 221140 -297830
rect 219540 -297920 221140 -297870
rect 219540 -297980 219560 -297920
rect 221120 -297980 221140 -297920
rect 219540 -298000 221140 -297980
rect 222540 -297830 224140 -297800
rect 222540 -297870 222560 -297830
rect 224120 -297870 224140 -297830
rect 222540 -297920 224140 -297870
rect 222540 -297980 222560 -297920
rect 224120 -297980 224140 -297920
rect 222540 -298000 224140 -297980
rect 225540 -297830 227140 -297800
rect 225540 -297870 225560 -297830
rect 227120 -297870 227140 -297830
rect 225540 -297920 227140 -297870
rect 225540 -297980 225560 -297920
rect 227120 -297980 227140 -297920
rect 225540 -298000 227140 -297980
rect 228540 -297830 230140 -297800
rect 228540 -297870 228560 -297830
rect 230120 -297870 230140 -297830
rect 228540 -297920 230140 -297870
rect 228540 -297980 228560 -297920
rect 230120 -297980 230140 -297920
rect 228540 -298000 230140 -297980
rect 231540 -297830 233140 -297800
rect 231540 -297870 231560 -297830
rect 233120 -297870 233140 -297830
rect 231540 -297920 233140 -297870
rect 231540 -297980 231560 -297920
rect 233120 -297980 233140 -297920
rect 231540 -298000 233140 -297980
rect 234540 -297830 236140 -297800
rect 234540 -297870 234560 -297830
rect 236120 -297870 236140 -297830
rect 234540 -297920 236140 -297870
rect 234540 -297980 234560 -297920
rect 236120 -297980 236140 -297920
rect 234540 -298000 236140 -297980
rect 237540 -297830 239140 -297800
rect 237540 -297870 237560 -297830
rect 239120 -297870 239140 -297830
rect 237540 -297920 239140 -297870
rect 237540 -297980 237560 -297920
rect 239120 -297980 239140 -297920
rect 237540 -298000 239140 -297980
rect 240540 -297830 242140 -297800
rect 240540 -297870 240560 -297830
rect 242120 -297870 242140 -297830
rect 240540 -297920 242140 -297870
rect 240540 -297980 240560 -297920
rect 242120 -297980 242140 -297920
rect 240540 -298000 242140 -297980
rect 243540 -297830 245140 -297800
rect 243540 -297870 243560 -297830
rect 245120 -297870 245140 -297830
rect 243540 -297920 245140 -297870
rect 243540 -297980 243560 -297920
rect 245120 -297980 245140 -297920
rect 243540 -298000 245140 -297980
rect 246540 -297830 248140 -297800
rect 246540 -297870 246560 -297830
rect 248120 -297870 248140 -297830
rect 246540 -297920 248140 -297870
rect 246540 -297980 246560 -297920
rect 248120 -297980 248140 -297920
rect 246540 -298000 248140 -297980
rect 249540 -297830 251140 -297800
rect 249540 -297870 249560 -297830
rect 251120 -297870 251140 -297830
rect 249540 -297920 251140 -297870
rect 249540 -297980 249560 -297920
rect 251120 -297980 251140 -297920
rect 249540 -298000 251140 -297980
rect 252540 -297830 254140 -297800
rect 252540 -297870 252560 -297830
rect 254120 -297870 254140 -297830
rect 252540 -297920 254140 -297870
rect 252540 -297980 252560 -297920
rect 254120 -297980 254140 -297920
rect 252540 -298000 254140 -297980
rect 255540 -297830 257140 -297800
rect 255540 -297870 255560 -297830
rect 257120 -297870 257140 -297830
rect 255540 -297920 257140 -297870
rect 255540 -297980 255560 -297920
rect 257120 -297980 257140 -297920
rect 255540 -298000 257140 -297980
rect 258540 -297830 260140 -297800
rect 258540 -297870 258560 -297830
rect 260120 -297870 260140 -297830
rect 258540 -297920 260140 -297870
rect 258540 -297980 258560 -297920
rect 260120 -297980 260140 -297920
rect 258540 -298000 260140 -297980
rect 261540 -297830 263140 -297800
rect 261540 -297870 261560 -297830
rect 263120 -297870 263140 -297830
rect 261540 -297920 263140 -297870
rect 261540 -297980 261560 -297920
rect 263120 -297980 263140 -297920
rect 261540 -298000 263140 -297980
rect 264540 -297830 266140 -297800
rect 264540 -297870 264560 -297830
rect 266120 -297870 266140 -297830
rect 264540 -297920 266140 -297870
rect 264540 -297980 264560 -297920
rect 266120 -297980 266140 -297920
rect 264540 -298000 266140 -297980
rect 267540 -297830 269140 -297800
rect 267540 -297870 267560 -297830
rect 269120 -297870 269140 -297830
rect 267540 -297920 269140 -297870
rect 267540 -297980 267560 -297920
rect 269120 -297980 269140 -297920
rect 267540 -298000 269140 -297980
rect 270540 -297830 272140 -297800
rect 270540 -297870 270560 -297830
rect 272120 -297870 272140 -297830
rect 270540 -297920 272140 -297870
rect 270540 -297980 270560 -297920
rect 272120 -297980 272140 -297920
rect 270540 -298000 272140 -297980
rect 273540 -297830 275140 -297800
rect 273540 -297870 273560 -297830
rect 275120 -297870 275140 -297830
rect 273540 -297920 275140 -297870
rect 273540 -297980 273560 -297920
rect 275120 -297980 275140 -297920
rect 273540 -298000 275140 -297980
rect 276540 -297830 278140 -297800
rect 276540 -297870 276560 -297830
rect 278120 -297870 278140 -297830
rect 276540 -297920 278140 -297870
rect 276540 -297980 276560 -297920
rect 278120 -297980 278140 -297920
rect 276540 -298000 278140 -297980
rect 279540 -297830 281140 -297800
rect 279540 -297870 279560 -297830
rect 281120 -297870 281140 -297830
rect 279540 -297920 281140 -297870
rect 279540 -297980 279560 -297920
rect 281120 -297980 281140 -297920
rect 279540 -298000 281140 -297980
rect 282540 -297830 284140 -297800
rect 282540 -297870 282560 -297830
rect 284120 -297870 284140 -297830
rect 282540 -297920 284140 -297870
rect 282540 -297980 282560 -297920
rect 284120 -297980 284140 -297920
rect 282540 -298000 284140 -297980
rect 285540 -297830 287140 -297800
rect 285540 -297870 285560 -297830
rect 287120 -297870 287140 -297830
rect 285540 -297920 287140 -297870
rect 285540 -297980 285560 -297920
rect 287120 -297980 287140 -297920
rect 285540 -298000 287140 -297980
rect 288540 -297830 290140 -297800
rect 288540 -297870 288560 -297830
rect 290120 -297870 290140 -297830
rect 288540 -297920 290140 -297870
rect 288540 -297980 288560 -297920
rect 290120 -297980 290140 -297920
rect 288540 -298000 290140 -297980
rect 291540 -297830 293140 -297800
rect 291540 -297870 291560 -297830
rect 293120 -297870 293140 -297830
rect 291540 -297920 293140 -297870
rect 291540 -297980 291560 -297920
rect 293120 -297980 293140 -297920
rect 291540 -298000 293140 -297980
rect 294540 -297830 296140 -297800
rect 294540 -297870 294560 -297830
rect 296120 -297870 296140 -297830
rect 294540 -297920 296140 -297870
rect 294540 -297980 294560 -297920
rect 296120 -297980 296140 -297920
rect 294540 -298000 296140 -297980
rect 297540 -297830 299140 -297800
rect 297540 -297870 297560 -297830
rect 299120 -297870 299140 -297830
rect 297540 -297920 299140 -297870
rect 297540 -297980 297560 -297920
rect 299120 -297980 299140 -297920
rect 297540 -298000 299140 -297980
<< viali >>
rect 560 -297290 2120 -297230
rect 3560 -297290 5120 -297230
rect 6560 -297290 8120 -297230
rect 9560 -297290 11120 -297230
rect 12560 -297290 14120 -297230
rect 15560 -297290 17120 -297230
rect 18560 -297290 20120 -297230
rect 21560 -297290 23120 -297230
rect 24560 -297290 26120 -297230
rect 27560 -297290 29120 -297230
rect 30560 -297290 32120 -297230
rect 33560 -297290 35120 -297230
rect 36560 -297290 38120 -297230
rect 39560 -297290 41120 -297230
rect 42560 -297290 44120 -297230
rect 45560 -297290 47120 -297230
rect 48560 -297290 50120 -297230
rect 51560 -297290 53120 -297230
rect 54560 -297290 56120 -297230
rect 57560 -297290 59120 -297230
rect 60560 -297290 62120 -297230
rect 63560 -297290 65120 -297230
rect 66560 -297290 68120 -297230
rect 69560 -297290 71120 -297230
rect 72560 -297290 74120 -297230
rect 75560 -297290 77120 -297230
rect 78560 -297290 80120 -297230
rect 81560 -297290 83120 -297230
rect 84560 -297290 86120 -297230
rect 87560 -297290 89120 -297230
rect 90560 -297290 92120 -297230
rect 93560 -297290 95120 -297230
rect 96560 -297290 98120 -297230
rect 99560 -297290 101120 -297230
rect 102560 -297290 104120 -297230
rect 105560 -297290 107120 -297230
rect 108560 -297290 110120 -297230
rect 111560 -297290 113120 -297230
rect 114560 -297290 116120 -297230
rect 117560 -297290 119120 -297230
rect 120560 -297290 122120 -297230
rect 123560 -297290 125120 -297230
rect 126560 -297290 128120 -297230
rect 129560 -297290 131120 -297230
rect 132560 -297290 134120 -297230
rect 135560 -297290 137120 -297230
rect 138560 -297290 140120 -297230
rect 141560 -297290 143120 -297230
rect 144560 -297290 146120 -297230
rect 147560 -297290 149120 -297230
rect 150560 -297290 152120 -297230
rect 153560 -297290 155120 -297230
rect 156560 -297290 158120 -297230
rect 159560 -297290 161120 -297230
rect 162560 -297290 164120 -297230
rect 165560 -297290 167120 -297230
rect 168560 -297290 170120 -297230
rect 171560 -297290 173120 -297230
rect 174560 -297290 176120 -297230
rect 177560 -297290 179120 -297230
rect 180560 -297290 182120 -297230
rect 183560 -297290 185120 -297230
rect 186560 -297290 188120 -297230
rect 189560 -297290 191120 -297230
rect 192560 -297290 194120 -297230
rect 195560 -297290 197120 -297230
rect 198560 -297290 200120 -297230
rect 201560 -297290 203120 -297230
rect 204560 -297290 206120 -297230
rect 207560 -297290 209120 -297230
rect 210560 -297290 212120 -297230
rect 213560 -297290 215120 -297230
rect 216560 -297290 218120 -297230
rect 219560 -297290 221120 -297230
rect 222560 -297290 224120 -297230
rect 225560 -297290 227120 -297230
rect 228560 -297290 230120 -297230
rect 231560 -297290 233120 -297230
rect 234560 -297290 236120 -297230
rect 237560 -297290 239120 -297230
rect 240560 -297290 242120 -297230
rect 243560 -297290 245120 -297230
rect 246560 -297290 248120 -297230
rect 249560 -297290 251120 -297230
rect 252560 -297290 254120 -297230
rect 255560 -297290 257120 -297230
rect 258560 -297290 260120 -297230
rect 261560 -297290 263120 -297230
rect 264560 -297290 266120 -297230
rect 267560 -297290 269120 -297230
rect 270560 -297290 272120 -297230
rect 273560 -297290 275120 -297230
rect 276560 -297290 278120 -297230
rect 279560 -297290 281120 -297230
rect 282560 -297290 284120 -297230
rect 285560 -297290 287120 -297230
rect 288560 -297290 290120 -297230
rect 291560 -297290 293120 -297230
rect 294560 -297290 296120 -297230
rect 297560 -297290 299120 -297230
rect 240 -297700 420 -297500
rect 3240 -297700 3420 -297500
rect 6240 -297700 6420 -297500
rect 9240 -297700 9420 -297500
rect 12240 -297700 12420 -297500
rect 15240 -297700 15420 -297500
rect 18240 -297700 18420 -297500
rect 21240 -297700 21420 -297500
rect 24240 -297700 24420 -297500
rect 27240 -297700 27420 -297500
rect 30240 -297700 30420 -297500
rect 33240 -297700 33420 -297500
rect 36240 -297700 36420 -297500
rect 39240 -297700 39420 -297500
rect 42240 -297700 42420 -297500
rect 45240 -297700 45420 -297500
rect 48240 -297700 48420 -297500
rect 51240 -297700 51420 -297500
rect 54240 -297700 54420 -297500
rect 57240 -297700 57420 -297500
rect 60240 -297700 60420 -297500
rect 63240 -297700 63420 -297500
rect 66240 -297700 66420 -297500
rect 69240 -297700 69420 -297500
rect 72240 -297700 72420 -297500
rect 75240 -297700 75420 -297500
rect 78240 -297700 78420 -297500
rect 81240 -297700 81420 -297500
rect 84240 -297700 84420 -297500
rect 87240 -297700 87420 -297500
rect 90240 -297700 90420 -297500
rect 93240 -297700 93420 -297500
rect 96240 -297700 96420 -297500
rect 99240 -297700 99420 -297500
rect 102240 -297700 102420 -297500
rect 105240 -297700 105420 -297500
rect 108240 -297700 108420 -297500
rect 111240 -297700 111420 -297500
rect 114240 -297700 114420 -297500
rect 117240 -297700 117420 -297500
rect 120240 -297700 120420 -297500
rect 123240 -297700 123420 -297500
rect 126240 -297700 126420 -297500
rect 129240 -297700 129420 -297500
rect 132240 -297700 132420 -297500
rect 135240 -297700 135420 -297500
rect 138240 -297700 138420 -297500
rect 141240 -297700 141420 -297500
rect 144240 -297700 144420 -297500
rect 147240 -297700 147420 -297500
rect 150240 -297700 150420 -297500
rect 153240 -297700 153420 -297500
rect 156240 -297700 156420 -297500
rect 159240 -297700 159420 -297500
rect 162240 -297700 162420 -297500
rect 165240 -297700 165420 -297500
rect 168240 -297700 168420 -297500
rect 171240 -297700 171420 -297500
rect 174240 -297700 174420 -297500
rect 177240 -297700 177420 -297500
rect 180240 -297700 180420 -297500
rect 183240 -297700 183420 -297500
rect 186240 -297700 186420 -297500
rect 189240 -297700 189420 -297500
rect 192240 -297700 192420 -297500
rect 195240 -297700 195420 -297500
rect 198240 -297700 198420 -297500
rect 201240 -297700 201420 -297500
rect 204240 -297700 204420 -297500
rect 207240 -297700 207420 -297500
rect 210240 -297700 210420 -297500
rect 213240 -297700 213420 -297500
rect 216240 -297700 216420 -297500
rect 219240 -297700 219420 -297500
rect 222240 -297700 222420 -297500
rect 225240 -297700 225420 -297500
rect 228240 -297700 228420 -297500
rect 231240 -297700 231420 -297500
rect 234240 -297700 234420 -297500
rect 237240 -297700 237420 -297500
rect 240240 -297700 240420 -297500
rect 243240 -297700 243420 -297500
rect 246240 -297700 246420 -297500
rect 249240 -297700 249420 -297500
rect 252240 -297700 252420 -297500
rect 255240 -297700 255420 -297500
rect 258240 -297700 258420 -297500
rect 261240 -297700 261420 -297500
rect 264240 -297700 264420 -297500
rect 267240 -297700 267420 -297500
rect 270240 -297700 270420 -297500
rect 273240 -297700 273420 -297500
rect 276240 -297700 276420 -297500
rect 279240 -297700 279420 -297500
rect 282240 -297700 282420 -297500
rect 285240 -297700 285420 -297500
rect 288240 -297700 288420 -297500
rect 291240 -297700 291420 -297500
rect 294240 -297700 294420 -297500
rect 297240 -297700 297420 -297500
rect 560 -297980 2120 -297920
rect 3560 -297980 5120 -297920
rect 6560 -297980 8120 -297920
rect 9560 -297980 11120 -297920
rect 12560 -297980 14120 -297920
rect 15560 -297980 17120 -297920
rect 18560 -297980 20120 -297920
rect 21560 -297980 23120 -297920
rect 24560 -297980 26120 -297920
rect 27560 -297980 29120 -297920
rect 30560 -297980 32120 -297920
rect 33560 -297980 35120 -297920
rect 36560 -297980 38120 -297920
rect 39560 -297980 41120 -297920
rect 42560 -297980 44120 -297920
rect 45560 -297980 47120 -297920
rect 48560 -297980 50120 -297920
rect 51560 -297980 53120 -297920
rect 54560 -297980 56120 -297920
rect 57560 -297980 59120 -297920
rect 60560 -297980 62120 -297920
rect 63560 -297980 65120 -297920
rect 66560 -297980 68120 -297920
rect 69560 -297980 71120 -297920
rect 72560 -297980 74120 -297920
rect 75560 -297980 77120 -297920
rect 78560 -297980 80120 -297920
rect 81560 -297980 83120 -297920
rect 84560 -297980 86120 -297920
rect 87560 -297980 89120 -297920
rect 90560 -297980 92120 -297920
rect 93560 -297980 95120 -297920
rect 96560 -297980 98120 -297920
rect 99560 -297980 101120 -297920
rect 102560 -297980 104120 -297920
rect 105560 -297980 107120 -297920
rect 108560 -297980 110120 -297920
rect 111560 -297980 113120 -297920
rect 114560 -297980 116120 -297920
rect 117560 -297980 119120 -297920
rect 120560 -297980 122120 -297920
rect 123560 -297980 125120 -297920
rect 126560 -297980 128120 -297920
rect 129560 -297980 131120 -297920
rect 132560 -297980 134120 -297920
rect 135560 -297980 137120 -297920
rect 138560 -297980 140120 -297920
rect 141560 -297980 143120 -297920
rect 144560 -297980 146120 -297920
rect 147560 -297980 149120 -297920
rect 150560 -297980 152120 -297920
rect 153560 -297980 155120 -297920
rect 156560 -297980 158120 -297920
rect 159560 -297980 161120 -297920
rect 162560 -297980 164120 -297920
rect 165560 -297980 167120 -297920
rect 168560 -297980 170120 -297920
rect 171560 -297980 173120 -297920
rect 174560 -297980 176120 -297920
rect 177560 -297980 179120 -297920
rect 180560 -297980 182120 -297920
rect 183560 -297980 185120 -297920
rect 186560 -297980 188120 -297920
rect 189560 -297980 191120 -297920
rect 192560 -297980 194120 -297920
rect 195560 -297980 197120 -297920
rect 198560 -297980 200120 -297920
rect 201560 -297980 203120 -297920
rect 204560 -297980 206120 -297920
rect 207560 -297980 209120 -297920
rect 210560 -297980 212120 -297920
rect 213560 -297980 215120 -297920
rect 216560 -297980 218120 -297920
rect 219560 -297980 221120 -297920
rect 222560 -297980 224120 -297920
rect 225560 -297980 227120 -297920
rect 228560 -297980 230120 -297920
rect 231560 -297980 233120 -297920
rect 234560 -297980 236120 -297920
rect 237560 -297980 239120 -297920
rect 240560 -297980 242120 -297920
rect 243560 -297980 245120 -297920
rect 246560 -297980 248120 -297920
rect 249560 -297980 251120 -297920
rect 252560 -297980 254120 -297920
rect 255560 -297980 257120 -297920
rect 258560 -297980 260120 -297920
rect 261560 -297980 263120 -297920
rect 264560 -297980 266120 -297920
rect 267560 -297980 269120 -297920
rect 270560 -297980 272120 -297920
rect 273560 -297980 275120 -297920
rect 276560 -297980 278120 -297920
rect 279560 -297980 281120 -297920
rect 282560 -297980 284120 -297920
rect 285560 -297980 287120 -297920
rect 288560 -297980 290120 -297920
rect 291560 -297980 293120 -297920
rect 294560 -297980 296120 -297920
rect 297560 -297980 299120 -297920
<< metal1 >>
rect -1940 3450 299000 3460
rect -1940 3360 -1920 3450
rect -900 3360 50 3450
rect 140 3360 3050 3450
rect 3140 3360 6050 3450
rect 6140 3360 9050 3450
rect 9140 3360 12050 3450
rect 12140 3360 15050 3450
rect 15140 3360 18050 3450
rect 18140 3360 21050 3450
rect 21140 3360 24050 3450
rect 24140 3360 27050 3450
rect 27140 3360 30050 3450
rect 30140 3360 33050 3450
rect 33140 3360 36050 3450
rect 36140 3360 39050 3450
rect 39140 3360 42050 3450
rect 42140 3360 45050 3450
rect 45140 3360 48050 3450
rect 48140 3360 51050 3450
rect 51140 3360 54050 3450
rect 54140 3360 57050 3450
rect 57140 3360 60050 3450
rect 60140 3360 63050 3450
rect 63140 3360 66050 3450
rect 66140 3360 69050 3450
rect 69140 3360 72050 3450
rect 72140 3360 75050 3450
rect 75140 3360 78050 3450
rect 78140 3360 81050 3450
rect 81140 3360 84050 3450
rect 84140 3360 87050 3450
rect 87140 3360 90050 3450
rect 90140 3360 93050 3450
rect 93140 3360 96050 3450
rect 96140 3360 99050 3450
rect 99140 3360 102050 3450
rect 102140 3360 105050 3450
rect 105140 3360 108050 3450
rect 108140 3360 111050 3450
rect 111140 3360 114050 3450
rect 114140 3360 117050 3450
rect 117140 3360 120050 3450
rect 120140 3360 123050 3450
rect 123140 3360 126050 3450
rect 126140 3360 129050 3450
rect 129140 3360 132050 3450
rect 132140 3360 135050 3450
rect 135140 3360 138050 3450
rect 138140 3360 141050 3450
rect 141140 3360 144050 3450
rect 144140 3360 147050 3450
rect 147140 3360 150050 3450
rect 150140 3360 153050 3450
rect 153140 3360 156050 3450
rect 156140 3360 159050 3450
rect 159140 3360 162050 3450
rect 162140 3360 165050 3450
rect 165140 3360 168050 3450
rect 168140 3360 171050 3450
rect 171140 3360 174050 3450
rect 174140 3360 177050 3450
rect 177140 3360 180050 3450
rect 180140 3360 183050 3450
rect 183140 3360 186050 3450
rect 186140 3360 189050 3450
rect 189140 3360 192050 3450
rect 192140 3360 195050 3450
rect 195140 3360 198050 3450
rect 198140 3360 201050 3450
rect 201140 3360 204050 3450
rect 204140 3360 207050 3450
rect 207140 3360 210050 3450
rect 210140 3360 213050 3450
rect 213140 3360 216050 3450
rect 216140 3360 219050 3450
rect 219140 3360 222050 3450
rect 222140 3360 225050 3450
rect 225140 3360 228050 3450
rect 228140 3360 231050 3450
rect 231140 3360 234050 3450
rect 234140 3360 237050 3450
rect 237140 3360 240050 3450
rect 240140 3360 243050 3450
rect 243140 3360 246050 3450
rect 246140 3360 249050 3450
rect 249140 3360 252050 3450
rect 252140 3360 255050 3450
rect 255140 3360 258050 3450
rect 258140 3360 261050 3450
rect 261140 3360 264050 3450
rect 264140 3360 267050 3450
rect 267140 3360 270050 3450
rect 270140 3360 273050 3450
rect 273140 3360 276050 3450
rect 276140 3360 279050 3450
rect 279140 3360 282050 3450
rect 282140 3360 285050 3450
rect 285140 3360 288050 3450
rect 288140 3360 291050 3450
rect 291140 3360 294050 3450
rect 294140 3360 297050 3450
rect 297140 3360 299000 3450
rect -1940 3350 299000 3360
rect -2000 2970 -1800 3000
rect -2000 2820 0 2970
rect -2000 -30 -1800 2820
rect -1600 1560 0 1570
rect -1600 1490 -1580 1560
rect -1180 1490 -540 1560
rect -260 1490 0 1560
rect -1600 1480 0 1490
rect 300400 180 300600 3030
rect 300000 30 300600 180
rect -2000 -180 0 -30
rect -2000 -3030 -1800 -180
rect -1600 -1440 0 -1430
rect -1600 -1510 -1580 -1440
rect -1180 -1510 -540 -1440
rect -260 -1510 0 -1440
rect -1600 -1520 0 -1510
rect 300400 -2820 300600 30
rect 300000 -2970 300600 -2820
rect -2000 -3180 0 -3030
rect -2000 -6030 -1800 -3180
rect -1600 -4440 0 -4430
rect -1600 -4510 -1580 -4440
rect -1180 -4510 -540 -4440
rect -260 -4510 0 -4440
rect -1600 -4520 0 -4510
rect 300400 -5820 300600 -2970
rect 300000 -5970 300600 -5820
rect -2000 -6180 0 -6030
rect -2000 -9030 -1800 -6180
rect -1600 -7440 0 -7430
rect -1600 -7510 -1580 -7440
rect -1180 -7510 -540 -7440
rect -260 -7510 0 -7440
rect -1600 -7520 0 -7510
rect 300400 -8820 300600 -5970
rect 300000 -8970 300600 -8820
rect -2000 -9180 0 -9030
rect -2000 -12030 -1800 -9180
rect -1600 -10440 0 -10430
rect -1600 -10510 -1580 -10440
rect -1180 -10510 -540 -10440
rect -260 -10510 0 -10440
rect -1600 -10520 0 -10510
rect 300400 -11820 300600 -8970
rect 300000 -11970 300600 -11820
rect -2000 -12180 0 -12030
rect -2000 -15030 -1800 -12180
rect -1600 -13440 0 -13430
rect -1600 -13510 -1580 -13440
rect -1180 -13510 -540 -13440
rect -260 -13510 0 -13440
rect -1600 -13520 0 -13510
rect 300400 -14820 300600 -11970
rect 300000 -14970 300600 -14820
rect -2000 -15180 0 -15030
rect -2000 -18030 -1800 -15180
rect -1600 -16440 0 -16430
rect -1600 -16510 -1580 -16440
rect -1180 -16510 -540 -16440
rect -260 -16510 0 -16440
rect -1600 -16520 0 -16510
rect 300400 -17820 300600 -14970
rect 300000 -17970 300600 -17820
rect -2000 -18180 0 -18030
rect -2000 -21030 -1800 -18180
rect -1600 -19440 0 -19430
rect -1600 -19510 -1580 -19440
rect -1180 -19510 -540 -19440
rect -260 -19510 0 -19440
rect -1600 -19520 0 -19510
rect 300400 -20820 300600 -17970
rect 300000 -20970 300600 -20820
rect -2000 -21180 0 -21030
rect -2000 -24030 -1800 -21180
rect -1600 -22440 0 -22430
rect -1600 -22510 -1580 -22440
rect -1180 -22510 -540 -22440
rect -260 -22510 0 -22440
rect -1600 -22520 0 -22510
rect 300400 -23820 300600 -20970
rect 300000 -23970 300600 -23820
rect -2000 -24180 0 -24030
rect -2000 -27030 -1800 -24180
rect -1600 -25440 0 -25430
rect -1600 -25510 -1580 -25440
rect -1180 -25510 -540 -25440
rect -260 -25510 0 -25440
rect -1600 -25520 0 -25510
rect 300400 -26820 300600 -23970
rect 300000 -26970 300600 -26820
rect -2000 -27180 0 -27030
rect -2000 -30030 -1800 -27180
rect -1600 -28440 0 -28430
rect -1600 -28510 -1580 -28440
rect -1180 -28510 -540 -28440
rect -260 -28510 0 -28440
rect -1600 -28520 0 -28510
rect 300400 -29820 300600 -26970
rect 300000 -29970 300600 -29820
rect -2000 -30180 0 -30030
rect -2000 -33030 -1800 -30180
rect -1600 -31440 0 -31430
rect -1600 -31510 -1580 -31440
rect -1180 -31510 -540 -31440
rect -260 -31510 0 -31440
rect -1600 -31520 0 -31510
rect 300400 -32820 300600 -29970
rect 300000 -32970 300600 -32820
rect -2000 -33180 0 -33030
rect -2000 -36030 -1800 -33180
rect -1600 -34440 0 -34430
rect -1600 -34510 -1580 -34440
rect -1180 -34510 -540 -34440
rect -260 -34510 0 -34440
rect -1600 -34520 0 -34510
rect 300400 -35820 300600 -32970
rect 300000 -35970 300600 -35820
rect -2000 -36180 0 -36030
rect -2000 -39030 -1800 -36180
rect -1600 -37440 0 -37430
rect -1600 -37510 -1580 -37440
rect -1180 -37510 -540 -37440
rect -260 -37510 0 -37440
rect -1600 -37520 0 -37510
rect 300400 -38820 300600 -35970
rect 300000 -38970 300600 -38820
rect -2000 -39180 0 -39030
rect -2000 -42030 -1800 -39180
rect -1600 -40440 0 -40430
rect -1600 -40510 -1580 -40440
rect -1180 -40510 -540 -40440
rect -260 -40510 0 -40440
rect -1600 -40520 0 -40510
rect 300400 -41820 300600 -38970
rect 300000 -41970 300600 -41820
rect -2000 -42180 0 -42030
rect -2000 -45030 -1800 -42180
rect -1600 -43440 0 -43430
rect -1600 -43510 -1580 -43440
rect -1180 -43510 -540 -43440
rect -260 -43510 0 -43440
rect -1600 -43520 0 -43510
rect 300400 -44820 300600 -41970
rect 300000 -44970 300600 -44820
rect -2000 -45180 0 -45030
rect -2000 -48030 -1800 -45180
rect -1600 -46440 0 -46430
rect -1600 -46510 -1580 -46440
rect -1180 -46510 -540 -46440
rect -260 -46510 0 -46440
rect -1600 -46520 0 -46510
rect 300400 -47820 300600 -44970
rect 300000 -47970 300600 -47820
rect -2000 -48180 0 -48030
rect -2000 -51030 -1800 -48180
rect -1600 -49440 0 -49430
rect -1600 -49510 -1580 -49440
rect -1180 -49510 -540 -49440
rect -260 -49510 0 -49440
rect -1600 -49520 0 -49510
rect 300400 -50820 300600 -47970
rect 300000 -50970 300600 -50820
rect -2000 -51180 0 -51030
rect -2000 -54030 -1800 -51180
rect -1600 -52440 0 -52430
rect -1600 -52510 -1580 -52440
rect -1180 -52510 -540 -52440
rect -260 -52510 0 -52440
rect -1600 -52520 0 -52510
rect 300400 -53820 300600 -50970
rect 300000 -53970 300600 -53820
rect -2000 -54180 0 -54030
rect -2000 -57030 -1800 -54180
rect -1600 -55440 0 -55430
rect -1600 -55510 -1580 -55440
rect -1180 -55510 -540 -55440
rect -260 -55510 0 -55440
rect -1600 -55520 0 -55510
rect 300400 -56820 300600 -53970
rect 300000 -56970 300600 -56820
rect -2000 -57180 0 -57030
rect -2000 -60030 -1800 -57180
rect -1600 -58440 0 -58430
rect -1600 -58510 -1580 -58440
rect -1180 -58510 -540 -58440
rect -260 -58510 0 -58440
rect -1600 -58520 0 -58510
rect 300400 -59820 300600 -56970
rect 300000 -59970 300600 -59820
rect -2000 -60180 0 -60030
rect -2000 -63030 -1800 -60180
rect -1600 -61440 0 -61430
rect -1600 -61510 -1580 -61440
rect -1180 -61510 -540 -61440
rect -260 -61510 0 -61440
rect -1600 -61520 0 -61510
rect 300400 -62820 300600 -59970
rect 300000 -62970 300600 -62820
rect -2000 -63180 0 -63030
rect -2000 -66030 -1800 -63180
rect -1600 -64440 0 -64430
rect -1600 -64510 -1580 -64440
rect -1180 -64510 -540 -64440
rect -260 -64510 0 -64440
rect -1600 -64520 0 -64510
rect 300400 -65820 300600 -62970
rect 300000 -65970 300600 -65820
rect -2000 -66180 0 -66030
rect -2000 -69030 -1800 -66180
rect -1600 -67440 0 -67430
rect -1600 -67510 -1580 -67440
rect -1180 -67510 -540 -67440
rect -260 -67510 0 -67440
rect -1600 -67520 0 -67510
rect 300400 -68820 300600 -65970
rect 300000 -68970 300600 -68820
rect -2000 -69180 0 -69030
rect -2000 -72030 -1800 -69180
rect -1600 -70440 0 -70430
rect -1600 -70510 -1580 -70440
rect -1180 -70510 -540 -70440
rect -260 -70510 0 -70440
rect -1600 -70520 0 -70510
rect 300400 -71820 300600 -68970
rect 300000 -71970 300600 -71820
rect -2000 -72180 0 -72030
rect -2000 -75030 -1800 -72180
rect -1600 -73440 0 -73430
rect -1600 -73510 -1580 -73440
rect -1180 -73510 -540 -73440
rect -260 -73510 0 -73440
rect -1600 -73520 0 -73510
rect 300400 -74820 300600 -71970
rect 300000 -74970 300600 -74820
rect -2000 -75180 0 -75030
rect -2000 -78030 -1800 -75180
rect -1600 -76440 0 -76430
rect -1600 -76510 -1580 -76440
rect -1180 -76510 -540 -76440
rect -260 -76510 0 -76440
rect -1600 -76520 0 -76510
rect 300400 -77820 300600 -74970
rect 300000 -77970 300600 -77820
rect -2000 -78180 0 -78030
rect -2000 -81030 -1800 -78180
rect -1600 -79440 0 -79430
rect -1600 -79510 -1580 -79440
rect -1180 -79510 -540 -79440
rect -260 -79510 0 -79440
rect -1600 -79520 0 -79510
rect 300400 -80820 300600 -77970
rect 300000 -80970 300600 -80820
rect -2000 -81180 0 -81030
rect -2000 -84030 -1800 -81180
rect -1600 -82440 0 -82430
rect -1600 -82510 -1580 -82440
rect -1180 -82510 -540 -82440
rect -260 -82510 0 -82440
rect -1600 -82520 0 -82510
rect 300400 -83820 300600 -80970
rect 300000 -83970 300600 -83820
rect -2000 -84180 0 -84030
rect -2000 -87030 -1800 -84180
rect -1600 -85440 0 -85430
rect -1600 -85510 -1580 -85440
rect -1180 -85510 -540 -85440
rect -260 -85510 0 -85440
rect -1600 -85520 0 -85510
rect 300400 -86820 300600 -83970
rect 300000 -86970 300600 -86820
rect -2000 -87180 0 -87030
rect -2000 -90030 -1800 -87180
rect -1600 -88440 0 -88430
rect -1600 -88510 -1580 -88440
rect -1180 -88510 -540 -88440
rect -260 -88510 0 -88440
rect -1600 -88520 0 -88510
rect 300400 -89820 300600 -86970
rect 300000 -89970 300600 -89820
rect -2000 -90180 0 -90030
rect -2000 -93030 -1800 -90180
rect -1600 -91440 0 -91430
rect -1600 -91510 -1580 -91440
rect -1180 -91510 -540 -91440
rect -260 -91510 0 -91440
rect -1600 -91520 0 -91510
rect 300400 -92820 300600 -89970
rect 300000 -92970 300600 -92820
rect -2000 -93180 0 -93030
rect -2000 -96030 -1800 -93180
rect -1600 -94440 0 -94430
rect -1600 -94510 -1580 -94440
rect -1180 -94510 -540 -94440
rect -260 -94510 0 -94440
rect -1600 -94520 0 -94510
rect 300400 -95820 300600 -92970
rect 300000 -95970 300600 -95820
rect -2000 -96180 0 -96030
rect -2000 -99030 -1800 -96180
rect -1600 -97440 0 -97430
rect -1600 -97510 -1580 -97440
rect -1180 -97510 -540 -97440
rect -260 -97510 0 -97440
rect -1600 -97520 0 -97510
rect 300400 -98820 300600 -95970
rect 300000 -98970 300600 -98820
rect -2000 -99180 0 -99030
rect -2000 -102030 -1800 -99180
rect -1600 -100440 0 -100430
rect -1600 -100510 -1580 -100440
rect -1180 -100510 -540 -100440
rect -260 -100510 0 -100440
rect -1600 -100520 0 -100510
rect 300400 -101820 300600 -98970
rect 300000 -101970 300600 -101820
rect -2000 -102180 0 -102030
rect -2000 -105030 -1800 -102180
rect -1600 -103440 0 -103430
rect -1600 -103510 -1580 -103440
rect -1180 -103510 -540 -103440
rect -260 -103510 0 -103440
rect -1600 -103520 0 -103510
rect 300400 -104820 300600 -101970
rect 300000 -104970 300600 -104820
rect -2000 -105180 0 -105030
rect -2000 -108030 -1800 -105180
rect -1600 -106440 0 -106430
rect -1600 -106510 -1580 -106440
rect -1180 -106510 -540 -106440
rect -260 -106510 0 -106440
rect -1600 -106520 0 -106510
rect 300400 -107820 300600 -104970
rect 300000 -107970 300600 -107820
rect -2000 -108180 0 -108030
rect -2000 -111030 -1800 -108180
rect -1600 -109440 0 -109430
rect -1600 -109510 -1580 -109440
rect -1180 -109510 -540 -109440
rect -260 -109510 0 -109440
rect -1600 -109520 0 -109510
rect 300400 -110820 300600 -107970
rect 300000 -110970 300600 -110820
rect -2000 -111180 0 -111030
rect -2000 -114030 -1800 -111180
rect -1600 -112440 0 -112430
rect -1600 -112510 -1580 -112440
rect -1180 -112510 -540 -112440
rect -260 -112510 0 -112440
rect -1600 -112520 0 -112510
rect 300400 -113820 300600 -110970
rect 300000 -113970 300600 -113820
rect -2000 -114180 0 -114030
rect -2000 -117030 -1800 -114180
rect -1600 -115440 0 -115430
rect -1600 -115510 -1580 -115440
rect -1180 -115510 -540 -115440
rect -260 -115510 0 -115440
rect -1600 -115520 0 -115510
rect 300400 -116820 300600 -113970
rect 300000 -116970 300600 -116820
rect -2000 -117180 0 -117030
rect -2000 -120030 -1800 -117180
rect -1600 -118440 0 -118430
rect -1600 -118510 -1580 -118440
rect -1180 -118510 -540 -118440
rect -260 -118510 0 -118440
rect -1600 -118520 0 -118510
rect 300400 -119820 300600 -116970
rect 300000 -119970 300600 -119820
rect -2000 -120180 0 -120030
rect -2000 -123030 -1800 -120180
rect -1600 -121440 0 -121430
rect -1600 -121510 -1580 -121440
rect -1180 -121510 -540 -121440
rect -260 -121510 0 -121440
rect -1600 -121520 0 -121510
rect 300400 -122820 300600 -119970
rect 300000 -122970 300600 -122820
rect -2000 -123180 0 -123030
rect -2000 -126030 -1800 -123180
rect -1600 -124440 0 -124430
rect -1600 -124510 -1580 -124440
rect -1180 -124510 -540 -124440
rect -260 -124510 0 -124440
rect -1600 -124520 0 -124510
rect 300400 -125820 300600 -122970
rect 300000 -125970 300600 -125820
rect -2000 -126180 0 -126030
rect -2000 -129030 -1800 -126180
rect -1600 -127440 0 -127430
rect -1600 -127510 -1580 -127440
rect -1180 -127510 -540 -127440
rect -260 -127510 0 -127440
rect -1600 -127520 0 -127510
rect 300400 -128820 300600 -125970
rect 300000 -128970 300600 -128820
rect -2000 -129180 0 -129030
rect -2000 -132030 -1800 -129180
rect -1600 -130440 0 -130430
rect -1600 -130510 -1580 -130440
rect -1180 -130510 -540 -130440
rect -260 -130510 0 -130440
rect -1600 -130520 0 -130510
rect 300400 -131820 300600 -128970
rect 300000 -131970 300600 -131820
rect -2000 -132180 0 -132030
rect -2000 -135030 -1800 -132180
rect -1600 -133440 0 -133430
rect -1600 -133510 -1580 -133440
rect -1180 -133510 -540 -133440
rect -260 -133510 0 -133440
rect -1600 -133520 0 -133510
rect 300400 -134820 300600 -131970
rect 300000 -134970 300600 -134820
rect -2000 -135180 0 -135030
rect -2000 -138030 -1800 -135180
rect -1600 -136440 0 -136430
rect -1600 -136510 -1580 -136440
rect -1180 -136510 -540 -136440
rect -260 -136510 0 -136440
rect -1600 -136520 0 -136510
rect 300400 -137820 300600 -134970
rect 300000 -137970 300600 -137820
rect -2000 -138180 0 -138030
rect -2000 -141030 -1800 -138180
rect -1600 -139440 0 -139430
rect -1600 -139510 -1580 -139440
rect -1180 -139510 -540 -139440
rect -260 -139510 0 -139440
rect -1600 -139520 0 -139510
rect 300400 -140820 300600 -137970
rect 300000 -140970 300600 -140820
rect -2000 -141180 0 -141030
rect -2000 -144030 -1800 -141180
rect -1600 -142440 0 -142430
rect -1600 -142510 -1580 -142440
rect -1180 -142510 -540 -142440
rect -260 -142510 0 -142440
rect -1600 -142520 0 -142510
rect 300400 -143820 300600 -140970
rect 300000 -143970 300600 -143820
rect -2000 -144180 0 -144030
rect -2000 -147030 -1800 -144180
rect -1600 -145440 0 -145430
rect -1600 -145510 -1580 -145440
rect -1180 -145510 -540 -145440
rect -260 -145510 0 -145440
rect -1600 -145520 0 -145510
rect 300400 -146820 300600 -143970
rect 300000 -146970 300600 -146820
rect -2000 -147180 0 -147030
rect -2000 -150030 -1800 -147180
rect -1600 -148440 0 -148430
rect -1600 -148510 -1580 -148440
rect -1180 -148510 -540 -148440
rect -260 -148510 0 -148440
rect -1600 -148520 0 -148510
rect 300400 -149820 300600 -146970
rect 300000 -149970 300600 -149820
rect -2000 -150180 0 -150030
rect -2000 -153030 -1800 -150180
rect -1600 -151440 0 -151430
rect -1600 -151510 -1580 -151440
rect -1180 -151510 -540 -151440
rect -260 -151510 0 -151440
rect -1600 -151520 0 -151510
rect 300400 -152820 300600 -149970
rect 300000 -152970 300600 -152820
rect -2000 -153180 0 -153030
rect -2000 -156030 -1800 -153180
rect -1600 -154440 0 -154430
rect -1600 -154510 -1580 -154440
rect -1180 -154510 -540 -154440
rect -260 -154510 0 -154440
rect -1600 -154520 0 -154510
rect 300400 -155820 300600 -152970
rect 300000 -155970 300600 -155820
rect -2000 -156180 0 -156030
rect -2000 -159030 -1800 -156180
rect -1600 -157440 0 -157430
rect -1600 -157510 -1580 -157440
rect -1180 -157510 -540 -157440
rect -260 -157510 0 -157440
rect -1600 -157520 0 -157510
rect 300400 -158820 300600 -155970
rect 300000 -158970 300600 -158820
rect -2000 -159180 0 -159030
rect -2000 -162030 -1800 -159180
rect -1600 -160440 0 -160430
rect -1600 -160510 -1580 -160440
rect -1180 -160510 -540 -160440
rect -260 -160510 0 -160440
rect -1600 -160520 0 -160510
rect 300400 -161820 300600 -158970
rect 300000 -161970 300600 -161820
rect -2000 -162180 0 -162030
rect -2000 -165030 -1800 -162180
rect -1600 -163440 0 -163430
rect -1600 -163510 -1580 -163440
rect -1180 -163510 -540 -163440
rect -260 -163510 0 -163440
rect -1600 -163520 0 -163510
rect 300400 -164820 300600 -161970
rect 300000 -164970 300600 -164820
rect -2000 -165180 0 -165030
rect -2000 -168030 -1800 -165180
rect -1600 -166440 0 -166430
rect -1600 -166510 -1580 -166440
rect -1180 -166510 -540 -166440
rect -260 -166510 0 -166440
rect -1600 -166520 0 -166510
rect 300400 -167820 300600 -164970
rect 300000 -167970 300600 -167820
rect -2000 -168180 0 -168030
rect -2000 -171030 -1800 -168180
rect -1600 -169440 0 -169430
rect -1600 -169510 -1580 -169440
rect -1180 -169510 -540 -169440
rect -260 -169510 0 -169440
rect -1600 -169520 0 -169510
rect 300400 -170820 300600 -167970
rect 300000 -170970 300600 -170820
rect -2000 -171180 0 -171030
rect -2000 -174030 -1800 -171180
rect -1600 -172440 0 -172430
rect -1600 -172510 -1580 -172440
rect -1180 -172510 -540 -172440
rect -260 -172510 0 -172440
rect -1600 -172520 0 -172510
rect 300400 -173820 300600 -170970
rect 300000 -173970 300600 -173820
rect -2000 -174180 0 -174030
rect -2000 -177030 -1800 -174180
rect -1600 -175440 0 -175430
rect -1600 -175510 -1580 -175440
rect -1180 -175510 -540 -175440
rect -260 -175510 0 -175440
rect -1600 -175520 0 -175510
rect 300400 -176820 300600 -173970
rect 300000 -176970 300600 -176820
rect -2000 -177180 0 -177030
rect -2000 -180030 -1800 -177180
rect -1600 -178440 0 -178430
rect -1600 -178510 -1580 -178440
rect -1180 -178510 -540 -178440
rect -260 -178510 0 -178440
rect -1600 -178520 0 -178510
rect 300400 -179820 300600 -176970
rect 300000 -179970 300600 -179820
rect -2000 -180180 0 -180030
rect -2000 -183030 -1800 -180180
rect -1600 -181440 0 -181430
rect -1600 -181510 -1580 -181440
rect -1180 -181510 -540 -181440
rect -260 -181510 0 -181440
rect -1600 -181520 0 -181510
rect 300400 -182820 300600 -179970
rect 300000 -182970 300600 -182820
rect -2000 -183180 0 -183030
rect -2000 -186030 -1800 -183180
rect -1600 -184440 0 -184430
rect -1600 -184510 -1580 -184440
rect -1180 -184510 -540 -184440
rect -260 -184510 0 -184440
rect -1600 -184520 0 -184510
rect 300400 -185820 300600 -182970
rect 300000 -185970 300600 -185820
rect -2000 -186180 0 -186030
rect -2000 -189030 -1800 -186180
rect -1600 -187440 0 -187430
rect -1600 -187510 -1580 -187440
rect -1180 -187510 -540 -187440
rect -260 -187510 0 -187440
rect -1600 -187520 0 -187510
rect 300400 -188820 300600 -185970
rect 300000 -188970 300600 -188820
rect -2000 -189180 0 -189030
rect -2000 -192030 -1800 -189180
rect -1600 -190440 0 -190430
rect -1600 -190510 -1580 -190440
rect -1180 -190510 -540 -190440
rect -260 -190510 0 -190440
rect -1600 -190520 0 -190510
rect 300400 -191820 300600 -188970
rect 300000 -191970 300600 -191820
rect -2000 -192180 0 -192030
rect -2000 -195030 -1800 -192180
rect -1600 -193440 0 -193430
rect -1600 -193510 -1580 -193440
rect -1180 -193510 -540 -193440
rect -260 -193510 0 -193440
rect -1600 -193520 0 -193510
rect 300400 -194820 300600 -191970
rect 300000 -194970 300600 -194820
rect -2000 -195180 0 -195030
rect -2000 -198030 -1800 -195180
rect -1600 -196440 0 -196430
rect -1600 -196510 -1580 -196440
rect -1180 -196510 -540 -196440
rect -260 -196510 0 -196440
rect -1600 -196520 0 -196510
rect 300400 -197820 300600 -194970
rect 300000 -197970 300600 -197820
rect -2000 -198180 0 -198030
rect -2000 -201030 -1800 -198180
rect -1600 -199440 0 -199430
rect -1600 -199510 -1580 -199440
rect -1180 -199510 -540 -199440
rect -260 -199510 0 -199440
rect -1600 -199520 0 -199510
rect 300400 -200820 300600 -197970
rect 300000 -200970 300600 -200820
rect -2000 -201180 0 -201030
rect -2000 -204030 -1800 -201180
rect -1600 -202440 0 -202430
rect -1600 -202510 -1580 -202440
rect -1180 -202510 -540 -202440
rect -260 -202510 0 -202440
rect -1600 -202520 0 -202510
rect 300400 -203820 300600 -200970
rect 300000 -203970 300600 -203820
rect -2000 -204180 0 -204030
rect -2000 -207030 -1800 -204180
rect -1600 -205440 0 -205430
rect -1600 -205510 -1580 -205440
rect -1180 -205510 -540 -205440
rect -260 -205510 0 -205440
rect -1600 -205520 0 -205510
rect 300400 -206820 300600 -203970
rect 300000 -206970 300600 -206820
rect -2000 -207180 0 -207030
rect -2000 -210030 -1800 -207180
rect -1600 -208440 0 -208430
rect -1600 -208510 -1580 -208440
rect -1180 -208510 -540 -208440
rect -260 -208510 0 -208440
rect -1600 -208520 0 -208510
rect 300400 -209820 300600 -206970
rect 300000 -209970 300600 -209820
rect -2000 -210180 0 -210030
rect -2000 -213030 -1800 -210180
rect -1600 -211440 0 -211430
rect -1600 -211510 -1580 -211440
rect -1180 -211510 -540 -211440
rect -260 -211510 0 -211440
rect -1600 -211520 0 -211510
rect 300400 -212820 300600 -209970
rect 300000 -212970 300600 -212820
rect -2000 -213180 0 -213030
rect -2000 -216030 -1800 -213180
rect -1600 -214440 0 -214430
rect -1600 -214510 -1580 -214440
rect -1180 -214510 -540 -214440
rect -260 -214510 0 -214440
rect -1600 -214520 0 -214510
rect 300400 -215820 300600 -212970
rect 300000 -215970 300600 -215820
rect -2000 -216180 0 -216030
rect -2000 -219030 -1800 -216180
rect -1600 -217440 0 -217430
rect -1600 -217510 -1580 -217440
rect -1180 -217510 -540 -217440
rect -260 -217510 0 -217440
rect -1600 -217520 0 -217510
rect 300400 -218820 300600 -215970
rect 300000 -218970 300600 -218820
rect -2000 -219180 0 -219030
rect -2000 -222030 -1800 -219180
rect -1600 -220440 0 -220430
rect -1600 -220510 -1580 -220440
rect -1180 -220510 -540 -220440
rect -260 -220510 0 -220440
rect -1600 -220520 0 -220510
rect 300400 -221820 300600 -218970
rect 300000 -221970 300600 -221820
rect -2000 -222180 0 -222030
rect -2000 -225030 -1800 -222180
rect -1600 -223440 0 -223430
rect -1600 -223510 -1580 -223440
rect -1180 -223510 -540 -223440
rect -260 -223510 0 -223440
rect -1600 -223520 0 -223510
rect 300400 -224820 300600 -221970
rect 300000 -224970 300600 -224820
rect -2000 -225180 0 -225030
rect -2000 -228030 -1800 -225180
rect -1600 -226440 0 -226430
rect -1600 -226510 -1580 -226440
rect -1180 -226510 -540 -226440
rect -260 -226510 0 -226440
rect -1600 -226520 0 -226510
rect 300400 -227820 300600 -224970
rect 300000 -227970 300600 -227820
rect -2000 -228180 0 -228030
rect -2000 -231030 -1800 -228180
rect -1600 -229440 0 -229430
rect -1600 -229510 -1580 -229440
rect -1180 -229510 -540 -229440
rect -260 -229510 0 -229440
rect -1600 -229520 0 -229510
rect 300400 -230820 300600 -227970
rect 300000 -230970 300600 -230820
rect -2000 -231180 0 -231030
rect -2000 -234030 -1800 -231180
rect -1600 -232440 0 -232430
rect -1600 -232510 -1580 -232440
rect -1180 -232510 -540 -232440
rect -260 -232510 0 -232440
rect -1600 -232520 0 -232510
rect 300400 -233820 300600 -230970
rect 300000 -233970 300600 -233820
rect -2000 -234180 0 -234030
rect -2000 -237030 -1800 -234180
rect -1600 -235440 0 -235430
rect -1600 -235510 -1580 -235440
rect -1180 -235510 -540 -235440
rect -260 -235510 0 -235440
rect -1600 -235520 0 -235510
rect 300400 -236820 300600 -233970
rect 300000 -236970 300600 -236820
rect -2000 -237180 0 -237030
rect -2000 -240030 -1800 -237180
rect -1600 -238440 0 -238430
rect -1600 -238510 -1580 -238440
rect -1180 -238510 -540 -238440
rect -260 -238510 0 -238440
rect -1600 -238520 0 -238510
rect 300400 -239820 300600 -236970
rect 300000 -239970 300600 -239820
rect -2000 -240180 0 -240030
rect -2000 -243030 -1800 -240180
rect -1600 -241440 0 -241430
rect -1600 -241510 -1580 -241440
rect -1180 -241510 -540 -241440
rect -260 -241510 0 -241440
rect -1600 -241520 0 -241510
rect 300400 -242820 300600 -239970
rect 300000 -242970 300600 -242820
rect -2000 -243180 0 -243030
rect -2000 -246030 -1800 -243180
rect -1600 -244440 0 -244430
rect -1600 -244510 -1580 -244440
rect -1180 -244510 -540 -244440
rect -260 -244510 0 -244440
rect -1600 -244520 0 -244510
rect 300400 -245820 300600 -242970
rect 300000 -245970 300600 -245820
rect -2000 -246180 0 -246030
rect -2000 -249030 -1800 -246180
rect -1600 -247440 0 -247430
rect -1600 -247510 -1580 -247440
rect -1180 -247510 -540 -247440
rect -260 -247510 0 -247440
rect -1600 -247520 0 -247510
rect 300400 -248820 300600 -245970
rect 300000 -248970 300600 -248820
rect -2000 -249180 0 -249030
rect -2000 -252030 -1800 -249180
rect -1600 -250440 0 -250430
rect -1600 -250510 -1580 -250440
rect -1180 -250510 -540 -250440
rect -260 -250510 0 -250440
rect -1600 -250520 0 -250510
rect 300400 -251820 300600 -248970
rect 300000 -251970 300600 -251820
rect -2000 -252180 0 -252030
rect -2000 -255030 -1800 -252180
rect -1600 -253440 0 -253430
rect -1600 -253510 -1580 -253440
rect -1180 -253510 -540 -253440
rect -260 -253510 0 -253440
rect -1600 -253520 0 -253510
rect 300400 -254820 300600 -251970
rect 300000 -254970 300600 -254820
rect -2000 -255180 0 -255030
rect -2000 -258030 -1800 -255180
rect -1600 -256440 0 -256430
rect -1600 -256510 -1580 -256440
rect -1180 -256510 -540 -256440
rect -260 -256510 0 -256440
rect -1600 -256520 0 -256510
rect 300400 -257820 300600 -254970
rect 300000 -257970 300600 -257820
rect -2000 -258180 0 -258030
rect -2000 -261030 -1800 -258180
rect -1600 -259440 0 -259430
rect -1600 -259510 -1580 -259440
rect -1180 -259510 -540 -259440
rect -260 -259510 0 -259440
rect -1600 -259520 0 -259510
rect 300400 -260820 300600 -257970
rect 300000 -260970 300600 -260820
rect -2000 -261180 0 -261030
rect -2000 -264030 -1800 -261180
rect -1600 -262440 0 -262430
rect -1600 -262510 -1580 -262440
rect -1180 -262510 -540 -262440
rect -260 -262510 0 -262440
rect -1600 -262520 0 -262510
rect 300400 -263820 300600 -260970
rect 300000 -263970 300600 -263820
rect -2000 -264180 0 -264030
rect -2000 -267030 -1800 -264180
rect -1600 -265440 0 -265430
rect -1600 -265510 -1580 -265440
rect -1180 -265510 -540 -265440
rect -260 -265510 0 -265440
rect -1600 -265520 0 -265510
rect 300400 -266820 300600 -263970
rect 300000 -266970 300600 -266820
rect -2000 -267180 0 -267030
rect -2000 -270030 -1800 -267180
rect -1600 -268440 0 -268430
rect -1600 -268510 -1580 -268440
rect -1180 -268510 -540 -268440
rect -260 -268510 0 -268440
rect -1600 -268520 0 -268510
rect 300400 -269820 300600 -266970
rect 300000 -269970 300600 -269820
rect -2000 -270180 0 -270030
rect -2000 -273030 -1800 -270180
rect -1600 -271440 0 -271430
rect -1600 -271510 -1580 -271440
rect -1180 -271510 -540 -271440
rect -260 -271510 0 -271440
rect -1600 -271520 0 -271510
rect 300400 -272820 300600 -269970
rect 300000 -272970 300600 -272820
rect -2000 -273180 0 -273030
rect -2000 -276030 -1800 -273180
rect -1600 -274440 0 -274430
rect -1600 -274510 -1580 -274440
rect -1180 -274510 -540 -274440
rect -260 -274510 0 -274440
rect -1600 -274520 0 -274510
rect 300400 -275820 300600 -272970
rect 300000 -275970 300600 -275820
rect -2000 -276180 0 -276030
rect -2000 -279030 -1800 -276180
rect -1600 -277440 0 -277430
rect -1600 -277510 -1580 -277440
rect -1180 -277510 -540 -277440
rect -260 -277510 0 -277440
rect -1600 -277520 0 -277510
rect 300400 -278820 300600 -275970
rect 300000 -278970 300600 -278820
rect -2000 -279180 0 -279030
rect -2000 -282030 -1800 -279180
rect -1600 -280440 0 -280430
rect -1600 -280510 -1580 -280440
rect -1180 -280510 -540 -280440
rect -260 -280510 0 -280440
rect -1600 -280520 0 -280510
rect 300400 -281820 300600 -278970
rect 300000 -281970 300600 -281820
rect -2000 -282180 0 -282030
rect -2000 -285030 -1800 -282180
rect -1600 -283440 0 -283430
rect -1600 -283510 -1580 -283440
rect -1180 -283510 -540 -283440
rect -260 -283510 0 -283440
rect -1600 -283520 0 -283510
rect 300400 -284820 300600 -281970
rect 300000 -284970 300600 -284820
rect -2000 -285180 0 -285030
rect -2000 -288030 -1800 -285180
rect -1600 -286440 0 -286430
rect -1600 -286510 -1580 -286440
rect -1180 -286510 -540 -286440
rect -260 -286510 0 -286440
rect -1600 -286520 0 -286510
rect 300400 -287820 300600 -284970
rect 300000 -287970 300600 -287820
rect -2000 -288180 0 -288030
rect -2000 -291030 -1800 -288180
rect -1600 -289440 0 -289430
rect -1600 -289510 -1580 -289440
rect -1180 -289510 -540 -289440
rect -260 -289510 0 -289440
rect -1600 -289520 0 -289510
rect 300400 -290820 300600 -287970
rect 300000 -290970 300600 -290820
rect -2000 -291180 0 -291030
rect -2000 -294030 -1800 -291180
rect -1600 -292440 0 -292430
rect -1600 -292510 -1580 -292440
rect -1180 -292510 -540 -292440
rect -260 -292510 0 -292440
rect -1600 -292520 0 -292510
rect 300400 -293820 300600 -290970
rect 300000 -293970 300600 -293820
rect -2000 -294180 0 -294030
rect -2000 -297000 -1800 -294180
rect -1600 -295440 0 -295430
rect -1600 -295510 -1580 -295440
rect -1180 -295510 -540 -295440
rect -260 -295510 0 -295440
rect -1600 -295520 0 -295510
rect 300400 -296820 300600 -293970
rect 300000 -296970 300600 -296820
rect 540 -297200 560 -297130
rect 2120 -297200 2140 -297130
rect 540 -297230 2140 -297200
rect 540 -297290 560 -297230
rect 2120 -297290 2140 -297230
rect 540 -297300 2140 -297290
rect 3540 -297200 3560 -297130
rect 5120 -297200 5140 -297130
rect 3540 -297230 5140 -297200
rect 3540 -297290 3560 -297230
rect 5120 -297290 5140 -297230
rect 3540 -297300 5140 -297290
rect 6540 -297200 6560 -297130
rect 8120 -297200 8140 -297130
rect 6540 -297230 8140 -297200
rect 6540 -297290 6560 -297230
rect 8120 -297290 8140 -297230
rect 6540 -297300 8140 -297290
rect 9540 -297200 9560 -297130
rect 11120 -297200 11140 -297130
rect 9540 -297230 11140 -297200
rect 9540 -297290 9560 -297230
rect 11120 -297290 11140 -297230
rect 9540 -297300 11140 -297290
rect 12540 -297200 12560 -297130
rect 14120 -297200 14140 -297130
rect 12540 -297230 14140 -297200
rect 12540 -297290 12560 -297230
rect 14120 -297290 14140 -297230
rect 12540 -297300 14140 -297290
rect 15540 -297200 15560 -297130
rect 17120 -297200 17140 -297130
rect 15540 -297230 17140 -297200
rect 15540 -297290 15560 -297230
rect 17120 -297290 17140 -297230
rect 15540 -297300 17140 -297290
rect 18540 -297200 18560 -297130
rect 20120 -297200 20140 -297130
rect 18540 -297230 20140 -297200
rect 18540 -297290 18560 -297230
rect 20120 -297290 20140 -297230
rect 18540 -297300 20140 -297290
rect 21540 -297200 21560 -297130
rect 23120 -297200 23140 -297130
rect 21540 -297230 23140 -297200
rect 21540 -297290 21560 -297230
rect 23120 -297290 23140 -297230
rect 21540 -297300 23140 -297290
rect 24540 -297200 24560 -297130
rect 26120 -297200 26140 -297130
rect 24540 -297230 26140 -297200
rect 24540 -297290 24560 -297230
rect 26120 -297290 26140 -297230
rect 24540 -297300 26140 -297290
rect 27540 -297200 27560 -297130
rect 29120 -297200 29140 -297130
rect 27540 -297230 29140 -297200
rect 27540 -297290 27560 -297230
rect 29120 -297290 29140 -297230
rect 27540 -297300 29140 -297290
rect 30540 -297200 30560 -297130
rect 32120 -297200 32140 -297130
rect 30540 -297230 32140 -297200
rect 30540 -297290 30560 -297230
rect 32120 -297290 32140 -297230
rect 30540 -297300 32140 -297290
rect 33540 -297200 33560 -297130
rect 35120 -297200 35140 -297130
rect 33540 -297230 35140 -297200
rect 33540 -297290 33560 -297230
rect 35120 -297290 35140 -297230
rect 33540 -297300 35140 -297290
rect 36540 -297200 36560 -297130
rect 38120 -297200 38140 -297130
rect 36540 -297230 38140 -297200
rect 36540 -297290 36560 -297230
rect 38120 -297290 38140 -297230
rect 36540 -297300 38140 -297290
rect 39540 -297200 39560 -297130
rect 41120 -297200 41140 -297130
rect 39540 -297230 41140 -297200
rect 39540 -297290 39560 -297230
rect 41120 -297290 41140 -297230
rect 39540 -297300 41140 -297290
rect 42540 -297200 42560 -297130
rect 44120 -297200 44140 -297130
rect 42540 -297230 44140 -297200
rect 42540 -297290 42560 -297230
rect 44120 -297290 44140 -297230
rect 42540 -297300 44140 -297290
rect 45540 -297200 45560 -297130
rect 47120 -297200 47140 -297130
rect 45540 -297230 47140 -297200
rect 45540 -297290 45560 -297230
rect 47120 -297290 47140 -297230
rect 45540 -297300 47140 -297290
rect 48540 -297200 48560 -297130
rect 50120 -297200 50140 -297130
rect 48540 -297230 50140 -297200
rect 48540 -297290 48560 -297230
rect 50120 -297290 50140 -297230
rect 48540 -297300 50140 -297290
rect 51540 -297200 51560 -297130
rect 53120 -297200 53140 -297130
rect 51540 -297230 53140 -297200
rect 51540 -297290 51560 -297230
rect 53120 -297290 53140 -297230
rect 51540 -297300 53140 -297290
rect 54540 -297200 54560 -297130
rect 56120 -297200 56140 -297130
rect 54540 -297230 56140 -297200
rect 54540 -297290 54560 -297230
rect 56120 -297290 56140 -297230
rect 54540 -297300 56140 -297290
rect 57540 -297200 57560 -297130
rect 59120 -297200 59140 -297130
rect 57540 -297230 59140 -297200
rect 57540 -297290 57560 -297230
rect 59120 -297290 59140 -297230
rect 57540 -297300 59140 -297290
rect 60540 -297200 60560 -297130
rect 62120 -297200 62140 -297130
rect 60540 -297230 62140 -297200
rect 60540 -297290 60560 -297230
rect 62120 -297290 62140 -297230
rect 60540 -297300 62140 -297290
rect 63540 -297200 63560 -297130
rect 65120 -297200 65140 -297130
rect 63540 -297230 65140 -297200
rect 63540 -297290 63560 -297230
rect 65120 -297290 65140 -297230
rect 63540 -297300 65140 -297290
rect 66540 -297200 66560 -297130
rect 68120 -297200 68140 -297130
rect 66540 -297230 68140 -297200
rect 66540 -297290 66560 -297230
rect 68120 -297290 68140 -297230
rect 66540 -297300 68140 -297290
rect 69540 -297200 69560 -297130
rect 71120 -297200 71140 -297130
rect 69540 -297230 71140 -297200
rect 69540 -297290 69560 -297230
rect 71120 -297290 71140 -297230
rect 69540 -297300 71140 -297290
rect 72540 -297200 72560 -297130
rect 74120 -297200 74140 -297130
rect 72540 -297230 74140 -297200
rect 72540 -297290 72560 -297230
rect 74120 -297290 74140 -297230
rect 72540 -297300 74140 -297290
rect 75540 -297200 75560 -297130
rect 77120 -297200 77140 -297130
rect 75540 -297230 77140 -297200
rect 75540 -297290 75560 -297230
rect 77120 -297290 77140 -297230
rect 75540 -297300 77140 -297290
rect 78540 -297200 78560 -297130
rect 80120 -297200 80140 -297130
rect 78540 -297230 80140 -297200
rect 78540 -297290 78560 -297230
rect 80120 -297290 80140 -297230
rect 78540 -297300 80140 -297290
rect 81540 -297200 81560 -297130
rect 83120 -297200 83140 -297130
rect 81540 -297230 83140 -297200
rect 81540 -297290 81560 -297230
rect 83120 -297290 83140 -297230
rect 81540 -297300 83140 -297290
rect 84540 -297200 84560 -297130
rect 86120 -297200 86140 -297130
rect 84540 -297230 86140 -297200
rect 84540 -297290 84560 -297230
rect 86120 -297290 86140 -297230
rect 84540 -297300 86140 -297290
rect 87540 -297200 87560 -297130
rect 89120 -297200 89140 -297130
rect 87540 -297230 89140 -297200
rect 87540 -297290 87560 -297230
rect 89120 -297290 89140 -297230
rect 87540 -297300 89140 -297290
rect 90540 -297200 90560 -297130
rect 92120 -297200 92140 -297130
rect 90540 -297230 92140 -297200
rect 90540 -297290 90560 -297230
rect 92120 -297290 92140 -297230
rect 90540 -297300 92140 -297290
rect 93540 -297200 93560 -297130
rect 95120 -297200 95140 -297130
rect 93540 -297230 95140 -297200
rect 93540 -297290 93560 -297230
rect 95120 -297290 95140 -297230
rect 93540 -297300 95140 -297290
rect 96540 -297200 96560 -297130
rect 98120 -297200 98140 -297130
rect 96540 -297230 98140 -297200
rect 96540 -297290 96560 -297230
rect 98120 -297290 98140 -297230
rect 96540 -297300 98140 -297290
rect 99540 -297200 99560 -297130
rect 101120 -297200 101140 -297130
rect 99540 -297230 101140 -297200
rect 99540 -297290 99560 -297230
rect 101120 -297290 101140 -297230
rect 99540 -297300 101140 -297290
rect 102540 -297200 102560 -297130
rect 104120 -297200 104140 -297130
rect 102540 -297230 104140 -297200
rect 102540 -297290 102560 -297230
rect 104120 -297290 104140 -297230
rect 102540 -297300 104140 -297290
rect 105540 -297200 105560 -297130
rect 107120 -297200 107140 -297130
rect 105540 -297230 107140 -297200
rect 105540 -297290 105560 -297230
rect 107120 -297290 107140 -297230
rect 105540 -297300 107140 -297290
rect 108540 -297200 108560 -297130
rect 110120 -297200 110140 -297130
rect 108540 -297230 110140 -297200
rect 108540 -297290 108560 -297230
rect 110120 -297290 110140 -297230
rect 108540 -297300 110140 -297290
rect 111540 -297200 111560 -297130
rect 113120 -297200 113140 -297130
rect 111540 -297230 113140 -297200
rect 111540 -297290 111560 -297230
rect 113120 -297290 113140 -297230
rect 111540 -297300 113140 -297290
rect 114540 -297200 114560 -297130
rect 116120 -297200 116140 -297130
rect 114540 -297230 116140 -297200
rect 114540 -297290 114560 -297230
rect 116120 -297290 116140 -297230
rect 114540 -297300 116140 -297290
rect 117540 -297200 117560 -297130
rect 119120 -297200 119140 -297130
rect 117540 -297230 119140 -297200
rect 117540 -297290 117560 -297230
rect 119120 -297290 119140 -297230
rect 117540 -297300 119140 -297290
rect 120540 -297200 120560 -297130
rect 122120 -297200 122140 -297130
rect 120540 -297230 122140 -297200
rect 120540 -297290 120560 -297230
rect 122120 -297290 122140 -297230
rect 120540 -297300 122140 -297290
rect 123540 -297200 123560 -297130
rect 125120 -297200 125140 -297130
rect 123540 -297230 125140 -297200
rect 123540 -297290 123560 -297230
rect 125120 -297290 125140 -297230
rect 123540 -297300 125140 -297290
rect 126540 -297200 126560 -297130
rect 128120 -297200 128140 -297130
rect 126540 -297230 128140 -297200
rect 126540 -297290 126560 -297230
rect 128120 -297290 128140 -297230
rect 126540 -297300 128140 -297290
rect 129540 -297200 129560 -297130
rect 131120 -297200 131140 -297130
rect 129540 -297230 131140 -297200
rect 129540 -297290 129560 -297230
rect 131120 -297290 131140 -297230
rect 129540 -297300 131140 -297290
rect 132540 -297200 132560 -297130
rect 134120 -297200 134140 -297130
rect 132540 -297230 134140 -297200
rect 132540 -297290 132560 -297230
rect 134120 -297290 134140 -297230
rect 132540 -297300 134140 -297290
rect 135540 -297200 135560 -297130
rect 137120 -297200 137140 -297130
rect 135540 -297230 137140 -297200
rect 135540 -297290 135560 -297230
rect 137120 -297290 137140 -297230
rect 135540 -297300 137140 -297290
rect 138540 -297200 138560 -297130
rect 140120 -297200 140140 -297130
rect 138540 -297230 140140 -297200
rect 138540 -297290 138560 -297230
rect 140120 -297290 140140 -297230
rect 138540 -297300 140140 -297290
rect 141540 -297200 141560 -297130
rect 143120 -297200 143140 -297130
rect 141540 -297230 143140 -297200
rect 141540 -297290 141560 -297230
rect 143120 -297290 143140 -297230
rect 141540 -297300 143140 -297290
rect 144540 -297200 144560 -297130
rect 146120 -297200 146140 -297130
rect 144540 -297230 146140 -297200
rect 144540 -297290 144560 -297230
rect 146120 -297290 146140 -297230
rect 144540 -297300 146140 -297290
rect 147540 -297200 147560 -297130
rect 149120 -297200 149140 -297130
rect 147540 -297230 149140 -297200
rect 147540 -297290 147560 -297230
rect 149120 -297290 149140 -297230
rect 147540 -297300 149140 -297290
rect 150540 -297200 150560 -297130
rect 152120 -297200 152140 -297130
rect 150540 -297230 152140 -297200
rect 150540 -297290 150560 -297230
rect 152120 -297290 152140 -297230
rect 150540 -297300 152140 -297290
rect 153540 -297200 153560 -297130
rect 155120 -297200 155140 -297130
rect 153540 -297230 155140 -297200
rect 153540 -297290 153560 -297230
rect 155120 -297290 155140 -297230
rect 153540 -297300 155140 -297290
rect 156540 -297200 156560 -297130
rect 158120 -297200 158140 -297130
rect 156540 -297230 158140 -297200
rect 156540 -297290 156560 -297230
rect 158120 -297290 158140 -297230
rect 156540 -297300 158140 -297290
rect 159540 -297200 159560 -297130
rect 161120 -297200 161140 -297130
rect 159540 -297230 161140 -297200
rect 159540 -297290 159560 -297230
rect 161120 -297290 161140 -297230
rect 159540 -297300 161140 -297290
rect 162540 -297200 162560 -297130
rect 164120 -297200 164140 -297130
rect 162540 -297230 164140 -297200
rect 162540 -297290 162560 -297230
rect 164120 -297290 164140 -297230
rect 162540 -297300 164140 -297290
rect 165540 -297200 165560 -297130
rect 167120 -297200 167140 -297130
rect 165540 -297230 167140 -297200
rect 165540 -297290 165560 -297230
rect 167120 -297290 167140 -297230
rect 165540 -297300 167140 -297290
rect 168540 -297200 168560 -297130
rect 170120 -297200 170140 -297130
rect 168540 -297230 170140 -297200
rect 168540 -297290 168560 -297230
rect 170120 -297290 170140 -297230
rect 168540 -297300 170140 -297290
rect 171540 -297200 171560 -297130
rect 173120 -297200 173140 -297130
rect 171540 -297230 173140 -297200
rect 171540 -297290 171560 -297230
rect 173120 -297290 173140 -297230
rect 171540 -297300 173140 -297290
rect 174540 -297200 174560 -297130
rect 176120 -297200 176140 -297130
rect 174540 -297230 176140 -297200
rect 174540 -297290 174560 -297230
rect 176120 -297290 176140 -297230
rect 174540 -297300 176140 -297290
rect 177540 -297200 177560 -297130
rect 179120 -297200 179140 -297130
rect 177540 -297230 179140 -297200
rect 177540 -297290 177560 -297230
rect 179120 -297290 179140 -297230
rect 177540 -297300 179140 -297290
rect 180540 -297200 180560 -297130
rect 182120 -297200 182140 -297130
rect 180540 -297230 182140 -297200
rect 180540 -297290 180560 -297230
rect 182120 -297290 182140 -297230
rect 180540 -297300 182140 -297290
rect 183540 -297200 183560 -297130
rect 185120 -297200 185140 -297130
rect 183540 -297230 185140 -297200
rect 183540 -297290 183560 -297230
rect 185120 -297290 185140 -297230
rect 183540 -297300 185140 -297290
rect 186540 -297200 186560 -297130
rect 188120 -297200 188140 -297130
rect 186540 -297230 188140 -297200
rect 186540 -297290 186560 -297230
rect 188120 -297290 188140 -297230
rect 186540 -297300 188140 -297290
rect 189540 -297200 189560 -297130
rect 191120 -297200 191140 -297130
rect 189540 -297230 191140 -297200
rect 189540 -297290 189560 -297230
rect 191120 -297290 191140 -297230
rect 189540 -297300 191140 -297290
rect 192540 -297200 192560 -297130
rect 194120 -297200 194140 -297130
rect 192540 -297230 194140 -297200
rect 192540 -297290 192560 -297230
rect 194120 -297290 194140 -297230
rect 192540 -297300 194140 -297290
rect 195540 -297200 195560 -297130
rect 197120 -297200 197140 -297130
rect 195540 -297230 197140 -297200
rect 195540 -297290 195560 -297230
rect 197120 -297290 197140 -297230
rect 195540 -297300 197140 -297290
rect 198540 -297200 198560 -297130
rect 200120 -297200 200140 -297130
rect 198540 -297230 200140 -297200
rect 198540 -297290 198560 -297230
rect 200120 -297290 200140 -297230
rect 198540 -297300 200140 -297290
rect 201540 -297200 201560 -297130
rect 203120 -297200 203140 -297130
rect 201540 -297230 203140 -297200
rect 201540 -297290 201560 -297230
rect 203120 -297290 203140 -297230
rect 201540 -297300 203140 -297290
rect 204540 -297200 204560 -297130
rect 206120 -297200 206140 -297130
rect 204540 -297230 206140 -297200
rect 204540 -297290 204560 -297230
rect 206120 -297290 206140 -297230
rect 204540 -297300 206140 -297290
rect 207540 -297200 207560 -297130
rect 209120 -297200 209140 -297130
rect 207540 -297230 209140 -297200
rect 207540 -297290 207560 -297230
rect 209120 -297290 209140 -297230
rect 207540 -297300 209140 -297290
rect 210540 -297200 210560 -297130
rect 212120 -297200 212140 -297130
rect 210540 -297230 212140 -297200
rect 210540 -297290 210560 -297230
rect 212120 -297290 212140 -297230
rect 210540 -297300 212140 -297290
rect 213540 -297200 213560 -297130
rect 215120 -297200 215140 -297130
rect 213540 -297230 215140 -297200
rect 213540 -297290 213560 -297230
rect 215120 -297290 215140 -297230
rect 213540 -297300 215140 -297290
rect 216540 -297200 216560 -297130
rect 218120 -297200 218140 -297130
rect 216540 -297230 218140 -297200
rect 216540 -297290 216560 -297230
rect 218120 -297290 218140 -297230
rect 216540 -297300 218140 -297290
rect 219540 -297200 219560 -297130
rect 221120 -297200 221140 -297130
rect 219540 -297230 221140 -297200
rect 219540 -297290 219560 -297230
rect 221120 -297290 221140 -297230
rect 219540 -297300 221140 -297290
rect 222540 -297200 222560 -297130
rect 224120 -297200 224140 -297130
rect 222540 -297230 224140 -297200
rect 222540 -297290 222560 -297230
rect 224120 -297290 224140 -297230
rect 222540 -297300 224140 -297290
rect 225540 -297200 225560 -297130
rect 227120 -297200 227140 -297130
rect 225540 -297230 227140 -297200
rect 225540 -297290 225560 -297230
rect 227120 -297290 227140 -297230
rect 225540 -297300 227140 -297290
rect 228540 -297200 228560 -297130
rect 230120 -297200 230140 -297130
rect 228540 -297230 230140 -297200
rect 228540 -297290 228560 -297230
rect 230120 -297290 230140 -297230
rect 228540 -297300 230140 -297290
rect 231540 -297200 231560 -297130
rect 233120 -297200 233140 -297130
rect 231540 -297230 233140 -297200
rect 231540 -297290 231560 -297230
rect 233120 -297290 233140 -297230
rect 231540 -297300 233140 -297290
rect 234540 -297200 234560 -297130
rect 236120 -297200 236140 -297130
rect 234540 -297230 236140 -297200
rect 234540 -297290 234560 -297230
rect 236120 -297290 236140 -297230
rect 234540 -297300 236140 -297290
rect 237540 -297200 237560 -297130
rect 239120 -297200 239140 -297130
rect 237540 -297230 239140 -297200
rect 237540 -297290 237560 -297230
rect 239120 -297290 239140 -297230
rect 237540 -297300 239140 -297290
rect 240540 -297200 240560 -297130
rect 242120 -297200 242140 -297130
rect 240540 -297230 242140 -297200
rect 240540 -297290 240560 -297230
rect 242120 -297290 242140 -297230
rect 240540 -297300 242140 -297290
rect 243540 -297200 243560 -297130
rect 245120 -297200 245140 -297130
rect 243540 -297230 245140 -297200
rect 243540 -297290 243560 -297230
rect 245120 -297290 245140 -297230
rect 243540 -297300 245140 -297290
rect 246540 -297200 246560 -297130
rect 248120 -297200 248140 -297130
rect 246540 -297230 248140 -297200
rect 246540 -297290 246560 -297230
rect 248120 -297290 248140 -297230
rect 246540 -297300 248140 -297290
rect 249540 -297200 249560 -297130
rect 251120 -297200 251140 -297130
rect 249540 -297230 251140 -297200
rect 249540 -297290 249560 -297230
rect 251120 -297290 251140 -297230
rect 249540 -297300 251140 -297290
rect 252540 -297200 252560 -297130
rect 254120 -297200 254140 -297130
rect 252540 -297230 254140 -297200
rect 252540 -297290 252560 -297230
rect 254120 -297290 254140 -297230
rect 252540 -297300 254140 -297290
rect 255540 -297200 255560 -297130
rect 257120 -297200 257140 -297130
rect 255540 -297230 257140 -297200
rect 255540 -297290 255560 -297230
rect 257120 -297290 257140 -297230
rect 255540 -297300 257140 -297290
rect 258540 -297200 258560 -297130
rect 260120 -297200 260140 -297130
rect 258540 -297230 260140 -297200
rect 258540 -297290 258560 -297230
rect 260120 -297290 260140 -297230
rect 258540 -297300 260140 -297290
rect 261540 -297200 261560 -297130
rect 263120 -297200 263140 -297130
rect 261540 -297230 263140 -297200
rect 261540 -297290 261560 -297230
rect 263120 -297290 263140 -297230
rect 261540 -297300 263140 -297290
rect 264540 -297200 264560 -297130
rect 266120 -297200 266140 -297130
rect 264540 -297230 266140 -297200
rect 264540 -297290 264560 -297230
rect 266120 -297290 266140 -297230
rect 264540 -297300 266140 -297290
rect 267540 -297200 267560 -297130
rect 269120 -297200 269140 -297130
rect 267540 -297230 269140 -297200
rect 267540 -297290 267560 -297230
rect 269120 -297290 269140 -297230
rect 267540 -297300 269140 -297290
rect 270540 -297200 270560 -297130
rect 272120 -297200 272140 -297130
rect 270540 -297230 272140 -297200
rect 270540 -297290 270560 -297230
rect 272120 -297290 272140 -297230
rect 270540 -297300 272140 -297290
rect 273540 -297200 273560 -297130
rect 275120 -297200 275140 -297130
rect 273540 -297230 275140 -297200
rect 273540 -297290 273560 -297230
rect 275120 -297290 275140 -297230
rect 273540 -297300 275140 -297290
rect 276540 -297200 276560 -297130
rect 278120 -297200 278140 -297130
rect 276540 -297230 278140 -297200
rect 276540 -297290 276560 -297230
rect 278120 -297290 278140 -297230
rect 276540 -297300 278140 -297290
rect 279540 -297200 279560 -297130
rect 281120 -297200 281140 -297130
rect 279540 -297230 281140 -297200
rect 279540 -297290 279560 -297230
rect 281120 -297290 281140 -297230
rect 279540 -297300 281140 -297290
rect 282540 -297200 282560 -297130
rect 284120 -297200 284140 -297130
rect 282540 -297230 284140 -297200
rect 282540 -297290 282560 -297230
rect 284120 -297290 284140 -297230
rect 282540 -297300 284140 -297290
rect 285540 -297200 285560 -297130
rect 287120 -297200 287140 -297130
rect 285540 -297230 287140 -297200
rect 285540 -297290 285560 -297230
rect 287120 -297290 287140 -297230
rect 285540 -297300 287140 -297290
rect 288540 -297200 288560 -297130
rect 290120 -297200 290140 -297130
rect 288540 -297230 290140 -297200
rect 288540 -297290 288560 -297230
rect 290120 -297290 290140 -297230
rect 288540 -297300 290140 -297290
rect 291540 -297200 291560 -297130
rect 293120 -297200 293140 -297130
rect 291540 -297230 293140 -297200
rect 291540 -297290 291560 -297230
rect 293120 -297290 293140 -297230
rect 291540 -297300 293140 -297290
rect 294540 -297200 294560 -297130
rect 296120 -297200 296140 -297130
rect 294540 -297230 296140 -297200
rect 294540 -297290 294560 -297230
rect 296120 -297290 296140 -297230
rect 294540 -297300 296140 -297290
rect 297540 -297200 297560 -297130
rect 299120 -297200 299140 -297130
rect 297540 -297230 299140 -297200
rect 297540 -297290 297560 -297230
rect 299120 -297290 299140 -297230
rect 297540 -297300 299140 -297290
rect 220 -297500 440 -297490
rect 220 -297700 240 -297500
rect 420 -297700 440 -297500
rect 220 -297710 440 -297700
rect 3220 -297500 3440 -297490
rect 3220 -297700 3240 -297500
rect 3420 -297700 3440 -297500
rect 3220 -297710 3440 -297700
rect 6220 -297500 6440 -297490
rect 6220 -297700 6240 -297500
rect 6420 -297700 6440 -297500
rect 6220 -297710 6440 -297700
rect 9220 -297500 9440 -297490
rect 9220 -297700 9240 -297500
rect 9420 -297700 9440 -297500
rect 9220 -297710 9440 -297700
rect 12220 -297500 12440 -297490
rect 12220 -297700 12240 -297500
rect 12420 -297700 12440 -297500
rect 12220 -297710 12440 -297700
rect 15220 -297500 15440 -297490
rect 15220 -297700 15240 -297500
rect 15420 -297700 15440 -297500
rect 15220 -297710 15440 -297700
rect 18220 -297500 18440 -297490
rect 18220 -297700 18240 -297500
rect 18420 -297700 18440 -297500
rect 18220 -297710 18440 -297700
rect 21220 -297500 21440 -297490
rect 21220 -297700 21240 -297500
rect 21420 -297700 21440 -297500
rect 21220 -297710 21440 -297700
rect 24220 -297500 24440 -297490
rect 24220 -297700 24240 -297500
rect 24420 -297700 24440 -297500
rect 24220 -297710 24440 -297700
rect 27220 -297500 27440 -297490
rect 27220 -297700 27240 -297500
rect 27420 -297700 27440 -297500
rect 27220 -297710 27440 -297700
rect 30220 -297500 30440 -297490
rect 30220 -297700 30240 -297500
rect 30420 -297700 30440 -297500
rect 30220 -297710 30440 -297700
rect 33220 -297500 33440 -297490
rect 33220 -297700 33240 -297500
rect 33420 -297700 33440 -297500
rect 33220 -297710 33440 -297700
rect 36220 -297500 36440 -297490
rect 36220 -297700 36240 -297500
rect 36420 -297700 36440 -297500
rect 36220 -297710 36440 -297700
rect 39220 -297500 39440 -297490
rect 39220 -297700 39240 -297500
rect 39420 -297700 39440 -297500
rect 39220 -297710 39440 -297700
rect 42220 -297500 42440 -297490
rect 42220 -297700 42240 -297500
rect 42420 -297700 42440 -297500
rect 42220 -297710 42440 -297700
rect 45220 -297500 45440 -297490
rect 45220 -297700 45240 -297500
rect 45420 -297700 45440 -297500
rect 45220 -297710 45440 -297700
rect 48220 -297500 48440 -297490
rect 48220 -297700 48240 -297500
rect 48420 -297700 48440 -297500
rect 48220 -297710 48440 -297700
rect 51220 -297500 51440 -297490
rect 51220 -297700 51240 -297500
rect 51420 -297700 51440 -297500
rect 51220 -297710 51440 -297700
rect 54220 -297500 54440 -297490
rect 54220 -297700 54240 -297500
rect 54420 -297700 54440 -297500
rect 54220 -297710 54440 -297700
rect 57220 -297500 57440 -297490
rect 57220 -297700 57240 -297500
rect 57420 -297700 57440 -297500
rect 57220 -297710 57440 -297700
rect 60220 -297500 60440 -297490
rect 60220 -297700 60240 -297500
rect 60420 -297700 60440 -297500
rect 60220 -297710 60440 -297700
rect 63220 -297500 63440 -297490
rect 63220 -297700 63240 -297500
rect 63420 -297700 63440 -297500
rect 63220 -297710 63440 -297700
rect 66220 -297500 66440 -297490
rect 66220 -297700 66240 -297500
rect 66420 -297700 66440 -297500
rect 66220 -297710 66440 -297700
rect 69220 -297500 69440 -297490
rect 69220 -297700 69240 -297500
rect 69420 -297700 69440 -297500
rect 69220 -297710 69440 -297700
rect 72220 -297500 72440 -297490
rect 72220 -297700 72240 -297500
rect 72420 -297700 72440 -297500
rect 72220 -297710 72440 -297700
rect 75220 -297500 75440 -297490
rect 75220 -297700 75240 -297500
rect 75420 -297700 75440 -297500
rect 75220 -297710 75440 -297700
rect 78220 -297500 78440 -297490
rect 78220 -297700 78240 -297500
rect 78420 -297700 78440 -297500
rect 78220 -297710 78440 -297700
rect 81220 -297500 81440 -297490
rect 81220 -297700 81240 -297500
rect 81420 -297700 81440 -297500
rect 81220 -297710 81440 -297700
rect 84220 -297500 84440 -297490
rect 84220 -297700 84240 -297500
rect 84420 -297700 84440 -297500
rect 84220 -297710 84440 -297700
rect 87220 -297500 87440 -297490
rect 87220 -297700 87240 -297500
rect 87420 -297700 87440 -297500
rect 87220 -297710 87440 -297700
rect 90220 -297500 90440 -297490
rect 90220 -297700 90240 -297500
rect 90420 -297700 90440 -297500
rect 90220 -297710 90440 -297700
rect 93220 -297500 93440 -297490
rect 93220 -297700 93240 -297500
rect 93420 -297700 93440 -297500
rect 93220 -297710 93440 -297700
rect 96220 -297500 96440 -297490
rect 96220 -297700 96240 -297500
rect 96420 -297700 96440 -297500
rect 96220 -297710 96440 -297700
rect 99220 -297500 99440 -297490
rect 99220 -297700 99240 -297500
rect 99420 -297700 99440 -297500
rect 99220 -297710 99440 -297700
rect 102220 -297500 102440 -297490
rect 102220 -297700 102240 -297500
rect 102420 -297700 102440 -297500
rect 102220 -297710 102440 -297700
rect 105220 -297500 105440 -297490
rect 105220 -297700 105240 -297500
rect 105420 -297700 105440 -297500
rect 105220 -297710 105440 -297700
rect 108220 -297500 108440 -297490
rect 108220 -297700 108240 -297500
rect 108420 -297700 108440 -297500
rect 108220 -297710 108440 -297700
rect 111220 -297500 111440 -297490
rect 111220 -297700 111240 -297500
rect 111420 -297700 111440 -297500
rect 111220 -297710 111440 -297700
rect 114220 -297500 114440 -297490
rect 114220 -297700 114240 -297500
rect 114420 -297700 114440 -297500
rect 114220 -297710 114440 -297700
rect 117220 -297500 117440 -297490
rect 117220 -297700 117240 -297500
rect 117420 -297700 117440 -297500
rect 117220 -297710 117440 -297700
rect 120220 -297500 120440 -297490
rect 120220 -297700 120240 -297500
rect 120420 -297700 120440 -297500
rect 120220 -297710 120440 -297700
rect 123220 -297500 123440 -297490
rect 123220 -297700 123240 -297500
rect 123420 -297700 123440 -297500
rect 123220 -297710 123440 -297700
rect 126220 -297500 126440 -297490
rect 126220 -297700 126240 -297500
rect 126420 -297700 126440 -297500
rect 126220 -297710 126440 -297700
rect 129220 -297500 129440 -297490
rect 129220 -297700 129240 -297500
rect 129420 -297700 129440 -297500
rect 129220 -297710 129440 -297700
rect 132220 -297500 132440 -297490
rect 132220 -297700 132240 -297500
rect 132420 -297700 132440 -297500
rect 132220 -297710 132440 -297700
rect 135220 -297500 135440 -297490
rect 135220 -297700 135240 -297500
rect 135420 -297700 135440 -297500
rect 135220 -297710 135440 -297700
rect 138220 -297500 138440 -297490
rect 138220 -297700 138240 -297500
rect 138420 -297700 138440 -297500
rect 138220 -297710 138440 -297700
rect 141220 -297500 141440 -297490
rect 141220 -297700 141240 -297500
rect 141420 -297700 141440 -297500
rect 141220 -297710 141440 -297700
rect 144220 -297500 144440 -297490
rect 144220 -297700 144240 -297500
rect 144420 -297700 144440 -297500
rect 144220 -297710 144440 -297700
rect 147220 -297500 147440 -297490
rect 147220 -297700 147240 -297500
rect 147420 -297700 147440 -297500
rect 147220 -297710 147440 -297700
rect 150220 -297500 150440 -297490
rect 150220 -297700 150240 -297500
rect 150420 -297700 150440 -297500
rect 150220 -297710 150440 -297700
rect 153220 -297500 153440 -297490
rect 153220 -297700 153240 -297500
rect 153420 -297700 153440 -297500
rect 153220 -297710 153440 -297700
rect 156220 -297500 156440 -297490
rect 156220 -297700 156240 -297500
rect 156420 -297700 156440 -297500
rect 156220 -297710 156440 -297700
rect 159220 -297500 159440 -297490
rect 159220 -297700 159240 -297500
rect 159420 -297700 159440 -297500
rect 159220 -297710 159440 -297700
rect 162220 -297500 162440 -297490
rect 162220 -297700 162240 -297500
rect 162420 -297700 162440 -297500
rect 162220 -297710 162440 -297700
rect 165220 -297500 165440 -297490
rect 165220 -297700 165240 -297500
rect 165420 -297700 165440 -297500
rect 165220 -297710 165440 -297700
rect 168220 -297500 168440 -297490
rect 168220 -297700 168240 -297500
rect 168420 -297700 168440 -297500
rect 168220 -297710 168440 -297700
rect 171220 -297500 171440 -297490
rect 171220 -297700 171240 -297500
rect 171420 -297700 171440 -297500
rect 171220 -297710 171440 -297700
rect 174220 -297500 174440 -297490
rect 174220 -297700 174240 -297500
rect 174420 -297700 174440 -297500
rect 174220 -297710 174440 -297700
rect 177220 -297500 177440 -297490
rect 177220 -297700 177240 -297500
rect 177420 -297700 177440 -297500
rect 177220 -297710 177440 -297700
rect 180220 -297500 180440 -297490
rect 180220 -297700 180240 -297500
rect 180420 -297700 180440 -297500
rect 180220 -297710 180440 -297700
rect 183220 -297500 183440 -297490
rect 183220 -297700 183240 -297500
rect 183420 -297700 183440 -297500
rect 183220 -297710 183440 -297700
rect 186220 -297500 186440 -297490
rect 186220 -297700 186240 -297500
rect 186420 -297700 186440 -297500
rect 186220 -297710 186440 -297700
rect 189220 -297500 189440 -297490
rect 189220 -297700 189240 -297500
rect 189420 -297700 189440 -297500
rect 189220 -297710 189440 -297700
rect 192220 -297500 192440 -297490
rect 192220 -297700 192240 -297500
rect 192420 -297700 192440 -297500
rect 192220 -297710 192440 -297700
rect 195220 -297500 195440 -297490
rect 195220 -297700 195240 -297500
rect 195420 -297700 195440 -297500
rect 195220 -297710 195440 -297700
rect 198220 -297500 198440 -297490
rect 198220 -297700 198240 -297500
rect 198420 -297700 198440 -297500
rect 198220 -297710 198440 -297700
rect 201220 -297500 201440 -297490
rect 201220 -297700 201240 -297500
rect 201420 -297700 201440 -297500
rect 201220 -297710 201440 -297700
rect 204220 -297500 204440 -297490
rect 204220 -297700 204240 -297500
rect 204420 -297700 204440 -297500
rect 204220 -297710 204440 -297700
rect 207220 -297500 207440 -297490
rect 207220 -297700 207240 -297500
rect 207420 -297700 207440 -297500
rect 207220 -297710 207440 -297700
rect 210220 -297500 210440 -297490
rect 210220 -297700 210240 -297500
rect 210420 -297700 210440 -297500
rect 210220 -297710 210440 -297700
rect 213220 -297500 213440 -297490
rect 213220 -297700 213240 -297500
rect 213420 -297700 213440 -297500
rect 213220 -297710 213440 -297700
rect 216220 -297500 216440 -297490
rect 216220 -297700 216240 -297500
rect 216420 -297700 216440 -297500
rect 216220 -297710 216440 -297700
rect 219220 -297500 219440 -297490
rect 219220 -297700 219240 -297500
rect 219420 -297700 219440 -297500
rect 219220 -297710 219440 -297700
rect 222220 -297500 222440 -297490
rect 222220 -297700 222240 -297500
rect 222420 -297700 222440 -297500
rect 222220 -297710 222440 -297700
rect 225220 -297500 225440 -297490
rect 225220 -297700 225240 -297500
rect 225420 -297700 225440 -297500
rect 225220 -297710 225440 -297700
rect 228220 -297500 228440 -297490
rect 228220 -297700 228240 -297500
rect 228420 -297700 228440 -297500
rect 228220 -297710 228440 -297700
rect 231220 -297500 231440 -297490
rect 231220 -297700 231240 -297500
rect 231420 -297700 231440 -297500
rect 231220 -297710 231440 -297700
rect 234220 -297500 234440 -297490
rect 234220 -297700 234240 -297500
rect 234420 -297700 234440 -297500
rect 234220 -297710 234440 -297700
rect 237220 -297500 237440 -297490
rect 237220 -297700 237240 -297500
rect 237420 -297700 237440 -297500
rect 237220 -297710 237440 -297700
rect 240220 -297500 240440 -297490
rect 240220 -297700 240240 -297500
rect 240420 -297700 240440 -297500
rect 240220 -297710 240440 -297700
rect 243220 -297500 243440 -297490
rect 243220 -297700 243240 -297500
rect 243420 -297700 243440 -297500
rect 243220 -297710 243440 -297700
rect 246220 -297500 246440 -297490
rect 246220 -297700 246240 -297500
rect 246420 -297700 246440 -297500
rect 246220 -297710 246440 -297700
rect 249220 -297500 249440 -297490
rect 249220 -297700 249240 -297500
rect 249420 -297700 249440 -297500
rect 249220 -297710 249440 -297700
rect 252220 -297500 252440 -297490
rect 252220 -297700 252240 -297500
rect 252420 -297700 252440 -297500
rect 252220 -297710 252440 -297700
rect 255220 -297500 255440 -297490
rect 255220 -297700 255240 -297500
rect 255420 -297700 255440 -297500
rect 255220 -297710 255440 -297700
rect 258220 -297500 258440 -297490
rect 258220 -297700 258240 -297500
rect 258420 -297700 258440 -297500
rect 258220 -297710 258440 -297700
rect 261220 -297500 261440 -297490
rect 261220 -297700 261240 -297500
rect 261420 -297700 261440 -297500
rect 261220 -297710 261440 -297700
rect 264220 -297500 264440 -297490
rect 264220 -297700 264240 -297500
rect 264420 -297700 264440 -297500
rect 264220 -297710 264440 -297700
rect 267220 -297500 267440 -297490
rect 267220 -297700 267240 -297500
rect 267420 -297700 267440 -297500
rect 267220 -297710 267440 -297700
rect 270220 -297500 270440 -297490
rect 270220 -297700 270240 -297500
rect 270420 -297700 270440 -297500
rect 270220 -297710 270440 -297700
rect 273220 -297500 273440 -297490
rect 273220 -297700 273240 -297500
rect 273420 -297700 273440 -297500
rect 273220 -297710 273440 -297700
rect 276220 -297500 276440 -297490
rect 276220 -297700 276240 -297500
rect 276420 -297700 276440 -297500
rect 276220 -297710 276440 -297700
rect 279220 -297500 279440 -297490
rect 279220 -297700 279240 -297500
rect 279420 -297700 279440 -297500
rect 279220 -297710 279440 -297700
rect 282220 -297500 282440 -297490
rect 282220 -297700 282240 -297500
rect 282420 -297700 282440 -297500
rect 282220 -297710 282440 -297700
rect 285220 -297500 285440 -297490
rect 285220 -297700 285240 -297500
rect 285420 -297700 285440 -297500
rect 285220 -297710 285440 -297700
rect 288220 -297500 288440 -297490
rect 288220 -297700 288240 -297500
rect 288420 -297700 288440 -297500
rect 288220 -297710 288440 -297700
rect 291220 -297500 291440 -297490
rect 291220 -297700 291240 -297500
rect 291420 -297700 291440 -297500
rect 291220 -297710 291440 -297700
rect 294220 -297500 294440 -297490
rect 294220 -297700 294240 -297500
rect 294420 -297700 294440 -297500
rect 294220 -297710 294440 -297700
rect 297220 -297500 297440 -297490
rect 297220 -297700 297240 -297500
rect 297420 -297700 297440 -297500
rect 297220 -297710 297440 -297700
rect 540 -297920 300740 -297900
rect 540 -298080 560 -297920
rect 540 -298100 300740 -298080
<< via1 >>
rect -1920 3360 -900 3450
rect 50 3360 140 3450
rect 3050 3360 3140 3450
rect 6050 3360 6140 3450
rect 9050 3360 9140 3450
rect 12050 3360 12140 3450
rect 15050 3360 15140 3450
rect 18050 3360 18140 3450
rect 21050 3360 21140 3450
rect 24050 3360 24140 3450
rect 27050 3360 27140 3450
rect 30050 3360 30140 3450
rect 33050 3360 33140 3450
rect 36050 3360 36140 3450
rect 39050 3360 39140 3450
rect 42050 3360 42140 3450
rect 45050 3360 45140 3450
rect 48050 3360 48140 3450
rect 51050 3360 51140 3450
rect 54050 3360 54140 3450
rect 57050 3360 57140 3450
rect 60050 3360 60140 3450
rect 63050 3360 63140 3450
rect 66050 3360 66140 3450
rect 69050 3360 69140 3450
rect 72050 3360 72140 3450
rect 75050 3360 75140 3450
rect 78050 3360 78140 3450
rect 81050 3360 81140 3450
rect 84050 3360 84140 3450
rect 87050 3360 87140 3450
rect 90050 3360 90140 3450
rect 93050 3360 93140 3450
rect 96050 3360 96140 3450
rect 99050 3360 99140 3450
rect 102050 3360 102140 3450
rect 105050 3360 105140 3450
rect 108050 3360 108140 3450
rect 111050 3360 111140 3450
rect 114050 3360 114140 3450
rect 117050 3360 117140 3450
rect 120050 3360 120140 3450
rect 123050 3360 123140 3450
rect 126050 3360 126140 3450
rect 129050 3360 129140 3450
rect 132050 3360 132140 3450
rect 135050 3360 135140 3450
rect 138050 3360 138140 3450
rect 141050 3360 141140 3450
rect 144050 3360 144140 3450
rect 147050 3360 147140 3450
rect 150050 3360 150140 3450
rect 153050 3360 153140 3450
rect 156050 3360 156140 3450
rect 159050 3360 159140 3450
rect 162050 3360 162140 3450
rect 165050 3360 165140 3450
rect 168050 3360 168140 3450
rect 171050 3360 171140 3450
rect 174050 3360 174140 3450
rect 177050 3360 177140 3450
rect 180050 3360 180140 3450
rect 183050 3360 183140 3450
rect 186050 3360 186140 3450
rect 189050 3360 189140 3450
rect 192050 3360 192140 3450
rect 195050 3360 195140 3450
rect 198050 3360 198140 3450
rect 201050 3360 201140 3450
rect 204050 3360 204140 3450
rect 207050 3360 207140 3450
rect 210050 3360 210140 3450
rect 213050 3360 213140 3450
rect 216050 3360 216140 3450
rect 219050 3360 219140 3450
rect 222050 3360 222140 3450
rect 225050 3360 225140 3450
rect 228050 3360 228140 3450
rect 231050 3360 231140 3450
rect 234050 3360 234140 3450
rect 237050 3360 237140 3450
rect 240050 3360 240140 3450
rect 243050 3360 243140 3450
rect 246050 3360 246140 3450
rect 249050 3360 249140 3450
rect 252050 3360 252140 3450
rect 255050 3360 255140 3450
rect 258050 3360 258140 3450
rect 261050 3360 261140 3450
rect 264050 3360 264140 3450
rect 267050 3360 267140 3450
rect 270050 3360 270140 3450
rect 273050 3360 273140 3450
rect 276050 3360 276140 3450
rect 279050 3360 279140 3450
rect 282050 3360 282140 3450
rect 285050 3360 285140 3450
rect 288050 3360 288140 3450
rect 291050 3360 291140 3450
rect 294050 3360 294140 3450
rect 297050 3360 297140 3450
rect -1580 1490 -1180 1560
rect -540 1490 -260 1560
rect -1580 -1510 -1180 -1440
rect -540 -1510 -260 -1440
rect -1580 -4510 -1180 -4440
rect -540 -4510 -260 -4440
rect -1580 -7510 -1180 -7440
rect -540 -7510 -260 -7440
rect -1580 -10510 -1180 -10440
rect -540 -10510 -260 -10440
rect -1580 -13510 -1180 -13440
rect -540 -13510 -260 -13440
rect -1580 -16510 -1180 -16440
rect -540 -16510 -260 -16440
rect -1580 -19510 -1180 -19440
rect -540 -19510 -260 -19440
rect -1580 -22510 -1180 -22440
rect -540 -22510 -260 -22440
rect -1580 -25510 -1180 -25440
rect -540 -25510 -260 -25440
rect -1580 -28510 -1180 -28440
rect -540 -28510 -260 -28440
rect -1580 -31510 -1180 -31440
rect -540 -31510 -260 -31440
rect -1580 -34510 -1180 -34440
rect -540 -34510 -260 -34440
rect -1580 -37510 -1180 -37440
rect -540 -37510 -260 -37440
rect -1580 -40510 -1180 -40440
rect -540 -40510 -260 -40440
rect -1580 -43510 -1180 -43440
rect -540 -43510 -260 -43440
rect -1580 -46510 -1180 -46440
rect -540 -46510 -260 -46440
rect -1580 -49510 -1180 -49440
rect -540 -49510 -260 -49440
rect -1580 -52510 -1180 -52440
rect -540 -52510 -260 -52440
rect -1580 -55510 -1180 -55440
rect -540 -55510 -260 -55440
rect -1580 -58510 -1180 -58440
rect -540 -58510 -260 -58440
rect -1580 -61510 -1180 -61440
rect -540 -61510 -260 -61440
rect -1580 -64510 -1180 -64440
rect -540 -64510 -260 -64440
rect -1580 -67510 -1180 -67440
rect -540 -67510 -260 -67440
rect -1580 -70510 -1180 -70440
rect -540 -70510 -260 -70440
rect -1580 -73510 -1180 -73440
rect -540 -73510 -260 -73440
rect -1580 -76510 -1180 -76440
rect -540 -76510 -260 -76440
rect -1580 -79510 -1180 -79440
rect -540 -79510 -260 -79440
rect -1580 -82510 -1180 -82440
rect -540 -82510 -260 -82440
rect -1580 -85510 -1180 -85440
rect -540 -85510 -260 -85440
rect -1580 -88510 -1180 -88440
rect -540 -88510 -260 -88440
rect -1580 -91510 -1180 -91440
rect -540 -91510 -260 -91440
rect -1580 -94510 -1180 -94440
rect -540 -94510 -260 -94440
rect -1580 -97510 -1180 -97440
rect -540 -97510 -260 -97440
rect -1580 -100510 -1180 -100440
rect -540 -100510 -260 -100440
rect -1580 -103510 -1180 -103440
rect -540 -103510 -260 -103440
rect -1580 -106510 -1180 -106440
rect -540 -106510 -260 -106440
rect -1580 -109510 -1180 -109440
rect -540 -109510 -260 -109440
rect -1580 -112510 -1180 -112440
rect -540 -112510 -260 -112440
rect -1580 -115510 -1180 -115440
rect -540 -115510 -260 -115440
rect -1580 -118510 -1180 -118440
rect -540 -118510 -260 -118440
rect -1580 -121510 -1180 -121440
rect -540 -121510 -260 -121440
rect -1580 -124510 -1180 -124440
rect -540 -124510 -260 -124440
rect -1580 -127510 -1180 -127440
rect -540 -127510 -260 -127440
rect -1580 -130510 -1180 -130440
rect -540 -130510 -260 -130440
rect -1580 -133510 -1180 -133440
rect -540 -133510 -260 -133440
rect -1580 -136510 -1180 -136440
rect -540 -136510 -260 -136440
rect -1580 -139510 -1180 -139440
rect -540 -139510 -260 -139440
rect -1580 -142510 -1180 -142440
rect -540 -142510 -260 -142440
rect -1580 -145510 -1180 -145440
rect -540 -145510 -260 -145440
rect -1580 -148510 -1180 -148440
rect -540 -148510 -260 -148440
rect -1580 -151510 -1180 -151440
rect -540 -151510 -260 -151440
rect -1580 -154510 -1180 -154440
rect -540 -154510 -260 -154440
rect -1580 -157510 -1180 -157440
rect -540 -157510 -260 -157440
rect -1580 -160510 -1180 -160440
rect -540 -160510 -260 -160440
rect -1580 -163510 -1180 -163440
rect -540 -163510 -260 -163440
rect -1580 -166510 -1180 -166440
rect -540 -166510 -260 -166440
rect -1580 -169510 -1180 -169440
rect -540 -169510 -260 -169440
rect -1580 -172510 -1180 -172440
rect -540 -172510 -260 -172440
rect -1580 -175510 -1180 -175440
rect -540 -175510 -260 -175440
rect -1580 -178510 -1180 -178440
rect -540 -178510 -260 -178440
rect -1580 -181510 -1180 -181440
rect -540 -181510 -260 -181440
rect -1580 -184510 -1180 -184440
rect -540 -184510 -260 -184440
rect -1580 -187510 -1180 -187440
rect -540 -187510 -260 -187440
rect -1580 -190510 -1180 -190440
rect -540 -190510 -260 -190440
rect -1580 -193510 -1180 -193440
rect -540 -193510 -260 -193440
rect -1580 -196510 -1180 -196440
rect -540 -196510 -260 -196440
rect -1580 -199510 -1180 -199440
rect -540 -199510 -260 -199440
rect -1580 -202510 -1180 -202440
rect -540 -202510 -260 -202440
rect -1580 -205510 -1180 -205440
rect -540 -205510 -260 -205440
rect -1580 -208510 -1180 -208440
rect -540 -208510 -260 -208440
rect -1580 -211510 -1180 -211440
rect -540 -211510 -260 -211440
rect -1580 -214510 -1180 -214440
rect -540 -214510 -260 -214440
rect -1580 -217510 -1180 -217440
rect -540 -217510 -260 -217440
rect -1580 -220510 -1180 -220440
rect -540 -220510 -260 -220440
rect -1580 -223510 -1180 -223440
rect -540 -223510 -260 -223440
rect -1580 -226510 -1180 -226440
rect -540 -226510 -260 -226440
rect -1580 -229510 -1180 -229440
rect -540 -229510 -260 -229440
rect -1580 -232510 -1180 -232440
rect -540 -232510 -260 -232440
rect -1580 -235510 -1180 -235440
rect -540 -235510 -260 -235440
rect -1580 -238510 -1180 -238440
rect -540 -238510 -260 -238440
rect -1580 -241510 -1180 -241440
rect -540 -241510 -260 -241440
rect -1580 -244510 -1180 -244440
rect -540 -244510 -260 -244440
rect -1580 -247510 -1180 -247440
rect -540 -247510 -260 -247440
rect -1580 -250510 -1180 -250440
rect -540 -250510 -260 -250440
rect -1580 -253510 -1180 -253440
rect -540 -253510 -260 -253440
rect -1580 -256510 -1180 -256440
rect -540 -256510 -260 -256440
rect -1580 -259510 -1180 -259440
rect -540 -259510 -260 -259440
rect -1580 -262510 -1180 -262440
rect -540 -262510 -260 -262440
rect -1580 -265510 -1180 -265440
rect -540 -265510 -260 -265440
rect -1580 -268510 -1180 -268440
rect -540 -268510 -260 -268440
rect -1580 -271510 -1180 -271440
rect -540 -271510 -260 -271440
rect -1580 -274510 -1180 -274440
rect -540 -274510 -260 -274440
rect -1580 -277510 -1180 -277440
rect -540 -277510 -260 -277440
rect -1580 -280510 -1180 -280440
rect -540 -280510 -260 -280440
rect -1580 -283510 -1180 -283440
rect -540 -283510 -260 -283440
rect -1580 -286510 -1180 -286440
rect -540 -286510 -260 -286440
rect -1580 -289510 -1180 -289440
rect -540 -289510 -260 -289440
rect -1580 -292510 -1180 -292440
rect -540 -292510 -260 -292440
rect -1580 -295510 -1180 -295440
rect -540 -295510 -260 -295440
rect 560 -297200 2120 -297130
rect 3560 -297200 5120 -297130
rect 6560 -297200 8120 -297130
rect 9560 -297200 11120 -297130
rect 12560 -297200 14120 -297130
rect 15560 -297200 17120 -297130
rect 18560 -297200 20120 -297130
rect 21560 -297200 23120 -297130
rect 24560 -297200 26120 -297130
rect 27560 -297200 29120 -297130
rect 30560 -297200 32120 -297130
rect 33560 -297200 35120 -297130
rect 36560 -297200 38120 -297130
rect 39560 -297200 41120 -297130
rect 42560 -297200 44120 -297130
rect 45560 -297200 47120 -297130
rect 48560 -297200 50120 -297130
rect 51560 -297200 53120 -297130
rect 54560 -297200 56120 -297130
rect 57560 -297200 59120 -297130
rect 60560 -297200 62120 -297130
rect 63560 -297200 65120 -297130
rect 66560 -297200 68120 -297130
rect 69560 -297200 71120 -297130
rect 72560 -297200 74120 -297130
rect 75560 -297200 77120 -297130
rect 78560 -297200 80120 -297130
rect 81560 -297200 83120 -297130
rect 84560 -297200 86120 -297130
rect 87560 -297200 89120 -297130
rect 90560 -297200 92120 -297130
rect 93560 -297200 95120 -297130
rect 96560 -297200 98120 -297130
rect 99560 -297200 101120 -297130
rect 102560 -297200 104120 -297130
rect 105560 -297200 107120 -297130
rect 108560 -297200 110120 -297130
rect 111560 -297200 113120 -297130
rect 114560 -297200 116120 -297130
rect 117560 -297200 119120 -297130
rect 120560 -297200 122120 -297130
rect 123560 -297200 125120 -297130
rect 126560 -297200 128120 -297130
rect 129560 -297200 131120 -297130
rect 132560 -297200 134120 -297130
rect 135560 -297200 137120 -297130
rect 138560 -297200 140120 -297130
rect 141560 -297200 143120 -297130
rect 144560 -297200 146120 -297130
rect 147560 -297200 149120 -297130
rect 150560 -297200 152120 -297130
rect 153560 -297200 155120 -297130
rect 156560 -297200 158120 -297130
rect 159560 -297200 161120 -297130
rect 162560 -297200 164120 -297130
rect 165560 -297200 167120 -297130
rect 168560 -297200 170120 -297130
rect 171560 -297200 173120 -297130
rect 174560 -297200 176120 -297130
rect 177560 -297200 179120 -297130
rect 180560 -297200 182120 -297130
rect 183560 -297200 185120 -297130
rect 186560 -297200 188120 -297130
rect 189560 -297200 191120 -297130
rect 192560 -297200 194120 -297130
rect 195560 -297200 197120 -297130
rect 198560 -297200 200120 -297130
rect 201560 -297200 203120 -297130
rect 204560 -297200 206120 -297130
rect 207560 -297200 209120 -297130
rect 210560 -297200 212120 -297130
rect 213560 -297200 215120 -297130
rect 216560 -297200 218120 -297130
rect 219560 -297200 221120 -297130
rect 222560 -297200 224120 -297130
rect 225560 -297200 227120 -297130
rect 228560 -297200 230120 -297130
rect 231560 -297200 233120 -297130
rect 234560 -297200 236120 -297130
rect 237560 -297200 239120 -297130
rect 240560 -297200 242120 -297130
rect 243560 -297200 245120 -297130
rect 246560 -297200 248120 -297130
rect 249560 -297200 251120 -297130
rect 252560 -297200 254120 -297130
rect 255560 -297200 257120 -297130
rect 258560 -297200 260120 -297130
rect 261560 -297200 263120 -297130
rect 264560 -297200 266120 -297130
rect 267560 -297200 269120 -297130
rect 270560 -297200 272120 -297130
rect 273560 -297200 275120 -297130
rect 276560 -297200 278120 -297130
rect 279560 -297200 281120 -297130
rect 282560 -297200 284120 -297130
rect 285560 -297200 287120 -297130
rect 288560 -297200 290120 -297130
rect 291560 -297200 293120 -297130
rect 294560 -297200 296120 -297130
rect 297560 -297200 299120 -297130
rect 240 -297700 420 -297500
rect 3240 -297700 3420 -297500
rect 6240 -297700 6420 -297500
rect 9240 -297700 9420 -297500
rect 12240 -297700 12420 -297500
rect 15240 -297700 15420 -297500
rect 18240 -297700 18420 -297500
rect 21240 -297700 21420 -297500
rect 24240 -297700 24420 -297500
rect 27240 -297700 27420 -297500
rect 30240 -297700 30420 -297500
rect 33240 -297700 33420 -297500
rect 36240 -297700 36420 -297500
rect 39240 -297700 39420 -297500
rect 42240 -297700 42420 -297500
rect 45240 -297700 45420 -297500
rect 48240 -297700 48420 -297500
rect 51240 -297700 51420 -297500
rect 54240 -297700 54420 -297500
rect 57240 -297700 57420 -297500
rect 60240 -297700 60420 -297500
rect 63240 -297700 63420 -297500
rect 66240 -297700 66420 -297500
rect 69240 -297700 69420 -297500
rect 72240 -297700 72420 -297500
rect 75240 -297700 75420 -297500
rect 78240 -297700 78420 -297500
rect 81240 -297700 81420 -297500
rect 84240 -297700 84420 -297500
rect 87240 -297700 87420 -297500
rect 90240 -297700 90420 -297500
rect 93240 -297700 93420 -297500
rect 96240 -297700 96420 -297500
rect 99240 -297700 99420 -297500
rect 102240 -297700 102420 -297500
rect 105240 -297700 105420 -297500
rect 108240 -297700 108420 -297500
rect 111240 -297700 111420 -297500
rect 114240 -297700 114420 -297500
rect 117240 -297700 117420 -297500
rect 120240 -297700 120420 -297500
rect 123240 -297700 123420 -297500
rect 126240 -297700 126420 -297500
rect 129240 -297700 129420 -297500
rect 132240 -297700 132420 -297500
rect 135240 -297700 135420 -297500
rect 138240 -297700 138420 -297500
rect 141240 -297700 141420 -297500
rect 144240 -297700 144420 -297500
rect 147240 -297700 147420 -297500
rect 150240 -297700 150420 -297500
rect 153240 -297700 153420 -297500
rect 156240 -297700 156420 -297500
rect 159240 -297700 159420 -297500
rect 162240 -297700 162420 -297500
rect 165240 -297700 165420 -297500
rect 168240 -297700 168420 -297500
rect 171240 -297700 171420 -297500
rect 174240 -297700 174420 -297500
rect 177240 -297700 177420 -297500
rect 180240 -297700 180420 -297500
rect 183240 -297700 183420 -297500
rect 186240 -297700 186420 -297500
rect 189240 -297700 189420 -297500
rect 192240 -297700 192420 -297500
rect 195240 -297700 195420 -297500
rect 198240 -297700 198420 -297500
rect 201240 -297700 201420 -297500
rect 204240 -297700 204420 -297500
rect 207240 -297700 207420 -297500
rect 210240 -297700 210420 -297500
rect 213240 -297700 213420 -297500
rect 216240 -297700 216420 -297500
rect 219240 -297700 219420 -297500
rect 222240 -297700 222420 -297500
rect 225240 -297700 225420 -297500
rect 228240 -297700 228420 -297500
rect 231240 -297700 231420 -297500
rect 234240 -297700 234420 -297500
rect 237240 -297700 237420 -297500
rect 240240 -297700 240420 -297500
rect 243240 -297700 243420 -297500
rect 246240 -297700 246420 -297500
rect 249240 -297700 249420 -297500
rect 252240 -297700 252420 -297500
rect 255240 -297700 255420 -297500
rect 258240 -297700 258420 -297500
rect 261240 -297700 261420 -297500
rect 264240 -297700 264420 -297500
rect 267240 -297700 267420 -297500
rect 270240 -297700 270420 -297500
rect 273240 -297700 273420 -297500
rect 276240 -297700 276420 -297500
rect 279240 -297700 279420 -297500
rect 282240 -297700 282420 -297500
rect 285240 -297700 285420 -297500
rect 288240 -297700 288420 -297500
rect 291240 -297700 291420 -297500
rect 294240 -297700 294420 -297500
rect 297240 -297700 297420 -297500
rect 560 -297980 2120 -297920
rect 2120 -297980 3560 -297920
rect 3560 -297980 5120 -297920
rect 5120 -297980 6560 -297920
rect 6560 -297980 8120 -297920
rect 8120 -297980 9560 -297920
rect 9560 -297980 11120 -297920
rect 11120 -297980 12560 -297920
rect 12560 -297980 14120 -297920
rect 14120 -297980 15560 -297920
rect 15560 -297980 17120 -297920
rect 17120 -297980 18560 -297920
rect 18560 -297980 20120 -297920
rect 20120 -297980 21560 -297920
rect 21560 -297980 23120 -297920
rect 23120 -297980 24560 -297920
rect 24560 -297980 26120 -297920
rect 26120 -297980 27560 -297920
rect 27560 -297980 29120 -297920
rect 29120 -297980 30560 -297920
rect 30560 -297980 32120 -297920
rect 32120 -297980 33560 -297920
rect 33560 -297980 35120 -297920
rect 35120 -297980 36560 -297920
rect 36560 -297980 38120 -297920
rect 38120 -297980 39560 -297920
rect 39560 -297980 41120 -297920
rect 41120 -297980 42560 -297920
rect 42560 -297980 44120 -297920
rect 44120 -297980 45560 -297920
rect 45560 -297980 47120 -297920
rect 47120 -297980 48560 -297920
rect 48560 -297980 50120 -297920
rect 50120 -297980 51560 -297920
rect 51560 -297980 53120 -297920
rect 53120 -297980 54560 -297920
rect 54560 -297980 56120 -297920
rect 56120 -297980 57560 -297920
rect 57560 -297980 59120 -297920
rect 59120 -297980 60560 -297920
rect 60560 -297980 62120 -297920
rect 62120 -297980 63560 -297920
rect 63560 -297980 65120 -297920
rect 65120 -297980 66560 -297920
rect 66560 -297980 68120 -297920
rect 68120 -297980 69560 -297920
rect 69560 -297980 71120 -297920
rect 71120 -297980 72560 -297920
rect 72560 -297980 74120 -297920
rect 74120 -297980 75560 -297920
rect 75560 -297980 77120 -297920
rect 77120 -297980 78560 -297920
rect 78560 -297980 80120 -297920
rect 80120 -297980 81560 -297920
rect 81560 -297980 83120 -297920
rect 83120 -297980 84560 -297920
rect 84560 -297980 86120 -297920
rect 86120 -297980 87560 -297920
rect 87560 -297980 89120 -297920
rect 89120 -297980 90560 -297920
rect 90560 -297980 92120 -297920
rect 92120 -297980 93560 -297920
rect 93560 -297980 95120 -297920
rect 95120 -297980 96560 -297920
rect 96560 -297980 98120 -297920
rect 98120 -297980 99560 -297920
rect 99560 -297980 101120 -297920
rect 101120 -297980 102560 -297920
rect 102560 -297980 104120 -297920
rect 104120 -297980 105560 -297920
rect 105560 -297980 107120 -297920
rect 107120 -297980 108560 -297920
rect 108560 -297980 110120 -297920
rect 110120 -297980 111560 -297920
rect 111560 -297980 113120 -297920
rect 113120 -297980 114560 -297920
rect 114560 -297980 116120 -297920
rect 116120 -297980 117560 -297920
rect 117560 -297980 119120 -297920
rect 119120 -297980 120560 -297920
rect 120560 -297980 122120 -297920
rect 122120 -297980 123560 -297920
rect 123560 -297980 125120 -297920
rect 125120 -297980 126560 -297920
rect 126560 -297980 128120 -297920
rect 128120 -297980 129560 -297920
rect 129560 -297980 131120 -297920
rect 131120 -297980 132560 -297920
rect 132560 -297980 134120 -297920
rect 134120 -297980 135560 -297920
rect 135560 -297980 137120 -297920
rect 137120 -297980 138560 -297920
rect 138560 -297980 140120 -297920
rect 140120 -297980 141560 -297920
rect 141560 -297980 143120 -297920
rect 143120 -297980 144560 -297920
rect 144560 -297980 146120 -297920
rect 146120 -297980 147560 -297920
rect 147560 -297980 149120 -297920
rect 149120 -297980 150560 -297920
rect 150560 -297980 152120 -297920
rect 152120 -297980 153560 -297920
rect 153560 -297980 155120 -297920
rect 155120 -297980 156560 -297920
rect 156560 -297980 158120 -297920
rect 158120 -297980 159560 -297920
rect 159560 -297980 161120 -297920
rect 161120 -297980 162560 -297920
rect 162560 -297980 164120 -297920
rect 164120 -297980 165560 -297920
rect 165560 -297980 167120 -297920
rect 167120 -297980 168560 -297920
rect 168560 -297980 170120 -297920
rect 170120 -297980 171560 -297920
rect 171560 -297980 173120 -297920
rect 173120 -297980 174560 -297920
rect 174560 -297980 176120 -297920
rect 176120 -297980 177560 -297920
rect 177560 -297980 179120 -297920
rect 179120 -297980 180560 -297920
rect 180560 -297980 182120 -297920
rect 182120 -297980 183560 -297920
rect 183560 -297980 185120 -297920
rect 185120 -297980 186560 -297920
rect 186560 -297980 188120 -297920
rect 188120 -297980 189560 -297920
rect 189560 -297980 191120 -297920
rect 191120 -297980 192560 -297920
rect 192560 -297980 194120 -297920
rect 194120 -297980 195560 -297920
rect 195560 -297980 197120 -297920
rect 197120 -297980 198560 -297920
rect 198560 -297980 200120 -297920
rect 200120 -297980 201560 -297920
rect 201560 -297980 203120 -297920
rect 203120 -297980 204560 -297920
rect 204560 -297980 206120 -297920
rect 206120 -297980 207560 -297920
rect 207560 -297980 209120 -297920
rect 209120 -297980 210560 -297920
rect 210560 -297980 212120 -297920
rect 212120 -297980 213560 -297920
rect 213560 -297980 215120 -297920
rect 215120 -297980 216560 -297920
rect 216560 -297980 218120 -297920
rect 218120 -297980 219560 -297920
rect 219560 -297980 221120 -297920
rect 221120 -297980 222560 -297920
rect 222560 -297980 224120 -297920
rect 224120 -297980 225560 -297920
rect 225560 -297980 227120 -297920
rect 227120 -297980 228560 -297920
rect 228560 -297980 230120 -297920
rect 230120 -297980 231560 -297920
rect 231560 -297980 233120 -297920
rect 233120 -297980 234560 -297920
rect 234560 -297980 236120 -297920
rect 236120 -297980 237560 -297920
rect 237560 -297980 239120 -297920
rect 239120 -297980 240560 -297920
rect 240560 -297980 242120 -297920
rect 242120 -297980 243560 -297920
rect 243560 -297980 245120 -297920
rect 245120 -297980 246560 -297920
rect 246560 -297980 248120 -297920
rect 248120 -297980 249560 -297920
rect 249560 -297980 251120 -297920
rect 251120 -297980 252560 -297920
rect 252560 -297980 254120 -297920
rect 254120 -297980 255560 -297920
rect 255560 -297980 257120 -297920
rect 257120 -297980 258560 -297920
rect 258560 -297980 260120 -297920
rect 260120 -297980 261560 -297920
rect 261560 -297980 263120 -297920
rect 263120 -297980 264560 -297920
rect 264560 -297980 266120 -297920
rect 266120 -297980 267560 -297920
rect 267560 -297980 269120 -297920
rect 269120 -297980 270560 -297920
rect 270560 -297980 272120 -297920
rect 272120 -297980 273560 -297920
rect 273560 -297980 275120 -297920
rect 275120 -297980 276560 -297920
rect 276560 -297980 278120 -297920
rect 278120 -297980 279560 -297920
rect 279560 -297980 281120 -297920
rect 281120 -297980 282560 -297920
rect 282560 -297980 284120 -297920
rect 284120 -297980 285560 -297920
rect 285560 -297980 287120 -297920
rect 287120 -297980 288560 -297920
rect 288560 -297980 290120 -297920
rect 290120 -297980 291560 -297920
rect 291560 -297980 293120 -297920
rect 293120 -297980 294560 -297920
rect 294560 -297980 296120 -297920
rect 296120 -297980 297560 -297920
rect 297560 -297980 299120 -297920
rect 299120 -297980 300740 -297920
rect 560 -298080 300740 -297980
<< metal2 >>
rect 0 4040 300000 4150
rect -3000 3450 -890 3460
rect -3000 3360 -1920 3450
rect -900 3360 -890 3450
rect -3000 3350 -890 3360
rect -3000 1560 -1000 1570
rect -3000 1490 -1580 1560
rect -1180 1490 -1000 1560
rect -3000 1480 -1000 1490
rect -750 230 -640 4000
rect 480 3650 590 3660
rect 480 3560 490 3650
rect 580 3560 590 3650
rect 480 3550 590 3560
rect 40 3450 150 3460
rect 40 3360 50 3450
rect 140 3360 150 3450
rect 40 3350 150 3360
rect 60 3000 130 3350
rect 500 3000 570 3550
rect 1020 3000 1090 4040
rect 3480 3650 3590 3660
rect 3480 3560 3490 3650
rect 3580 3560 3590 3650
rect 3480 3550 3590 3560
rect 3040 3450 3150 3460
rect 3040 3360 3050 3450
rect 3140 3360 3150 3450
rect 3040 3350 3150 3360
rect 3060 3000 3130 3350
rect 3500 3000 3570 3550
rect 4020 3000 4090 4040
rect 6480 3650 6590 3660
rect 6480 3560 6490 3650
rect 6580 3560 6590 3650
rect 6480 3550 6590 3560
rect 6040 3450 6150 3460
rect 6040 3360 6050 3450
rect 6140 3360 6150 3450
rect 6040 3350 6150 3360
rect 6060 3000 6130 3350
rect 6500 3000 6570 3550
rect 7020 3000 7090 4040
rect 9480 3650 9590 3660
rect 9480 3560 9490 3650
rect 9580 3560 9590 3650
rect 9480 3550 9590 3560
rect 9040 3450 9150 3460
rect 9040 3360 9050 3450
rect 9140 3360 9150 3450
rect 9040 3350 9150 3360
rect 9060 3000 9130 3350
rect 9500 3000 9570 3550
rect 10020 3000 10090 4040
rect 12480 3650 12590 3660
rect 12480 3560 12490 3650
rect 12580 3560 12590 3650
rect 12480 3550 12590 3560
rect 12040 3450 12150 3460
rect 12040 3360 12050 3450
rect 12140 3360 12150 3450
rect 12040 3350 12150 3360
rect 12060 3000 12130 3350
rect 12500 3000 12570 3550
rect 13020 3000 13090 4040
rect 15480 3650 15590 3660
rect 15480 3560 15490 3650
rect 15580 3560 15590 3650
rect 15480 3550 15590 3560
rect 15040 3450 15150 3460
rect 15040 3360 15050 3450
rect 15140 3360 15150 3450
rect 15040 3350 15150 3360
rect 15060 3000 15130 3350
rect 15500 3000 15570 3550
rect 16020 3000 16090 4040
rect 18480 3650 18590 3660
rect 18480 3560 18490 3650
rect 18580 3560 18590 3650
rect 18480 3550 18590 3560
rect 18040 3450 18150 3460
rect 18040 3360 18050 3450
rect 18140 3360 18150 3450
rect 18040 3350 18150 3360
rect 18060 3000 18130 3350
rect 18500 3000 18570 3550
rect 19020 3000 19090 4040
rect 21480 3650 21590 3660
rect 21480 3560 21490 3650
rect 21580 3560 21590 3650
rect 21480 3550 21590 3560
rect 21040 3450 21150 3460
rect 21040 3360 21050 3450
rect 21140 3360 21150 3450
rect 21040 3350 21150 3360
rect 21060 3000 21130 3350
rect 21500 3000 21570 3550
rect 22020 3000 22090 4040
rect 24480 3650 24590 3660
rect 24480 3560 24490 3650
rect 24580 3560 24590 3650
rect 24480 3550 24590 3560
rect 24040 3450 24150 3460
rect 24040 3360 24050 3450
rect 24140 3360 24150 3450
rect 24040 3350 24150 3360
rect 24060 3000 24130 3350
rect 24500 3000 24570 3550
rect 25020 3000 25090 4040
rect 27480 3650 27590 3660
rect 27480 3560 27490 3650
rect 27580 3560 27590 3650
rect 27480 3550 27590 3560
rect 27040 3450 27150 3460
rect 27040 3360 27050 3450
rect 27140 3360 27150 3450
rect 27040 3350 27150 3360
rect 27060 3000 27130 3350
rect 27500 3000 27570 3550
rect 28020 3000 28090 4040
rect 30480 3650 30590 3660
rect 30480 3560 30490 3650
rect 30580 3560 30590 3650
rect 30480 3550 30590 3560
rect 30040 3450 30150 3460
rect 30040 3360 30050 3450
rect 30140 3360 30150 3450
rect 30040 3350 30150 3360
rect 30060 3000 30130 3350
rect 30500 3000 30570 3550
rect 31020 3000 31090 4040
rect 33480 3650 33590 3660
rect 33480 3560 33490 3650
rect 33580 3560 33590 3650
rect 33480 3550 33590 3560
rect 33040 3450 33150 3460
rect 33040 3360 33050 3450
rect 33140 3360 33150 3450
rect 33040 3350 33150 3360
rect 33060 3000 33130 3350
rect 33500 3000 33570 3550
rect 34020 3000 34090 4040
rect 36480 3650 36590 3660
rect 36480 3560 36490 3650
rect 36580 3560 36590 3650
rect 36480 3550 36590 3560
rect 36040 3450 36150 3460
rect 36040 3360 36050 3450
rect 36140 3360 36150 3450
rect 36040 3350 36150 3360
rect 36060 3000 36130 3350
rect 36500 3000 36570 3550
rect 37020 3000 37090 4040
rect 39480 3650 39590 3660
rect 39480 3560 39490 3650
rect 39580 3560 39590 3650
rect 39480 3550 39590 3560
rect 39040 3450 39150 3460
rect 39040 3360 39050 3450
rect 39140 3360 39150 3450
rect 39040 3350 39150 3360
rect 39060 3000 39130 3350
rect 39500 3000 39570 3550
rect 40020 3000 40090 4040
rect 42480 3650 42590 3660
rect 42480 3560 42490 3650
rect 42580 3560 42590 3650
rect 42480 3550 42590 3560
rect 42040 3450 42150 3460
rect 42040 3360 42050 3450
rect 42140 3360 42150 3450
rect 42040 3350 42150 3360
rect 42060 3000 42130 3350
rect 42500 3000 42570 3550
rect 43020 3000 43090 4040
rect 45480 3650 45590 3660
rect 45480 3560 45490 3650
rect 45580 3560 45590 3650
rect 45480 3550 45590 3560
rect 45040 3450 45150 3460
rect 45040 3360 45050 3450
rect 45140 3360 45150 3450
rect 45040 3350 45150 3360
rect 45060 3000 45130 3350
rect 45500 3000 45570 3550
rect 46020 3000 46090 4040
rect 48480 3650 48590 3660
rect 48480 3560 48490 3650
rect 48580 3560 48590 3650
rect 48480 3550 48590 3560
rect 48040 3450 48150 3460
rect 48040 3360 48050 3450
rect 48140 3360 48150 3450
rect 48040 3350 48150 3360
rect 48060 3000 48130 3350
rect 48500 3000 48570 3550
rect 49020 3000 49090 4040
rect 51480 3650 51590 3660
rect 51480 3560 51490 3650
rect 51580 3560 51590 3650
rect 51480 3550 51590 3560
rect 51040 3450 51150 3460
rect 51040 3360 51050 3450
rect 51140 3360 51150 3450
rect 51040 3350 51150 3360
rect 51060 3000 51130 3350
rect 51500 3000 51570 3550
rect 52020 3000 52090 4040
rect 54480 3650 54590 3660
rect 54480 3560 54490 3650
rect 54580 3560 54590 3650
rect 54480 3550 54590 3560
rect 54040 3450 54150 3460
rect 54040 3360 54050 3450
rect 54140 3360 54150 3450
rect 54040 3350 54150 3360
rect 54060 3000 54130 3350
rect 54500 3000 54570 3550
rect 55020 3000 55090 4040
rect 57480 3650 57590 3660
rect 57480 3560 57490 3650
rect 57580 3560 57590 3650
rect 57480 3550 57590 3560
rect 57040 3450 57150 3460
rect 57040 3360 57050 3450
rect 57140 3360 57150 3450
rect 57040 3350 57150 3360
rect 57060 3000 57130 3350
rect 57500 3000 57570 3550
rect 58020 3000 58090 4040
rect 60480 3650 60590 3660
rect 60480 3560 60490 3650
rect 60580 3560 60590 3650
rect 60480 3550 60590 3560
rect 60040 3450 60150 3460
rect 60040 3360 60050 3450
rect 60140 3360 60150 3450
rect 60040 3350 60150 3360
rect 60060 3000 60130 3350
rect 60500 3000 60570 3550
rect 61020 3000 61090 4040
rect 63480 3650 63590 3660
rect 63480 3560 63490 3650
rect 63580 3560 63590 3650
rect 63480 3550 63590 3560
rect 63040 3450 63150 3460
rect 63040 3360 63050 3450
rect 63140 3360 63150 3450
rect 63040 3350 63150 3360
rect 63060 3000 63130 3350
rect 63500 3000 63570 3550
rect 64020 3000 64090 4040
rect 66480 3650 66590 3660
rect 66480 3560 66490 3650
rect 66580 3560 66590 3650
rect 66480 3550 66590 3560
rect 66040 3450 66150 3460
rect 66040 3360 66050 3450
rect 66140 3360 66150 3450
rect 66040 3350 66150 3360
rect 66060 3000 66130 3350
rect 66500 3000 66570 3550
rect 67020 3000 67090 4040
rect 69480 3650 69590 3660
rect 69480 3560 69490 3650
rect 69580 3560 69590 3650
rect 69480 3550 69590 3560
rect 69040 3450 69150 3460
rect 69040 3360 69050 3450
rect 69140 3360 69150 3450
rect 69040 3350 69150 3360
rect 69060 3000 69130 3350
rect 69500 3000 69570 3550
rect 70020 3000 70090 4040
rect 72480 3650 72590 3660
rect 72480 3560 72490 3650
rect 72580 3560 72590 3650
rect 72480 3550 72590 3560
rect 72040 3450 72150 3460
rect 72040 3360 72050 3450
rect 72140 3360 72150 3450
rect 72040 3350 72150 3360
rect 72060 3000 72130 3350
rect 72500 3000 72570 3550
rect 73020 3000 73090 4040
rect 75480 3650 75590 3660
rect 75480 3560 75490 3650
rect 75580 3560 75590 3650
rect 75480 3550 75590 3560
rect 75040 3450 75150 3460
rect 75040 3360 75050 3450
rect 75140 3360 75150 3450
rect 75040 3350 75150 3360
rect 75060 3000 75130 3350
rect 75500 3000 75570 3550
rect 76020 3000 76090 4040
rect 78480 3650 78590 3660
rect 78480 3560 78490 3650
rect 78580 3560 78590 3650
rect 78480 3550 78590 3560
rect 78040 3450 78150 3460
rect 78040 3360 78050 3450
rect 78140 3360 78150 3450
rect 78040 3350 78150 3360
rect 78060 3000 78130 3350
rect 78500 3000 78570 3550
rect 79020 3000 79090 4040
rect 81480 3650 81590 3660
rect 81480 3560 81490 3650
rect 81580 3560 81590 3650
rect 81480 3550 81590 3560
rect 81040 3450 81150 3460
rect 81040 3360 81050 3450
rect 81140 3360 81150 3450
rect 81040 3350 81150 3360
rect 81060 3000 81130 3350
rect 81500 3000 81570 3550
rect 82020 3000 82090 4040
rect 84480 3650 84590 3660
rect 84480 3560 84490 3650
rect 84580 3560 84590 3650
rect 84480 3550 84590 3560
rect 84040 3450 84150 3460
rect 84040 3360 84050 3450
rect 84140 3360 84150 3450
rect 84040 3350 84150 3360
rect 84060 3000 84130 3350
rect 84500 3000 84570 3550
rect 85020 3000 85090 4040
rect 87480 3650 87590 3660
rect 87480 3560 87490 3650
rect 87580 3560 87590 3650
rect 87480 3550 87590 3560
rect 87040 3450 87150 3460
rect 87040 3360 87050 3450
rect 87140 3360 87150 3450
rect 87040 3350 87150 3360
rect 87060 3000 87130 3350
rect 87500 3000 87570 3550
rect 88020 3000 88090 4040
rect 90480 3650 90590 3660
rect 90480 3560 90490 3650
rect 90580 3560 90590 3650
rect 90480 3550 90590 3560
rect 90040 3450 90150 3460
rect 90040 3360 90050 3450
rect 90140 3360 90150 3450
rect 90040 3350 90150 3360
rect 90060 3000 90130 3350
rect 90500 3000 90570 3550
rect 91020 3000 91090 4040
rect 93480 3650 93590 3660
rect 93480 3560 93490 3650
rect 93580 3560 93590 3650
rect 93480 3550 93590 3560
rect 93040 3450 93150 3460
rect 93040 3360 93050 3450
rect 93140 3360 93150 3450
rect 93040 3350 93150 3360
rect 93060 3000 93130 3350
rect 93500 3000 93570 3550
rect 94020 3000 94090 4040
rect 96480 3650 96590 3660
rect 96480 3560 96490 3650
rect 96580 3560 96590 3650
rect 96480 3550 96590 3560
rect 96040 3450 96150 3460
rect 96040 3360 96050 3450
rect 96140 3360 96150 3450
rect 96040 3350 96150 3360
rect 96060 3000 96130 3350
rect 96500 3000 96570 3550
rect 97020 3000 97090 4040
rect 99480 3650 99590 3660
rect 99480 3560 99490 3650
rect 99580 3560 99590 3650
rect 99480 3550 99590 3560
rect 99040 3450 99150 3460
rect 99040 3360 99050 3450
rect 99140 3360 99150 3450
rect 99040 3350 99150 3360
rect 99060 3000 99130 3350
rect 99500 3000 99570 3550
rect 100020 3000 100090 4040
rect 102480 3650 102590 3660
rect 102480 3560 102490 3650
rect 102580 3560 102590 3650
rect 102480 3550 102590 3560
rect 102040 3450 102150 3460
rect 102040 3360 102050 3450
rect 102140 3360 102150 3450
rect 102040 3350 102150 3360
rect 102060 3000 102130 3350
rect 102500 3000 102570 3550
rect 103020 3000 103090 4040
rect 105480 3650 105590 3660
rect 105480 3560 105490 3650
rect 105580 3560 105590 3650
rect 105480 3550 105590 3560
rect 105040 3450 105150 3460
rect 105040 3360 105050 3450
rect 105140 3360 105150 3450
rect 105040 3350 105150 3360
rect 105060 3000 105130 3350
rect 105500 3000 105570 3550
rect 106020 3000 106090 4040
rect 108480 3650 108590 3660
rect 108480 3560 108490 3650
rect 108580 3560 108590 3650
rect 108480 3550 108590 3560
rect 108040 3450 108150 3460
rect 108040 3360 108050 3450
rect 108140 3360 108150 3450
rect 108040 3350 108150 3360
rect 108060 3000 108130 3350
rect 108500 3000 108570 3550
rect 109020 3000 109090 4040
rect 111480 3650 111590 3660
rect 111480 3560 111490 3650
rect 111580 3560 111590 3650
rect 111480 3550 111590 3560
rect 111040 3450 111150 3460
rect 111040 3360 111050 3450
rect 111140 3360 111150 3450
rect 111040 3350 111150 3360
rect 111060 3000 111130 3350
rect 111500 3000 111570 3550
rect 112020 3000 112090 4040
rect 114480 3650 114590 3660
rect 114480 3560 114490 3650
rect 114580 3560 114590 3650
rect 114480 3550 114590 3560
rect 114040 3450 114150 3460
rect 114040 3360 114050 3450
rect 114140 3360 114150 3450
rect 114040 3350 114150 3360
rect 114060 3000 114130 3350
rect 114500 3000 114570 3550
rect 115020 3000 115090 4040
rect 117480 3650 117590 3660
rect 117480 3560 117490 3650
rect 117580 3560 117590 3650
rect 117480 3550 117590 3560
rect 117040 3450 117150 3460
rect 117040 3360 117050 3450
rect 117140 3360 117150 3450
rect 117040 3350 117150 3360
rect 117060 3000 117130 3350
rect 117500 3000 117570 3550
rect 118020 3000 118090 4040
rect 120480 3650 120590 3660
rect 120480 3560 120490 3650
rect 120580 3560 120590 3650
rect 120480 3550 120590 3560
rect 120040 3450 120150 3460
rect 120040 3360 120050 3450
rect 120140 3360 120150 3450
rect 120040 3350 120150 3360
rect 120060 3000 120130 3350
rect 120500 3000 120570 3550
rect 121020 3000 121090 4040
rect 123480 3650 123590 3660
rect 123480 3560 123490 3650
rect 123580 3560 123590 3650
rect 123480 3550 123590 3560
rect 123040 3450 123150 3460
rect 123040 3360 123050 3450
rect 123140 3360 123150 3450
rect 123040 3350 123150 3360
rect 123060 3000 123130 3350
rect 123500 3000 123570 3550
rect 124020 3000 124090 4040
rect 126480 3650 126590 3660
rect 126480 3560 126490 3650
rect 126580 3560 126590 3650
rect 126480 3550 126590 3560
rect 126040 3450 126150 3460
rect 126040 3360 126050 3450
rect 126140 3360 126150 3450
rect 126040 3350 126150 3360
rect 126060 3000 126130 3350
rect 126500 3000 126570 3550
rect 127020 3000 127090 4040
rect 129480 3650 129590 3660
rect 129480 3560 129490 3650
rect 129580 3560 129590 3650
rect 129480 3550 129590 3560
rect 129040 3450 129150 3460
rect 129040 3360 129050 3450
rect 129140 3360 129150 3450
rect 129040 3350 129150 3360
rect 129060 3000 129130 3350
rect 129500 3000 129570 3550
rect 130020 3000 130090 4040
rect 132480 3650 132590 3660
rect 132480 3560 132490 3650
rect 132580 3560 132590 3650
rect 132480 3550 132590 3560
rect 132040 3450 132150 3460
rect 132040 3360 132050 3450
rect 132140 3360 132150 3450
rect 132040 3350 132150 3360
rect 132060 3000 132130 3350
rect 132500 3000 132570 3550
rect 133020 3000 133090 4040
rect 135480 3650 135590 3660
rect 135480 3560 135490 3650
rect 135580 3560 135590 3650
rect 135480 3550 135590 3560
rect 135040 3450 135150 3460
rect 135040 3360 135050 3450
rect 135140 3360 135150 3450
rect 135040 3350 135150 3360
rect 135060 3000 135130 3350
rect 135500 3000 135570 3550
rect 136020 3000 136090 4040
rect 138480 3650 138590 3660
rect 138480 3560 138490 3650
rect 138580 3560 138590 3650
rect 138480 3550 138590 3560
rect 138040 3450 138150 3460
rect 138040 3360 138050 3450
rect 138140 3360 138150 3450
rect 138040 3350 138150 3360
rect 138060 3000 138130 3350
rect 138500 3000 138570 3550
rect 139020 3000 139090 4040
rect 141480 3650 141590 3660
rect 141480 3560 141490 3650
rect 141580 3560 141590 3650
rect 141480 3550 141590 3560
rect 141040 3450 141150 3460
rect 141040 3360 141050 3450
rect 141140 3360 141150 3450
rect 141040 3350 141150 3360
rect 141060 3000 141130 3350
rect 141500 3000 141570 3550
rect 142020 3000 142090 4040
rect 144480 3650 144590 3660
rect 144480 3560 144490 3650
rect 144580 3560 144590 3650
rect 144480 3550 144590 3560
rect 144040 3450 144150 3460
rect 144040 3360 144050 3450
rect 144140 3360 144150 3450
rect 144040 3350 144150 3360
rect 144060 3000 144130 3350
rect 144500 3000 144570 3550
rect 145020 3000 145090 4040
rect 147480 3650 147590 3660
rect 147480 3560 147490 3650
rect 147580 3560 147590 3650
rect 147480 3550 147590 3560
rect 147040 3450 147150 3460
rect 147040 3360 147050 3450
rect 147140 3360 147150 3450
rect 147040 3350 147150 3360
rect 147060 3000 147130 3350
rect 147500 3000 147570 3550
rect 148020 3000 148090 4040
rect 150480 3650 150590 3660
rect 150480 3560 150490 3650
rect 150580 3560 150590 3650
rect 150480 3550 150590 3560
rect 150040 3450 150150 3460
rect 150040 3360 150050 3450
rect 150140 3360 150150 3450
rect 150040 3350 150150 3360
rect 150060 3000 150130 3350
rect 150500 3000 150570 3550
rect 151020 3000 151090 4040
rect 153480 3650 153590 3660
rect 153480 3560 153490 3650
rect 153580 3560 153590 3650
rect 153480 3550 153590 3560
rect 153040 3450 153150 3460
rect 153040 3360 153050 3450
rect 153140 3360 153150 3450
rect 153040 3350 153150 3360
rect 153060 3000 153130 3350
rect 153500 3000 153570 3550
rect 154020 3000 154090 4040
rect 156480 3650 156590 3660
rect 156480 3560 156490 3650
rect 156580 3560 156590 3650
rect 156480 3550 156590 3560
rect 156040 3450 156150 3460
rect 156040 3360 156050 3450
rect 156140 3360 156150 3450
rect 156040 3350 156150 3360
rect 156060 3000 156130 3350
rect 156500 3000 156570 3550
rect 157020 3000 157090 4040
rect 159480 3650 159590 3660
rect 159480 3560 159490 3650
rect 159580 3560 159590 3650
rect 159480 3550 159590 3560
rect 159040 3450 159150 3460
rect 159040 3360 159050 3450
rect 159140 3360 159150 3450
rect 159040 3350 159150 3360
rect 159060 3000 159130 3350
rect 159500 3000 159570 3550
rect 160020 3000 160090 4040
rect 162480 3650 162590 3660
rect 162480 3560 162490 3650
rect 162580 3560 162590 3650
rect 162480 3550 162590 3560
rect 162040 3450 162150 3460
rect 162040 3360 162050 3450
rect 162140 3360 162150 3450
rect 162040 3350 162150 3360
rect 162060 3000 162130 3350
rect 162500 3000 162570 3550
rect 163020 3000 163090 4040
rect 165480 3650 165590 3660
rect 165480 3560 165490 3650
rect 165580 3560 165590 3650
rect 165480 3550 165590 3560
rect 165040 3450 165150 3460
rect 165040 3360 165050 3450
rect 165140 3360 165150 3450
rect 165040 3350 165150 3360
rect 165060 3000 165130 3350
rect 165500 3000 165570 3550
rect 166020 3000 166090 4040
rect 168480 3650 168590 3660
rect 168480 3560 168490 3650
rect 168580 3560 168590 3650
rect 168480 3550 168590 3560
rect 168040 3450 168150 3460
rect 168040 3360 168050 3450
rect 168140 3360 168150 3450
rect 168040 3350 168150 3360
rect 168060 3000 168130 3350
rect 168500 3000 168570 3550
rect 169020 3000 169090 4040
rect 171480 3650 171590 3660
rect 171480 3560 171490 3650
rect 171580 3560 171590 3650
rect 171480 3550 171590 3560
rect 171040 3450 171150 3460
rect 171040 3360 171050 3450
rect 171140 3360 171150 3450
rect 171040 3350 171150 3360
rect 171060 3000 171130 3350
rect 171500 3000 171570 3550
rect 172020 3000 172090 4040
rect 174480 3650 174590 3660
rect 174480 3560 174490 3650
rect 174580 3560 174590 3650
rect 174480 3550 174590 3560
rect 174040 3450 174150 3460
rect 174040 3360 174050 3450
rect 174140 3360 174150 3450
rect 174040 3350 174150 3360
rect 174060 3000 174130 3350
rect 174500 3000 174570 3550
rect 175020 3000 175090 4040
rect 177480 3650 177590 3660
rect 177480 3560 177490 3650
rect 177580 3560 177590 3650
rect 177480 3550 177590 3560
rect 177040 3450 177150 3460
rect 177040 3360 177050 3450
rect 177140 3360 177150 3450
rect 177040 3350 177150 3360
rect 177060 3000 177130 3350
rect 177500 3000 177570 3550
rect 178020 3000 178090 4040
rect 180480 3650 180590 3660
rect 180480 3560 180490 3650
rect 180580 3560 180590 3650
rect 180480 3550 180590 3560
rect 180040 3450 180150 3460
rect 180040 3360 180050 3450
rect 180140 3360 180150 3450
rect 180040 3350 180150 3360
rect 180060 3000 180130 3350
rect 180500 3000 180570 3550
rect 181020 3000 181090 4040
rect 183480 3650 183590 3660
rect 183480 3560 183490 3650
rect 183580 3560 183590 3650
rect 183480 3550 183590 3560
rect 183040 3450 183150 3460
rect 183040 3360 183050 3450
rect 183140 3360 183150 3450
rect 183040 3350 183150 3360
rect 183060 3000 183130 3350
rect 183500 3000 183570 3550
rect 184020 3000 184090 4040
rect 186480 3650 186590 3660
rect 186480 3560 186490 3650
rect 186580 3560 186590 3650
rect 186480 3550 186590 3560
rect 186040 3450 186150 3460
rect 186040 3360 186050 3450
rect 186140 3360 186150 3450
rect 186040 3350 186150 3360
rect 186060 3000 186130 3350
rect 186500 3000 186570 3550
rect 187020 3000 187090 4040
rect 189480 3650 189590 3660
rect 189480 3560 189490 3650
rect 189580 3560 189590 3650
rect 189480 3550 189590 3560
rect 189040 3450 189150 3460
rect 189040 3360 189050 3450
rect 189140 3360 189150 3450
rect 189040 3350 189150 3360
rect 189060 3000 189130 3350
rect 189500 3000 189570 3550
rect 190020 3000 190090 4040
rect 192480 3650 192590 3660
rect 192480 3560 192490 3650
rect 192580 3560 192590 3650
rect 192480 3550 192590 3560
rect 192040 3450 192150 3460
rect 192040 3360 192050 3450
rect 192140 3360 192150 3450
rect 192040 3350 192150 3360
rect 192060 3000 192130 3350
rect 192500 3000 192570 3550
rect 193020 3000 193090 4040
rect 195480 3650 195590 3660
rect 195480 3560 195490 3650
rect 195580 3560 195590 3650
rect 195480 3550 195590 3560
rect 195040 3450 195150 3460
rect 195040 3360 195050 3450
rect 195140 3360 195150 3450
rect 195040 3350 195150 3360
rect 195060 3000 195130 3350
rect 195500 3000 195570 3550
rect 196020 3000 196090 4040
rect 198480 3650 198590 3660
rect 198480 3560 198490 3650
rect 198580 3560 198590 3650
rect 198480 3550 198590 3560
rect 198040 3450 198150 3460
rect 198040 3360 198050 3450
rect 198140 3360 198150 3450
rect 198040 3350 198150 3360
rect 198060 3000 198130 3350
rect 198500 3000 198570 3550
rect 199020 3000 199090 4040
rect 201480 3650 201590 3660
rect 201480 3560 201490 3650
rect 201580 3560 201590 3650
rect 201480 3550 201590 3560
rect 201040 3450 201150 3460
rect 201040 3360 201050 3450
rect 201140 3360 201150 3450
rect 201040 3350 201150 3360
rect 201060 3000 201130 3350
rect 201500 3000 201570 3550
rect 202020 3000 202090 4040
rect 204480 3650 204590 3660
rect 204480 3560 204490 3650
rect 204580 3560 204590 3650
rect 204480 3550 204590 3560
rect 204040 3450 204150 3460
rect 204040 3360 204050 3450
rect 204140 3360 204150 3450
rect 204040 3350 204150 3360
rect 204060 3000 204130 3350
rect 204500 3000 204570 3550
rect 205020 3000 205090 4040
rect 207480 3650 207590 3660
rect 207480 3560 207490 3650
rect 207580 3560 207590 3650
rect 207480 3550 207590 3560
rect 207040 3450 207150 3460
rect 207040 3360 207050 3450
rect 207140 3360 207150 3450
rect 207040 3350 207150 3360
rect 207060 3000 207130 3350
rect 207500 3000 207570 3550
rect 208020 3000 208090 4040
rect 210480 3650 210590 3660
rect 210480 3560 210490 3650
rect 210580 3560 210590 3650
rect 210480 3550 210590 3560
rect 210040 3450 210150 3460
rect 210040 3360 210050 3450
rect 210140 3360 210150 3450
rect 210040 3350 210150 3360
rect 210060 3000 210130 3350
rect 210500 3000 210570 3550
rect 211020 3000 211090 4040
rect 213480 3650 213590 3660
rect 213480 3560 213490 3650
rect 213580 3560 213590 3650
rect 213480 3550 213590 3560
rect 213040 3450 213150 3460
rect 213040 3360 213050 3450
rect 213140 3360 213150 3450
rect 213040 3350 213150 3360
rect 213060 3000 213130 3350
rect 213500 3000 213570 3550
rect 214020 3000 214090 4040
rect 216480 3650 216590 3660
rect 216480 3560 216490 3650
rect 216580 3560 216590 3650
rect 216480 3550 216590 3560
rect 216040 3450 216150 3460
rect 216040 3360 216050 3450
rect 216140 3360 216150 3450
rect 216040 3350 216150 3360
rect 216060 3000 216130 3350
rect 216500 3000 216570 3550
rect 217020 3000 217090 4040
rect 219480 3650 219590 3660
rect 219480 3560 219490 3650
rect 219580 3560 219590 3650
rect 219480 3550 219590 3560
rect 219040 3450 219150 3460
rect 219040 3360 219050 3450
rect 219140 3360 219150 3450
rect 219040 3350 219150 3360
rect 219060 3000 219130 3350
rect 219500 3000 219570 3550
rect 220020 3000 220090 4040
rect 222480 3650 222590 3660
rect 222480 3560 222490 3650
rect 222580 3560 222590 3650
rect 222480 3550 222590 3560
rect 222040 3450 222150 3460
rect 222040 3360 222050 3450
rect 222140 3360 222150 3450
rect 222040 3350 222150 3360
rect 222060 3000 222130 3350
rect 222500 3000 222570 3550
rect 223020 3000 223090 4040
rect 225480 3650 225590 3660
rect 225480 3560 225490 3650
rect 225580 3560 225590 3650
rect 225480 3550 225590 3560
rect 225040 3450 225150 3460
rect 225040 3360 225050 3450
rect 225140 3360 225150 3450
rect 225040 3350 225150 3360
rect 225060 3000 225130 3350
rect 225500 3000 225570 3550
rect 226020 3000 226090 4040
rect 228480 3650 228590 3660
rect 228480 3560 228490 3650
rect 228580 3560 228590 3650
rect 228480 3550 228590 3560
rect 228040 3450 228150 3460
rect 228040 3360 228050 3450
rect 228140 3360 228150 3450
rect 228040 3350 228150 3360
rect 228060 3000 228130 3350
rect 228500 3000 228570 3550
rect 229020 3000 229090 4040
rect 231480 3650 231590 3660
rect 231480 3560 231490 3650
rect 231580 3560 231590 3650
rect 231480 3550 231590 3560
rect 231040 3450 231150 3460
rect 231040 3360 231050 3450
rect 231140 3360 231150 3450
rect 231040 3350 231150 3360
rect 231060 3000 231130 3350
rect 231500 3000 231570 3550
rect 232020 3000 232090 4040
rect 234480 3650 234590 3660
rect 234480 3560 234490 3650
rect 234580 3560 234590 3650
rect 234480 3550 234590 3560
rect 234040 3450 234150 3460
rect 234040 3360 234050 3450
rect 234140 3360 234150 3450
rect 234040 3350 234150 3360
rect 234060 3000 234130 3350
rect 234500 3000 234570 3550
rect 235020 3000 235090 4040
rect 237480 3650 237590 3660
rect 237480 3560 237490 3650
rect 237580 3560 237590 3650
rect 237480 3550 237590 3560
rect 237040 3450 237150 3460
rect 237040 3360 237050 3450
rect 237140 3360 237150 3450
rect 237040 3350 237150 3360
rect 237060 3000 237130 3350
rect 237500 3000 237570 3550
rect 238020 3000 238090 4040
rect 240480 3650 240590 3660
rect 240480 3560 240490 3650
rect 240580 3560 240590 3650
rect 240480 3550 240590 3560
rect 240040 3450 240150 3460
rect 240040 3360 240050 3450
rect 240140 3360 240150 3450
rect 240040 3350 240150 3360
rect 240060 3000 240130 3350
rect 240500 3000 240570 3550
rect 241020 3000 241090 4040
rect 243480 3650 243590 3660
rect 243480 3560 243490 3650
rect 243580 3560 243590 3650
rect 243480 3550 243590 3560
rect 243040 3450 243150 3460
rect 243040 3360 243050 3450
rect 243140 3360 243150 3450
rect 243040 3350 243150 3360
rect 243060 3000 243130 3350
rect 243500 3000 243570 3550
rect 244020 3000 244090 4040
rect 246480 3650 246590 3660
rect 246480 3560 246490 3650
rect 246580 3560 246590 3650
rect 246480 3550 246590 3560
rect 246040 3450 246150 3460
rect 246040 3360 246050 3450
rect 246140 3360 246150 3450
rect 246040 3350 246150 3360
rect 246060 3000 246130 3350
rect 246500 3000 246570 3550
rect 247020 3000 247090 4040
rect 249480 3650 249590 3660
rect 249480 3560 249490 3650
rect 249580 3560 249590 3650
rect 249480 3550 249590 3560
rect 249040 3450 249150 3460
rect 249040 3360 249050 3450
rect 249140 3360 249150 3450
rect 249040 3350 249150 3360
rect 249060 3000 249130 3350
rect 249500 3000 249570 3550
rect 250020 3000 250090 4040
rect 252480 3650 252590 3660
rect 252480 3560 252490 3650
rect 252580 3560 252590 3650
rect 252480 3550 252590 3560
rect 252040 3450 252150 3460
rect 252040 3360 252050 3450
rect 252140 3360 252150 3450
rect 252040 3350 252150 3360
rect 252060 3000 252130 3350
rect 252500 3000 252570 3550
rect 253020 3000 253090 4040
rect 255480 3650 255590 3660
rect 255480 3560 255490 3650
rect 255580 3560 255590 3650
rect 255480 3550 255590 3560
rect 255040 3450 255150 3460
rect 255040 3360 255050 3450
rect 255140 3360 255150 3450
rect 255040 3350 255150 3360
rect 255060 3000 255130 3350
rect 255500 3000 255570 3550
rect 256020 3000 256090 4040
rect 258480 3650 258590 3660
rect 258480 3560 258490 3650
rect 258580 3560 258590 3650
rect 258480 3550 258590 3560
rect 258040 3450 258150 3460
rect 258040 3360 258050 3450
rect 258140 3360 258150 3450
rect 258040 3350 258150 3360
rect 258060 3000 258130 3350
rect 258500 3000 258570 3550
rect 259020 3000 259090 4040
rect 261480 3650 261590 3660
rect 261480 3560 261490 3650
rect 261580 3560 261590 3650
rect 261480 3550 261590 3560
rect 261040 3450 261150 3460
rect 261040 3360 261050 3450
rect 261140 3360 261150 3450
rect 261040 3350 261150 3360
rect 261060 3000 261130 3350
rect 261500 3000 261570 3550
rect 262020 3000 262090 4040
rect 264480 3650 264590 3660
rect 264480 3560 264490 3650
rect 264580 3560 264590 3650
rect 264480 3550 264590 3560
rect 264040 3450 264150 3460
rect 264040 3360 264050 3450
rect 264140 3360 264150 3450
rect 264040 3350 264150 3360
rect 264060 3000 264130 3350
rect 264500 3000 264570 3550
rect 265020 3000 265090 4040
rect 267480 3650 267590 3660
rect 267480 3560 267490 3650
rect 267580 3560 267590 3650
rect 267480 3550 267590 3560
rect 267040 3450 267150 3460
rect 267040 3360 267050 3450
rect 267140 3360 267150 3450
rect 267040 3350 267150 3360
rect 267060 3000 267130 3350
rect 267500 3000 267570 3550
rect 268020 3000 268090 4040
rect 270480 3650 270590 3660
rect 270480 3560 270490 3650
rect 270580 3560 270590 3650
rect 270480 3550 270590 3560
rect 270040 3450 270150 3460
rect 270040 3360 270050 3450
rect 270140 3360 270150 3450
rect 270040 3350 270150 3360
rect 270060 3000 270130 3350
rect 270500 3000 270570 3550
rect 271020 3000 271090 4040
rect 273480 3650 273590 3660
rect 273480 3560 273490 3650
rect 273580 3560 273590 3650
rect 273480 3550 273590 3560
rect 273040 3450 273150 3460
rect 273040 3360 273050 3450
rect 273140 3360 273150 3450
rect 273040 3350 273150 3360
rect 273060 3000 273130 3350
rect 273500 3000 273570 3550
rect 274020 3000 274090 4040
rect 276480 3650 276590 3660
rect 276480 3560 276490 3650
rect 276580 3560 276590 3650
rect 276480 3550 276590 3560
rect 276040 3450 276150 3460
rect 276040 3360 276050 3450
rect 276140 3360 276150 3450
rect 276040 3350 276150 3360
rect 276060 3000 276130 3350
rect 276500 3000 276570 3550
rect 277020 3000 277090 4040
rect 279480 3650 279590 3660
rect 279480 3560 279490 3650
rect 279580 3560 279590 3650
rect 279480 3550 279590 3560
rect 279040 3450 279150 3460
rect 279040 3360 279050 3450
rect 279140 3360 279150 3450
rect 279040 3350 279150 3360
rect 279060 3000 279130 3350
rect 279500 3000 279570 3550
rect 280020 3000 280090 4040
rect 282480 3650 282590 3660
rect 282480 3560 282490 3650
rect 282580 3560 282590 3650
rect 282480 3550 282590 3560
rect 282040 3450 282150 3460
rect 282040 3360 282050 3450
rect 282140 3360 282150 3450
rect 282040 3350 282150 3360
rect 282060 3000 282130 3350
rect 282500 3000 282570 3550
rect 283020 3000 283090 4040
rect 285480 3650 285590 3660
rect 285480 3560 285490 3650
rect 285580 3560 285590 3650
rect 285480 3550 285590 3560
rect 285040 3450 285150 3460
rect 285040 3360 285050 3450
rect 285140 3360 285150 3450
rect 285040 3350 285150 3360
rect 285060 3000 285130 3350
rect 285500 3000 285570 3550
rect 286020 3000 286090 4040
rect 288480 3650 288590 3660
rect 288480 3560 288490 3650
rect 288580 3560 288590 3650
rect 288480 3550 288590 3560
rect 288040 3450 288150 3460
rect 288040 3360 288050 3450
rect 288140 3360 288150 3450
rect 288040 3350 288150 3360
rect 288060 3000 288130 3350
rect 288500 3000 288570 3550
rect 289020 3000 289090 4040
rect 291480 3650 291590 3660
rect 291480 3560 291490 3650
rect 291580 3560 291590 3650
rect 291480 3550 291590 3560
rect 291040 3450 291150 3460
rect 291040 3360 291050 3450
rect 291140 3360 291150 3450
rect 291040 3350 291150 3360
rect 291060 3000 291130 3350
rect 291500 3000 291570 3550
rect 292020 3000 292090 4040
rect 294480 3650 294590 3660
rect 294480 3560 294490 3650
rect 294580 3560 294590 3650
rect 294480 3550 294590 3560
rect 294040 3450 294150 3460
rect 294040 3360 294050 3450
rect 294140 3360 294150 3450
rect 294040 3350 294150 3360
rect 294060 3000 294130 3350
rect 294500 3000 294570 3550
rect 295020 3000 295090 4040
rect 297480 3650 297590 3660
rect 297480 3560 297490 3650
rect 297580 3560 297590 3650
rect 297480 3550 297590 3560
rect 297040 3450 297150 3460
rect 297040 3360 297050 3450
rect 297140 3360 297150 3450
rect 297040 3350 297150 3360
rect 297060 3000 297130 3350
rect 297500 3000 297570 3550
rect 298020 3000 298090 4040
rect -560 1560 -260 1570
rect -560 1490 -540 1560
rect -560 1480 -260 1490
rect -750 160 -740 230
rect -650 160 -640 230
rect -3000 -1440 -1000 -1430
rect -3000 -1510 -1580 -1440
rect -1180 -1510 -1000 -1440
rect -3000 -1520 -1000 -1510
rect -750 -2770 -640 160
rect -560 -1440 -260 -1430
rect -560 -1510 -540 -1440
rect -560 -1520 -260 -1510
rect -750 -2840 -740 -2770
rect -650 -2840 -640 -2770
rect -3000 -4440 -1000 -4430
rect -3000 -4510 -1580 -4440
rect -1180 -4510 -1000 -4440
rect -3000 -4520 -1000 -4510
rect -750 -5770 -640 -2840
rect -560 -4440 -260 -4430
rect -560 -4510 -540 -4440
rect -560 -4520 -260 -4510
rect -750 -5840 -740 -5770
rect -650 -5840 -640 -5770
rect -3000 -7440 -1000 -7430
rect -3000 -7510 -1580 -7440
rect -1180 -7510 -1000 -7440
rect -3000 -7520 -1000 -7510
rect -750 -8770 -640 -5840
rect -560 -7440 -260 -7430
rect -560 -7510 -540 -7440
rect -560 -7520 -260 -7510
rect -750 -8840 -740 -8770
rect -650 -8840 -640 -8770
rect -3000 -10440 -1000 -10430
rect -3000 -10510 -1580 -10440
rect -1180 -10510 -1000 -10440
rect -3000 -10520 -1000 -10510
rect -750 -11770 -640 -8840
rect -560 -10440 -260 -10430
rect -560 -10510 -540 -10440
rect -560 -10520 -260 -10510
rect -750 -11840 -740 -11770
rect -650 -11840 -640 -11770
rect -3000 -13440 -1000 -13430
rect -3000 -13510 -1580 -13440
rect -1180 -13510 -1000 -13440
rect -3000 -13520 -1000 -13510
rect -750 -14770 -640 -11840
rect -560 -13440 -260 -13430
rect -560 -13510 -540 -13440
rect -560 -13520 -260 -13510
rect -750 -14840 -740 -14770
rect -650 -14840 -640 -14770
rect -3000 -16440 -1000 -16430
rect -3000 -16510 -1580 -16440
rect -1180 -16510 -1000 -16440
rect -3000 -16520 -1000 -16510
rect -750 -17770 -640 -14840
rect -560 -16440 -260 -16430
rect -560 -16510 -540 -16440
rect -560 -16520 -260 -16510
rect -750 -17840 -740 -17770
rect -650 -17840 -640 -17770
rect -3000 -19440 -1000 -19430
rect -3000 -19510 -1580 -19440
rect -1180 -19510 -1000 -19440
rect -3000 -19520 -1000 -19510
rect -750 -20770 -640 -17840
rect -560 -19440 -260 -19430
rect -560 -19510 -540 -19440
rect -560 -19520 -260 -19510
rect -750 -20840 -740 -20770
rect -650 -20840 -640 -20770
rect -3000 -22440 -1000 -22430
rect -3000 -22510 -1580 -22440
rect -1180 -22510 -1000 -22440
rect -3000 -22520 -1000 -22510
rect -750 -23770 -640 -20840
rect -560 -22440 -260 -22430
rect -560 -22510 -540 -22440
rect -560 -22520 -260 -22510
rect -750 -23840 -740 -23770
rect -650 -23840 -640 -23770
rect -3000 -25440 -1000 -25430
rect -3000 -25510 -1580 -25440
rect -1180 -25510 -1000 -25440
rect -3000 -25520 -1000 -25510
rect -750 -26770 -640 -23840
rect -560 -25440 -260 -25430
rect -560 -25510 -540 -25440
rect -560 -25520 -260 -25510
rect -750 -26840 -740 -26770
rect -650 -26840 -640 -26770
rect -3000 -28440 -1000 -28430
rect -3000 -28510 -1580 -28440
rect -1180 -28510 -1000 -28440
rect -3000 -28520 -1000 -28510
rect -750 -29770 -640 -26840
rect -560 -28440 -260 -28430
rect -560 -28510 -540 -28440
rect -560 -28520 -260 -28510
rect -750 -29840 -740 -29770
rect -650 -29840 -640 -29770
rect -3000 -31440 -1000 -31430
rect -3000 -31510 -1580 -31440
rect -1180 -31510 -1000 -31440
rect -3000 -31520 -1000 -31510
rect -750 -32770 -640 -29840
rect -560 -31440 -260 -31430
rect -560 -31510 -540 -31440
rect -560 -31520 -260 -31510
rect -750 -32840 -740 -32770
rect -650 -32840 -640 -32770
rect -3000 -34440 -1000 -34430
rect -3000 -34510 -1580 -34440
rect -1180 -34510 -1000 -34440
rect -3000 -34520 -1000 -34510
rect -750 -35770 -640 -32840
rect -560 -34440 -260 -34430
rect -560 -34510 -540 -34440
rect -560 -34520 -260 -34510
rect -750 -35840 -740 -35770
rect -650 -35840 -640 -35770
rect -3000 -37440 -1000 -37430
rect -3000 -37510 -1580 -37440
rect -1180 -37510 -1000 -37440
rect -3000 -37520 -1000 -37510
rect -750 -38770 -640 -35840
rect -560 -37440 -260 -37430
rect -560 -37510 -540 -37440
rect -560 -37520 -260 -37510
rect -750 -38840 -740 -38770
rect -650 -38840 -640 -38770
rect -3000 -40440 -1000 -40430
rect -3000 -40510 -1580 -40440
rect -1180 -40510 -1000 -40440
rect -3000 -40520 -1000 -40510
rect -750 -41770 -640 -38840
rect -560 -40440 -260 -40430
rect -560 -40510 -540 -40440
rect -560 -40520 -260 -40510
rect -750 -41840 -740 -41770
rect -650 -41840 -640 -41770
rect -3000 -43440 -1000 -43430
rect -3000 -43510 -1580 -43440
rect -1180 -43510 -1000 -43440
rect -3000 -43520 -1000 -43510
rect -750 -44770 -640 -41840
rect -560 -43440 -260 -43430
rect -560 -43510 -540 -43440
rect -560 -43520 -260 -43510
rect -750 -44840 -740 -44770
rect -650 -44840 -640 -44770
rect -3000 -46440 -1000 -46430
rect -3000 -46510 -1580 -46440
rect -1180 -46510 -1000 -46440
rect -3000 -46520 -1000 -46510
rect -750 -47770 -640 -44840
rect -560 -46440 -260 -46430
rect -560 -46510 -540 -46440
rect -560 -46520 -260 -46510
rect -750 -47840 -740 -47770
rect -650 -47840 -640 -47770
rect -3000 -49440 -1000 -49430
rect -3000 -49510 -1580 -49440
rect -1180 -49510 -1000 -49440
rect -3000 -49520 -1000 -49510
rect -750 -50770 -640 -47840
rect -560 -49440 -260 -49430
rect -560 -49510 -540 -49440
rect -560 -49520 -260 -49510
rect -750 -50840 -740 -50770
rect -650 -50840 -640 -50770
rect -3000 -52440 -1000 -52430
rect -3000 -52510 -1580 -52440
rect -1180 -52510 -1000 -52440
rect -3000 -52520 -1000 -52510
rect -750 -53770 -640 -50840
rect -560 -52440 -260 -52430
rect -560 -52510 -540 -52440
rect -560 -52520 -260 -52510
rect -750 -53840 -740 -53770
rect -650 -53840 -640 -53770
rect -3000 -55440 -1000 -55430
rect -3000 -55510 -1580 -55440
rect -1180 -55510 -1000 -55440
rect -3000 -55520 -1000 -55510
rect -750 -56770 -640 -53840
rect -560 -55440 -260 -55430
rect -560 -55510 -540 -55440
rect -560 -55520 -260 -55510
rect -750 -56840 -740 -56770
rect -650 -56840 -640 -56770
rect -3000 -58440 -1000 -58430
rect -3000 -58510 -1580 -58440
rect -1180 -58510 -1000 -58440
rect -3000 -58520 -1000 -58510
rect -750 -59770 -640 -56840
rect -560 -58440 -260 -58430
rect -560 -58510 -540 -58440
rect -560 -58520 -260 -58510
rect -750 -59840 -740 -59770
rect -650 -59840 -640 -59770
rect -3000 -61440 -1000 -61430
rect -3000 -61510 -1580 -61440
rect -1180 -61510 -1000 -61440
rect -3000 -61520 -1000 -61510
rect -750 -62770 -640 -59840
rect -560 -61440 -260 -61430
rect -560 -61510 -540 -61440
rect -560 -61520 -260 -61510
rect -750 -62840 -740 -62770
rect -650 -62840 -640 -62770
rect -3000 -64440 -1000 -64430
rect -3000 -64510 -1580 -64440
rect -1180 -64510 -1000 -64440
rect -3000 -64520 -1000 -64510
rect -750 -65770 -640 -62840
rect -560 -64440 -260 -64430
rect -560 -64510 -540 -64440
rect -560 -64520 -260 -64510
rect -750 -65840 -740 -65770
rect -650 -65840 -640 -65770
rect -3000 -67440 -1000 -67430
rect -3000 -67510 -1580 -67440
rect -1180 -67510 -1000 -67440
rect -3000 -67520 -1000 -67510
rect -750 -68770 -640 -65840
rect -560 -67440 -260 -67430
rect -560 -67510 -540 -67440
rect -560 -67520 -260 -67510
rect -750 -68840 -740 -68770
rect -650 -68840 -640 -68770
rect -3000 -70440 -1000 -70430
rect -3000 -70510 -1580 -70440
rect -1180 -70510 -1000 -70440
rect -3000 -70520 -1000 -70510
rect -750 -71770 -640 -68840
rect -560 -70440 -260 -70430
rect -560 -70510 -540 -70440
rect -560 -70520 -260 -70510
rect -750 -71840 -740 -71770
rect -650 -71840 -640 -71770
rect -3000 -73440 -1000 -73430
rect -3000 -73510 -1580 -73440
rect -1180 -73510 -1000 -73440
rect -3000 -73520 -1000 -73510
rect -750 -74770 -640 -71840
rect -560 -73440 -260 -73430
rect -560 -73510 -540 -73440
rect -560 -73520 -260 -73510
rect -750 -74840 -740 -74770
rect -650 -74840 -640 -74770
rect -3000 -76440 -1000 -76430
rect -3000 -76510 -1580 -76440
rect -1180 -76510 -1000 -76440
rect -3000 -76520 -1000 -76510
rect -750 -77770 -640 -74840
rect -560 -76440 -260 -76430
rect -560 -76510 -540 -76440
rect -560 -76520 -260 -76510
rect -750 -77840 -740 -77770
rect -650 -77840 -640 -77770
rect -3000 -79440 -1000 -79430
rect -3000 -79510 -1580 -79440
rect -1180 -79510 -1000 -79440
rect -3000 -79520 -1000 -79510
rect -750 -80770 -640 -77840
rect -560 -79440 -260 -79430
rect -560 -79510 -540 -79440
rect -560 -79520 -260 -79510
rect -750 -80840 -740 -80770
rect -650 -80840 -640 -80770
rect -3000 -82440 -1000 -82430
rect -3000 -82510 -1580 -82440
rect -1180 -82510 -1000 -82440
rect -3000 -82520 -1000 -82510
rect -750 -83770 -640 -80840
rect -560 -82440 -260 -82430
rect -560 -82510 -540 -82440
rect -560 -82520 -260 -82510
rect -750 -83840 -740 -83770
rect -650 -83840 -640 -83770
rect -3000 -85440 -1000 -85430
rect -3000 -85510 -1580 -85440
rect -1180 -85510 -1000 -85440
rect -3000 -85520 -1000 -85510
rect -750 -86770 -640 -83840
rect -560 -85440 -260 -85430
rect -560 -85510 -540 -85440
rect -560 -85520 -260 -85510
rect -750 -86840 -740 -86770
rect -650 -86840 -640 -86770
rect -3000 -88440 -1000 -88430
rect -3000 -88510 -1580 -88440
rect -1180 -88510 -1000 -88440
rect -3000 -88520 -1000 -88510
rect -750 -89770 -640 -86840
rect -560 -88440 -260 -88430
rect -560 -88510 -540 -88440
rect -560 -88520 -260 -88510
rect -750 -89840 -740 -89770
rect -650 -89840 -640 -89770
rect -3000 -91440 -1000 -91430
rect -3000 -91510 -1580 -91440
rect -1180 -91510 -1000 -91440
rect -3000 -91520 -1000 -91510
rect -750 -92770 -640 -89840
rect -560 -91440 -260 -91430
rect -560 -91510 -540 -91440
rect -560 -91520 -260 -91510
rect -750 -92840 -740 -92770
rect -650 -92840 -640 -92770
rect -3000 -94440 -1000 -94430
rect -3000 -94510 -1580 -94440
rect -1180 -94510 -1000 -94440
rect -3000 -94520 -1000 -94510
rect -750 -95770 -640 -92840
rect -560 -94440 -260 -94430
rect -560 -94510 -540 -94440
rect -560 -94520 -260 -94510
rect -750 -95840 -740 -95770
rect -650 -95840 -640 -95770
rect -3000 -97440 -1000 -97430
rect -3000 -97510 -1580 -97440
rect -1180 -97510 -1000 -97440
rect -3000 -97520 -1000 -97510
rect -750 -98770 -640 -95840
rect -560 -97440 -260 -97430
rect -560 -97510 -540 -97440
rect -560 -97520 -260 -97510
rect -750 -98840 -740 -98770
rect -650 -98840 -640 -98770
rect -3000 -100440 -1000 -100430
rect -3000 -100510 -1580 -100440
rect -1180 -100510 -1000 -100440
rect -3000 -100520 -1000 -100510
rect -750 -101770 -640 -98840
rect -560 -100440 -260 -100430
rect -560 -100510 -540 -100440
rect -560 -100520 -260 -100510
rect -750 -101840 -740 -101770
rect -650 -101840 -640 -101770
rect -3000 -103440 -1000 -103430
rect -3000 -103510 -1580 -103440
rect -1180 -103510 -1000 -103440
rect -3000 -103520 -1000 -103510
rect -750 -104770 -640 -101840
rect -560 -103440 -260 -103430
rect -560 -103510 -540 -103440
rect -560 -103520 -260 -103510
rect -750 -104840 -740 -104770
rect -650 -104840 -640 -104770
rect -3000 -106440 -1000 -106430
rect -3000 -106510 -1580 -106440
rect -1180 -106510 -1000 -106440
rect -3000 -106520 -1000 -106510
rect -750 -107770 -640 -104840
rect -560 -106440 -260 -106430
rect -560 -106510 -540 -106440
rect -560 -106520 -260 -106510
rect -750 -107840 -740 -107770
rect -650 -107840 -640 -107770
rect -3000 -109440 -1000 -109430
rect -3000 -109510 -1580 -109440
rect -1180 -109510 -1000 -109440
rect -3000 -109520 -1000 -109510
rect -750 -110770 -640 -107840
rect -560 -109440 -260 -109430
rect -560 -109510 -540 -109440
rect -560 -109520 -260 -109510
rect -750 -110840 -740 -110770
rect -650 -110840 -640 -110770
rect -3000 -112440 -1000 -112430
rect -3000 -112510 -1580 -112440
rect -1180 -112510 -1000 -112440
rect -3000 -112520 -1000 -112510
rect -750 -113770 -640 -110840
rect -560 -112440 -260 -112430
rect -560 -112510 -540 -112440
rect -560 -112520 -260 -112510
rect -750 -113840 -740 -113770
rect -650 -113840 -640 -113770
rect -3000 -115440 -1000 -115430
rect -3000 -115510 -1580 -115440
rect -1180 -115510 -1000 -115440
rect -3000 -115520 -1000 -115510
rect -750 -116770 -640 -113840
rect -560 -115440 -260 -115430
rect -560 -115510 -540 -115440
rect -560 -115520 -260 -115510
rect -750 -116840 -740 -116770
rect -650 -116840 -640 -116770
rect -3000 -118440 -1000 -118430
rect -3000 -118510 -1580 -118440
rect -1180 -118510 -1000 -118440
rect -3000 -118520 -1000 -118510
rect -750 -119770 -640 -116840
rect -560 -118440 -260 -118430
rect -560 -118510 -540 -118440
rect -560 -118520 -260 -118510
rect -750 -119840 -740 -119770
rect -650 -119840 -640 -119770
rect -3000 -121440 -1000 -121430
rect -3000 -121510 -1580 -121440
rect -1180 -121510 -1000 -121440
rect -3000 -121520 -1000 -121510
rect -750 -122770 -640 -119840
rect -560 -121440 -260 -121430
rect -560 -121510 -540 -121440
rect -560 -121520 -260 -121510
rect -750 -122840 -740 -122770
rect -650 -122840 -640 -122770
rect -3000 -124440 -1000 -124430
rect -3000 -124510 -1580 -124440
rect -1180 -124510 -1000 -124440
rect -3000 -124520 -1000 -124510
rect -750 -125770 -640 -122840
rect -560 -124440 -260 -124430
rect -560 -124510 -540 -124440
rect -560 -124520 -260 -124510
rect -750 -125840 -740 -125770
rect -650 -125840 -640 -125770
rect -3000 -127440 -1000 -127430
rect -3000 -127510 -1580 -127440
rect -1180 -127510 -1000 -127440
rect -3000 -127520 -1000 -127510
rect -750 -128770 -640 -125840
rect -560 -127440 -260 -127430
rect -560 -127510 -540 -127440
rect -560 -127520 -260 -127510
rect -750 -128840 -740 -128770
rect -650 -128840 -640 -128770
rect -3000 -130440 -1000 -130430
rect -3000 -130510 -1580 -130440
rect -1180 -130510 -1000 -130440
rect -3000 -130520 -1000 -130510
rect -750 -131770 -640 -128840
rect -560 -130440 -260 -130430
rect -560 -130510 -540 -130440
rect -560 -130520 -260 -130510
rect -750 -131840 -740 -131770
rect -650 -131840 -640 -131770
rect -3000 -133440 -1000 -133430
rect -3000 -133510 -1580 -133440
rect -1180 -133510 -1000 -133440
rect -3000 -133520 -1000 -133510
rect -750 -134770 -640 -131840
rect -560 -133440 -260 -133430
rect -560 -133510 -540 -133440
rect -560 -133520 -260 -133510
rect -750 -134840 -740 -134770
rect -650 -134840 -640 -134770
rect -3000 -136440 -1000 -136430
rect -3000 -136510 -1580 -136440
rect -1180 -136510 -1000 -136440
rect -3000 -136520 -1000 -136510
rect -750 -137770 -640 -134840
rect -560 -136440 -260 -136430
rect -560 -136510 -540 -136440
rect -560 -136520 -260 -136510
rect -750 -137840 -740 -137770
rect -650 -137840 -640 -137770
rect -3000 -139440 -1000 -139430
rect -3000 -139510 -1580 -139440
rect -1180 -139510 -1000 -139440
rect -3000 -139520 -1000 -139510
rect -750 -140770 -640 -137840
rect -560 -139440 -260 -139430
rect -560 -139510 -540 -139440
rect -560 -139520 -260 -139510
rect -750 -140840 -740 -140770
rect -650 -140840 -640 -140770
rect -3000 -142440 -1000 -142430
rect -3000 -142510 -1580 -142440
rect -1180 -142510 -1000 -142440
rect -3000 -142520 -1000 -142510
rect -750 -143770 -640 -140840
rect -560 -142440 -260 -142430
rect -560 -142510 -540 -142440
rect -560 -142520 -260 -142510
rect -750 -143840 -740 -143770
rect -650 -143840 -640 -143770
rect -3000 -145440 -1000 -145430
rect -3000 -145510 -1580 -145440
rect -1180 -145510 -1000 -145440
rect -3000 -145520 -1000 -145510
rect -750 -146770 -640 -143840
rect -560 -145440 -260 -145430
rect -560 -145510 -540 -145440
rect -560 -145520 -260 -145510
rect -750 -146840 -740 -146770
rect -650 -146840 -640 -146770
rect -3000 -148440 -1000 -148430
rect -3000 -148510 -1580 -148440
rect -1180 -148510 -1000 -148440
rect -3000 -148520 -1000 -148510
rect -750 -149770 -640 -146840
rect -560 -148440 -260 -148430
rect -560 -148510 -540 -148440
rect -560 -148520 -260 -148510
rect -750 -149840 -740 -149770
rect -650 -149840 -640 -149770
rect -3000 -151440 -1000 -151430
rect -3000 -151510 -1580 -151440
rect -1180 -151510 -1000 -151440
rect -3000 -151520 -1000 -151510
rect -750 -152770 -640 -149840
rect -560 -151440 -260 -151430
rect -560 -151510 -540 -151440
rect -560 -151520 -260 -151510
rect -750 -152840 -740 -152770
rect -650 -152840 -640 -152770
rect -3000 -154440 -1000 -154430
rect -3000 -154510 -1580 -154440
rect -1180 -154510 -1000 -154440
rect -3000 -154520 -1000 -154510
rect -750 -155770 -640 -152840
rect -560 -154440 -260 -154430
rect -560 -154510 -540 -154440
rect -560 -154520 -260 -154510
rect -750 -155840 -740 -155770
rect -650 -155840 -640 -155770
rect -3000 -157440 -1000 -157430
rect -3000 -157510 -1580 -157440
rect -1180 -157510 -1000 -157440
rect -3000 -157520 -1000 -157510
rect -750 -158770 -640 -155840
rect -560 -157440 -260 -157430
rect -560 -157510 -540 -157440
rect -560 -157520 -260 -157510
rect -750 -158840 -740 -158770
rect -650 -158840 -640 -158770
rect -3000 -160440 -1000 -160430
rect -3000 -160510 -1580 -160440
rect -1180 -160510 -1000 -160440
rect -3000 -160520 -1000 -160510
rect -750 -161770 -640 -158840
rect -560 -160440 -260 -160430
rect -560 -160510 -540 -160440
rect -560 -160520 -260 -160510
rect -750 -161840 -740 -161770
rect -650 -161840 -640 -161770
rect -3000 -163440 -1000 -163430
rect -3000 -163510 -1580 -163440
rect -1180 -163510 -1000 -163440
rect -3000 -163520 -1000 -163510
rect -750 -164770 -640 -161840
rect -560 -163440 -260 -163430
rect -560 -163510 -540 -163440
rect -560 -163520 -260 -163510
rect -750 -164840 -740 -164770
rect -650 -164840 -640 -164770
rect -3000 -166440 -1000 -166430
rect -3000 -166510 -1580 -166440
rect -1180 -166510 -1000 -166440
rect -3000 -166520 -1000 -166510
rect -750 -167770 -640 -164840
rect -560 -166440 -260 -166430
rect -560 -166510 -540 -166440
rect -560 -166520 -260 -166510
rect -750 -167840 -740 -167770
rect -650 -167840 -640 -167770
rect -3000 -169440 -1000 -169430
rect -3000 -169510 -1580 -169440
rect -1180 -169510 -1000 -169440
rect -3000 -169520 -1000 -169510
rect -750 -170770 -640 -167840
rect -560 -169440 -260 -169430
rect -560 -169510 -540 -169440
rect -560 -169520 -260 -169510
rect -750 -170840 -740 -170770
rect -650 -170840 -640 -170770
rect -3000 -172440 -1000 -172430
rect -3000 -172510 -1580 -172440
rect -1180 -172510 -1000 -172440
rect -3000 -172520 -1000 -172510
rect -750 -173770 -640 -170840
rect -560 -172440 -260 -172430
rect -560 -172510 -540 -172440
rect -560 -172520 -260 -172510
rect -750 -173840 -740 -173770
rect -650 -173840 -640 -173770
rect -3000 -175440 -1000 -175430
rect -3000 -175510 -1580 -175440
rect -1180 -175510 -1000 -175440
rect -3000 -175520 -1000 -175510
rect -750 -176770 -640 -173840
rect -560 -175440 -260 -175430
rect -560 -175510 -540 -175440
rect -560 -175520 -260 -175510
rect -750 -176840 -740 -176770
rect -650 -176840 -640 -176770
rect -3000 -178440 -1000 -178430
rect -3000 -178510 -1580 -178440
rect -1180 -178510 -1000 -178440
rect -3000 -178520 -1000 -178510
rect -750 -179770 -640 -176840
rect -560 -178440 -260 -178430
rect -560 -178510 -540 -178440
rect -560 -178520 -260 -178510
rect -750 -179840 -740 -179770
rect -650 -179840 -640 -179770
rect -3000 -181440 -1000 -181430
rect -3000 -181510 -1580 -181440
rect -1180 -181510 -1000 -181440
rect -3000 -181520 -1000 -181510
rect -750 -182770 -640 -179840
rect -560 -181440 -260 -181430
rect -560 -181510 -540 -181440
rect -560 -181520 -260 -181510
rect -750 -182840 -740 -182770
rect -650 -182840 -640 -182770
rect -3000 -184440 -1000 -184430
rect -3000 -184510 -1580 -184440
rect -1180 -184510 -1000 -184440
rect -3000 -184520 -1000 -184510
rect -750 -185770 -640 -182840
rect -560 -184440 -260 -184430
rect -560 -184510 -540 -184440
rect -560 -184520 -260 -184510
rect -750 -185840 -740 -185770
rect -650 -185840 -640 -185770
rect -3000 -187440 -1000 -187430
rect -3000 -187510 -1580 -187440
rect -1180 -187510 -1000 -187440
rect -3000 -187520 -1000 -187510
rect -750 -188770 -640 -185840
rect -560 -187440 -260 -187430
rect -560 -187510 -540 -187440
rect -560 -187520 -260 -187510
rect -750 -188840 -740 -188770
rect -650 -188840 -640 -188770
rect -3000 -190440 -1000 -190430
rect -3000 -190510 -1580 -190440
rect -1180 -190510 -1000 -190440
rect -3000 -190520 -1000 -190510
rect -750 -191770 -640 -188840
rect -560 -190440 -260 -190430
rect -560 -190510 -540 -190440
rect -560 -190520 -260 -190510
rect -750 -191840 -740 -191770
rect -650 -191840 -640 -191770
rect -3000 -193440 -1000 -193430
rect -3000 -193510 -1580 -193440
rect -1180 -193510 -1000 -193440
rect -3000 -193520 -1000 -193510
rect -750 -194770 -640 -191840
rect -560 -193440 -260 -193430
rect -560 -193510 -540 -193440
rect -560 -193520 -260 -193510
rect -750 -194840 -740 -194770
rect -650 -194840 -640 -194770
rect -3000 -196440 -1000 -196430
rect -3000 -196510 -1580 -196440
rect -1180 -196510 -1000 -196440
rect -3000 -196520 -1000 -196510
rect -750 -197770 -640 -194840
rect -560 -196440 -260 -196430
rect -560 -196510 -540 -196440
rect -560 -196520 -260 -196510
rect -750 -197840 -740 -197770
rect -650 -197840 -640 -197770
rect -3000 -199440 -1000 -199430
rect -3000 -199510 -1580 -199440
rect -1180 -199510 -1000 -199440
rect -3000 -199520 -1000 -199510
rect -750 -200770 -640 -197840
rect -560 -199440 -260 -199430
rect -560 -199510 -540 -199440
rect -560 -199520 -260 -199510
rect -750 -200840 -740 -200770
rect -650 -200840 -640 -200770
rect -3000 -202440 -1000 -202430
rect -3000 -202510 -1580 -202440
rect -1180 -202510 -1000 -202440
rect -3000 -202520 -1000 -202510
rect -750 -203770 -640 -200840
rect -560 -202440 -260 -202430
rect -560 -202510 -540 -202440
rect -560 -202520 -260 -202510
rect -750 -203840 -740 -203770
rect -650 -203840 -640 -203770
rect -3000 -205440 -1000 -205430
rect -3000 -205510 -1580 -205440
rect -1180 -205510 -1000 -205440
rect -3000 -205520 -1000 -205510
rect -750 -206770 -640 -203840
rect -560 -205440 -260 -205430
rect -560 -205510 -540 -205440
rect -560 -205520 -260 -205510
rect -750 -206840 -740 -206770
rect -650 -206840 -640 -206770
rect -3000 -208440 -1000 -208430
rect -3000 -208510 -1580 -208440
rect -1180 -208510 -1000 -208440
rect -3000 -208520 -1000 -208510
rect -750 -209770 -640 -206840
rect -560 -208440 -260 -208430
rect -560 -208510 -540 -208440
rect -560 -208520 -260 -208510
rect -750 -209840 -740 -209770
rect -650 -209840 -640 -209770
rect -3000 -211440 -1000 -211430
rect -3000 -211510 -1580 -211440
rect -1180 -211510 -1000 -211440
rect -3000 -211520 -1000 -211510
rect -750 -212770 -640 -209840
rect -560 -211440 -260 -211430
rect -560 -211510 -540 -211440
rect -560 -211520 -260 -211510
rect -750 -212840 -740 -212770
rect -650 -212840 -640 -212770
rect -3000 -214440 -1000 -214430
rect -3000 -214510 -1580 -214440
rect -1180 -214510 -1000 -214440
rect -3000 -214520 -1000 -214510
rect -750 -215770 -640 -212840
rect -560 -214440 -260 -214430
rect -560 -214510 -540 -214440
rect -560 -214520 -260 -214510
rect -750 -215840 -740 -215770
rect -650 -215840 -640 -215770
rect -3000 -217440 -1000 -217430
rect -3000 -217510 -1580 -217440
rect -1180 -217510 -1000 -217440
rect -3000 -217520 -1000 -217510
rect -750 -218770 -640 -215840
rect -560 -217440 -260 -217430
rect -560 -217510 -540 -217440
rect -560 -217520 -260 -217510
rect -750 -218840 -740 -218770
rect -650 -218840 -640 -218770
rect -3000 -220440 -1000 -220430
rect -3000 -220510 -1580 -220440
rect -1180 -220510 -1000 -220440
rect -3000 -220520 -1000 -220510
rect -750 -221770 -640 -218840
rect -560 -220440 -260 -220430
rect -560 -220510 -540 -220440
rect -560 -220520 -260 -220510
rect -750 -221840 -740 -221770
rect -650 -221840 -640 -221770
rect -3000 -223440 -1000 -223430
rect -3000 -223510 -1580 -223440
rect -1180 -223510 -1000 -223440
rect -3000 -223520 -1000 -223510
rect -750 -224770 -640 -221840
rect -560 -223440 -260 -223430
rect -560 -223510 -540 -223440
rect -560 -223520 -260 -223510
rect -750 -224840 -740 -224770
rect -650 -224840 -640 -224770
rect -3000 -226440 -1000 -226430
rect -3000 -226510 -1580 -226440
rect -1180 -226510 -1000 -226440
rect -3000 -226520 -1000 -226510
rect -750 -227770 -640 -224840
rect -560 -226440 -260 -226430
rect -560 -226510 -540 -226440
rect -560 -226520 -260 -226510
rect -750 -227840 -740 -227770
rect -650 -227840 -640 -227770
rect -3000 -229440 -1000 -229430
rect -3000 -229510 -1580 -229440
rect -1180 -229510 -1000 -229440
rect -3000 -229520 -1000 -229510
rect -750 -230770 -640 -227840
rect -560 -229440 -260 -229430
rect -560 -229510 -540 -229440
rect -560 -229520 -260 -229510
rect -750 -230840 -740 -230770
rect -650 -230840 -640 -230770
rect -3000 -232440 -1000 -232430
rect -3000 -232510 -1580 -232440
rect -1180 -232510 -1000 -232440
rect -3000 -232520 -1000 -232510
rect -750 -233770 -640 -230840
rect -560 -232440 -260 -232430
rect -560 -232510 -540 -232440
rect -560 -232520 -260 -232510
rect -750 -233840 -740 -233770
rect -650 -233840 -640 -233770
rect -3000 -235440 -1000 -235430
rect -3000 -235510 -1580 -235440
rect -1180 -235510 -1000 -235440
rect -3000 -235520 -1000 -235510
rect -750 -236770 -640 -233840
rect -560 -235440 -260 -235430
rect -560 -235510 -540 -235440
rect -560 -235520 -260 -235510
rect -750 -236840 -740 -236770
rect -650 -236840 -640 -236770
rect -3000 -238440 -1000 -238430
rect -3000 -238510 -1580 -238440
rect -1180 -238510 -1000 -238440
rect -3000 -238520 -1000 -238510
rect -750 -239770 -640 -236840
rect -560 -238440 -260 -238430
rect -560 -238510 -540 -238440
rect -560 -238520 -260 -238510
rect -750 -239840 -740 -239770
rect -650 -239840 -640 -239770
rect -3000 -241440 -1000 -241430
rect -3000 -241510 -1580 -241440
rect -1180 -241510 -1000 -241440
rect -3000 -241520 -1000 -241510
rect -750 -242770 -640 -239840
rect -560 -241440 -260 -241430
rect -560 -241510 -540 -241440
rect -560 -241520 -260 -241510
rect -750 -242840 -740 -242770
rect -650 -242840 -640 -242770
rect -3000 -244440 -1000 -244430
rect -3000 -244510 -1580 -244440
rect -1180 -244510 -1000 -244440
rect -3000 -244520 -1000 -244510
rect -750 -245770 -640 -242840
rect -560 -244440 -260 -244430
rect -560 -244510 -540 -244440
rect -560 -244520 -260 -244510
rect -750 -245840 -740 -245770
rect -650 -245840 -640 -245770
rect -3000 -247440 -1000 -247430
rect -3000 -247510 -1580 -247440
rect -1180 -247510 -1000 -247440
rect -3000 -247520 -1000 -247510
rect -750 -248770 -640 -245840
rect -560 -247440 -260 -247430
rect -560 -247510 -540 -247440
rect -560 -247520 -260 -247510
rect -750 -248840 -740 -248770
rect -650 -248840 -640 -248770
rect -3000 -250440 -1000 -250430
rect -3000 -250510 -1580 -250440
rect -1180 -250510 -1000 -250440
rect -3000 -250520 -1000 -250510
rect -750 -251770 -640 -248840
rect -560 -250440 -260 -250430
rect -560 -250510 -540 -250440
rect -560 -250520 -260 -250510
rect -750 -251840 -740 -251770
rect -650 -251840 -640 -251770
rect -3000 -253440 -1000 -253430
rect -3000 -253510 -1580 -253440
rect -1180 -253510 -1000 -253440
rect -3000 -253520 -1000 -253510
rect -750 -254770 -640 -251840
rect -560 -253440 -260 -253430
rect -560 -253510 -540 -253440
rect -560 -253520 -260 -253510
rect -750 -254840 -740 -254770
rect -650 -254840 -640 -254770
rect -3000 -256440 -1000 -256430
rect -3000 -256510 -1580 -256440
rect -1180 -256510 -1000 -256440
rect -3000 -256520 -1000 -256510
rect -750 -257770 -640 -254840
rect -560 -256440 -260 -256430
rect -560 -256510 -540 -256440
rect -560 -256520 -260 -256510
rect -750 -257840 -740 -257770
rect -650 -257840 -640 -257770
rect -3000 -259440 -1000 -259430
rect -3000 -259510 -1580 -259440
rect -1180 -259510 -1000 -259440
rect -3000 -259520 -1000 -259510
rect -750 -260770 -640 -257840
rect -560 -259440 -260 -259430
rect -560 -259510 -540 -259440
rect -560 -259520 -260 -259510
rect -750 -260840 -740 -260770
rect -650 -260840 -640 -260770
rect -3000 -262440 -1000 -262430
rect -3000 -262510 -1580 -262440
rect -1180 -262510 -1000 -262440
rect -3000 -262520 -1000 -262510
rect -750 -263770 -640 -260840
rect -560 -262440 -260 -262430
rect -560 -262510 -540 -262440
rect -560 -262520 -260 -262510
rect -750 -263840 -740 -263770
rect -650 -263840 -640 -263770
rect -3000 -265440 -1000 -265430
rect -3000 -265510 -1580 -265440
rect -1180 -265510 -1000 -265440
rect -3000 -265520 -1000 -265510
rect -750 -266770 -640 -263840
rect -560 -265440 -260 -265430
rect -560 -265510 -540 -265440
rect -560 -265520 -260 -265510
rect -750 -266840 -740 -266770
rect -650 -266840 -640 -266770
rect -3000 -268440 -1000 -268430
rect -3000 -268510 -1580 -268440
rect -1180 -268510 -1000 -268440
rect -3000 -268520 -1000 -268510
rect -750 -269770 -640 -266840
rect -560 -268440 -260 -268430
rect -560 -268510 -540 -268440
rect -560 -268520 -260 -268510
rect -750 -269840 -740 -269770
rect -650 -269840 -640 -269770
rect -3000 -271440 -1000 -271430
rect -3000 -271510 -1580 -271440
rect -1180 -271510 -1000 -271440
rect -3000 -271520 -1000 -271510
rect -750 -272770 -640 -269840
rect -560 -271440 -260 -271430
rect -560 -271510 -540 -271440
rect -560 -271520 -260 -271510
rect -750 -272840 -740 -272770
rect -650 -272840 -640 -272770
rect -3000 -274440 -1000 -274430
rect -3000 -274510 -1580 -274440
rect -1180 -274510 -1000 -274440
rect -3000 -274520 -1000 -274510
rect -750 -275770 -640 -272840
rect -560 -274440 -260 -274430
rect -560 -274510 -540 -274440
rect -560 -274520 -260 -274510
rect -750 -275840 -740 -275770
rect -650 -275840 -640 -275770
rect -3000 -277440 -1000 -277430
rect -3000 -277510 -1580 -277440
rect -1180 -277510 -1000 -277440
rect -3000 -277520 -1000 -277510
rect -750 -278770 -640 -275840
rect -560 -277440 -260 -277430
rect -560 -277510 -540 -277440
rect -560 -277520 -260 -277510
rect -750 -278840 -740 -278770
rect -650 -278840 -640 -278770
rect -3000 -280440 -1000 -280430
rect -3000 -280510 -1580 -280440
rect -1180 -280510 -1000 -280440
rect -3000 -280520 -1000 -280510
rect -750 -281770 -640 -278840
rect -560 -280440 -260 -280430
rect -560 -280510 -540 -280440
rect -560 -280520 -260 -280510
rect -750 -281840 -740 -281770
rect -650 -281840 -640 -281770
rect -3000 -283440 -1000 -283430
rect -3000 -283510 -1580 -283440
rect -1180 -283510 -1000 -283440
rect -3000 -283520 -1000 -283510
rect -750 -284770 -640 -281840
rect -560 -283440 -260 -283430
rect -560 -283510 -540 -283440
rect -560 -283520 -260 -283510
rect -750 -284840 -740 -284770
rect -650 -284840 -640 -284770
rect -3000 -286440 -1000 -286430
rect -3000 -286510 -1580 -286440
rect -1180 -286510 -1000 -286440
rect -3000 -286520 -1000 -286510
rect -750 -287770 -640 -284840
rect -560 -286440 -260 -286430
rect -560 -286510 -540 -286440
rect -560 -286520 -260 -286510
rect -750 -287840 -740 -287770
rect -650 -287840 -640 -287770
rect -3000 -289440 -1000 -289430
rect -3000 -289510 -1580 -289440
rect -1180 -289510 -1000 -289440
rect -3000 -289520 -1000 -289510
rect -750 -290770 -640 -287840
rect -560 -289440 -260 -289430
rect -560 -289510 -540 -289440
rect -560 -289520 -260 -289510
rect -750 -290840 -740 -290770
rect -650 -290840 -640 -290770
rect -3000 -292440 -1000 -292430
rect -3000 -292510 -1580 -292440
rect -1180 -292510 -1000 -292440
rect -3000 -292520 -1000 -292510
rect -750 -293770 -640 -290840
rect -560 -292440 -260 -292430
rect -560 -292510 -540 -292440
rect -560 -292520 -260 -292510
rect -750 -293840 -740 -293770
rect -650 -293840 -640 -293770
rect -3000 -295440 -1000 -295430
rect -3000 -295510 -1580 -295440
rect -1180 -295510 -1000 -295440
rect -3000 -295520 -1000 -295510
rect -750 -296770 -640 -293840
rect -560 -295440 -260 -295430
rect -560 -295510 -540 -295440
rect -560 -295520 -260 -295510
rect -750 -296840 -740 -296770
rect -650 -296840 -640 -296770
rect -750 -297000 -640 -296840
rect 540 -297080 2780 -297060
rect 540 -297200 560 -297080
rect 2760 -297180 2780 -297080
rect 2120 -297200 2780 -297180
rect 3540 -297080 5780 -297060
rect 3540 -297200 3560 -297080
rect 5760 -297180 5780 -297080
rect 5120 -297200 5780 -297180
rect 6540 -297080 8780 -297060
rect 6540 -297200 6560 -297080
rect 8760 -297180 8780 -297080
rect 8120 -297200 8780 -297180
rect 9540 -297080 11780 -297060
rect 9540 -297200 9560 -297080
rect 11760 -297180 11780 -297080
rect 11120 -297200 11780 -297180
rect 12540 -297080 14780 -297060
rect 12540 -297200 12560 -297080
rect 14760 -297180 14780 -297080
rect 14120 -297200 14780 -297180
rect 15540 -297080 17780 -297060
rect 15540 -297200 15560 -297080
rect 17760 -297180 17780 -297080
rect 17120 -297200 17780 -297180
rect 18540 -297080 20780 -297060
rect 18540 -297200 18560 -297080
rect 20760 -297180 20780 -297080
rect 20120 -297200 20780 -297180
rect 21540 -297080 23780 -297060
rect 21540 -297200 21560 -297080
rect 23760 -297180 23780 -297080
rect 23120 -297200 23780 -297180
rect 24540 -297080 26780 -297060
rect 24540 -297200 24560 -297080
rect 26760 -297180 26780 -297080
rect 26120 -297200 26780 -297180
rect 27540 -297080 29780 -297060
rect 27540 -297200 27560 -297080
rect 29760 -297180 29780 -297080
rect 29120 -297200 29780 -297180
rect 30540 -297080 32780 -297060
rect 30540 -297200 30560 -297080
rect 32760 -297180 32780 -297080
rect 32120 -297200 32780 -297180
rect 33540 -297080 35780 -297060
rect 33540 -297200 33560 -297080
rect 35760 -297180 35780 -297080
rect 35120 -297200 35780 -297180
rect 36540 -297080 38780 -297060
rect 36540 -297200 36560 -297080
rect 38760 -297180 38780 -297080
rect 38120 -297200 38780 -297180
rect 39540 -297080 41780 -297060
rect 39540 -297200 39560 -297080
rect 41760 -297180 41780 -297080
rect 41120 -297200 41780 -297180
rect 42540 -297080 44780 -297060
rect 42540 -297200 42560 -297080
rect 44760 -297180 44780 -297080
rect 44120 -297200 44780 -297180
rect 45540 -297080 47780 -297060
rect 45540 -297200 45560 -297080
rect 47760 -297180 47780 -297080
rect 47120 -297200 47780 -297180
rect 48540 -297080 50780 -297060
rect 48540 -297200 48560 -297080
rect 50760 -297180 50780 -297080
rect 50120 -297200 50780 -297180
rect 51540 -297080 53780 -297060
rect 51540 -297200 51560 -297080
rect 53760 -297180 53780 -297080
rect 53120 -297200 53780 -297180
rect 54540 -297080 56780 -297060
rect 54540 -297200 54560 -297080
rect 56760 -297180 56780 -297080
rect 56120 -297200 56780 -297180
rect 57540 -297080 59780 -297060
rect 57540 -297200 57560 -297080
rect 59760 -297180 59780 -297080
rect 59120 -297200 59780 -297180
rect 60540 -297080 62780 -297060
rect 60540 -297200 60560 -297080
rect 62760 -297180 62780 -297080
rect 62120 -297200 62780 -297180
rect 63540 -297080 65780 -297060
rect 63540 -297200 63560 -297080
rect 65760 -297180 65780 -297080
rect 65120 -297200 65780 -297180
rect 66540 -297080 68780 -297060
rect 66540 -297200 66560 -297080
rect 68760 -297180 68780 -297080
rect 68120 -297200 68780 -297180
rect 69540 -297080 71780 -297060
rect 69540 -297200 69560 -297080
rect 71760 -297180 71780 -297080
rect 71120 -297200 71780 -297180
rect 72540 -297080 74780 -297060
rect 72540 -297200 72560 -297080
rect 74760 -297180 74780 -297080
rect 74120 -297200 74780 -297180
rect 75540 -297080 77780 -297060
rect 75540 -297200 75560 -297080
rect 77760 -297180 77780 -297080
rect 77120 -297200 77780 -297180
rect 78540 -297080 80780 -297060
rect 78540 -297200 78560 -297080
rect 80760 -297180 80780 -297080
rect 80120 -297200 80780 -297180
rect 81540 -297080 83780 -297060
rect 81540 -297200 81560 -297080
rect 83760 -297180 83780 -297080
rect 83120 -297200 83780 -297180
rect 84540 -297080 86780 -297060
rect 84540 -297200 84560 -297080
rect 86760 -297180 86780 -297080
rect 86120 -297200 86780 -297180
rect 87540 -297080 89780 -297060
rect 87540 -297200 87560 -297080
rect 89760 -297180 89780 -297080
rect 89120 -297200 89780 -297180
rect 90540 -297080 92780 -297060
rect 90540 -297200 90560 -297080
rect 92760 -297180 92780 -297080
rect 92120 -297200 92780 -297180
rect 93540 -297080 95780 -297060
rect 93540 -297200 93560 -297080
rect 95760 -297180 95780 -297080
rect 95120 -297200 95780 -297180
rect 96540 -297080 98780 -297060
rect 96540 -297200 96560 -297080
rect 98760 -297180 98780 -297080
rect 98120 -297200 98780 -297180
rect 99540 -297080 101780 -297060
rect 99540 -297200 99560 -297080
rect 101760 -297180 101780 -297080
rect 101120 -297200 101780 -297180
rect 102540 -297080 104780 -297060
rect 102540 -297200 102560 -297080
rect 104760 -297180 104780 -297080
rect 104120 -297200 104780 -297180
rect 105540 -297080 107780 -297060
rect 105540 -297200 105560 -297080
rect 107760 -297180 107780 -297080
rect 107120 -297200 107780 -297180
rect 108540 -297080 110780 -297060
rect 108540 -297200 108560 -297080
rect 110760 -297180 110780 -297080
rect 110120 -297200 110780 -297180
rect 111540 -297080 113780 -297060
rect 111540 -297200 111560 -297080
rect 113760 -297180 113780 -297080
rect 113120 -297200 113780 -297180
rect 114540 -297080 116780 -297060
rect 114540 -297200 114560 -297080
rect 116760 -297180 116780 -297080
rect 116120 -297200 116780 -297180
rect 117540 -297080 119780 -297060
rect 117540 -297200 117560 -297080
rect 119760 -297180 119780 -297080
rect 119120 -297200 119780 -297180
rect 120540 -297080 122780 -297060
rect 120540 -297200 120560 -297080
rect 122760 -297180 122780 -297080
rect 122120 -297200 122780 -297180
rect 123540 -297080 125780 -297060
rect 123540 -297200 123560 -297080
rect 125760 -297180 125780 -297080
rect 125120 -297200 125780 -297180
rect 126540 -297080 128780 -297060
rect 126540 -297200 126560 -297080
rect 128760 -297180 128780 -297080
rect 128120 -297200 128780 -297180
rect 129540 -297080 131780 -297060
rect 129540 -297200 129560 -297080
rect 131760 -297180 131780 -297080
rect 131120 -297200 131780 -297180
rect 132540 -297080 134780 -297060
rect 132540 -297200 132560 -297080
rect 134760 -297180 134780 -297080
rect 134120 -297200 134780 -297180
rect 135540 -297080 137780 -297060
rect 135540 -297200 135560 -297080
rect 137760 -297180 137780 -297080
rect 137120 -297200 137780 -297180
rect 138540 -297080 140780 -297060
rect 138540 -297200 138560 -297080
rect 140760 -297180 140780 -297080
rect 140120 -297200 140780 -297180
rect 141540 -297080 143780 -297060
rect 141540 -297200 141560 -297080
rect 143760 -297180 143780 -297080
rect 143120 -297200 143780 -297180
rect 144540 -297080 146780 -297060
rect 144540 -297200 144560 -297080
rect 146760 -297180 146780 -297080
rect 146120 -297200 146780 -297180
rect 147540 -297080 149780 -297060
rect 147540 -297200 147560 -297080
rect 149760 -297180 149780 -297080
rect 149120 -297200 149780 -297180
rect 150540 -297080 152780 -297060
rect 150540 -297200 150560 -297080
rect 152760 -297180 152780 -297080
rect 152120 -297200 152780 -297180
rect 153540 -297080 155780 -297060
rect 153540 -297200 153560 -297080
rect 155760 -297180 155780 -297080
rect 155120 -297200 155780 -297180
rect 156540 -297080 158780 -297060
rect 156540 -297200 156560 -297080
rect 158760 -297180 158780 -297080
rect 158120 -297200 158780 -297180
rect 159540 -297080 161780 -297060
rect 159540 -297200 159560 -297080
rect 161760 -297180 161780 -297080
rect 161120 -297200 161780 -297180
rect 162540 -297080 164780 -297060
rect 162540 -297200 162560 -297080
rect 164760 -297180 164780 -297080
rect 164120 -297200 164780 -297180
rect 165540 -297080 167780 -297060
rect 165540 -297200 165560 -297080
rect 167760 -297180 167780 -297080
rect 167120 -297200 167780 -297180
rect 168540 -297080 170780 -297060
rect 168540 -297200 168560 -297080
rect 170760 -297180 170780 -297080
rect 170120 -297200 170780 -297180
rect 171540 -297080 173780 -297060
rect 171540 -297200 171560 -297080
rect 173760 -297180 173780 -297080
rect 173120 -297200 173780 -297180
rect 174540 -297080 176780 -297060
rect 174540 -297200 174560 -297080
rect 176760 -297180 176780 -297080
rect 176120 -297200 176780 -297180
rect 177540 -297080 179780 -297060
rect 177540 -297200 177560 -297080
rect 179760 -297180 179780 -297080
rect 179120 -297200 179780 -297180
rect 180540 -297080 182780 -297060
rect 180540 -297200 180560 -297080
rect 182760 -297180 182780 -297080
rect 182120 -297200 182780 -297180
rect 183540 -297080 185780 -297060
rect 183540 -297200 183560 -297080
rect 185760 -297180 185780 -297080
rect 185120 -297200 185780 -297180
rect 186540 -297080 188780 -297060
rect 186540 -297200 186560 -297080
rect 188760 -297180 188780 -297080
rect 188120 -297200 188780 -297180
rect 189540 -297080 191780 -297060
rect 189540 -297200 189560 -297080
rect 191760 -297180 191780 -297080
rect 191120 -297200 191780 -297180
rect 192540 -297080 194780 -297060
rect 192540 -297200 192560 -297080
rect 194760 -297180 194780 -297080
rect 194120 -297200 194780 -297180
rect 195540 -297080 197780 -297060
rect 195540 -297200 195560 -297080
rect 197760 -297180 197780 -297080
rect 197120 -297200 197780 -297180
rect 198540 -297080 200780 -297060
rect 198540 -297200 198560 -297080
rect 200760 -297180 200780 -297080
rect 200120 -297200 200780 -297180
rect 201540 -297080 203780 -297060
rect 201540 -297200 201560 -297080
rect 203760 -297180 203780 -297080
rect 203120 -297200 203780 -297180
rect 204540 -297080 206780 -297060
rect 204540 -297200 204560 -297080
rect 206760 -297180 206780 -297080
rect 206120 -297200 206780 -297180
rect 207540 -297080 209780 -297060
rect 207540 -297200 207560 -297080
rect 209760 -297180 209780 -297080
rect 209120 -297200 209780 -297180
rect 210540 -297080 212780 -297060
rect 210540 -297200 210560 -297080
rect 212760 -297180 212780 -297080
rect 212120 -297200 212780 -297180
rect 213540 -297080 215780 -297060
rect 213540 -297200 213560 -297080
rect 215760 -297180 215780 -297080
rect 215120 -297200 215780 -297180
rect 216540 -297080 218780 -297060
rect 216540 -297200 216560 -297080
rect 218760 -297180 218780 -297080
rect 218120 -297200 218780 -297180
rect 219540 -297080 221780 -297060
rect 219540 -297200 219560 -297080
rect 221760 -297180 221780 -297080
rect 221120 -297200 221780 -297180
rect 222540 -297080 224780 -297060
rect 222540 -297200 222560 -297080
rect 224760 -297180 224780 -297080
rect 224120 -297200 224780 -297180
rect 225540 -297080 227780 -297060
rect 225540 -297200 225560 -297080
rect 227760 -297180 227780 -297080
rect 227120 -297200 227780 -297180
rect 228540 -297080 230780 -297060
rect 228540 -297200 228560 -297080
rect 230760 -297180 230780 -297080
rect 230120 -297200 230780 -297180
rect 231540 -297080 233780 -297060
rect 231540 -297200 231560 -297080
rect 233760 -297180 233780 -297080
rect 233120 -297200 233780 -297180
rect 234540 -297080 236780 -297060
rect 234540 -297200 234560 -297080
rect 236760 -297180 236780 -297080
rect 236120 -297200 236780 -297180
rect 237540 -297080 239780 -297060
rect 237540 -297200 237560 -297080
rect 239760 -297180 239780 -297080
rect 239120 -297200 239780 -297180
rect 240540 -297080 242780 -297060
rect 240540 -297200 240560 -297080
rect 242760 -297180 242780 -297080
rect 242120 -297200 242780 -297180
rect 243540 -297080 245780 -297060
rect 243540 -297200 243560 -297080
rect 245760 -297180 245780 -297080
rect 245120 -297200 245780 -297180
rect 246540 -297080 248780 -297060
rect 246540 -297200 246560 -297080
rect 248760 -297180 248780 -297080
rect 248120 -297200 248780 -297180
rect 249540 -297080 251780 -297060
rect 249540 -297200 249560 -297080
rect 251760 -297180 251780 -297080
rect 251120 -297200 251780 -297180
rect 252540 -297080 254780 -297060
rect 252540 -297200 252560 -297080
rect 254760 -297180 254780 -297080
rect 254120 -297200 254780 -297180
rect 255540 -297080 257780 -297060
rect 255540 -297200 255560 -297080
rect 257760 -297180 257780 -297080
rect 257120 -297200 257780 -297180
rect 258540 -297080 260780 -297060
rect 258540 -297200 258560 -297080
rect 260760 -297180 260780 -297080
rect 260120 -297200 260780 -297180
rect 261540 -297080 263780 -297060
rect 261540 -297200 261560 -297080
rect 263760 -297180 263780 -297080
rect 263120 -297200 263780 -297180
rect 264540 -297080 266780 -297060
rect 264540 -297200 264560 -297080
rect 266760 -297180 266780 -297080
rect 266120 -297200 266780 -297180
rect 267540 -297080 269780 -297060
rect 267540 -297200 267560 -297080
rect 269760 -297180 269780 -297080
rect 269120 -297200 269780 -297180
rect 270540 -297080 272780 -297060
rect 270540 -297200 270560 -297080
rect 272760 -297180 272780 -297080
rect 272120 -297200 272780 -297180
rect 273540 -297080 275780 -297060
rect 273540 -297200 273560 -297080
rect 275760 -297180 275780 -297080
rect 275120 -297200 275780 -297180
rect 276540 -297080 278780 -297060
rect 276540 -297200 276560 -297080
rect 278760 -297180 278780 -297080
rect 278120 -297200 278780 -297180
rect 279540 -297080 281780 -297060
rect 279540 -297200 279560 -297080
rect 281760 -297180 281780 -297080
rect 281120 -297200 281780 -297180
rect 282540 -297080 284780 -297060
rect 282540 -297200 282560 -297080
rect 284760 -297180 284780 -297080
rect 284120 -297200 284780 -297180
rect 285540 -297080 287780 -297060
rect 285540 -297200 285560 -297080
rect 287760 -297180 287780 -297080
rect 287120 -297200 287780 -297180
rect 288540 -297080 290780 -297060
rect 288540 -297200 288560 -297080
rect 290760 -297180 290780 -297080
rect 290120 -297200 290780 -297180
rect 291540 -297080 293780 -297060
rect 291540 -297200 291560 -297080
rect 293760 -297180 293780 -297080
rect 293120 -297200 293780 -297180
rect 294540 -297080 296780 -297060
rect 294540 -297200 294560 -297080
rect 296760 -297180 296780 -297080
rect 296120 -297200 296780 -297180
rect 297540 -297080 299780 -297060
rect 297540 -297200 297560 -297080
rect 299760 -297180 299780 -297080
rect 299120 -297200 299780 -297180
rect 220 -297500 440 -297490
rect 220 -297700 240 -297500
rect 420 -297700 440 -297500
rect 220 -297710 440 -297700
rect 3220 -297500 3440 -297490
rect 3220 -297700 3240 -297500
rect 3420 -297700 3440 -297500
rect 3220 -297710 3440 -297700
rect 6220 -297500 6440 -297490
rect 6220 -297700 6240 -297500
rect 6420 -297700 6440 -297500
rect 6220 -297710 6440 -297700
rect 9220 -297500 9440 -297490
rect 9220 -297700 9240 -297500
rect 9420 -297700 9440 -297500
rect 9220 -297710 9440 -297700
rect 12220 -297500 12440 -297490
rect 12220 -297700 12240 -297500
rect 12420 -297700 12440 -297500
rect 12220 -297710 12440 -297700
rect 15220 -297500 15440 -297490
rect 15220 -297700 15240 -297500
rect 15420 -297700 15440 -297500
rect 15220 -297710 15440 -297700
rect 18220 -297500 18440 -297490
rect 18220 -297700 18240 -297500
rect 18420 -297700 18440 -297500
rect 18220 -297710 18440 -297700
rect 21220 -297500 21440 -297490
rect 21220 -297700 21240 -297500
rect 21420 -297700 21440 -297500
rect 21220 -297710 21440 -297700
rect 24220 -297500 24440 -297490
rect 24220 -297700 24240 -297500
rect 24420 -297700 24440 -297500
rect 24220 -297710 24440 -297700
rect 27220 -297500 27440 -297490
rect 27220 -297700 27240 -297500
rect 27420 -297700 27440 -297500
rect 27220 -297710 27440 -297700
rect 30220 -297500 30440 -297490
rect 30220 -297700 30240 -297500
rect 30420 -297700 30440 -297500
rect 30220 -297710 30440 -297700
rect 33220 -297500 33440 -297490
rect 33220 -297700 33240 -297500
rect 33420 -297700 33440 -297500
rect 33220 -297710 33440 -297700
rect 36220 -297500 36440 -297490
rect 36220 -297700 36240 -297500
rect 36420 -297700 36440 -297500
rect 36220 -297710 36440 -297700
rect 39220 -297500 39440 -297490
rect 39220 -297700 39240 -297500
rect 39420 -297700 39440 -297500
rect 39220 -297710 39440 -297700
rect 42220 -297500 42440 -297490
rect 42220 -297700 42240 -297500
rect 42420 -297700 42440 -297500
rect 42220 -297710 42440 -297700
rect 45220 -297500 45440 -297490
rect 45220 -297700 45240 -297500
rect 45420 -297700 45440 -297500
rect 45220 -297710 45440 -297700
rect 48220 -297500 48440 -297490
rect 48220 -297700 48240 -297500
rect 48420 -297700 48440 -297500
rect 48220 -297710 48440 -297700
rect 51220 -297500 51440 -297490
rect 51220 -297700 51240 -297500
rect 51420 -297700 51440 -297500
rect 51220 -297710 51440 -297700
rect 54220 -297500 54440 -297490
rect 54220 -297700 54240 -297500
rect 54420 -297700 54440 -297500
rect 54220 -297710 54440 -297700
rect 57220 -297500 57440 -297490
rect 57220 -297700 57240 -297500
rect 57420 -297700 57440 -297500
rect 57220 -297710 57440 -297700
rect 60220 -297500 60440 -297490
rect 60220 -297700 60240 -297500
rect 60420 -297700 60440 -297500
rect 60220 -297710 60440 -297700
rect 63220 -297500 63440 -297490
rect 63220 -297700 63240 -297500
rect 63420 -297700 63440 -297500
rect 63220 -297710 63440 -297700
rect 66220 -297500 66440 -297490
rect 66220 -297700 66240 -297500
rect 66420 -297700 66440 -297500
rect 66220 -297710 66440 -297700
rect 69220 -297500 69440 -297490
rect 69220 -297700 69240 -297500
rect 69420 -297700 69440 -297500
rect 69220 -297710 69440 -297700
rect 72220 -297500 72440 -297490
rect 72220 -297700 72240 -297500
rect 72420 -297700 72440 -297500
rect 72220 -297710 72440 -297700
rect 75220 -297500 75440 -297490
rect 75220 -297700 75240 -297500
rect 75420 -297700 75440 -297500
rect 75220 -297710 75440 -297700
rect 78220 -297500 78440 -297490
rect 78220 -297700 78240 -297500
rect 78420 -297700 78440 -297500
rect 78220 -297710 78440 -297700
rect 81220 -297500 81440 -297490
rect 81220 -297700 81240 -297500
rect 81420 -297700 81440 -297500
rect 81220 -297710 81440 -297700
rect 84220 -297500 84440 -297490
rect 84220 -297700 84240 -297500
rect 84420 -297700 84440 -297500
rect 84220 -297710 84440 -297700
rect 87220 -297500 87440 -297490
rect 87220 -297700 87240 -297500
rect 87420 -297700 87440 -297500
rect 87220 -297710 87440 -297700
rect 90220 -297500 90440 -297490
rect 90220 -297700 90240 -297500
rect 90420 -297700 90440 -297500
rect 90220 -297710 90440 -297700
rect 93220 -297500 93440 -297490
rect 93220 -297700 93240 -297500
rect 93420 -297700 93440 -297500
rect 93220 -297710 93440 -297700
rect 96220 -297500 96440 -297490
rect 96220 -297700 96240 -297500
rect 96420 -297700 96440 -297500
rect 96220 -297710 96440 -297700
rect 99220 -297500 99440 -297490
rect 99220 -297700 99240 -297500
rect 99420 -297700 99440 -297500
rect 99220 -297710 99440 -297700
rect 102220 -297500 102440 -297490
rect 102220 -297700 102240 -297500
rect 102420 -297700 102440 -297500
rect 102220 -297710 102440 -297700
rect 105220 -297500 105440 -297490
rect 105220 -297700 105240 -297500
rect 105420 -297700 105440 -297500
rect 105220 -297710 105440 -297700
rect 108220 -297500 108440 -297490
rect 108220 -297700 108240 -297500
rect 108420 -297700 108440 -297500
rect 108220 -297710 108440 -297700
rect 111220 -297500 111440 -297490
rect 111220 -297700 111240 -297500
rect 111420 -297700 111440 -297500
rect 111220 -297710 111440 -297700
rect 114220 -297500 114440 -297490
rect 114220 -297700 114240 -297500
rect 114420 -297700 114440 -297500
rect 114220 -297710 114440 -297700
rect 117220 -297500 117440 -297490
rect 117220 -297700 117240 -297500
rect 117420 -297700 117440 -297500
rect 117220 -297710 117440 -297700
rect 120220 -297500 120440 -297490
rect 120220 -297700 120240 -297500
rect 120420 -297700 120440 -297500
rect 120220 -297710 120440 -297700
rect 123220 -297500 123440 -297490
rect 123220 -297700 123240 -297500
rect 123420 -297700 123440 -297500
rect 123220 -297710 123440 -297700
rect 126220 -297500 126440 -297490
rect 126220 -297700 126240 -297500
rect 126420 -297700 126440 -297500
rect 126220 -297710 126440 -297700
rect 129220 -297500 129440 -297490
rect 129220 -297700 129240 -297500
rect 129420 -297700 129440 -297500
rect 129220 -297710 129440 -297700
rect 132220 -297500 132440 -297490
rect 132220 -297700 132240 -297500
rect 132420 -297700 132440 -297500
rect 132220 -297710 132440 -297700
rect 135220 -297500 135440 -297490
rect 135220 -297700 135240 -297500
rect 135420 -297700 135440 -297500
rect 135220 -297710 135440 -297700
rect 138220 -297500 138440 -297490
rect 138220 -297700 138240 -297500
rect 138420 -297700 138440 -297500
rect 138220 -297710 138440 -297700
rect 141220 -297500 141440 -297490
rect 141220 -297700 141240 -297500
rect 141420 -297700 141440 -297500
rect 141220 -297710 141440 -297700
rect 144220 -297500 144440 -297490
rect 144220 -297700 144240 -297500
rect 144420 -297700 144440 -297500
rect 144220 -297710 144440 -297700
rect 147220 -297500 147440 -297490
rect 147220 -297700 147240 -297500
rect 147420 -297700 147440 -297500
rect 147220 -297710 147440 -297700
rect 150220 -297500 150440 -297490
rect 150220 -297700 150240 -297500
rect 150420 -297700 150440 -297500
rect 150220 -297710 150440 -297700
rect 153220 -297500 153440 -297490
rect 153220 -297700 153240 -297500
rect 153420 -297700 153440 -297500
rect 153220 -297710 153440 -297700
rect 156220 -297500 156440 -297490
rect 156220 -297700 156240 -297500
rect 156420 -297700 156440 -297500
rect 156220 -297710 156440 -297700
rect 159220 -297500 159440 -297490
rect 159220 -297700 159240 -297500
rect 159420 -297700 159440 -297500
rect 159220 -297710 159440 -297700
rect 162220 -297500 162440 -297490
rect 162220 -297700 162240 -297500
rect 162420 -297700 162440 -297500
rect 162220 -297710 162440 -297700
rect 165220 -297500 165440 -297490
rect 165220 -297700 165240 -297500
rect 165420 -297700 165440 -297500
rect 165220 -297710 165440 -297700
rect 168220 -297500 168440 -297490
rect 168220 -297700 168240 -297500
rect 168420 -297700 168440 -297500
rect 168220 -297710 168440 -297700
rect 171220 -297500 171440 -297490
rect 171220 -297700 171240 -297500
rect 171420 -297700 171440 -297500
rect 171220 -297710 171440 -297700
rect 174220 -297500 174440 -297490
rect 174220 -297700 174240 -297500
rect 174420 -297700 174440 -297500
rect 174220 -297710 174440 -297700
rect 177220 -297500 177440 -297490
rect 177220 -297700 177240 -297500
rect 177420 -297700 177440 -297500
rect 177220 -297710 177440 -297700
rect 180220 -297500 180440 -297490
rect 180220 -297700 180240 -297500
rect 180420 -297700 180440 -297500
rect 180220 -297710 180440 -297700
rect 183220 -297500 183440 -297490
rect 183220 -297700 183240 -297500
rect 183420 -297700 183440 -297500
rect 183220 -297710 183440 -297700
rect 186220 -297500 186440 -297490
rect 186220 -297700 186240 -297500
rect 186420 -297700 186440 -297500
rect 186220 -297710 186440 -297700
rect 189220 -297500 189440 -297490
rect 189220 -297700 189240 -297500
rect 189420 -297700 189440 -297500
rect 189220 -297710 189440 -297700
rect 192220 -297500 192440 -297490
rect 192220 -297700 192240 -297500
rect 192420 -297700 192440 -297500
rect 192220 -297710 192440 -297700
rect 195220 -297500 195440 -297490
rect 195220 -297700 195240 -297500
rect 195420 -297700 195440 -297500
rect 195220 -297710 195440 -297700
rect 198220 -297500 198440 -297490
rect 198220 -297700 198240 -297500
rect 198420 -297700 198440 -297500
rect 198220 -297710 198440 -297700
rect 201220 -297500 201440 -297490
rect 201220 -297700 201240 -297500
rect 201420 -297700 201440 -297500
rect 201220 -297710 201440 -297700
rect 204220 -297500 204440 -297490
rect 204220 -297700 204240 -297500
rect 204420 -297700 204440 -297500
rect 204220 -297710 204440 -297700
rect 207220 -297500 207440 -297490
rect 207220 -297700 207240 -297500
rect 207420 -297700 207440 -297500
rect 207220 -297710 207440 -297700
rect 210220 -297500 210440 -297490
rect 210220 -297700 210240 -297500
rect 210420 -297700 210440 -297500
rect 210220 -297710 210440 -297700
rect 213220 -297500 213440 -297490
rect 213220 -297700 213240 -297500
rect 213420 -297700 213440 -297500
rect 213220 -297710 213440 -297700
rect 216220 -297500 216440 -297490
rect 216220 -297700 216240 -297500
rect 216420 -297700 216440 -297500
rect 216220 -297710 216440 -297700
rect 219220 -297500 219440 -297490
rect 219220 -297700 219240 -297500
rect 219420 -297700 219440 -297500
rect 219220 -297710 219440 -297700
rect 222220 -297500 222440 -297490
rect 222220 -297700 222240 -297500
rect 222420 -297700 222440 -297500
rect 222220 -297710 222440 -297700
rect 225220 -297500 225440 -297490
rect 225220 -297700 225240 -297500
rect 225420 -297700 225440 -297500
rect 225220 -297710 225440 -297700
rect 228220 -297500 228440 -297490
rect 228220 -297700 228240 -297500
rect 228420 -297700 228440 -297500
rect 228220 -297710 228440 -297700
rect 231220 -297500 231440 -297490
rect 231220 -297700 231240 -297500
rect 231420 -297700 231440 -297500
rect 231220 -297710 231440 -297700
rect 234220 -297500 234440 -297490
rect 234220 -297700 234240 -297500
rect 234420 -297700 234440 -297500
rect 234220 -297710 234440 -297700
rect 237220 -297500 237440 -297490
rect 237220 -297700 237240 -297500
rect 237420 -297700 237440 -297500
rect 237220 -297710 237440 -297700
rect 240220 -297500 240440 -297490
rect 240220 -297700 240240 -297500
rect 240420 -297700 240440 -297500
rect 240220 -297710 240440 -297700
rect 243220 -297500 243440 -297490
rect 243220 -297700 243240 -297500
rect 243420 -297700 243440 -297500
rect 243220 -297710 243440 -297700
rect 246220 -297500 246440 -297490
rect 246220 -297700 246240 -297500
rect 246420 -297700 246440 -297500
rect 246220 -297710 246440 -297700
rect 249220 -297500 249440 -297490
rect 249220 -297700 249240 -297500
rect 249420 -297700 249440 -297500
rect 249220 -297710 249440 -297700
rect 252220 -297500 252440 -297490
rect 252220 -297700 252240 -297500
rect 252420 -297700 252440 -297500
rect 252220 -297710 252440 -297700
rect 255220 -297500 255440 -297490
rect 255220 -297700 255240 -297500
rect 255420 -297700 255440 -297500
rect 255220 -297710 255440 -297700
rect 258220 -297500 258440 -297490
rect 258220 -297700 258240 -297500
rect 258420 -297700 258440 -297500
rect 258220 -297710 258440 -297700
rect 261220 -297500 261440 -297490
rect 261220 -297700 261240 -297500
rect 261420 -297700 261440 -297500
rect 261220 -297710 261440 -297700
rect 264220 -297500 264440 -297490
rect 264220 -297700 264240 -297500
rect 264420 -297700 264440 -297500
rect 264220 -297710 264440 -297700
rect 267220 -297500 267440 -297490
rect 267220 -297700 267240 -297500
rect 267420 -297700 267440 -297500
rect 267220 -297710 267440 -297700
rect 270220 -297500 270440 -297490
rect 270220 -297700 270240 -297500
rect 270420 -297700 270440 -297500
rect 270220 -297710 270440 -297700
rect 273220 -297500 273440 -297490
rect 273220 -297700 273240 -297500
rect 273420 -297700 273440 -297500
rect 273220 -297710 273440 -297700
rect 276220 -297500 276440 -297490
rect 276220 -297700 276240 -297500
rect 276420 -297700 276440 -297500
rect 276220 -297710 276440 -297700
rect 279220 -297500 279440 -297490
rect 279220 -297700 279240 -297500
rect 279420 -297700 279440 -297500
rect 279220 -297710 279440 -297700
rect 282220 -297500 282440 -297490
rect 282220 -297700 282240 -297500
rect 282420 -297700 282440 -297500
rect 282220 -297710 282440 -297700
rect 285220 -297500 285440 -297490
rect 285220 -297700 285240 -297500
rect 285420 -297700 285440 -297500
rect 285220 -297710 285440 -297700
rect 288220 -297500 288440 -297490
rect 288220 -297700 288240 -297500
rect 288420 -297700 288440 -297500
rect 288220 -297710 288440 -297700
rect 291220 -297500 291440 -297490
rect 291220 -297700 291240 -297500
rect 291420 -297700 291440 -297500
rect 291220 -297710 291440 -297700
rect 294220 -297500 294440 -297490
rect 294220 -297700 294240 -297500
rect 294420 -297700 294440 -297500
rect 294220 -297710 294440 -297700
rect 297220 -297500 297440 -297490
rect 297220 -297700 297240 -297500
rect 297420 -297700 297440 -297500
rect 297220 -297710 297440 -297700
rect 540 -297920 300740 -297900
rect 540 -298080 560 -297920
rect 540 -298100 300740 -298080
<< via2 >>
rect 490 3560 580 3650
rect 3490 3560 3580 3650
rect 6490 3560 6580 3650
rect 9490 3560 9580 3650
rect 12490 3560 12580 3650
rect 15490 3560 15580 3650
rect 18490 3560 18580 3650
rect 21490 3560 21580 3650
rect 24490 3560 24580 3650
rect 27490 3560 27580 3650
rect 30490 3560 30580 3650
rect 33490 3560 33580 3650
rect 36490 3560 36580 3650
rect 39490 3560 39580 3650
rect 42490 3560 42580 3650
rect 45490 3560 45580 3650
rect 48490 3560 48580 3650
rect 51490 3560 51580 3650
rect 54490 3560 54580 3650
rect 57490 3560 57580 3650
rect 60490 3560 60580 3650
rect 63490 3560 63580 3650
rect 66490 3560 66580 3650
rect 69490 3560 69580 3650
rect 72490 3560 72580 3650
rect 75490 3560 75580 3650
rect 78490 3560 78580 3650
rect 81490 3560 81580 3650
rect 84490 3560 84580 3650
rect 87490 3560 87580 3650
rect 90490 3560 90580 3650
rect 93490 3560 93580 3650
rect 96490 3560 96580 3650
rect 99490 3560 99580 3650
rect 102490 3560 102580 3650
rect 105490 3560 105580 3650
rect 108490 3560 108580 3650
rect 111490 3560 111580 3650
rect 114490 3560 114580 3650
rect 117490 3560 117580 3650
rect 120490 3560 120580 3650
rect 123490 3560 123580 3650
rect 126490 3560 126580 3650
rect 129490 3560 129580 3650
rect 132490 3560 132580 3650
rect 135490 3560 135580 3650
rect 138490 3560 138580 3650
rect 141490 3560 141580 3650
rect 144490 3560 144580 3650
rect 147490 3560 147580 3650
rect 150490 3560 150580 3650
rect 153490 3560 153580 3650
rect 156490 3560 156580 3650
rect 159490 3560 159580 3650
rect 162490 3560 162580 3650
rect 165490 3560 165580 3650
rect 168490 3560 168580 3650
rect 171490 3560 171580 3650
rect 174490 3560 174580 3650
rect 177490 3560 177580 3650
rect 180490 3560 180580 3650
rect 183490 3560 183580 3650
rect 186490 3560 186580 3650
rect 189490 3560 189580 3650
rect 192490 3560 192580 3650
rect 195490 3560 195580 3650
rect 198490 3560 198580 3650
rect 201490 3560 201580 3650
rect 204490 3560 204580 3650
rect 207490 3560 207580 3650
rect 210490 3560 210580 3650
rect 213490 3560 213580 3650
rect 216490 3560 216580 3650
rect 219490 3560 219580 3650
rect 222490 3560 222580 3650
rect 225490 3560 225580 3650
rect 228490 3560 228580 3650
rect 231490 3560 231580 3650
rect 234490 3560 234580 3650
rect 237490 3560 237580 3650
rect 240490 3560 240580 3650
rect 243490 3560 243580 3650
rect 246490 3560 246580 3650
rect 249490 3560 249580 3650
rect 252490 3560 252580 3650
rect 255490 3560 255580 3650
rect 258490 3560 258580 3650
rect 261490 3560 261580 3650
rect 264490 3560 264580 3650
rect 267490 3560 267580 3650
rect 270490 3560 270580 3650
rect 273490 3560 273580 3650
rect 276490 3560 276580 3650
rect 279490 3560 279580 3650
rect 282490 3560 282580 3650
rect 285490 3560 285580 3650
rect 288490 3560 288580 3650
rect 291490 3560 291580 3650
rect 294490 3560 294580 3650
rect 297490 3560 297580 3650
rect -540 1490 -260 1560
rect -740 160 -650 230
rect -540 -1510 -260 -1440
rect -740 -2840 -650 -2770
rect -540 -4510 -260 -4440
rect -740 -5840 -650 -5770
rect -540 -7510 -260 -7440
rect -740 -8840 -650 -8770
rect -540 -10510 -260 -10440
rect -740 -11840 -650 -11770
rect -540 -13510 -260 -13440
rect -740 -14840 -650 -14770
rect -540 -16510 -260 -16440
rect -740 -17840 -650 -17770
rect -540 -19510 -260 -19440
rect -740 -20840 -650 -20770
rect -540 -22510 -260 -22440
rect -740 -23840 -650 -23770
rect -540 -25510 -260 -25440
rect -740 -26840 -650 -26770
rect -540 -28510 -260 -28440
rect -740 -29840 -650 -29770
rect -540 -31510 -260 -31440
rect -740 -32840 -650 -32770
rect -540 -34510 -260 -34440
rect -740 -35840 -650 -35770
rect -540 -37510 -260 -37440
rect -740 -38840 -650 -38770
rect -540 -40510 -260 -40440
rect -740 -41840 -650 -41770
rect -540 -43510 -260 -43440
rect -740 -44840 -650 -44770
rect -540 -46510 -260 -46440
rect -740 -47840 -650 -47770
rect -540 -49510 -260 -49440
rect -740 -50840 -650 -50770
rect -540 -52510 -260 -52440
rect -740 -53840 -650 -53770
rect -540 -55510 -260 -55440
rect -740 -56840 -650 -56770
rect -540 -58510 -260 -58440
rect -740 -59840 -650 -59770
rect -540 -61510 -260 -61440
rect -740 -62840 -650 -62770
rect -540 -64510 -260 -64440
rect -740 -65840 -650 -65770
rect -540 -67510 -260 -67440
rect -740 -68840 -650 -68770
rect -540 -70510 -260 -70440
rect -740 -71840 -650 -71770
rect -540 -73510 -260 -73440
rect -740 -74840 -650 -74770
rect -540 -76510 -260 -76440
rect -740 -77840 -650 -77770
rect -540 -79510 -260 -79440
rect -740 -80840 -650 -80770
rect -540 -82510 -260 -82440
rect -740 -83840 -650 -83770
rect -540 -85510 -260 -85440
rect -740 -86840 -650 -86770
rect -540 -88510 -260 -88440
rect -740 -89840 -650 -89770
rect -540 -91510 -260 -91440
rect -740 -92840 -650 -92770
rect -540 -94510 -260 -94440
rect -740 -95840 -650 -95770
rect -540 -97510 -260 -97440
rect -740 -98840 -650 -98770
rect -540 -100510 -260 -100440
rect -740 -101840 -650 -101770
rect -540 -103510 -260 -103440
rect -740 -104840 -650 -104770
rect -540 -106510 -260 -106440
rect -740 -107840 -650 -107770
rect -540 -109510 -260 -109440
rect -740 -110840 -650 -110770
rect -540 -112510 -260 -112440
rect -740 -113840 -650 -113770
rect -540 -115510 -260 -115440
rect -740 -116840 -650 -116770
rect -540 -118510 -260 -118440
rect -740 -119840 -650 -119770
rect -540 -121510 -260 -121440
rect -740 -122840 -650 -122770
rect -540 -124510 -260 -124440
rect -740 -125840 -650 -125770
rect -540 -127510 -260 -127440
rect -740 -128840 -650 -128770
rect -540 -130510 -260 -130440
rect -740 -131840 -650 -131770
rect -540 -133510 -260 -133440
rect -740 -134840 -650 -134770
rect -540 -136510 -260 -136440
rect -740 -137840 -650 -137770
rect -540 -139510 -260 -139440
rect -740 -140840 -650 -140770
rect -540 -142510 -260 -142440
rect -740 -143840 -650 -143770
rect -540 -145510 -260 -145440
rect -740 -146840 -650 -146770
rect -540 -148510 -260 -148440
rect -740 -149840 -650 -149770
rect -540 -151510 -260 -151440
rect -740 -152840 -650 -152770
rect -540 -154510 -260 -154440
rect -740 -155840 -650 -155770
rect -540 -157510 -260 -157440
rect -740 -158840 -650 -158770
rect -540 -160510 -260 -160440
rect -740 -161840 -650 -161770
rect -540 -163510 -260 -163440
rect -740 -164840 -650 -164770
rect -540 -166510 -260 -166440
rect -740 -167840 -650 -167770
rect -540 -169510 -260 -169440
rect -740 -170840 -650 -170770
rect -540 -172510 -260 -172440
rect -740 -173840 -650 -173770
rect -540 -175510 -260 -175440
rect -740 -176840 -650 -176770
rect -540 -178510 -260 -178440
rect -740 -179840 -650 -179770
rect -540 -181510 -260 -181440
rect -740 -182840 -650 -182770
rect -540 -184510 -260 -184440
rect -740 -185840 -650 -185770
rect -540 -187510 -260 -187440
rect -740 -188840 -650 -188770
rect -540 -190510 -260 -190440
rect -740 -191840 -650 -191770
rect -540 -193510 -260 -193440
rect -740 -194840 -650 -194770
rect -540 -196510 -260 -196440
rect -740 -197840 -650 -197770
rect -540 -199510 -260 -199440
rect -740 -200840 -650 -200770
rect -540 -202510 -260 -202440
rect -740 -203840 -650 -203770
rect -540 -205510 -260 -205440
rect -740 -206840 -650 -206770
rect -540 -208510 -260 -208440
rect -740 -209840 -650 -209770
rect -540 -211510 -260 -211440
rect -740 -212840 -650 -212770
rect -540 -214510 -260 -214440
rect -740 -215840 -650 -215770
rect -540 -217510 -260 -217440
rect -740 -218840 -650 -218770
rect -540 -220510 -260 -220440
rect -740 -221840 -650 -221770
rect -540 -223510 -260 -223440
rect -740 -224840 -650 -224770
rect -540 -226510 -260 -226440
rect -740 -227840 -650 -227770
rect -540 -229510 -260 -229440
rect -740 -230840 -650 -230770
rect -540 -232510 -260 -232440
rect -740 -233840 -650 -233770
rect -540 -235510 -260 -235440
rect -740 -236840 -650 -236770
rect -540 -238510 -260 -238440
rect -740 -239840 -650 -239770
rect -540 -241510 -260 -241440
rect -740 -242840 -650 -242770
rect -540 -244510 -260 -244440
rect -740 -245840 -650 -245770
rect -540 -247510 -260 -247440
rect -740 -248840 -650 -248770
rect -540 -250510 -260 -250440
rect -740 -251840 -650 -251770
rect -540 -253510 -260 -253440
rect -740 -254840 -650 -254770
rect -540 -256510 -260 -256440
rect -740 -257840 -650 -257770
rect -540 -259510 -260 -259440
rect -740 -260840 -650 -260770
rect -540 -262510 -260 -262440
rect -740 -263840 -650 -263770
rect -540 -265510 -260 -265440
rect -740 -266840 -650 -266770
rect -540 -268510 -260 -268440
rect -740 -269840 -650 -269770
rect -540 -271510 -260 -271440
rect -740 -272840 -650 -272770
rect -540 -274510 -260 -274440
rect -740 -275840 -650 -275770
rect -540 -277510 -260 -277440
rect -740 -278840 -650 -278770
rect -540 -280510 -260 -280440
rect -740 -281840 -650 -281770
rect -540 -283510 -260 -283440
rect -740 -284840 -650 -284770
rect -540 -286510 -260 -286440
rect -740 -287840 -650 -287770
rect -540 -289510 -260 -289440
rect -740 -290840 -650 -290770
rect -540 -292510 -260 -292440
rect -740 -293840 -650 -293770
rect -540 -295510 -260 -295440
rect -740 -296840 -650 -296770
rect 560 -297130 2760 -297080
rect 560 -297180 2120 -297130
rect 2120 -297180 2760 -297130
rect 3560 -297130 5760 -297080
rect 3560 -297180 5120 -297130
rect 5120 -297180 5760 -297130
rect 6560 -297130 8760 -297080
rect 6560 -297180 8120 -297130
rect 8120 -297180 8760 -297130
rect 9560 -297130 11760 -297080
rect 9560 -297180 11120 -297130
rect 11120 -297180 11760 -297130
rect 12560 -297130 14760 -297080
rect 12560 -297180 14120 -297130
rect 14120 -297180 14760 -297130
rect 15560 -297130 17760 -297080
rect 15560 -297180 17120 -297130
rect 17120 -297180 17760 -297130
rect 18560 -297130 20760 -297080
rect 18560 -297180 20120 -297130
rect 20120 -297180 20760 -297130
rect 21560 -297130 23760 -297080
rect 21560 -297180 23120 -297130
rect 23120 -297180 23760 -297130
rect 24560 -297130 26760 -297080
rect 24560 -297180 26120 -297130
rect 26120 -297180 26760 -297130
rect 27560 -297130 29760 -297080
rect 27560 -297180 29120 -297130
rect 29120 -297180 29760 -297130
rect 30560 -297130 32760 -297080
rect 30560 -297180 32120 -297130
rect 32120 -297180 32760 -297130
rect 33560 -297130 35760 -297080
rect 33560 -297180 35120 -297130
rect 35120 -297180 35760 -297130
rect 36560 -297130 38760 -297080
rect 36560 -297180 38120 -297130
rect 38120 -297180 38760 -297130
rect 39560 -297130 41760 -297080
rect 39560 -297180 41120 -297130
rect 41120 -297180 41760 -297130
rect 42560 -297130 44760 -297080
rect 42560 -297180 44120 -297130
rect 44120 -297180 44760 -297130
rect 45560 -297130 47760 -297080
rect 45560 -297180 47120 -297130
rect 47120 -297180 47760 -297130
rect 48560 -297130 50760 -297080
rect 48560 -297180 50120 -297130
rect 50120 -297180 50760 -297130
rect 51560 -297130 53760 -297080
rect 51560 -297180 53120 -297130
rect 53120 -297180 53760 -297130
rect 54560 -297130 56760 -297080
rect 54560 -297180 56120 -297130
rect 56120 -297180 56760 -297130
rect 57560 -297130 59760 -297080
rect 57560 -297180 59120 -297130
rect 59120 -297180 59760 -297130
rect 60560 -297130 62760 -297080
rect 60560 -297180 62120 -297130
rect 62120 -297180 62760 -297130
rect 63560 -297130 65760 -297080
rect 63560 -297180 65120 -297130
rect 65120 -297180 65760 -297130
rect 66560 -297130 68760 -297080
rect 66560 -297180 68120 -297130
rect 68120 -297180 68760 -297130
rect 69560 -297130 71760 -297080
rect 69560 -297180 71120 -297130
rect 71120 -297180 71760 -297130
rect 72560 -297130 74760 -297080
rect 72560 -297180 74120 -297130
rect 74120 -297180 74760 -297130
rect 75560 -297130 77760 -297080
rect 75560 -297180 77120 -297130
rect 77120 -297180 77760 -297130
rect 78560 -297130 80760 -297080
rect 78560 -297180 80120 -297130
rect 80120 -297180 80760 -297130
rect 81560 -297130 83760 -297080
rect 81560 -297180 83120 -297130
rect 83120 -297180 83760 -297130
rect 84560 -297130 86760 -297080
rect 84560 -297180 86120 -297130
rect 86120 -297180 86760 -297130
rect 87560 -297130 89760 -297080
rect 87560 -297180 89120 -297130
rect 89120 -297180 89760 -297130
rect 90560 -297130 92760 -297080
rect 90560 -297180 92120 -297130
rect 92120 -297180 92760 -297130
rect 93560 -297130 95760 -297080
rect 93560 -297180 95120 -297130
rect 95120 -297180 95760 -297130
rect 96560 -297130 98760 -297080
rect 96560 -297180 98120 -297130
rect 98120 -297180 98760 -297130
rect 99560 -297130 101760 -297080
rect 99560 -297180 101120 -297130
rect 101120 -297180 101760 -297130
rect 102560 -297130 104760 -297080
rect 102560 -297180 104120 -297130
rect 104120 -297180 104760 -297130
rect 105560 -297130 107760 -297080
rect 105560 -297180 107120 -297130
rect 107120 -297180 107760 -297130
rect 108560 -297130 110760 -297080
rect 108560 -297180 110120 -297130
rect 110120 -297180 110760 -297130
rect 111560 -297130 113760 -297080
rect 111560 -297180 113120 -297130
rect 113120 -297180 113760 -297130
rect 114560 -297130 116760 -297080
rect 114560 -297180 116120 -297130
rect 116120 -297180 116760 -297130
rect 117560 -297130 119760 -297080
rect 117560 -297180 119120 -297130
rect 119120 -297180 119760 -297130
rect 120560 -297130 122760 -297080
rect 120560 -297180 122120 -297130
rect 122120 -297180 122760 -297130
rect 123560 -297130 125760 -297080
rect 123560 -297180 125120 -297130
rect 125120 -297180 125760 -297130
rect 126560 -297130 128760 -297080
rect 126560 -297180 128120 -297130
rect 128120 -297180 128760 -297130
rect 129560 -297130 131760 -297080
rect 129560 -297180 131120 -297130
rect 131120 -297180 131760 -297130
rect 132560 -297130 134760 -297080
rect 132560 -297180 134120 -297130
rect 134120 -297180 134760 -297130
rect 135560 -297130 137760 -297080
rect 135560 -297180 137120 -297130
rect 137120 -297180 137760 -297130
rect 138560 -297130 140760 -297080
rect 138560 -297180 140120 -297130
rect 140120 -297180 140760 -297130
rect 141560 -297130 143760 -297080
rect 141560 -297180 143120 -297130
rect 143120 -297180 143760 -297130
rect 144560 -297130 146760 -297080
rect 144560 -297180 146120 -297130
rect 146120 -297180 146760 -297130
rect 147560 -297130 149760 -297080
rect 147560 -297180 149120 -297130
rect 149120 -297180 149760 -297130
rect 150560 -297130 152760 -297080
rect 150560 -297180 152120 -297130
rect 152120 -297180 152760 -297130
rect 153560 -297130 155760 -297080
rect 153560 -297180 155120 -297130
rect 155120 -297180 155760 -297130
rect 156560 -297130 158760 -297080
rect 156560 -297180 158120 -297130
rect 158120 -297180 158760 -297130
rect 159560 -297130 161760 -297080
rect 159560 -297180 161120 -297130
rect 161120 -297180 161760 -297130
rect 162560 -297130 164760 -297080
rect 162560 -297180 164120 -297130
rect 164120 -297180 164760 -297130
rect 165560 -297130 167760 -297080
rect 165560 -297180 167120 -297130
rect 167120 -297180 167760 -297130
rect 168560 -297130 170760 -297080
rect 168560 -297180 170120 -297130
rect 170120 -297180 170760 -297130
rect 171560 -297130 173760 -297080
rect 171560 -297180 173120 -297130
rect 173120 -297180 173760 -297130
rect 174560 -297130 176760 -297080
rect 174560 -297180 176120 -297130
rect 176120 -297180 176760 -297130
rect 177560 -297130 179760 -297080
rect 177560 -297180 179120 -297130
rect 179120 -297180 179760 -297130
rect 180560 -297130 182760 -297080
rect 180560 -297180 182120 -297130
rect 182120 -297180 182760 -297130
rect 183560 -297130 185760 -297080
rect 183560 -297180 185120 -297130
rect 185120 -297180 185760 -297130
rect 186560 -297130 188760 -297080
rect 186560 -297180 188120 -297130
rect 188120 -297180 188760 -297130
rect 189560 -297130 191760 -297080
rect 189560 -297180 191120 -297130
rect 191120 -297180 191760 -297130
rect 192560 -297130 194760 -297080
rect 192560 -297180 194120 -297130
rect 194120 -297180 194760 -297130
rect 195560 -297130 197760 -297080
rect 195560 -297180 197120 -297130
rect 197120 -297180 197760 -297130
rect 198560 -297130 200760 -297080
rect 198560 -297180 200120 -297130
rect 200120 -297180 200760 -297130
rect 201560 -297130 203760 -297080
rect 201560 -297180 203120 -297130
rect 203120 -297180 203760 -297130
rect 204560 -297130 206760 -297080
rect 204560 -297180 206120 -297130
rect 206120 -297180 206760 -297130
rect 207560 -297130 209760 -297080
rect 207560 -297180 209120 -297130
rect 209120 -297180 209760 -297130
rect 210560 -297130 212760 -297080
rect 210560 -297180 212120 -297130
rect 212120 -297180 212760 -297130
rect 213560 -297130 215760 -297080
rect 213560 -297180 215120 -297130
rect 215120 -297180 215760 -297130
rect 216560 -297130 218760 -297080
rect 216560 -297180 218120 -297130
rect 218120 -297180 218760 -297130
rect 219560 -297130 221760 -297080
rect 219560 -297180 221120 -297130
rect 221120 -297180 221760 -297130
rect 222560 -297130 224760 -297080
rect 222560 -297180 224120 -297130
rect 224120 -297180 224760 -297130
rect 225560 -297130 227760 -297080
rect 225560 -297180 227120 -297130
rect 227120 -297180 227760 -297130
rect 228560 -297130 230760 -297080
rect 228560 -297180 230120 -297130
rect 230120 -297180 230760 -297130
rect 231560 -297130 233760 -297080
rect 231560 -297180 233120 -297130
rect 233120 -297180 233760 -297130
rect 234560 -297130 236760 -297080
rect 234560 -297180 236120 -297130
rect 236120 -297180 236760 -297130
rect 237560 -297130 239760 -297080
rect 237560 -297180 239120 -297130
rect 239120 -297180 239760 -297130
rect 240560 -297130 242760 -297080
rect 240560 -297180 242120 -297130
rect 242120 -297180 242760 -297130
rect 243560 -297130 245760 -297080
rect 243560 -297180 245120 -297130
rect 245120 -297180 245760 -297130
rect 246560 -297130 248760 -297080
rect 246560 -297180 248120 -297130
rect 248120 -297180 248760 -297130
rect 249560 -297130 251760 -297080
rect 249560 -297180 251120 -297130
rect 251120 -297180 251760 -297130
rect 252560 -297130 254760 -297080
rect 252560 -297180 254120 -297130
rect 254120 -297180 254760 -297130
rect 255560 -297130 257760 -297080
rect 255560 -297180 257120 -297130
rect 257120 -297180 257760 -297130
rect 258560 -297130 260760 -297080
rect 258560 -297180 260120 -297130
rect 260120 -297180 260760 -297130
rect 261560 -297130 263760 -297080
rect 261560 -297180 263120 -297130
rect 263120 -297180 263760 -297130
rect 264560 -297130 266760 -297080
rect 264560 -297180 266120 -297130
rect 266120 -297180 266760 -297130
rect 267560 -297130 269760 -297080
rect 267560 -297180 269120 -297130
rect 269120 -297180 269760 -297130
rect 270560 -297130 272760 -297080
rect 270560 -297180 272120 -297130
rect 272120 -297180 272760 -297130
rect 273560 -297130 275760 -297080
rect 273560 -297180 275120 -297130
rect 275120 -297180 275760 -297130
rect 276560 -297130 278760 -297080
rect 276560 -297180 278120 -297130
rect 278120 -297180 278760 -297130
rect 279560 -297130 281760 -297080
rect 279560 -297180 281120 -297130
rect 281120 -297180 281760 -297130
rect 282560 -297130 284760 -297080
rect 282560 -297180 284120 -297130
rect 284120 -297180 284760 -297130
rect 285560 -297130 287760 -297080
rect 285560 -297180 287120 -297130
rect 287120 -297180 287760 -297130
rect 288560 -297130 290760 -297080
rect 288560 -297180 290120 -297130
rect 290120 -297180 290760 -297130
rect 291560 -297130 293760 -297080
rect 291560 -297180 293120 -297130
rect 293120 -297180 293760 -297130
rect 294560 -297130 296760 -297080
rect 294560 -297180 296120 -297130
rect 296120 -297180 296760 -297130
rect 297560 -297130 299760 -297080
rect 297560 -297180 299120 -297130
rect 299120 -297180 299760 -297130
rect 240 -297700 420 -297500
rect 3240 -297700 3420 -297500
rect 6240 -297700 6420 -297500
rect 9240 -297700 9420 -297500
rect 12240 -297700 12420 -297500
rect 15240 -297700 15420 -297500
rect 18240 -297700 18420 -297500
rect 21240 -297700 21420 -297500
rect 24240 -297700 24420 -297500
rect 27240 -297700 27420 -297500
rect 30240 -297700 30420 -297500
rect 33240 -297700 33420 -297500
rect 36240 -297700 36420 -297500
rect 39240 -297700 39420 -297500
rect 42240 -297700 42420 -297500
rect 45240 -297700 45420 -297500
rect 48240 -297700 48420 -297500
rect 51240 -297700 51420 -297500
rect 54240 -297700 54420 -297500
rect 57240 -297700 57420 -297500
rect 60240 -297700 60420 -297500
rect 63240 -297700 63420 -297500
rect 66240 -297700 66420 -297500
rect 69240 -297700 69420 -297500
rect 72240 -297700 72420 -297500
rect 75240 -297700 75420 -297500
rect 78240 -297700 78420 -297500
rect 81240 -297700 81420 -297500
rect 84240 -297700 84420 -297500
rect 87240 -297700 87420 -297500
rect 90240 -297700 90420 -297500
rect 93240 -297700 93420 -297500
rect 96240 -297700 96420 -297500
rect 99240 -297700 99420 -297500
rect 102240 -297700 102420 -297500
rect 105240 -297700 105420 -297500
rect 108240 -297700 108420 -297500
rect 111240 -297700 111420 -297500
rect 114240 -297700 114420 -297500
rect 117240 -297700 117420 -297500
rect 120240 -297700 120420 -297500
rect 123240 -297700 123420 -297500
rect 126240 -297700 126420 -297500
rect 129240 -297700 129420 -297500
rect 132240 -297700 132420 -297500
rect 135240 -297700 135420 -297500
rect 138240 -297700 138420 -297500
rect 141240 -297700 141420 -297500
rect 144240 -297700 144420 -297500
rect 147240 -297700 147420 -297500
rect 150240 -297700 150420 -297500
rect 153240 -297700 153420 -297500
rect 156240 -297700 156420 -297500
rect 159240 -297700 159420 -297500
rect 162240 -297700 162420 -297500
rect 165240 -297700 165420 -297500
rect 168240 -297700 168420 -297500
rect 171240 -297700 171420 -297500
rect 174240 -297700 174420 -297500
rect 177240 -297700 177420 -297500
rect 180240 -297700 180420 -297500
rect 183240 -297700 183420 -297500
rect 186240 -297700 186420 -297500
rect 189240 -297700 189420 -297500
rect 192240 -297700 192420 -297500
rect 195240 -297700 195420 -297500
rect 198240 -297700 198420 -297500
rect 201240 -297700 201420 -297500
rect 204240 -297700 204420 -297500
rect 207240 -297700 207420 -297500
rect 210240 -297700 210420 -297500
rect 213240 -297700 213420 -297500
rect 216240 -297700 216420 -297500
rect 219240 -297700 219420 -297500
rect 222240 -297700 222420 -297500
rect 225240 -297700 225420 -297500
rect 228240 -297700 228420 -297500
rect 231240 -297700 231420 -297500
rect 234240 -297700 234420 -297500
rect 237240 -297700 237420 -297500
rect 240240 -297700 240420 -297500
rect 243240 -297700 243420 -297500
rect 246240 -297700 246420 -297500
rect 249240 -297700 249420 -297500
rect 252240 -297700 252420 -297500
rect 255240 -297700 255420 -297500
rect 258240 -297700 258420 -297500
rect 261240 -297700 261420 -297500
rect 264240 -297700 264420 -297500
rect 267240 -297700 267420 -297500
rect 270240 -297700 270420 -297500
rect 273240 -297700 273420 -297500
rect 276240 -297700 276420 -297500
rect 279240 -297700 279420 -297500
rect 282240 -297700 282420 -297500
rect 285240 -297700 285420 -297500
rect 288240 -297700 288420 -297500
rect 291240 -297700 291420 -297500
rect 294240 -297700 294420 -297500
rect 297240 -297700 297420 -297500
<< metal3 >>
rect -1200 2840 -1110 5000
rect 480 3650 590 3660
rect 480 3560 490 3650
rect 580 3560 590 3650
rect 480 3550 590 3560
rect 3480 3650 3590 3660
rect 3480 3560 3490 3650
rect 3580 3560 3590 3650
rect 3480 3550 3590 3560
rect 6480 3650 6590 3660
rect 6480 3560 6490 3650
rect 6580 3560 6590 3650
rect 6480 3550 6590 3560
rect 9480 3650 9590 3660
rect 9480 3560 9490 3650
rect 9580 3560 9590 3650
rect 9480 3550 9590 3560
rect 12480 3650 12590 3660
rect 12480 3560 12490 3650
rect 12580 3560 12590 3650
rect 12480 3550 12590 3560
rect 15480 3650 15590 3660
rect 15480 3560 15490 3650
rect 15580 3560 15590 3650
rect 15480 3550 15590 3560
rect 18480 3650 18590 3660
rect 18480 3560 18490 3650
rect 18580 3560 18590 3650
rect 18480 3550 18590 3560
rect 21480 3650 21590 3660
rect 21480 3560 21490 3650
rect 21580 3560 21590 3650
rect 21480 3550 21590 3560
rect 24480 3650 24590 3660
rect 24480 3560 24490 3650
rect 24580 3560 24590 3650
rect 24480 3550 24590 3560
rect 27480 3650 27590 3660
rect 27480 3560 27490 3650
rect 27580 3560 27590 3650
rect 27480 3550 27590 3560
rect 30480 3650 30590 3660
rect 30480 3560 30490 3650
rect 30580 3560 30590 3650
rect 30480 3550 30590 3560
rect 33480 3650 33590 3660
rect 33480 3560 33490 3650
rect 33580 3560 33590 3650
rect 33480 3550 33590 3560
rect 36480 3650 36590 3660
rect 36480 3560 36490 3650
rect 36580 3560 36590 3650
rect 36480 3550 36590 3560
rect 39480 3650 39590 3660
rect 39480 3560 39490 3650
rect 39580 3560 39590 3650
rect 39480 3550 39590 3560
rect 42480 3650 42590 3660
rect 42480 3560 42490 3650
rect 42580 3560 42590 3650
rect 42480 3550 42590 3560
rect 45480 3650 45590 3660
rect 45480 3560 45490 3650
rect 45580 3560 45590 3650
rect 45480 3550 45590 3560
rect 48480 3650 48590 3660
rect 48480 3560 48490 3650
rect 48580 3560 48590 3650
rect 48480 3550 48590 3560
rect 51480 3650 51590 3660
rect 51480 3560 51490 3650
rect 51580 3560 51590 3650
rect 51480 3550 51590 3560
rect 54480 3650 54590 3660
rect 54480 3560 54490 3650
rect 54580 3560 54590 3650
rect 54480 3550 54590 3560
rect 57480 3650 57590 3660
rect 57480 3560 57490 3650
rect 57580 3560 57590 3650
rect 57480 3550 57590 3560
rect 60480 3650 60590 3660
rect 60480 3560 60490 3650
rect 60580 3560 60590 3650
rect 60480 3550 60590 3560
rect 63480 3650 63590 3660
rect 63480 3560 63490 3650
rect 63580 3560 63590 3650
rect 63480 3550 63590 3560
rect 66480 3650 66590 3660
rect 66480 3560 66490 3650
rect 66580 3560 66590 3650
rect 66480 3550 66590 3560
rect 69480 3650 69590 3660
rect 69480 3560 69490 3650
rect 69580 3560 69590 3650
rect 69480 3550 69590 3560
rect 72480 3650 72590 3660
rect 72480 3560 72490 3650
rect 72580 3560 72590 3650
rect 72480 3550 72590 3560
rect 75480 3650 75590 3660
rect 75480 3560 75490 3650
rect 75580 3560 75590 3650
rect 75480 3550 75590 3560
rect 78480 3650 78590 3660
rect 78480 3560 78490 3650
rect 78580 3560 78590 3650
rect 78480 3550 78590 3560
rect 81480 3650 81590 3660
rect 81480 3560 81490 3650
rect 81580 3560 81590 3650
rect 81480 3550 81590 3560
rect 84480 3650 84590 3660
rect 84480 3560 84490 3650
rect 84580 3560 84590 3650
rect 84480 3550 84590 3560
rect 87480 3650 87590 3660
rect 87480 3560 87490 3650
rect 87580 3560 87590 3650
rect 87480 3550 87590 3560
rect 90480 3650 90590 3660
rect 90480 3560 90490 3650
rect 90580 3560 90590 3650
rect 90480 3550 90590 3560
rect 93480 3650 93590 3660
rect 93480 3560 93490 3650
rect 93580 3560 93590 3650
rect 93480 3550 93590 3560
rect 96480 3650 96590 3660
rect 96480 3560 96490 3650
rect 96580 3560 96590 3650
rect 96480 3550 96590 3560
rect 99480 3650 99590 3660
rect 99480 3560 99490 3650
rect 99580 3560 99590 3650
rect 99480 3550 99590 3560
rect 102480 3650 102590 3660
rect 102480 3560 102490 3650
rect 102580 3560 102590 3650
rect 102480 3550 102590 3560
rect 105480 3650 105590 3660
rect 105480 3560 105490 3650
rect 105580 3560 105590 3650
rect 105480 3550 105590 3560
rect 108480 3650 108590 3660
rect 108480 3560 108490 3650
rect 108580 3560 108590 3650
rect 108480 3550 108590 3560
rect 111480 3650 111590 3660
rect 111480 3560 111490 3650
rect 111580 3560 111590 3650
rect 111480 3550 111590 3560
rect 114480 3650 114590 3660
rect 114480 3560 114490 3650
rect 114580 3560 114590 3650
rect 114480 3550 114590 3560
rect 117480 3650 117590 3660
rect 117480 3560 117490 3650
rect 117580 3560 117590 3650
rect 117480 3550 117590 3560
rect 120480 3650 120590 3660
rect 120480 3560 120490 3650
rect 120580 3560 120590 3650
rect 120480 3550 120590 3560
rect 123480 3650 123590 3660
rect 123480 3560 123490 3650
rect 123580 3560 123590 3650
rect 123480 3550 123590 3560
rect 126480 3650 126590 3660
rect 126480 3560 126490 3650
rect 126580 3560 126590 3650
rect 126480 3550 126590 3560
rect 129480 3650 129590 3660
rect 129480 3560 129490 3650
rect 129580 3560 129590 3650
rect 129480 3550 129590 3560
rect 132480 3650 132590 3660
rect 132480 3560 132490 3650
rect 132580 3560 132590 3650
rect 132480 3550 132590 3560
rect 135480 3650 135590 3660
rect 135480 3560 135490 3650
rect 135580 3560 135590 3650
rect 135480 3550 135590 3560
rect 138480 3650 138590 3660
rect 138480 3560 138490 3650
rect 138580 3560 138590 3650
rect 138480 3550 138590 3560
rect 141480 3650 141590 3660
rect 141480 3560 141490 3650
rect 141580 3560 141590 3650
rect 141480 3550 141590 3560
rect 144480 3650 144590 3660
rect 144480 3560 144490 3650
rect 144580 3560 144590 3650
rect 144480 3550 144590 3560
rect 147480 3650 147590 3660
rect 147480 3560 147490 3650
rect 147580 3560 147590 3650
rect 147480 3550 147590 3560
rect 150480 3650 150590 3660
rect 150480 3560 150490 3650
rect 150580 3560 150590 3650
rect 150480 3550 150590 3560
rect 153480 3650 153590 3660
rect 153480 3560 153490 3650
rect 153580 3560 153590 3650
rect 153480 3550 153590 3560
rect 156480 3650 156590 3660
rect 156480 3560 156490 3650
rect 156580 3560 156590 3650
rect 156480 3550 156590 3560
rect 159480 3650 159590 3660
rect 159480 3560 159490 3650
rect 159580 3560 159590 3650
rect 159480 3550 159590 3560
rect 162480 3650 162590 3660
rect 162480 3560 162490 3650
rect 162580 3560 162590 3650
rect 162480 3550 162590 3560
rect 165480 3650 165590 3660
rect 165480 3560 165490 3650
rect 165580 3560 165590 3650
rect 165480 3550 165590 3560
rect 168480 3650 168590 3660
rect 168480 3560 168490 3650
rect 168580 3560 168590 3650
rect 168480 3550 168590 3560
rect 171480 3650 171590 3660
rect 171480 3560 171490 3650
rect 171580 3560 171590 3650
rect 171480 3550 171590 3560
rect 174480 3650 174590 3660
rect 174480 3560 174490 3650
rect 174580 3560 174590 3650
rect 174480 3550 174590 3560
rect 177480 3650 177590 3660
rect 177480 3560 177490 3650
rect 177580 3560 177590 3650
rect 177480 3550 177590 3560
rect 180480 3650 180590 3660
rect 180480 3560 180490 3650
rect 180580 3560 180590 3650
rect 180480 3550 180590 3560
rect 183480 3650 183590 3660
rect 183480 3560 183490 3650
rect 183580 3560 183590 3650
rect 183480 3550 183590 3560
rect 186480 3650 186590 3660
rect 186480 3560 186490 3650
rect 186580 3560 186590 3650
rect 186480 3550 186590 3560
rect 189480 3650 189590 3660
rect 189480 3560 189490 3650
rect 189580 3560 189590 3650
rect 189480 3550 189590 3560
rect 192480 3650 192590 3660
rect 192480 3560 192490 3650
rect 192580 3560 192590 3650
rect 192480 3550 192590 3560
rect 195480 3650 195590 3660
rect 195480 3560 195490 3650
rect 195580 3560 195590 3650
rect 195480 3550 195590 3560
rect 198480 3650 198590 3660
rect 198480 3560 198490 3650
rect 198580 3560 198590 3650
rect 198480 3550 198590 3560
rect 201480 3650 201590 3660
rect 201480 3560 201490 3650
rect 201580 3560 201590 3650
rect 201480 3550 201590 3560
rect 204480 3650 204590 3660
rect 204480 3560 204490 3650
rect 204580 3560 204590 3650
rect 204480 3550 204590 3560
rect 207480 3650 207590 3660
rect 207480 3560 207490 3650
rect 207580 3560 207590 3650
rect 207480 3550 207590 3560
rect 210480 3650 210590 3660
rect 210480 3560 210490 3650
rect 210580 3560 210590 3650
rect 210480 3550 210590 3560
rect 213480 3650 213590 3660
rect 213480 3560 213490 3650
rect 213580 3560 213590 3650
rect 213480 3550 213590 3560
rect 216480 3650 216590 3660
rect 216480 3560 216490 3650
rect 216580 3560 216590 3650
rect 216480 3550 216590 3560
rect 219480 3650 219590 3660
rect 219480 3560 219490 3650
rect 219580 3560 219590 3650
rect 219480 3550 219590 3560
rect 222480 3650 222590 3660
rect 222480 3560 222490 3650
rect 222580 3560 222590 3650
rect 222480 3550 222590 3560
rect 225480 3650 225590 3660
rect 225480 3560 225490 3650
rect 225580 3560 225590 3650
rect 225480 3550 225590 3560
rect 228480 3650 228590 3660
rect 228480 3560 228490 3650
rect 228580 3560 228590 3650
rect 228480 3550 228590 3560
rect 231480 3650 231590 3660
rect 231480 3560 231490 3650
rect 231580 3560 231590 3650
rect 231480 3550 231590 3560
rect 234480 3650 234590 3660
rect 234480 3560 234490 3650
rect 234580 3560 234590 3650
rect 234480 3550 234590 3560
rect 237480 3650 237590 3660
rect 237480 3560 237490 3650
rect 237580 3560 237590 3650
rect 237480 3550 237590 3560
rect 240480 3650 240590 3660
rect 240480 3560 240490 3650
rect 240580 3560 240590 3650
rect 240480 3550 240590 3560
rect 243480 3650 243590 3660
rect 243480 3560 243490 3650
rect 243580 3560 243590 3650
rect 243480 3550 243590 3560
rect 246480 3650 246590 3660
rect 246480 3560 246490 3650
rect 246580 3560 246590 3650
rect 246480 3550 246590 3560
rect 249480 3650 249590 3660
rect 249480 3560 249490 3650
rect 249580 3560 249590 3650
rect 249480 3550 249590 3560
rect 252480 3650 252590 3660
rect 252480 3560 252490 3650
rect 252580 3560 252590 3650
rect 252480 3550 252590 3560
rect 255480 3650 255590 3660
rect 255480 3560 255490 3650
rect 255580 3560 255590 3650
rect 255480 3550 255590 3560
rect 258480 3650 258590 3660
rect 258480 3560 258490 3650
rect 258580 3560 258590 3650
rect 258480 3550 258590 3560
rect 261480 3650 261590 3660
rect 261480 3560 261490 3650
rect 261580 3560 261590 3650
rect 261480 3550 261590 3560
rect 264480 3650 264590 3660
rect 264480 3560 264490 3650
rect 264580 3560 264590 3650
rect 264480 3550 264590 3560
rect 267480 3650 267590 3660
rect 267480 3560 267490 3650
rect 267580 3560 267590 3650
rect 267480 3550 267590 3560
rect 270480 3650 270590 3660
rect 270480 3560 270490 3650
rect 270580 3560 270590 3650
rect 270480 3550 270590 3560
rect 273480 3650 273590 3660
rect 273480 3560 273490 3650
rect 273580 3560 273590 3650
rect 273480 3550 273590 3560
rect 276480 3650 276590 3660
rect 276480 3560 276490 3650
rect 276580 3560 276590 3650
rect 276480 3550 276590 3560
rect 279480 3650 279590 3660
rect 279480 3560 279490 3650
rect 279580 3560 279590 3650
rect 279480 3550 279590 3560
rect 282480 3650 282590 3660
rect 282480 3560 282490 3650
rect 282580 3560 282590 3650
rect 282480 3550 282590 3560
rect 285480 3650 285590 3660
rect 285480 3560 285490 3650
rect 285580 3560 285590 3650
rect 285480 3550 285590 3560
rect 288480 3650 288590 3660
rect 288480 3560 288490 3650
rect 288580 3560 288590 3650
rect 288480 3550 288590 3560
rect 291480 3650 291590 3660
rect 291480 3560 291490 3650
rect 291580 3560 291590 3650
rect 291480 3550 291590 3560
rect 294480 3650 294590 3660
rect 294480 3560 294490 3650
rect 294580 3560 294590 3650
rect 294480 3550 294590 3560
rect 297480 3650 297590 3660
rect 297480 3560 297490 3650
rect 297580 3560 297590 3650
rect 297480 3550 297590 3560
rect -1200 2750 200 2840
rect -1200 -160 -1110 2750
rect -480 2550 -370 2560
rect -480 2540 520 2550
rect -480 2470 -470 2540
rect -380 2470 520 2540
rect -480 2460 520 2470
rect -480 2450 -370 2460
rect -560 1560 440 1570
rect -560 1490 -540 1560
rect -260 1490 440 1560
rect -560 1480 440 1490
rect -760 230 40 250
rect -760 160 -740 230
rect -650 160 40 230
rect -750 140 -640 160
rect -1200 -250 200 -160
rect -1200 -3160 -1110 -250
rect -480 -450 -370 -440
rect -480 -460 520 -450
rect -480 -530 -470 -460
rect -380 -530 520 -460
rect -480 -540 520 -530
rect -480 -550 -370 -540
rect -560 -1440 440 -1430
rect -560 -1510 -540 -1440
rect -260 -1510 440 -1440
rect -560 -1520 440 -1510
rect -760 -2770 40 -2750
rect -760 -2840 -740 -2770
rect -650 -2840 40 -2770
rect -750 -2860 -640 -2840
rect -1200 -3250 200 -3160
rect -1200 -6160 -1110 -3250
rect -480 -3450 -370 -3440
rect -480 -3460 520 -3450
rect -480 -3530 -470 -3460
rect -380 -3530 520 -3460
rect -480 -3540 520 -3530
rect -480 -3550 -370 -3540
rect -560 -4440 440 -4430
rect -560 -4510 -540 -4440
rect -260 -4510 440 -4440
rect -560 -4520 440 -4510
rect -760 -5770 40 -5750
rect -760 -5840 -740 -5770
rect -650 -5840 40 -5770
rect -750 -5860 -640 -5840
rect -1200 -6250 200 -6160
rect -1200 -9160 -1110 -6250
rect -480 -6450 -370 -6440
rect -480 -6460 520 -6450
rect -480 -6530 -470 -6460
rect -380 -6530 520 -6460
rect -480 -6540 520 -6530
rect -480 -6550 -370 -6540
rect -560 -7440 440 -7430
rect -560 -7510 -540 -7440
rect -260 -7510 440 -7440
rect -560 -7520 440 -7510
rect -760 -8770 40 -8750
rect -760 -8840 -740 -8770
rect -650 -8840 40 -8770
rect -750 -8860 -640 -8840
rect -1200 -9250 200 -9160
rect -1200 -12160 -1110 -9250
rect -480 -9450 -370 -9440
rect -480 -9460 520 -9450
rect -480 -9530 -470 -9460
rect -380 -9530 520 -9460
rect -480 -9540 520 -9530
rect -480 -9550 -370 -9540
rect -560 -10440 440 -10430
rect -560 -10510 -540 -10440
rect -260 -10510 440 -10440
rect -560 -10520 440 -10510
rect -760 -11770 40 -11750
rect -760 -11840 -740 -11770
rect -650 -11840 40 -11770
rect -750 -11860 -640 -11840
rect -1200 -12250 200 -12160
rect -1200 -15160 -1110 -12250
rect -480 -12450 -370 -12440
rect -480 -12460 520 -12450
rect -480 -12530 -470 -12460
rect -380 -12530 520 -12460
rect -480 -12540 520 -12530
rect -480 -12550 -370 -12540
rect -560 -13440 440 -13430
rect -560 -13510 -540 -13440
rect -260 -13510 440 -13440
rect -560 -13520 440 -13510
rect -760 -14770 40 -14750
rect -760 -14840 -740 -14770
rect -650 -14840 40 -14770
rect -750 -14860 -640 -14840
rect -1200 -15250 200 -15160
rect -1200 -18160 -1110 -15250
rect -480 -15450 -370 -15440
rect -480 -15460 520 -15450
rect -480 -15530 -470 -15460
rect -380 -15530 520 -15460
rect -480 -15540 520 -15530
rect -480 -15550 -370 -15540
rect -560 -16440 440 -16430
rect -560 -16510 -540 -16440
rect -260 -16510 440 -16440
rect -560 -16520 440 -16510
rect -760 -17770 40 -17750
rect -760 -17840 -740 -17770
rect -650 -17840 40 -17770
rect -750 -17860 -640 -17840
rect -1200 -18250 200 -18160
rect -1200 -21160 -1110 -18250
rect -480 -18450 -370 -18440
rect -480 -18460 520 -18450
rect -480 -18530 -470 -18460
rect -380 -18530 520 -18460
rect -480 -18540 520 -18530
rect -480 -18550 -370 -18540
rect -560 -19440 440 -19430
rect -560 -19510 -540 -19440
rect -260 -19510 440 -19440
rect -560 -19520 440 -19510
rect -760 -20770 40 -20750
rect -760 -20840 -740 -20770
rect -650 -20840 40 -20770
rect -750 -20860 -640 -20840
rect -1200 -21250 200 -21160
rect -1200 -24160 -1110 -21250
rect -480 -21450 -370 -21440
rect -480 -21460 520 -21450
rect -480 -21530 -470 -21460
rect -380 -21530 520 -21460
rect -480 -21540 520 -21530
rect -480 -21550 -370 -21540
rect -560 -22440 440 -22430
rect -560 -22510 -540 -22440
rect -260 -22510 440 -22440
rect -560 -22520 440 -22510
rect -760 -23770 40 -23750
rect -760 -23840 -740 -23770
rect -650 -23840 40 -23770
rect -750 -23860 -640 -23840
rect -1200 -24250 200 -24160
rect -1200 -27160 -1110 -24250
rect -480 -24450 -370 -24440
rect -480 -24460 520 -24450
rect -480 -24530 -470 -24460
rect -380 -24530 520 -24460
rect -480 -24540 520 -24530
rect -480 -24550 -370 -24540
rect -560 -25440 440 -25430
rect -560 -25510 -540 -25440
rect -260 -25510 440 -25440
rect -560 -25520 440 -25510
rect -760 -26770 40 -26750
rect -760 -26840 -740 -26770
rect -650 -26840 40 -26770
rect -750 -26860 -640 -26840
rect -1200 -27250 200 -27160
rect -1200 -30160 -1110 -27250
rect -480 -27450 -370 -27440
rect -480 -27460 520 -27450
rect -480 -27530 -470 -27460
rect -380 -27530 520 -27460
rect -480 -27540 520 -27530
rect -480 -27550 -370 -27540
rect -560 -28440 440 -28430
rect -560 -28510 -540 -28440
rect -260 -28510 440 -28440
rect -560 -28520 440 -28510
rect -760 -29770 40 -29750
rect -760 -29840 -740 -29770
rect -650 -29840 40 -29770
rect -750 -29860 -640 -29840
rect -1200 -30250 200 -30160
rect -1200 -33160 -1110 -30250
rect -480 -30450 -370 -30440
rect -480 -30460 520 -30450
rect -480 -30530 -470 -30460
rect -380 -30530 520 -30460
rect -480 -30540 520 -30530
rect -480 -30550 -370 -30540
rect -560 -31440 440 -31430
rect -560 -31510 -540 -31440
rect -260 -31510 440 -31440
rect -560 -31520 440 -31510
rect -760 -32770 40 -32750
rect -760 -32840 -740 -32770
rect -650 -32840 40 -32770
rect -750 -32860 -640 -32840
rect -1200 -33250 200 -33160
rect -1200 -36160 -1110 -33250
rect -480 -33450 -370 -33440
rect -480 -33460 520 -33450
rect -480 -33530 -470 -33460
rect -380 -33530 520 -33460
rect -480 -33540 520 -33530
rect -480 -33550 -370 -33540
rect -560 -34440 440 -34430
rect -560 -34510 -540 -34440
rect -260 -34510 440 -34440
rect -560 -34520 440 -34510
rect -760 -35770 40 -35750
rect -760 -35840 -740 -35770
rect -650 -35840 40 -35770
rect -750 -35860 -640 -35840
rect -1200 -36250 200 -36160
rect -1200 -39160 -1110 -36250
rect -480 -36450 -370 -36440
rect -480 -36460 520 -36450
rect -480 -36530 -470 -36460
rect -380 -36530 520 -36460
rect -480 -36540 520 -36530
rect -480 -36550 -370 -36540
rect -560 -37440 440 -37430
rect -560 -37510 -540 -37440
rect -260 -37510 440 -37440
rect -560 -37520 440 -37510
rect -760 -38770 40 -38750
rect -760 -38840 -740 -38770
rect -650 -38840 40 -38770
rect -750 -38860 -640 -38840
rect -1200 -39250 200 -39160
rect -1200 -42160 -1110 -39250
rect -480 -39450 -370 -39440
rect -480 -39460 520 -39450
rect -480 -39530 -470 -39460
rect -380 -39530 520 -39460
rect -480 -39540 520 -39530
rect -480 -39550 -370 -39540
rect -560 -40440 440 -40430
rect -560 -40510 -540 -40440
rect -260 -40510 440 -40440
rect -560 -40520 440 -40510
rect -760 -41770 40 -41750
rect -760 -41840 -740 -41770
rect -650 -41840 40 -41770
rect -750 -41860 -640 -41840
rect -1200 -42250 200 -42160
rect -1200 -45160 -1110 -42250
rect -480 -42450 -370 -42440
rect -480 -42460 520 -42450
rect -480 -42530 -470 -42460
rect -380 -42530 520 -42460
rect -480 -42540 520 -42530
rect -480 -42550 -370 -42540
rect -560 -43440 440 -43430
rect -560 -43510 -540 -43440
rect -260 -43510 440 -43440
rect -560 -43520 440 -43510
rect -760 -44770 40 -44750
rect -760 -44840 -740 -44770
rect -650 -44840 40 -44770
rect -750 -44860 -640 -44840
rect -1200 -45250 200 -45160
rect -1200 -48160 -1110 -45250
rect -480 -45450 -370 -45440
rect -480 -45460 520 -45450
rect -480 -45530 -470 -45460
rect -380 -45530 520 -45460
rect -480 -45540 520 -45530
rect -480 -45550 -370 -45540
rect -560 -46440 440 -46430
rect -560 -46510 -540 -46440
rect -260 -46510 440 -46440
rect -560 -46520 440 -46510
rect -760 -47770 40 -47750
rect -760 -47840 -740 -47770
rect -650 -47840 40 -47770
rect -750 -47860 -640 -47840
rect -1200 -48250 200 -48160
rect -1200 -51160 -1110 -48250
rect -480 -48450 -370 -48440
rect -480 -48460 520 -48450
rect -480 -48530 -470 -48460
rect -380 -48530 520 -48460
rect -480 -48540 520 -48530
rect -480 -48550 -370 -48540
rect -560 -49440 440 -49430
rect -560 -49510 -540 -49440
rect -260 -49510 440 -49440
rect -560 -49520 440 -49510
rect -760 -50770 40 -50750
rect -760 -50840 -740 -50770
rect -650 -50840 40 -50770
rect -750 -50860 -640 -50840
rect -1200 -51250 200 -51160
rect -1200 -54160 -1110 -51250
rect -480 -51450 -370 -51440
rect -480 -51460 520 -51450
rect -480 -51530 -470 -51460
rect -380 -51530 520 -51460
rect -480 -51540 520 -51530
rect -480 -51550 -370 -51540
rect -560 -52440 440 -52430
rect -560 -52510 -540 -52440
rect -260 -52510 440 -52440
rect -560 -52520 440 -52510
rect -760 -53770 40 -53750
rect -760 -53840 -740 -53770
rect -650 -53840 40 -53770
rect -750 -53860 -640 -53840
rect -1200 -54250 200 -54160
rect -1200 -57160 -1110 -54250
rect -480 -54450 -370 -54440
rect -480 -54460 520 -54450
rect -480 -54530 -470 -54460
rect -380 -54530 520 -54460
rect -480 -54540 520 -54530
rect -480 -54550 -370 -54540
rect -560 -55440 440 -55430
rect -560 -55510 -540 -55440
rect -260 -55510 440 -55440
rect -560 -55520 440 -55510
rect -760 -56770 40 -56750
rect -760 -56840 -740 -56770
rect -650 -56840 40 -56770
rect -750 -56860 -640 -56840
rect -1200 -57250 200 -57160
rect -1200 -60160 -1110 -57250
rect -480 -57450 -370 -57440
rect -480 -57460 520 -57450
rect -480 -57530 -470 -57460
rect -380 -57530 520 -57460
rect -480 -57540 520 -57530
rect -480 -57550 -370 -57540
rect -560 -58440 440 -58430
rect -560 -58510 -540 -58440
rect -260 -58510 440 -58440
rect -560 -58520 440 -58510
rect -760 -59770 40 -59750
rect -760 -59840 -740 -59770
rect -650 -59840 40 -59770
rect -750 -59860 -640 -59840
rect -1200 -60250 200 -60160
rect -1200 -63160 -1110 -60250
rect -480 -60450 -370 -60440
rect -480 -60460 520 -60450
rect -480 -60530 -470 -60460
rect -380 -60530 520 -60460
rect -480 -60540 520 -60530
rect -480 -60550 -370 -60540
rect -560 -61440 440 -61430
rect -560 -61510 -540 -61440
rect -260 -61510 440 -61440
rect -560 -61520 440 -61510
rect -760 -62770 40 -62750
rect -760 -62840 -740 -62770
rect -650 -62840 40 -62770
rect -750 -62860 -640 -62840
rect -1200 -63250 200 -63160
rect -1200 -66160 -1110 -63250
rect -480 -63450 -370 -63440
rect -480 -63460 520 -63450
rect -480 -63530 -470 -63460
rect -380 -63530 520 -63460
rect -480 -63540 520 -63530
rect -480 -63550 -370 -63540
rect -560 -64440 440 -64430
rect -560 -64510 -540 -64440
rect -260 -64510 440 -64440
rect -560 -64520 440 -64510
rect -760 -65770 40 -65750
rect -760 -65840 -740 -65770
rect -650 -65840 40 -65770
rect -750 -65860 -640 -65840
rect -1200 -66250 200 -66160
rect -1200 -69160 -1110 -66250
rect -480 -66450 -370 -66440
rect -480 -66460 520 -66450
rect -480 -66530 -470 -66460
rect -380 -66530 520 -66460
rect -480 -66540 520 -66530
rect -480 -66550 -370 -66540
rect -560 -67440 440 -67430
rect -560 -67510 -540 -67440
rect -260 -67510 440 -67440
rect -560 -67520 440 -67510
rect -760 -68770 40 -68750
rect -760 -68840 -740 -68770
rect -650 -68840 40 -68770
rect -750 -68860 -640 -68840
rect -1200 -69250 200 -69160
rect -1200 -72160 -1110 -69250
rect -480 -69450 -370 -69440
rect -480 -69460 520 -69450
rect -480 -69530 -470 -69460
rect -380 -69530 520 -69460
rect -480 -69540 520 -69530
rect -480 -69550 -370 -69540
rect -560 -70440 440 -70430
rect -560 -70510 -540 -70440
rect -260 -70510 440 -70440
rect -560 -70520 440 -70510
rect -760 -71770 40 -71750
rect -760 -71840 -740 -71770
rect -650 -71840 40 -71770
rect -750 -71860 -640 -71840
rect -1200 -72250 200 -72160
rect -1200 -75160 -1110 -72250
rect -480 -72450 -370 -72440
rect -480 -72460 520 -72450
rect -480 -72530 -470 -72460
rect -380 -72530 520 -72460
rect -480 -72540 520 -72530
rect -480 -72550 -370 -72540
rect -560 -73440 440 -73430
rect -560 -73510 -540 -73440
rect -260 -73510 440 -73440
rect -560 -73520 440 -73510
rect -760 -74770 40 -74750
rect -760 -74840 -740 -74770
rect -650 -74840 40 -74770
rect -750 -74860 -640 -74840
rect -1200 -75250 200 -75160
rect -1200 -78160 -1110 -75250
rect -480 -75450 -370 -75440
rect -480 -75460 520 -75450
rect -480 -75530 -470 -75460
rect -380 -75530 520 -75460
rect -480 -75540 520 -75530
rect -480 -75550 -370 -75540
rect -560 -76440 440 -76430
rect -560 -76510 -540 -76440
rect -260 -76510 440 -76440
rect -560 -76520 440 -76510
rect -760 -77770 40 -77750
rect -760 -77840 -740 -77770
rect -650 -77840 40 -77770
rect -750 -77860 -640 -77840
rect -1200 -78250 200 -78160
rect -1200 -81160 -1110 -78250
rect -480 -78450 -370 -78440
rect -480 -78460 520 -78450
rect -480 -78530 -470 -78460
rect -380 -78530 520 -78460
rect -480 -78540 520 -78530
rect -480 -78550 -370 -78540
rect -560 -79440 440 -79430
rect -560 -79510 -540 -79440
rect -260 -79510 440 -79440
rect -560 -79520 440 -79510
rect -760 -80770 40 -80750
rect -760 -80840 -740 -80770
rect -650 -80840 40 -80770
rect -750 -80860 -640 -80840
rect -1200 -81250 200 -81160
rect -1200 -84160 -1110 -81250
rect -480 -81450 -370 -81440
rect -480 -81460 520 -81450
rect -480 -81530 -470 -81460
rect -380 -81530 520 -81460
rect -480 -81540 520 -81530
rect -480 -81550 -370 -81540
rect -560 -82440 440 -82430
rect -560 -82510 -540 -82440
rect -260 -82510 440 -82440
rect -560 -82520 440 -82510
rect -760 -83770 40 -83750
rect -760 -83840 -740 -83770
rect -650 -83840 40 -83770
rect -750 -83860 -640 -83840
rect -1200 -84250 200 -84160
rect -1200 -87160 -1110 -84250
rect -480 -84450 -370 -84440
rect -480 -84460 520 -84450
rect -480 -84530 -470 -84460
rect -380 -84530 520 -84460
rect -480 -84540 520 -84530
rect -480 -84550 -370 -84540
rect -560 -85440 440 -85430
rect -560 -85510 -540 -85440
rect -260 -85510 440 -85440
rect -560 -85520 440 -85510
rect -760 -86770 40 -86750
rect -760 -86840 -740 -86770
rect -650 -86840 40 -86770
rect -750 -86860 -640 -86840
rect -1200 -87250 200 -87160
rect -1200 -90160 -1110 -87250
rect -480 -87450 -370 -87440
rect -480 -87460 520 -87450
rect -480 -87530 -470 -87460
rect -380 -87530 520 -87460
rect -480 -87540 520 -87530
rect -480 -87550 -370 -87540
rect -560 -88440 440 -88430
rect -560 -88510 -540 -88440
rect -260 -88510 440 -88440
rect -560 -88520 440 -88510
rect -760 -89770 40 -89750
rect -760 -89840 -740 -89770
rect -650 -89840 40 -89770
rect -750 -89860 -640 -89840
rect -1200 -90250 200 -90160
rect -1200 -93160 -1110 -90250
rect -480 -90450 -370 -90440
rect -480 -90460 520 -90450
rect -480 -90530 -470 -90460
rect -380 -90530 520 -90460
rect -480 -90540 520 -90530
rect -480 -90550 -370 -90540
rect -560 -91440 440 -91430
rect -560 -91510 -540 -91440
rect -260 -91510 440 -91440
rect -560 -91520 440 -91510
rect -760 -92770 40 -92750
rect -760 -92840 -740 -92770
rect -650 -92840 40 -92770
rect -750 -92860 -640 -92840
rect -1200 -93250 200 -93160
rect -1200 -96160 -1110 -93250
rect -480 -93450 -370 -93440
rect -480 -93460 520 -93450
rect -480 -93530 -470 -93460
rect -380 -93530 520 -93460
rect -480 -93540 520 -93530
rect -480 -93550 -370 -93540
rect -560 -94440 440 -94430
rect -560 -94510 -540 -94440
rect -260 -94510 440 -94440
rect -560 -94520 440 -94510
rect -760 -95770 40 -95750
rect -760 -95840 -740 -95770
rect -650 -95840 40 -95770
rect -750 -95860 -640 -95840
rect -1200 -96250 200 -96160
rect -1200 -99160 -1110 -96250
rect -480 -96450 -370 -96440
rect -480 -96460 520 -96450
rect -480 -96530 -470 -96460
rect -380 -96530 520 -96460
rect -480 -96540 520 -96530
rect -480 -96550 -370 -96540
rect -560 -97440 440 -97430
rect -560 -97510 -540 -97440
rect -260 -97510 440 -97440
rect -560 -97520 440 -97510
rect -760 -98770 40 -98750
rect -760 -98840 -740 -98770
rect -650 -98840 40 -98770
rect -750 -98860 -640 -98840
rect -1200 -99250 200 -99160
rect -1200 -102160 -1110 -99250
rect -480 -99450 -370 -99440
rect -480 -99460 520 -99450
rect -480 -99530 -470 -99460
rect -380 -99530 520 -99460
rect -480 -99540 520 -99530
rect -480 -99550 -370 -99540
rect -560 -100440 440 -100430
rect -560 -100510 -540 -100440
rect -260 -100510 440 -100440
rect -560 -100520 440 -100510
rect -760 -101770 40 -101750
rect -760 -101840 -740 -101770
rect -650 -101840 40 -101770
rect -750 -101860 -640 -101840
rect -1200 -102250 200 -102160
rect -1200 -105160 -1110 -102250
rect -480 -102450 -370 -102440
rect -480 -102460 520 -102450
rect -480 -102530 -470 -102460
rect -380 -102530 520 -102460
rect -480 -102540 520 -102530
rect -480 -102550 -370 -102540
rect -560 -103440 440 -103430
rect -560 -103510 -540 -103440
rect -260 -103510 440 -103440
rect -560 -103520 440 -103510
rect -760 -104770 40 -104750
rect -760 -104840 -740 -104770
rect -650 -104840 40 -104770
rect -750 -104860 -640 -104840
rect -1200 -105250 200 -105160
rect -1200 -108160 -1110 -105250
rect -480 -105450 -370 -105440
rect -480 -105460 520 -105450
rect -480 -105530 -470 -105460
rect -380 -105530 520 -105460
rect -480 -105540 520 -105530
rect -480 -105550 -370 -105540
rect -560 -106440 440 -106430
rect -560 -106510 -540 -106440
rect -260 -106510 440 -106440
rect -560 -106520 440 -106510
rect -760 -107770 40 -107750
rect -760 -107840 -740 -107770
rect -650 -107840 40 -107770
rect -750 -107860 -640 -107840
rect -1200 -108250 200 -108160
rect -1200 -111160 -1110 -108250
rect -480 -108450 -370 -108440
rect -480 -108460 520 -108450
rect -480 -108530 -470 -108460
rect -380 -108530 520 -108460
rect -480 -108540 520 -108530
rect -480 -108550 -370 -108540
rect -560 -109440 440 -109430
rect -560 -109510 -540 -109440
rect -260 -109510 440 -109440
rect -560 -109520 440 -109510
rect -760 -110770 40 -110750
rect -760 -110840 -740 -110770
rect -650 -110840 40 -110770
rect -750 -110860 -640 -110840
rect -1200 -111250 200 -111160
rect -1200 -114160 -1110 -111250
rect -480 -111450 -370 -111440
rect -480 -111460 520 -111450
rect -480 -111530 -470 -111460
rect -380 -111530 520 -111460
rect -480 -111540 520 -111530
rect -480 -111550 -370 -111540
rect -560 -112440 440 -112430
rect -560 -112510 -540 -112440
rect -260 -112510 440 -112440
rect -560 -112520 440 -112510
rect -760 -113770 40 -113750
rect -760 -113840 -740 -113770
rect -650 -113840 40 -113770
rect -750 -113860 -640 -113840
rect -1200 -114250 200 -114160
rect -1200 -117160 -1110 -114250
rect -480 -114450 -370 -114440
rect -480 -114460 520 -114450
rect -480 -114530 -470 -114460
rect -380 -114530 520 -114460
rect -480 -114540 520 -114530
rect -480 -114550 -370 -114540
rect -560 -115440 440 -115430
rect -560 -115510 -540 -115440
rect -260 -115510 440 -115440
rect -560 -115520 440 -115510
rect -760 -116770 40 -116750
rect -760 -116840 -740 -116770
rect -650 -116840 40 -116770
rect -750 -116860 -640 -116840
rect -1200 -117250 200 -117160
rect -1200 -120160 -1110 -117250
rect -480 -117450 -370 -117440
rect -480 -117460 520 -117450
rect -480 -117530 -470 -117460
rect -380 -117530 520 -117460
rect -480 -117540 520 -117530
rect -480 -117550 -370 -117540
rect -560 -118440 440 -118430
rect -560 -118510 -540 -118440
rect -260 -118510 440 -118440
rect -560 -118520 440 -118510
rect -760 -119770 40 -119750
rect -760 -119840 -740 -119770
rect -650 -119840 40 -119770
rect -750 -119860 -640 -119840
rect -1200 -120250 200 -120160
rect -1200 -123160 -1110 -120250
rect -480 -120450 -370 -120440
rect -480 -120460 520 -120450
rect -480 -120530 -470 -120460
rect -380 -120530 520 -120460
rect -480 -120540 520 -120530
rect -480 -120550 -370 -120540
rect -560 -121440 440 -121430
rect -560 -121510 -540 -121440
rect -260 -121510 440 -121440
rect -560 -121520 440 -121510
rect -760 -122770 40 -122750
rect -760 -122840 -740 -122770
rect -650 -122840 40 -122770
rect -750 -122860 -640 -122840
rect -1200 -123250 200 -123160
rect -1200 -126160 -1110 -123250
rect -480 -123450 -370 -123440
rect -480 -123460 520 -123450
rect -480 -123530 -470 -123460
rect -380 -123530 520 -123460
rect -480 -123540 520 -123530
rect -480 -123550 -370 -123540
rect -560 -124440 440 -124430
rect -560 -124510 -540 -124440
rect -260 -124510 440 -124440
rect -560 -124520 440 -124510
rect -760 -125770 40 -125750
rect -760 -125840 -740 -125770
rect -650 -125840 40 -125770
rect -750 -125860 -640 -125840
rect -1200 -126250 200 -126160
rect -1200 -129160 -1110 -126250
rect -480 -126450 -370 -126440
rect -480 -126460 520 -126450
rect -480 -126530 -470 -126460
rect -380 -126530 520 -126460
rect -480 -126540 520 -126530
rect -480 -126550 -370 -126540
rect -560 -127440 440 -127430
rect -560 -127510 -540 -127440
rect -260 -127510 440 -127440
rect -560 -127520 440 -127510
rect -760 -128770 40 -128750
rect -760 -128840 -740 -128770
rect -650 -128840 40 -128770
rect -750 -128860 -640 -128840
rect -1200 -129250 200 -129160
rect -1200 -132160 -1110 -129250
rect -480 -129450 -370 -129440
rect -480 -129460 520 -129450
rect -480 -129530 -470 -129460
rect -380 -129530 520 -129460
rect -480 -129540 520 -129530
rect -480 -129550 -370 -129540
rect -560 -130440 440 -130430
rect -560 -130510 -540 -130440
rect -260 -130510 440 -130440
rect -560 -130520 440 -130510
rect -760 -131770 40 -131750
rect -760 -131840 -740 -131770
rect -650 -131840 40 -131770
rect -750 -131860 -640 -131840
rect -1200 -132250 200 -132160
rect -1200 -135160 -1110 -132250
rect -480 -132450 -370 -132440
rect -480 -132460 520 -132450
rect -480 -132530 -470 -132460
rect -380 -132530 520 -132460
rect -480 -132540 520 -132530
rect -480 -132550 -370 -132540
rect -560 -133440 440 -133430
rect -560 -133510 -540 -133440
rect -260 -133510 440 -133440
rect -560 -133520 440 -133510
rect -760 -134770 40 -134750
rect -760 -134840 -740 -134770
rect -650 -134840 40 -134770
rect -750 -134860 -640 -134840
rect -1200 -135250 200 -135160
rect -1200 -138160 -1110 -135250
rect -480 -135450 -370 -135440
rect -480 -135460 520 -135450
rect -480 -135530 -470 -135460
rect -380 -135530 520 -135460
rect -480 -135540 520 -135530
rect -480 -135550 -370 -135540
rect -560 -136440 440 -136430
rect -560 -136510 -540 -136440
rect -260 -136510 440 -136440
rect -560 -136520 440 -136510
rect -760 -137770 40 -137750
rect -760 -137840 -740 -137770
rect -650 -137840 40 -137770
rect -750 -137860 -640 -137840
rect -1200 -138250 200 -138160
rect -1200 -141160 -1110 -138250
rect -480 -138450 -370 -138440
rect -480 -138460 520 -138450
rect -480 -138530 -470 -138460
rect -380 -138530 520 -138460
rect -480 -138540 520 -138530
rect -480 -138550 -370 -138540
rect -560 -139440 440 -139430
rect -560 -139510 -540 -139440
rect -260 -139510 440 -139440
rect -560 -139520 440 -139510
rect -760 -140770 40 -140750
rect -760 -140840 -740 -140770
rect -650 -140840 40 -140770
rect -750 -140860 -640 -140840
rect -1200 -141250 200 -141160
rect -1200 -144160 -1110 -141250
rect -480 -141450 -370 -141440
rect -480 -141460 520 -141450
rect -480 -141530 -470 -141460
rect -380 -141530 520 -141460
rect -480 -141540 520 -141530
rect -480 -141550 -370 -141540
rect -560 -142440 440 -142430
rect -560 -142510 -540 -142440
rect -260 -142510 440 -142440
rect -560 -142520 440 -142510
rect -760 -143770 40 -143750
rect -760 -143840 -740 -143770
rect -650 -143840 40 -143770
rect -750 -143860 -640 -143840
rect -1200 -144250 200 -144160
rect -1200 -147160 -1110 -144250
rect -480 -144450 -370 -144440
rect -480 -144460 520 -144450
rect -480 -144530 -470 -144460
rect -380 -144530 520 -144460
rect -480 -144540 520 -144530
rect -480 -144550 -370 -144540
rect -560 -145440 440 -145430
rect -560 -145510 -540 -145440
rect -260 -145510 440 -145440
rect -560 -145520 440 -145510
rect -760 -146770 40 -146750
rect -760 -146840 -740 -146770
rect -650 -146840 40 -146770
rect -750 -146860 -640 -146840
rect -1200 -147250 200 -147160
rect -1200 -150160 -1110 -147250
rect -480 -147450 -370 -147440
rect -480 -147460 520 -147450
rect -480 -147530 -470 -147460
rect -380 -147530 520 -147460
rect -480 -147540 520 -147530
rect -480 -147550 -370 -147540
rect -560 -148440 440 -148430
rect -560 -148510 -540 -148440
rect -260 -148510 440 -148440
rect -560 -148520 440 -148510
rect -760 -149770 40 -149750
rect -760 -149840 -740 -149770
rect -650 -149840 40 -149770
rect -750 -149860 -640 -149840
rect -1200 -150250 200 -150160
rect -1200 -153160 -1110 -150250
rect -480 -150450 -370 -150440
rect -480 -150460 520 -150450
rect -480 -150530 -470 -150460
rect -380 -150530 520 -150460
rect -480 -150540 520 -150530
rect -480 -150550 -370 -150540
rect -560 -151440 440 -151430
rect -560 -151510 -540 -151440
rect -260 -151510 440 -151440
rect -560 -151520 440 -151510
rect -760 -152770 40 -152750
rect -760 -152840 -740 -152770
rect -650 -152840 40 -152770
rect -750 -152860 -640 -152840
rect -1200 -153250 200 -153160
rect -1200 -156160 -1110 -153250
rect -480 -153450 -370 -153440
rect -480 -153460 520 -153450
rect -480 -153530 -470 -153460
rect -380 -153530 520 -153460
rect -480 -153540 520 -153530
rect -480 -153550 -370 -153540
rect -560 -154440 440 -154430
rect -560 -154510 -540 -154440
rect -260 -154510 440 -154440
rect -560 -154520 440 -154510
rect -760 -155770 40 -155750
rect -760 -155840 -740 -155770
rect -650 -155840 40 -155770
rect -750 -155860 -640 -155840
rect -1200 -156250 200 -156160
rect -1200 -159160 -1110 -156250
rect -480 -156450 -370 -156440
rect -480 -156460 520 -156450
rect -480 -156530 -470 -156460
rect -380 -156530 520 -156460
rect -480 -156540 520 -156530
rect -480 -156550 -370 -156540
rect -560 -157440 440 -157430
rect -560 -157510 -540 -157440
rect -260 -157510 440 -157440
rect -560 -157520 440 -157510
rect -760 -158770 40 -158750
rect -760 -158840 -740 -158770
rect -650 -158840 40 -158770
rect -750 -158860 -640 -158840
rect -1200 -159250 200 -159160
rect -1200 -162160 -1110 -159250
rect -480 -159450 -370 -159440
rect -480 -159460 520 -159450
rect -480 -159530 -470 -159460
rect -380 -159530 520 -159460
rect -480 -159540 520 -159530
rect -480 -159550 -370 -159540
rect -560 -160440 440 -160430
rect -560 -160510 -540 -160440
rect -260 -160510 440 -160440
rect -560 -160520 440 -160510
rect -760 -161770 40 -161750
rect -760 -161840 -740 -161770
rect -650 -161840 40 -161770
rect -750 -161860 -640 -161840
rect -1200 -162250 200 -162160
rect -1200 -165160 -1110 -162250
rect -480 -162450 -370 -162440
rect -480 -162460 520 -162450
rect -480 -162530 -470 -162460
rect -380 -162530 520 -162460
rect -480 -162540 520 -162530
rect -480 -162550 -370 -162540
rect -560 -163440 440 -163430
rect -560 -163510 -540 -163440
rect -260 -163510 440 -163440
rect -560 -163520 440 -163510
rect -760 -164770 40 -164750
rect -760 -164840 -740 -164770
rect -650 -164840 40 -164770
rect -750 -164860 -640 -164840
rect -1200 -165250 200 -165160
rect -1200 -168160 -1110 -165250
rect -480 -165450 -370 -165440
rect -480 -165460 520 -165450
rect -480 -165530 -470 -165460
rect -380 -165530 520 -165460
rect -480 -165540 520 -165530
rect -480 -165550 -370 -165540
rect -560 -166440 440 -166430
rect -560 -166510 -540 -166440
rect -260 -166510 440 -166440
rect -560 -166520 440 -166510
rect -760 -167770 40 -167750
rect -760 -167840 -740 -167770
rect -650 -167840 40 -167770
rect -750 -167860 -640 -167840
rect -1200 -168250 200 -168160
rect -1200 -171160 -1110 -168250
rect -480 -168450 -370 -168440
rect -480 -168460 520 -168450
rect -480 -168530 -470 -168460
rect -380 -168530 520 -168460
rect -480 -168540 520 -168530
rect -480 -168550 -370 -168540
rect -560 -169440 440 -169430
rect -560 -169510 -540 -169440
rect -260 -169510 440 -169440
rect -560 -169520 440 -169510
rect -760 -170770 40 -170750
rect -760 -170840 -740 -170770
rect -650 -170840 40 -170770
rect -750 -170860 -640 -170840
rect -1200 -171250 200 -171160
rect -1200 -174160 -1110 -171250
rect -480 -171450 -370 -171440
rect -480 -171460 520 -171450
rect -480 -171530 -470 -171460
rect -380 -171530 520 -171460
rect -480 -171540 520 -171530
rect -480 -171550 -370 -171540
rect -560 -172440 440 -172430
rect -560 -172510 -540 -172440
rect -260 -172510 440 -172440
rect -560 -172520 440 -172510
rect -760 -173770 40 -173750
rect -760 -173840 -740 -173770
rect -650 -173840 40 -173770
rect -750 -173860 -640 -173840
rect -1200 -174250 200 -174160
rect -1200 -177160 -1110 -174250
rect -480 -174450 -370 -174440
rect -480 -174460 520 -174450
rect -480 -174530 -470 -174460
rect -380 -174530 520 -174460
rect -480 -174540 520 -174530
rect -480 -174550 -370 -174540
rect -560 -175440 440 -175430
rect -560 -175510 -540 -175440
rect -260 -175510 440 -175440
rect -560 -175520 440 -175510
rect -760 -176770 40 -176750
rect -760 -176840 -740 -176770
rect -650 -176840 40 -176770
rect -750 -176860 -640 -176840
rect -1200 -177250 200 -177160
rect -1200 -180160 -1110 -177250
rect -480 -177450 -370 -177440
rect -480 -177460 520 -177450
rect -480 -177530 -470 -177460
rect -380 -177530 520 -177460
rect -480 -177540 520 -177530
rect -480 -177550 -370 -177540
rect -560 -178440 440 -178430
rect -560 -178510 -540 -178440
rect -260 -178510 440 -178440
rect -560 -178520 440 -178510
rect -760 -179770 40 -179750
rect -760 -179840 -740 -179770
rect -650 -179840 40 -179770
rect -750 -179860 -640 -179840
rect -1200 -180250 200 -180160
rect -1200 -183160 -1110 -180250
rect -480 -180450 -370 -180440
rect -480 -180460 520 -180450
rect -480 -180530 -470 -180460
rect -380 -180530 520 -180460
rect -480 -180540 520 -180530
rect -480 -180550 -370 -180540
rect -560 -181440 440 -181430
rect -560 -181510 -540 -181440
rect -260 -181510 440 -181440
rect -560 -181520 440 -181510
rect -760 -182770 40 -182750
rect -760 -182840 -740 -182770
rect -650 -182840 40 -182770
rect -750 -182860 -640 -182840
rect -1200 -183250 200 -183160
rect -1200 -186160 -1110 -183250
rect -480 -183450 -370 -183440
rect -480 -183460 520 -183450
rect -480 -183530 -470 -183460
rect -380 -183530 520 -183460
rect -480 -183540 520 -183530
rect -480 -183550 -370 -183540
rect -560 -184440 440 -184430
rect -560 -184510 -540 -184440
rect -260 -184510 440 -184440
rect -560 -184520 440 -184510
rect -760 -185770 40 -185750
rect -760 -185840 -740 -185770
rect -650 -185840 40 -185770
rect -750 -185860 -640 -185840
rect -1200 -186250 200 -186160
rect -1200 -189160 -1110 -186250
rect -480 -186450 -370 -186440
rect -480 -186460 520 -186450
rect -480 -186530 -470 -186460
rect -380 -186530 520 -186460
rect -480 -186540 520 -186530
rect -480 -186550 -370 -186540
rect -560 -187440 440 -187430
rect -560 -187510 -540 -187440
rect -260 -187510 440 -187440
rect -560 -187520 440 -187510
rect -760 -188770 40 -188750
rect -760 -188840 -740 -188770
rect -650 -188840 40 -188770
rect -750 -188860 -640 -188840
rect -1200 -189250 200 -189160
rect -1200 -192160 -1110 -189250
rect -480 -189450 -370 -189440
rect -480 -189460 520 -189450
rect -480 -189530 -470 -189460
rect -380 -189530 520 -189460
rect -480 -189540 520 -189530
rect -480 -189550 -370 -189540
rect -560 -190440 440 -190430
rect -560 -190510 -540 -190440
rect -260 -190510 440 -190440
rect -560 -190520 440 -190510
rect -760 -191770 40 -191750
rect -760 -191840 -740 -191770
rect -650 -191840 40 -191770
rect -750 -191860 -640 -191840
rect -1200 -192250 200 -192160
rect -1200 -195160 -1110 -192250
rect -480 -192450 -370 -192440
rect -480 -192460 520 -192450
rect -480 -192530 -470 -192460
rect -380 -192530 520 -192460
rect -480 -192540 520 -192530
rect -480 -192550 -370 -192540
rect -560 -193440 440 -193430
rect -560 -193510 -540 -193440
rect -260 -193510 440 -193440
rect -560 -193520 440 -193510
rect -760 -194770 40 -194750
rect -760 -194840 -740 -194770
rect -650 -194840 40 -194770
rect -750 -194860 -640 -194840
rect -1200 -195250 200 -195160
rect -1200 -198160 -1110 -195250
rect -480 -195450 -370 -195440
rect -480 -195460 520 -195450
rect -480 -195530 -470 -195460
rect -380 -195530 520 -195460
rect -480 -195540 520 -195530
rect -480 -195550 -370 -195540
rect -560 -196440 440 -196430
rect -560 -196510 -540 -196440
rect -260 -196510 440 -196440
rect -560 -196520 440 -196510
rect -760 -197770 40 -197750
rect -760 -197840 -740 -197770
rect -650 -197840 40 -197770
rect -750 -197860 -640 -197840
rect -1200 -198250 200 -198160
rect -1200 -201160 -1110 -198250
rect -480 -198450 -370 -198440
rect -480 -198460 520 -198450
rect -480 -198530 -470 -198460
rect -380 -198530 520 -198460
rect -480 -198540 520 -198530
rect -480 -198550 -370 -198540
rect -560 -199440 440 -199430
rect -560 -199510 -540 -199440
rect -260 -199510 440 -199440
rect -560 -199520 440 -199510
rect -760 -200770 40 -200750
rect -760 -200840 -740 -200770
rect -650 -200840 40 -200770
rect -750 -200860 -640 -200840
rect -1200 -201250 200 -201160
rect -1200 -204160 -1110 -201250
rect -480 -201450 -370 -201440
rect -480 -201460 520 -201450
rect -480 -201530 -470 -201460
rect -380 -201530 520 -201460
rect -480 -201540 520 -201530
rect -480 -201550 -370 -201540
rect -560 -202440 440 -202430
rect -560 -202510 -540 -202440
rect -260 -202510 440 -202440
rect -560 -202520 440 -202510
rect -760 -203770 40 -203750
rect -760 -203840 -740 -203770
rect -650 -203840 40 -203770
rect -750 -203860 -640 -203840
rect -1200 -204250 200 -204160
rect -1200 -207160 -1110 -204250
rect -480 -204450 -370 -204440
rect -480 -204460 520 -204450
rect -480 -204530 -470 -204460
rect -380 -204530 520 -204460
rect -480 -204540 520 -204530
rect -480 -204550 -370 -204540
rect -560 -205440 440 -205430
rect -560 -205510 -540 -205440
rect -260 -205510 440 -205440
rect -560 -205520 440 -205510
rect -760 -206770 40 -206750
rect -760 -206840 -740 -206770
rect -650 -206840 40 -206770
rect -750 -206860 -640 -206840
rect -1200 -207250 200 -207160
rect -1200 -210160 -1110 -207250
rect -480 -207450 -370 -207440
rect -480 -207460 520 -207450
rect -480 -207530 -470 -207460
rect -380 -207530 520 -207460
rect -480 -207540 520 -207530
rect -480 -207550 -370 -207540
rect -560 -208440 440 -208430
rect -560 -208510 -540 -208440
rect -260 -208510 440 -208440
rect -560 -208520 440 -208510
rect -760 -209770 40 -209750
rect -760 -209840 -740 -209770
rect -650 -209840 40 -209770
rect -750 -209860 -640 -209840
rect -1200 -210250 200 -210160
rect -1200 -213160 -1110 -210250
rect -480 -210450 -370 -210440
rect -480 -210460 520 -210450
rect -480 -210530 -470 -210460
rect -380 -210530 520 -210460
rect -480 -210540 520 -210530
rect -480 -210550 -370 -210540
rect -560 -211440 440 -211430
rect -560 -211510 -540 -211440
rect -260 -211510 440 -211440
rect -560 -211520 440 -211510
rect -760 -212770 40 -212750
rect -760 -212840 -740 -212770
rect -650 -212840 40 -212770
rect -750 -212860 -640 -212840
rect -1200 -213250 200 -213160
rect -1200 -216160 -1110 -213250
rect -480 -213450 -370 -213440
rect -480 -213460 520 -213450
rect -480 -213530 -470 -213460
rect -380 -213530 520 -213460
rect -480 -213540 520 -213530
rect -480 -213550 -370 -213540
rect -560 -214440 440 -214430
rect -560 -214510 -540 -214440
rect -260 -214510 440 -214440
rect -560 -214520 440 -214510
rect -760 -215770 40 -215750
rect -760 -215840 -740 -215770
rect -650 -215840 40 -215770
rect -750 -215860 -640 -215840
rect -1200 -216250 200 -216160
rect -1200 -219160 -1110 -216250
rect -480 -216450 -370 -216440
rect -480 -216460 520 -216450
rect -480 -216530 -470 -216460
rect -380 -216530 520 -216460
rect -480 -216540 520 -216530
rect -480 -216550 -370 -216540
rect -560 -217440 440 -217430
rect -560 -217510 -540 -217440
rect -260 -217510 440 -217440
rect -560 -217520 440 -217510
rect -760 -218770 40 -218750
rect -760 -218840 -740 -218770
rect -650 -218840 40 -218770
rect -750 -218860 -640 -218840
rect -1200 -219250 200 -219160
rect -1200 -222160 -1110 -219250
rect -480 -219450 -370 -219440
rect -480 -219460 520 -219450
rect -480 -219530 -470 -219460
rect -380 -219530 520 -219460
rect -480 -219540 520 -219530
rect -480 -219550 -370 -219540
rect -560 -220440 440 -220430
rect -560 -220510 -540 -220440
rect -260 -220510 440 -220440
rect -560 -220520 440 -220510
rect -760 -221770 40 -221750
rect -760 -221840 -740 -221770
rect -650 -221840 40 -221770
rect -750 -221860 -640 -221840
rect -1200 -222250 200 -222160
rect -1200 -225160 -1110 -222250
rect -480 -222450 -370 -222440
rect -480 -222460 520 -222450
rect -480 -222530 -470 -222460
rect -380 -222530 520 -222460
rect -480 -222540 520 -222530
rect -480 -222550 -370 -222540
rect -560 -223440 440 -223430
rect -560 -223510 -540 -223440
rect -260 -223510 440 -223440
rect -560 -223520 440 -223510
rect -760 -224770 40 -224750
rect -760 -224840 -740 -224770
rect -650 -224840 40 -224770
rect -750 -224860 -640 -224840
rect -1200 -225250 200 -225160
rect -1200 -228160 -1110 -225250
rect -480 -225450 -370 -225440
rect -480 -225460 520 -225450
rect -480 -225530 -470 -225460
rect -380 -225530 520 -225460
rect -480 -225540 520 -225530
rect -480 -225550 -370 -225540
rect -560 -226440 440 -226430
rect -560 -226510 -540 -226440
rect -260 -226510 440 -226440
rect -560 -226520 440 -226510
rect -760 -227770 40 -227750
rect -760 -227840 -740 -227770
rect -650 -227840 40 -227770
rect -750 -227860 -640 -227840
rect -1200 -228250 200 -228160
rect -1200 -231160 -1110 -228250
rect -480 -228450 -370 -228440
rect -480 -228460 520 -228450
rect -480 -228530 -470 -228460
rect -380 -228530 520 -228460
rect -480 -228540 520 -228530
rect -480 -228550 -370 -228540
rect -560 -229440 440 -229430
rect -560 -229510 -540 -229440
rect -260 -229510 440 -229440
rect -560 -229520 440 -229510
rect -760 -230770 40 -230750
rect -760 -230840 -740 -230770
rect -650 -230840 40 -230770
rect -750 -230860 -640 -230840
rect -1200 -231250 200 -231160
rect -1200 -234160 -1110 -231250
rect -480 -231450 -370 -231440
rect -480 -231460 520 -231450
rect -480 -231530 -470 -231460
rect -380 -231530 520 -231460
rect -480 -231540 520 -231530
rect -480 -231550 -370 -231540
rect -560 -232440 440 -232430
rect -560 -232510 -540 -232440
rect -260 -232510 440 -232440
rect -560 -232520 440 -232510
rect -760 -233770 40 -233750
rect -760 -233840 -740 -233770
rect -650 -233840 40 -233770
rect -750 -233860 -640 -233840
rect -1200 -234250 200 -234160
rect -1200 -237160 -1110 -234250
rect -480 -234450 -370 -234440
rect -480 -234460 520 -234450
rect -480 -234530 -470 -234460
rect -380 -234530 520 -234460
rect -480 -234540 520 -234530
rect -480 -234550 -370 -234540
rect -560 -235440 440 -235430
rect -560 -235510 -540 -235440
rect -260 -235510 440 -235440
rect -560 -235520 440 -235510
rect -760 -236770 40 -236750
rect -760 -236840 -740 -236770
rect -650 -236840 40 -236770
rect -750 -236860 -640 -236840
rect -1200 -237250 200 -237160
rect -1200 -240160 -1110 -237250
rect -480 -237450 -370 -237440
rect -480 -237460 520 -237450
rect -480 -237530 -470 -237460
rect -380 -237530 520 -237460
rect -480 -237540 520 -237530
rect -480 -237550 -370 -237540
rect -560 -238440 440 -238430
rect -560 -238510 -540 -238440
rect -260 -238510 440 -238440
rect -560 -238520 440 -238510
rect -760 -239770 40 -239750
rect -760 -239840 -740 -239770
rect -650 -239840 40 -239770
rect -750 -239860 -640 -239840
rect -1200 -240250 200 -240160
rect -1200 -243160 -1110 -240250
rect -480 -240450 -370 -240440
rect -480 -240460 520 -240450
rect -480 -240530 -470 -240460
rect -380 -240530 520 -240460
rect -480 -240540 520 -240530
rect -480 -240550 -370 -240540
rect -560 -241440 440 -241430
rect -560 -241510 -540 -241440
rect -260 -241510 440 -241440
rect -560 -241520 440 -241510
rect -760 -242770 40 -242750
rect -760 -242840 -740 -242770
rect -650 -242840 40 -242770
rect -750 -242860 -640 -242840
rect -1200 -243250 200 -243160
rect -1200 -246160 -1110 -243250
rect -480 -243450 -370 -243440
rect -480 -243460 520 -243450
rect -480 -243530 -470 -243460
rect -380 -243530 520 -243460
rect -480 -243540 520 -243530
rect -480 -243550 -370 -243540
rect -560 -244440 440 -244430
rect -560 -244510 -540 -244440
rect -260 -244510 440 -244440
rect -560 -244520 440 -244510
rect -760 -245770 40 -245750
rect -760 -245840 -740 -245770
rect -650 -245840 40 -245770
rect -750 -245860 -640 -245840
rect -1200 -246250 200 -246160
rect -1200 -249160 -1110 -246250
rect -480 -246450 -370 -246440
rect -480 -246460 520 -246450
rect -480 -246530 -470 -246460
rect -380 -246530 520 -246460
rect -480 -246540 520 -246530
rect -480 -246550 -370 -246540
rect -560 -247440 440 -247430
rect -560 -247510 -540 -247440
rect -260 -247510 440 -247440
rect -560 -247520 440 -247510
rect -760 -248770 40 -248750
rect -760 -248840 -740 -248770
rect -650 -248840 40 -248770
rect -750 -248860 -640 -248840
rect -1200 -249250 200 -249160
rect -1200 -252160 -1110 -249250
rect -480 -249450 -370 -249440
rect -480 -249460 520 -249450
rect -480 -249530 -470 -249460
rect -380 -249530 520 -249460
rect -480 -249540 520 -249530
rect -480 -249550 -370 -249540
rect -560 -250440 440 -250430
rect -560 -250510 -540 -250440
rect -260 -250510 440 -250440
rect -560 -250520 440 -250510
rect -760 -251770 40 -251750
rect -760 -251840 -740 -251770
rect -650 -251840 40 -251770
rect -750 -251860 -640 -251840
rect -1200 -252250 200 -252160
rect -1200 -255160 -1110 -252250
rect -480 -252450 -370 -252440
rect -480 -252460 520 -252450
rect -480 -252530 -470 -252460
rect -380 -252530 520 -252460
rect -480 -252540 520 -252530
rect -480 -252550 -370 -252540
rect -560 -253440 440 -253430
rect -560 -253510 -540 -253440
rect -260 -253510 440 -253440
rect -560 -253520 440 -253510
rect -760 -254770 40 -254750
rect -760 -254840 -740 -254770
rect -650 -254840 40 -254770
rect -750 -254860 -640 -254840
rect -1200 -255250 200 -255160
rect -1200 -258160 -1110 -255250
rect -480 -255450 -370 -255440
rect -480 -255460 520 -255450
rect -480 -255530 -470 -255460
rect -380 -255530 520 -255460
rect -480 -255540 520 -255530
rect -480 -255550 -370 -255540
rect -560 -256440 440 -256430
rect -560 -256510 -540 -256440
rect -260 -256510 440 -256440
rect -560 -256520 440 -256510
rect -760 -257770 40 -257750
rect -760 -257840 -740 -257770
rect -650 -257840 40 -257770
rect -750 -257860 -640 -257840
rect -1200 -258250 200 -258160
rect -1200 -261160 -1110 -258250
rect -480 -258450 -370 -258440
rect -480 -258460 520 -258450
rect -480 -258530 -470 -258460
rect -380 -258530 520 -258460
rect -480 -258540 520 -258530
rect -480 -258550 -370 -258540
rect -560 -259440 440 -259430
rect -560 -259510 -540 -259440
rect -260 -259510 440 -259440
rect -560 -259520 440 -259510
rect -760 -260770 40 -260750
rect -760 -260840 -740 -260770
rect -650 -260840 40 -260770
rect -750 -260860 -640 -260840
rect -1200 -261250 200 -261160
rect -1200 -264160 -1110 -261250
rect -480 -261450 -370 -261440
rect -480 -261460 520 -261450
rect -480 -261530 -470 -261460
rect -380 -261530 520 -261460
rect -480 -261540 520 -261530
rect -480 -261550 -370 -261540
rect -560 -262440 440 -262430
rect -560 -262510 -540 -262440
rect -260 -262510 440 -262440
rect -560 -262520 440 -262510
rect -760 -263770 40 -263750
rect -760 -263840 -740 -263770
rect -650 -263840 40 -263770
rect -750 -263860 -640 -263840
rect -1200 -264250 200 -264160
rect -1200 -267160 -1110 -264250
rect -480 -264450 -370 -264440
rect -480 -264460 520 -264450
rect -480 -264530 -470 -264460
rect -380 -264530 520 -264460
rect -480 -264540 520 -264530
rect -480 -264550 -370 -264540
rect -560 -265440 440 -265430
rect -560 -265510 -540 -265440
rect -260 -265510 440 -265440
rect -560 -265520 440 -265510
rect -760 -266770 40 -266750
rect -760 -266840 -740 -266770
rect -650 -266840 40 -266770
rect -750 -266860 -640 -266840
rect -1200 -267250 200 -267160
rect -1200 -270160 -1110 -267250
rect -480 -267450 -370 -267440
rect -480 -267460 520 -267450
rect -480 -267530 -470 -267460
rect -380 -267530 520 -267460
rect -480 -267540 520 -267530
rect -480 -267550 -370 -267540
rect -560 -268440 440 -268430
rect -560 -268510 -540 -268440
rect -260 -268510 440 -268440
rect -560 -268520 440 -268510
rect -760 -269770 40 -269750
rect -760 -269840 -740 -269770
rect -650 -269840 40 -269770
rect -750 -269860 -640 -269840
rect -1200 -270250 200 -270160
rect -1200 -273160 -1110 -270250
rect -480 -270450 -370 -270440
rect -480 -270460 520 -270450
rect -480 -270530 -470 -270460
rect -380 -270530 520 -270460
rect -480 -270540 520 -270530
rect -480 -270550 -370 -270540
rect -560 -271440 440 -271430
rect -560 -271510 -540 -271440
rect -260 -271510 440 -271440
rect -560 -271520 440 -271510
rect -760 -272770 40 -272750
rect -760 -272840 -740 -272770
rect -650 -272840 40 -272770
rect -750 -272860 -640 -272840
rect -1200 -273250 200 -273160
rect -1200 -276160 -1110 -273250
rect -480 -273450 -370 -273440
rect -480 -273460 520 -273450
rect -480 -273530 -470 -273460
rect -380 -273530 520 -273460
rect -480 -273540 520 -273530
rect -480 -273550 -370 -273540
rect -560 -274440 440 -274430
rect -560 -274510 -540 -274440
rect -260 -274510 440 -274440
rect -560 -274520 440 -274510
rect -760 -275770 40 -275750
rect -760 -275840 -740 -275770
rect -650 -275840 40 -275770
rect -750 -275860 -640 -275840
rect -1200 -276250 200 -276160
rect -1200 -279160 -1110 -276250
rect -480 -276450 -370 -276440
rect -480 -276460 520 -276450
rect -480 -276530 -470 -276460
rect -380 -276530 520 -276460
rect -480 -276540 520 -276530
rect -480 -276550 -370 -276540
rect -560 -277440 440 -277430
rect -560 -277510 -540 -277440
rect -260 -277510 440 -277440
rect -560 -277520 440 -277510
rect -760 -278770 40 -278750
rect -760 -278840 -740 -278770
rect -650 -278840 40 -278770
rect -750 -278860 -640 -278840
rect -1200 -279250 200 -279160
rect -1200 -282160 -1110 -279250
rect -480 -279450 -370 -279440
rect -480 -279460 520 -279450
rect -480 -279530 -470 -279460
rect -380 -279530 520 -279460
rect -480 -279540 520 -279530
rect -480 -279550 -370 -279540
rect -560 -280440 440 -280430
rect -560 -280510 -540 -280440
rect -260 -280510 440 -280440
rect -560 -280520 440 -280510
rect -760 -281770 40 -281750
rect -760 -281840 -740 -281770
rect -650 -281840 40 -281770
rect -750 -281860 -640 -281840
rect -1200 -282250 200 -282160
rect -1200 -285160 -1110 -282250
rect -480 -282450 -370 -282440
rect -480 -282460 520 -282450
rect -480 -282530 -470 -282460
rect -380 -282530 520 -282460
rect -480 -282540 520 -282530
rect -480 -282550 -370 -282540
rect -560 -283440 440 -283430
rect -560 -283510 -540 -283440
rect -260 -283510 440 -283440
rect -560 -283520 440 -283510
rect -760 -284770 40 -284750
rect -760 -284840 -740 -284770
rect -650 -284840 40 -284770
rect -750 -284860 -640 -284840
rect -1200 -285250 200 -285160
rect -1200 -288160 -1110 -285250
rect -480 -285450 -370 -285440
rect -480 -285460 520 -285450
rect -480 -285530 -470 -285460
rect -380 -285530 520 -285460
rect -480 -285540 520 -285530
rect -480 -285550 -370 -285540
rect -560 -286440 440 -286430
rect -560 -286510 -540 -286440
rect -260 -286510 440 -286440
rect -560 -286520 440 -286510
rect -760 -287770 40 -287750
rect -760 -287840 -740 -287770
rect -650 -287840 40 -287770
rect -750 -287860 -640 -287840
rect -1200 -288250 200 -288160
rect -1200 -291160 -1110 -288250
rect -480 -288450 -370 -288440
rect -480 -288460 520 -288450
rect -480 -288530 -470 -288460
rect -380 -288530 520 -288460
rect -480 -288540 520 -288530
rect -480 -288550 -370 -288540
rect -560 -289440 440 -289430
rect -560 -289510 -540 -289440
rect -260 -289510 440 -289440
rect -560 -289520 440 -289510
rect -760 -290770 40 -290750
rect -760 -290840 -740 -290770
rect -650 -290840 40 -290770
rect -750 -290860 -640 -290840
rect -1200 -291250 200 -291160
rect -1200 -294160 -1110 -291250
rect -480 -291450 -370 -291440
rect -480 -291460 520 -291450
rect -480 -291530 -470 -291460
rect -380 -291530 520 -291460
rect -480 -291540 520 -291530
rect -480 -291550 -370 -291540
rect -560 -292440 440 -292430
rect -560 -292510 -540 -292440
rect -260 -292510 440 -292440
rect -560 -292520 440 -292510
rect -760 -293770 40 -293750
rect -760 -293840 -740 -293770
rect -650 -293840 40 -293770
rect -750 -293860 -640 -293840
rect -1200 -294250 200 -294160
rect -1200 -295000 -1110 -294250
rect -480 -294450 -370 -294440
rect -480 -294460 520 -294450
rect -480 -294530 -470 -294460
rect -380 -294530 520 -294460
rect -480 -294540 520 -294530
rect -480 -294550 -370 -294540
rect -560 -295440 440 -295430
rect -560 -295510 -540 -295440
rect -260 -295510 440 -295440
rect -560 -295520 440 -295510
rect -760 -296770 40 -296750
rect -760 -296840 -740 -296770
rect -650 -296840 40 -296770
rect -750 -296860 -640 -296840
rect 540 -297080 2780 -297060
rect 540 -297180 560 -297080
rect 2760 -297180 2780 -297080
rect 540 -297200 2780 -297180
rect 3540 -297080 5780 -297060
rect 3540 -297180 3560 -297080
rect 5760 -297180 5780 -297080
rect 3540 -297200 5780 -297180
rect 6540 -297080 8780 -297060
rect 6540 -297180 6560 -297080
rect 8760 -297180 8780 -297080
rect 6540 -297200 8780 -297180
rect 9540 -297080 11780 -297060
rect 9540 -297180 9560 -297080
rect 11760 -297180 11780 -297080
rect 9540 -297200 11780 -297180
rect 12540 -297080 14780 -297060
rect 12540 -297180 12560 -297080
rect 14760 -297180 14780 -297080
rect 12540 -297200 14780 -297180
rect 15540 -297080 17780 -297060
rect 15540 -297180 15560 -297080
rect 17760 -297180 17780 -297080
rect 15540 -297200 17780 -297180
rect 18540 -297080 20780 -297060
rect 18540 -297180 18560 -297080
rect 20760 -297180 20780 -297080
rect 18540 -297200 20780 -297180
rect 21540 -297080 23780 -297060
rect 21540 -297180 21560 -297080
rect 23760 -297180 23780 -297080
rect 21540 -297200 23780 -297180
rect 24540 -297080 26780 -297060
rect 24540 -297180 24560 -297080
rect 26760 -297180 26780 -297080
rect 24540 -297200 26780 -297180
rect 27540 -297080 29780 -297060
rect 27540 -297180 27560 -297080
rect 29760 -297180 29780 -297080
rect 27540 -297200 29780 -297180
rect 30540 -297080 32780 -297060
rect 30540 -297180 30560 -297080
rect 32760 -297180 32780 -297080
rect 30540 -297200 32780 -297180
rect 33540 -297080 35780 -297060
rect 33540 -297180 33560 -297080
rect 35760 -297180 35780 -297080
rect 33540 -297200 35780 -297180
rect 36540 -297080 38780 -297060
rect 36540 -297180 36560 -297080
rect 38760 -297180 38780 -297080
rect 36540 -297200 38780 -297180
rect 39540 -297080 41780 -297060
rect 39540 -297180 39560 -297080
rect 41760 -297180 41780 -297080
rect 39540 -297200 41780 -297180
rect 42540 -297080 44780 -297060
rect 42540 -297180 42560 -297080
rect 44760 -297180 44780 -297080
rect 42540 -297200 44780 -297180
rect 45540 -297080 47780 -297060
rect 45540 -297180 45560 -297080
rect 47760 -297180 47780 -297080
rect 45540 -297200 47780 -297180
rect 48540 -297080 50780 -297060
rect 48540 -297180 48560 -297080
rect 50760 -297180 50780 -297080
rect 48540 -297200 50780 -297180
rect 51540 -297080 53780 -297060
rect 51540 -297180 51560 -297080
rect 53760 -297180 53780 -297080
rect 51540 -297200 53780 -297180
rect 54540 -297080 56780 -297060
rect 54540 -297180 54560 -297080
rect 56760 -297180 56780 -297080
rect 54540 -297200 56780 -297180
rect 57540 -297080 59780 -297060
rect 57540 -297180 57560 -297080
rect 59760 -297180 59780 -297080
rect 57540 -297200 59780 -297180
rect 60540 -297080 62780 -297060
rect 60540 -297180 60560 -297080
rect 62760 -297180 62780 -297080
rect 60540 -297200 62780 -297180
rect 63540 -297080 65780 -297060
rect 63540 -297180 63560 -297080
rect 65760 -297180 65780 -297080
rect 63540 -297200 65780 -297180
rect 66540 -297080 68780 -297060
rect 66540 -297180 66560 -297080
rect 68760 -297180 68780 -297080
rect 66540 -297200 68780 -297180
rect 69540 -297080 71780 -297060
rect 69540 -297180 69560 -297080
rect 71760 -297180 71780 -297080
rect 69540 -297200 71780 -297180
rect 72540 -297080 74780 -297060
rect 72540 -297180 72560 -297080
rect 74760 -297180 74780 -297080
rect 72540 -297200 74780 -297180
rect 75540 -297080 77780 -297060
rect 75540 -297180 75560 -297080
rect 77760 -297180 77780 -297080
rect 75540 -297200 77780 -297180
rect 78540 -297080 80780 -297060
rect 78540 -297180 78560 -297080
rect 80760 -297180 80780 -297080
rect 78540 -297200 80780 -297180
rect 81540 -297080 83780 -297060
rect 81540 -297180 81560 -297080
rect 83760 -297180 83780 -297080
rect 81540 -297200 83780 -297180
rect 84540 -297080 86780 -297060
rect 84540 -297180 84560 -297080
rect 86760 -297180 86780 -297080
rect 84540 -297200 86780 -297180
rect 87540 -297080 89780 -297060
rect 87540 -297180 87560 -297080
rect 89760 -297180 89780 -297080
rect 87540 -297200 89780 -297180
rect 90540 -297080 92780 -297060
rect 90540 -297180 90560 -297080
rect 92760 -297180 92780 -297080
rect 90540 -297200 92780 -297180
rect 93540 -297080 95780 -297060
rect 93540 -297180 93560 -297080
rect 95760 -297180 95780 -297080
rect 93540 -297200 95780 -297180
rect 96540 -297080 98780 -297060
rect 96540 -297180 96560 -297080
rect 98760 -297180 98780 -297080
rect 96540 -297200 98780 -297180
rect 99540 -297080 101780 -297060
rect 99540 -297180 99560 -297080
rect 101760 -297180 101780 -297080
rect 99540 -297200 101780 -297180
rect 102540 -297080 104780 -297060
rect 102540 -297180 102560 -297080
rect 104760 -297180 104780 -297080
rect 102540 -297200 104780 -297180
rect 105540 -297080 107780 -297060
rect 105540 -297180 105560 -297080
rect 107760 -297180 107780 -297080
rect 105540 -297200 107780 -297180
rect 108540 -297080 110780 -297060
rect 108540 -297180 108560 -297080
rect 110760 -297180 110780 -297080
rect 108540 -297200 110780 -297180
rect 111540 -297080 113780 -297060
rect 111540 -297180 111560 -297080
rect 113760 -297180 113780 -297080
rect 111540 -297200 113780 -297180
rect 114540 -297080 116780 -297060
rect 114540 -297180 114560 -297080
rect 116760 -297180 116780 -297080
rect 114540 -297200 116780 -297180
rect 117540 -297080 119780 -297060
rect 117540 -297180 117560 -297080
rect 119760 -297180 119780 -297080
rect 117540 -297200 119780 -297180
rect 120540 -297080 122780 -297060
rect 120540 -297180 120560 -297080
rect 122760 -297180 122780 -297080
rect 120540 -297200 122780 -297180
rect 123540 -297080 125780 -297060
rect 123540 -297180 123560 -297080
rect 125760 -297180 125780 -297080
rect 123540 -297200 125780 -297180
rect 126540 -297080 128780 -297060
rect 126540 -297180 126560 -297080
rect 128760 -297180 128780 -297080
rect 126540 -297200 128780 -297180
rect 129540 -297080 131780 -297060
rect 129540 -297180 129560 -297080
rect 131760 -297180 131780 -297080
rect 129540 -297200 131780 -297180
rect 132540 -297080 134780 -297060
rect 132540 -297180 132560 -297080
rect 134760 -297180 134780 -297080
rect 132540 -297200 134780 -297180
rect 135540 -297080 137780 -297060
rect 135540 -297180 135560 -297080
rect 137760 -297180 137780 -297080
rect 135540 -297200 137780 -297180
rect 138540 -297080 140780 -297060
rect 138540 -297180 138560 -297080
rect 140760 -297180 140780 -297080
rect 138540 -297200 140780 -297180
rect 141540 -297080 143780 -297060
rect 141540 -297180 141560 -297080
rect 143760 -297180 143780 -297080
rect 141540 -297200 143780 -297180
rect 144540 -297080 146780 -297060
rect 144540 -297180 144560 -297080
rect 146760 -297180 146780 -297080
rect 144540 -297200 146780 -297180
rect 147540 -297080 149780 -297060
rect 147540 -297180 147560 -297080
rect 149760 -297180 149780 -297080
rect 147540 -297200 149780 -297180
rect 150540 -297080 152780 -297060
rect 150540 -297180 150560 -297080
rect 152760 -297180 152780 -297080
rect 150540 -297200 152780 -297180
rect 153540 -297080 155780 -297060
rect 153540 -297180 153560 -297080
rect 155760 -297180 155780 -297080
rect 153540 -297200 155780 -297180
rect 156540 -297080 158780 -297060
rect 156540 -297180 156560 -297080
rect 158760 -297180 158780 -297080
rect 156540 -297200 158780 -297180
rect 159540 -297080 161780 -297060
rect 159540 -297180 159560 -297080
rect 161760 -297180 161780 -297080
rect 159540 -297200 161780 -297180
rect 162540 -297080 164780 -297060
rect 162540 -297180 162560 -297080
rect 164760 -297180 164780 -297080
rect 162540 -297200 164780 -297180
rect 165540 -297080 167780 -297060
rect 165540 -297180 165560 -297080
rect 167760 -297180 167780 -297080
rect 165540 -297200 167780 -297180
rect 168540 -297080 170780 -297060
rect 168540 -297180 168560 -297080
rect 170760 -297180 170780 -297080
rect 168540 -297200 170780 -297180
rect 171540 -297080 173780 -297060
rect 171540 -297180 171560 -297080
rect 173760 -297180 173780 -297080
rect 171540 -297200 173780 -297180
rect 174540 -297080 176780 -297060
rect 174540 -297180 174560 -297080
rect 176760 -297180 176780 -297080
rect 174540 -297200 176780 -297180
rect 177540 -297080 179780 -297060
rect 177540 -297180 177560 -297080
rect 179760 -297180 179780 -297080
rect 177540 -297200 179780 -297180
rect 180540 -297080 182780 -297060
rect 180540 -297180 180560 -297080
rect 182760 -297180 182780 -297080
rect 180540 -297200 182780 -297180
rect 183540 -297080 185780 -297060
rect 183540 -297180 183560 -297080
rect 185760 -297180 185780 -297080
rect 183540 -297200 185780 -297180
rect 186540 -297080 188780 -297060
rect 186540 -297180 186560 -297080
rect 188760 -297180 188780 -297080
rect 186540 -297200 188780 -297180
rect 189540 -297080 191780 -297060
rect 189540 -297180 189560 -297080
rect 191760 -297180 191780 -297080
rect 189540 -297200 191780 -297180
rect 192540 -297080 194780 -297060
rect 192540 -297180 192560 -297080
rect 194760 -297180 194780 -297080
rect 192540 -297200 194780 -297180
rect 195540 -297080 197780 -297060
rect 195540 -297180 195560 -297080
rect 197760 -297180 197780 -297080
rect 195540 -297200 197780 -297180
rect 198540 -297080 200780 -297060
rect 198540 -297180 198560 -297080
rect 200760 -297180 200780 -297080
rect 198540 -297200 200780 -297180
rect 201540 -297080 203780 -297060
rect 201540 -297180 201560 -297080
rect 203760 -297180 203780 -297080
rect 201540 -297200 203780 -297180
rect 204540 -297080 206780 -297060
rect 204540 -297180 204560 -297080
rect 206760 -297180 206780 -297080
rect 204540 -297200 206780 -297180
rect 207540 -297080 209780 -297060
rect 207540 -297180 207560 -297080
rect 209760 -297180 209780 -297080
rect 207540 -297200 209780 -297180
rect 210540 -297080 212780 -297060
rect 210540 -297180 210560 -297080
rect 212760 -297180 212780 -297080
rect 210540 -297200 212780 -297180
rect 213540 -297080 215780 -297060
rect 213540 -297180 213560 -297080
rect 215760 -297180 215780 -297080
rect 213540 -297200 215780 -297180
rect 216540 -297080 218780 -297060
rect 216540 -297180 216560 -297080
rect 218760 -297180 218780 -297080
rect 216540 -297200 218780 -297180
rect 219540 -297080 221780 -297060
rect 219540 -297180 219560 -297080
rect 221760 -297180 221780 -297080
rect 219540 -297200 221780 -297180
rect 222540 -297080 224780 -297060
rect 222540 -297180 222560 -297080
rect 224760 -297180 224780 -297080
rect 222540 -297200 224780 -297180
rect 225540 -297080 227780 -297060
rect 225540 -297180 225560 -297080
rect 227760 -297180 227780 -297080
rect 225540 -297200 227780 -297180
rect 228540 -297080 230780 -297060
rect 228540 -297180 228560 -297080
rect 230760 -297180 230780 -297080
rect 228540 -297200 230780 -297180
rect 231540 -297080 233780 -297060
rect 231540 -297180 231560 -297080
rect 233760 -297180 233780 -297080
rect 231540 -297200 233780 -297180
rect 234540 -297080 236780 -297060
rect 234540 -297180 234560 -297080
rect 236760 -297180 236780 -297080
rect 234540 -297200 236780 -297180
rect 237540 -297080 239780 -297060
rect 237540 -297180 237560 -297080
rect 239760 -297180 239780 -297080
rect 237540 -297200 239780 -297180
rect 240540 -297080 242780 -297060
rect 240540 -297180 240560 -297080
rect 242760 -297180 242780 -297080
rect 240540 -297200 242780 -297180
rect 243540 -297080 245780 -297060
rect 243540 -297180 243560 -297080
rect 245760 -297180 245780 -297080
rect 243540 -297200 245780 -297180
rect 246540 -297080 248780 -297060
rect 246540 -297180 246560 -297080
rect 248760 -297180 248780 -297080
rect 246540 -297200 248780 -297180
rect 249540 -297080 251780 -297060
rect 249540 -297180 249560 -297080
rect 251760 -297180 251780 -297080
rect 249540 -297200 251780 -297180
rect 252540 -297080 254780 -297060
rect 252540 -297180 252560 -297080
rect 254760 -297180 254780 -297080
rect 252540 -297200 254780 -297180
rect 255540 -297080 257780 -297060
rect 255540 -297180 255560 -297080
rect 257760 -297180 257780 -297080
rect 255540 -297200 257780 -297180
rect 258540 -297080 260780 -297060
rect 258540 -297180 258560 -297080
rect 260760 -297180 260780 -297080
rect 258540 -297200 260780 -297180
rect 261540 -297080 263780 -297060
rect 261540 -297180 261560 -297080
rect 263760 -297180 263780 -297080
rect 261540 -297200 263780 -297180
rect 264540 -297080 266780 -297060
rect 264540 -297180 264560 -297080
rect 266760 -297180 266780 -297080
rect 264540 -297200 266780 -297180
rect 267540 -297080 269780 -297060
rect 267540 -297180 267560 -297080
rect 269760 -297180 269780 -297080
rect 267540 -297200 269780 -297180
rect 270540 -297080 272780 -297060
rect 270540 -297180 270560 -297080
rect 272760 -297180 272780 -297080
rect 270540 -297200 272780 -297180
rect 273540 -297080 275780 -297060
rect 273540 -297180 273560 -297080
rect 275760 -297180 275780 -297080
rect 273540 -297200 275780 -297180
rect 276540 -297080 278780 -297060
rect 276540 -297180 276560 -297080
rect 278760 -297180 278780 -297080
rect 276540 -297200 278780 -297180
rect 279540 -297080 281780 -297060
rect 279540 -297180 279560 -297080
rect 281760 -297180 281780 -297080
rect 279540 -297200 281780 -297180
rect 282540 -297080 284780 -297060
rect 282540 -297180 282560 -297080
rect 284760 -297180 284780 -297080
rect 282540 -297200 284780 -297180
rect 285540 -297080 287780 -297060
rect 285540 -297180 285560 -297080
rect 287760 -297180 287780 -297080
rect 285540 -297200 287780 -297180
rect 288540 -297080 290780 -297060
rect 288540 -297180 288560 -297080
rect 290760 -297180 290780 -297080
rect 288540 -297200 290780 -297180
rect 291540 -297080 293780 -297060
rect 291540 -297180 291560 -297080
rect 293760 -297180 293780 -297080
rect 291540 -297200 293780 -297180
rect 294540 -297080 296780 -297060
rect 294540 -297180 294560 -297080
rect 296760 -297180 296780 -297080
rect 294540 -297200 296780 -297180
rect 297540 -297080 299780 -297060
rect 297540 -297180 297560 -297080
rect 299760 -297180 299780 -297080
rect 297540 -297200 299780 -297180
rect 220 -297500 440 -297490
rect 220 -297700 240 -297500
rect 420 -297700 440 -297500
rect 220 -297710 440 -297700
rect 3220 -297500 3440 -297490
rect 3220 -297700 3240 -297500
rect 3420 -297700 3440 -297500
rect 3220 -297710 3440 -297700
rect 6220 -297500 6440 -297490
rect 6220 -297700 6240 -297500
rect 6420 -297700 6440 -297500
rect 6220 -297710 6440 -297700
rect 9220 -297500 9440 -297490
rect 9220 -297700 9240 -297500
rect 9420 -297700 9440 -297500
rect 9220 -297710 9440 -297700
rect 12220 -297500 12440 -297490
rect 12220 -297700 12240 -297500
rect 12420 -297700 12440 -297500
rect 12220 -297710 12440 -297700
rect 15220 -297500 15440 -297490
rect 15220 -297700 15240 -297500
rect 15420 -297700 15440 -297500
rect 15220 -297710 15440 -297700
rect 18220 -297500 18440 -297490
rect 18220 -297700 18240 -297500
rect 18420 -297700 18440 -297500
rect 18220 -297710 18440 -297700
rect 21220 -297500 21440 -297490
rect 21220 -297700 21240 -297500
rect 21420 -297700 21440 -297500
rect 21220 -297710 21440 -297700
rect 24220 -297500 24440 -297490
rect 24220 -297700 24240 -297500
rect 24420 -297700 24440 -297500
rect 24220 -297710 24440 -297700
rect 27220 -297500 27440 -297490
rect 27220 -297700 27240 -297500
rect 27420 -297700 27440 -297500
rect 27220 -297710 27440 -297700
rect 30220 -297500 30440 -297490
rect 30220 -297700 30240 -297500
rect 30420 -297700 30440 -297500
rect 30220 -297710 30440 -297700
rect 33220 -297500 33440 -297490
rect 33220 -297700 33240 -297500
rect 33420 -297700 33440 -297500
rect 33220 -297710 33440 -297700
rect 36220 -297500 36440 -297490
rect 36220 -297700 36240 -297500
rect 36420 -297700 36440 -297500
rect 36220 -297710 36440 -297700
rect 39220 -297500 39440 -297490
rect 39220 -297700 39240 -297500
rect 39420 -297700 39440 -297500
rect 39220 -297710 39440 -297700
rect 42220 -297500 42440 -297490
rect 42220 -297700 42240 -297500
rect 42420 -297700 42440 -297500
rect 42220 -297710 42440 -297700
rect 45220 -297500 45440 -297490
rect 45220 -297700 45240 -297500
rect 45420 -297700 45440 -297500
rect 45220 -297710 45440 -297700
rect 48220 -297500 48440 -297490
rect 48220 -297700 48240 -297500
rect 48420 -297700 48440 -297500
rect 48220 -297710 48440 -297700
rect 51220 -297500 51440 -297490
rect 51220 -297700 51240 -297500
rect 51420 -297700 51440 -297500
rect 51220 -297710 51440 -297700
rect 54220 -297500 54440 -297490
rect 54220 -297700 54240 -297500
rect 54420 -297700 54440 -297500
rect 54220 -297710 54440 -297700
rect 57220 -297500 57440 -297490
rect 57220 -297700 57240 -297500
rect 57420 -297700 57440 -297500
rect 57220 -297710 57440 -297700
rect 60220 -297500 60440 -297490
rect 60220 -297700 60240 -297500
rect 60420 -297700 60440 -297500
rect 60220 -297710 60440 -297700
rect 63220 -297500 63440 -297490
rect 63220 -297700 63240 -297500
rect 63420 -297700 63440 -297500
rect 63220 -297710 63440 -297700
rect 66220 -297500 66440 -297490
rect 66220 -297700 66240 -297500
rect 66420 -297700 66440 -297500
rect 66220 -297710 66440 -297700
rect 69220 -297500 69440 -297490
rect 69220 -297700 69240 -297500
rect 69420 -297700 69440 -297500
rect 69220 -297710 69440 -297700
rect 72220 -297500 72440 -297490
rect 72220 -297700 72240 -297500
rect 72420 -297700 72440 -297500
rect 72220 -297710 72440 -297700
rect 75220 -297500 75440 -297490
rect 75220 -297700 75240 -297500
rect 75420 -297700 75440 -297500
rect 75220 -297710 75440 -297700
rect 78220 -297500 78440 -297490
rect 78220 -297700 78240 -297500
rect 78420 -297700 78440 -297500
rect 78220 -297710 78440 -297700
rect 81220 -297500 81440 -297490
rect 81220 -297700 81240 -297500
rect 81420 -297700 81440 -297500
rect 81220 -297710 81440 -297700
rect 84220 -297500 84440 -297490
rect 84220 -297700 84240 -297500
rect 84420 -297700 84440 -297500
rect 84220 -297710 84440 -297700
rect 87220 -297500 87440 -297490
rect 87220 -297700 87240 -297500
rect 87420 -297700 87440 -297500
rect 87220 -297710 87440 -297700
rect 90220 -297500 90440 -297490
rect 90220 -297700 90240 -297500
rect 90420 -297700 90440 -297500
rect 90220 -297710 90440 -297700
rect 93220 -297500 93440 -297490
rect 93220 -297700 93240 -297500
rect 93420 -297700 93440 -297500
rect 93220 -297710 93440 -297700
rect 96220 -297500 96440 -297490
rect 96220 -297700 96240 -297500
rect 96420 -297700 96440 -297500
rect 96220 -297710 96440 -297700
rect 99220 -297500 99440 -297490
rect 99220 -297700 99240 -297500
rect 99420 -297700 99440 -297500
rect 99220 -297710 99440 -297700
rect 102220 -297500 102440 -297490
rect 102220 -297700 102240 -297500
rect 102420 -297700 102440 -297500
rect 102220 -297710 102440 -297700
rect 105220 -297500 105440 -297490
rect 105220 -297700 105240 -297500
rect 105420 -297700 105440 -297500
rect 105220 -297710 105440 -297700
rect 108220 -297500 108440 -297490
rect 108220 -297700 108240 -297500
rect 108420 -297700 108440 -297500
rect 108220 -297710 108440 -297700
rect 111220 -297500 111440 -297490
rect 111220 -297700 111240 -297500
rect 111420 -297700 111440 -297500
rect 111220 -297710 111440 -297700
rect 114220 -297500 114440 -297490
rect 114220 -297700 114240 -297500
rect 114420 -297700 114440 -297500
rect 114220 -297710 114440 -297700
rect 117220 -297500 117440 -297490
rect 117220 -297700 117240 -297500
rect 117420 -297700 117440 -297500
rect 117220 -297710 117440 -297700
rect 120220 -297500 120440 -297490
rect 120220 -297700 120240 -297500
rect 120420 -297700 120440 -297500
rect 120220 -297710 120440 -297700
rect 123220 -297500 123440 -297490
rect 123220 -297700 123240 -297500
rect 123420 -297700 123440 -297500
rect 123220 -297710 123440 -297700
rect 126220 -297500 126440 -297490
rect 126220 -297700 126240 -297500
rect 126420 -297700 126440 -297500
rect 126220 -297710 126440 -297700
rect 129220 -297500 129440 -297490
rect 129220 -297700 129240 -297500
rect 129420 -297700 129440 -297500
rect 129220 -297710 129440 -297700
rect 132220 -297500 132440 -297490
rect 132220 -297700 132240 -297500
rect 132420 -297700 132440 -297500
rect 132220 -297710 132440 -297700
rect 135220 -297500 135440 -297490
rect 135220 -297700 135240 -297500
rect 135420 -297700 135440 -297500
rect 135220 -297710 135440 -297700
rect 138220 -297500 138440 -297490
rect 138220 -297700 138240 -297500
rect 138420 -297700 138440 -297500
rect 138220 -297710 138440 -297700
rect 141220 -297500 141440 -297490
rect 141220 -297700 141240 -297500
rect 141420 -297700 141440 -297500
rect 141220 -297710 141440 -297700
rect 144220 -297500 144440 -297490
rect 144220 -297700 144240 -297500
rect 144420 -297700 144440 -297500
rect 144220 -297710 144440 -297700
rect 147220 -297500 147440 -297490
rect 147220 -297700 147240 -297500
rect 147420 -297700 147440 -297500
rect 147220 -297710 147440 -297700
rect 150220 -297500 150440 -297490
rect 150220 -297700 150240 -297500
rect 150420 -297700 150440 -297500
rect 150220 -297710 150440 -297700
rect 153220 -297500 153440 -297490
rect 153220 -297700 153240 -297500
rect 153420 -297700 153440 -297500
rect 153220 -297710 153440 -297700
rect 156220 -297500 156440 -297490
rect 156220 -297700 156240 -297500
rect 156420 -297700 156440 -297500
rect 156220 -297710 156440 -297700
rect 159220 -297500 159440 -297490
rect 159220 -297700 159240 -297500
rect 159420 -297700 159440 -297500
rect 159220 -297710 159440 -297700
rect 162220 -297500 162440 -297490
rect 162220 -297700 162240 -297500
rect 162420 -297700 162440 -297500
rect 162220 -297710 162440 -297700
rect 165220 -297500 165440 -297490
rect 165220 -297700 165240 -297500
rect 165420 -297700 165440 -297500
rect 165220 -297710 165440 -297700
rect 168220 -297500 168440 -297490
rect 168220 -297700 168240 -297500
rect 168420 -297700 168440 -297500
rect 168220 -297710 168440 -297700
rect 171220 -297500 171440 -297490
rect 171220 -297700 171240 -297500
rect 171420 -297700 171440 -297500
rect 171220 -297710 171440 -297700
rect 174220 -297500 174440 -297490
rect 174220 -297700 174240 -297500
rect 174420 -297700 174440 -297500
rect 174220 -297710 174440 -297700
rect 177220 -297500 177440 -297490
rect 177220 -297700 177240 -297500
rect 177420 -297700 177440 -297500
rect 177220 -297710 177440 -297700
rect 180220 -297500 180440 -297490
rect 180220 -297700 180240 -297500
rect 180420 -297700 180440 -297500
rect 180220 -297710 180440 -297700
rect 183220 -297500 183440 -297490
rect 183220 -297700 183240 -297500
rect 183420 -297700 183440 -297500
rect 183220 -297710 183440 -297700
rect 186220 -297500 186440 -297490
rect 186220 -297700 186240 -297500
rect 186420 -297700 186440 -297500
rect 186220 -297710 186440 -297700
rect 189220 -297500 189440 -297490
rect 189220 -297700 189240 -297500
rect 189420 -297700 189440 -297500
rect 189220 -297710 189440 -297700
rect 192220 -297500 192440 -297490
rect 192220 -297700 192240 -297500
rect 192420 -297700 192440 -297500
rect 192220 -297710 192440 -297700
rect 195220 -297500 195440 -297490
rect 195220 -297700 195240 -297500
rect 195420 -297700 195440 -297500
rect 195220 -297710 195440 -297700
rect 198220 -297500 198440 -297490
rect 198220 -297700 198240 -297500
rect 198420 -297700 198440 -297500
rect 198220 -297710 198440 -297700
rect 201220 -297500 201440 -297490
rect 201220 -297700 201240 -297500
rect 201420 -297700 201440 -297500
rect 201220 -297710 201440 -297700
rect 204220 -297500 204440 -297490
rect 204220 -297700 204240 -297500
rect 204420 -297700 204440 -297500
rect 204220 -297710 204440 -297700
rect 207220 -297500 207440 -297490
rect 207220 -297700 207240 -297500
rect 207420 -297700 207440 -297500
rect 207220 -297710 207440 -297700
rect 210220 -297500 210440 -297490
rect 210220 -297700 210240 -297500
rect 210420 -297700 210440 -297500
rect 210220 -297710 210440 -297700
rect 213220 -297500 213440 -297490
rect 213220 -297700 213240 -297500
rect 213420 -297700 213440 -297500
rect 213220 -297710 213440 -297700
rect 216220 -297500 216440 -297490
rect 216220 -297700 216240 -297500
rect 216420 -297700 216440 -297500
rect 216220 -297710 216440 -297700
rect 219220 -297500 219440 -297490
rect 219220 -297700 219240 -297500
rect 219420 -297700 219440 -297500
rect 219220 -297710 219440 -297700
rect 222220 -297500 222440 -297490
rect 222220 -297700 222240 -297500
rect 222420 -297700 222440 -297500
rect 222220 -297710 222440 -297700
rect 225220 -297500 225440 -297490
rect 225220 -297700 225240 -297500
rect 225420 -297700 225440 -297500
rect 225220 -297710 225440 -297700
rect 228220 -297500 228440 -297490
rect 228220 -297700 228240 -297500
rect 228420 -297700 228440 -297500
rect 228220 -297710 228440 -297700
rect 231220 -297500 231440 -297490
rect 231220 -297700 231240 -297500
rect 231420 -297700 231440 -297500
rect 231220 -297710 231440 -297700
rect 234220 -297500 234440 -297490
rect 234220 -297700 234240 -297500
rect 234420 -297700 234440 -297500
rect 234220 -297710 234440 -297700
rect 237220 -297500 237440 -297490
rect 237220 -297700 237240 -297500
rect 237420 -297700 237440 -297500
rect 237220 -297710 237440 -297700
rect 240220 -297500 240440 -297490
rect 240220 -297700 240240 -297500
rect 240420 -297700 240440 -297500
rect 240220 -297710 240440 -297700
rect 243220 -297500 243440 -297490
rect 243220 -297700 243240 -297500
rect 243420 -297700 243440 -297500
rect 243220 -297710 243440 -297700
rect 246220 -297500 246440 -297490
rect 246220 -297700 246240 -297500
rect 246420 -297700 246440 -297500
rect 246220 -297710 246440 -297700
rect 249220 -297500 249440 -297490
rect 249220 -297700 249240 -297500
rect 249420 -297700 249440 -297500
rect 249220 -297710 249440 -297700
rect 252220 -297500 252440 -297490
rect 252220 -297700 252240 -297500
rect 252420 -297700 252440 -297500
rect 252220 -297710 252440 -297700
rect 255220 -297500 255440 -297490
rect 255220 -297700 255240 -297500
rect 255420 -297700 255440 -297500
rect 255220 -297710 255440 -297700
rect 258220 -297500 258440 -297490
rect 258220 -297700 258240 -297500
rect 258420 -297700 258440 -297500
rect 258220 -297710 258440 -297700
rect 261220 -297500 261440 -297490
rect 261220 -297700 261240 -297500
rect 261420 -297700 261440 -297500
rect 261220 -297710 261440 -297700
rect 264220 -297500 264440 -297490
rect 264220 -297700 264240 -297500
rect 264420 -297700 264440 -297500
rect 264220 -297710 264440 -297700
rect 267220 -297500 267440 -297490
rect 267220 -297700 267240 -297500
rect 267420 -297700 267440 -297500
rect 267220 -297710 267440 -297700
rect 270220 -297500 270440 -297490
rect 270220 -297700 270240 -297500
rect 270420 -297700 270440 -297500
rect 270220 -297710 270440 -297700
rect 273220 -297500 273440 -297490
rect 273220 -297700 273240 -297500
rect 273420 -297700 273440 -297500
rect 273220 -297710 273440 -297700
rect 276220 -297500 276440 -297490
rect 276220 -297700 276240 -297500
rect 276420 -297700 276440 -297500
rect 276220 -297710 276440 -297700
rect 279220 -297500 279440 -297490
rect 279220 -297700 279240 -297500
rect 279420 -297700 279440 -297500
rect 279220 -297710 279440 -297700
rect 282220 -297500 282440 -297490
rect 282220 -297700 282240 -297500
rect 282420 -297700 282440 -297500
rect 282220 -297710 282440 -297700
rect 285220 -297500 285440 -297490
rect 285220 -297700 285240 -297500
rect 285420 -297700 285440 -297500
rect 285220 -297710 285440 -297700
rect 288220 -297500 288440 -297490
rect 288220 -297700 288240 -297500
rect 288420 -297700 288440 -297500
rect 288220 -297710 288440 -297700
rect 291220 -297500 291440 -297490
rect 291220 -297700 291240 -297500
rect 291420 -297700 291440 -297500
rect 291220 -297710 291440 -297700
rect 294220 -297500 294440 -297490
rect 294220 -297700 294240 -297500
rect 294420 -297700 294440 -297500
rect 294220 -297710 294440 -297700
rect 297220 -297500 297440 -297490
rect 297220 -297700 297240 -297500
rect 297420 -297700 297440 -297500
rect 297220 -297710 297440 -297700
<< via3 >>
rect 490 3560 580 3650
rect 3490 3560 3580 3650
rect 6490 3560 6580 3650
rect 9490 3560 9580 3650
rect 12490 3560 12580 3650
rect 15490 3560 15580 3650
rect 18490 3560 18580 3650
rect 21490 3560 21580 3650
rect 24490 3560 24580 3650
rect 27490 3560 27580 3650
rect 30490 3560 30580 3650
rect 33490 3560 33580 3650
rect 36490 3560 36580 3650
rect 39490 3560 39580 3650
rect 42490 3560 42580 3650
rect 45490 3560 45580 3650
rect 48490 3560 48580 3650
rect 51490 3560 51580 3650
rect 54490 3560 54580 3650
rect 57490 3560 57580 3650
rect 60490 3560 60580 3650
rect 63490 3560 63580 3650
rect 66490 3560 66580 3650
rect 69490 3560 69580 3650
rect 72490 3560 72580 3650
rect 75490 3560 75580 3650
rect 78490 3560 78580 3650
rect 81490 3560 81580 3650
rect 84490 3560 84580 3650
rect 87490 3560 87580 3650
rect 90490 3560 90580 3650
rect 93490 3560 93580 3650
rect 96490 3560 96580 3650
rect 99490 3560 99580 3650
rect 102490 3560 102580 3650
rect 105490 3560 105580 3650
rect 108490 3560 108580 3650
rect 111490 3560 111580 3650
rect 114490 3560 114580 3650
rect 117490 3560 117580 3650
rect 120490 3560 120580 3650
rect 123490 3560 123580 3650
rect 126490 3560 126580 3650
rect 129490 3560 129580 3650
rect 132490 3560 132580 3650
rect 135490 3560 135580 3650
rect 138490 3560 138580 3650
rect 141490 3560 141580 3650
rect 144490 3560 144580 3650
rect 147490 3560 147580 3650
rect 150490 3560 150580 3650
rect 153490 3560 153580 3650
rect 156490 3560 156580 3650
rect 159490 3560 159580 3650
rect 162490 3560 162580 3650
rect 165490 3560 165580 3650
rect 168490 3560 168580 3650
rect 171490 3560 171580 3650
rect 174490 3560 174580 3650
rect 177490 3560 177580 3650
rect 180490 3560 180580 3650
rect 183490 3560 183580 3650
rect 186490 3560 186580 3650
rect 189490 3560 189580 3650
rect 192490 3560 192580 3650
rect 195490 3560 195580 3650
rect 198490 3560 198580 3650
rect 201490 3560 201580 3650
rect 204490 3560 204580 3650
rect 207490 3560 207580 3650
rect 210490 3560 210580 3650
rect 213490 3560 213580 3650
rect 216490 3560 216580 3650
rect 219490 3560 219580 3650
rect 222490 3560 222580 3650
rect 225490 3560 225580 3650
rect 228490 3560 228580 3650
rect 231490 3560 231580 3650
rect 234490 3560 234580 3650
rect 237490 3560 237580 3650
rect 240490 3560 240580 3650
rect 243490 3560 243580 3650
rect 246490 3560 246580 3650
rect 249490 3560 249580 3650
rect 252490 3560 252580 3650
rect 255490 3560 255580 3650
rect 258490 3560 258580 3650
rect 261490 3560 261580 3650
rect 264490 3560 264580 3650
rect 267490 3560 267580 3650
rect 270490 3560 270580 3650
rect 273490 3560 273580 3650
rect 276490 3560 276580 3650
rect 279490 3560 279580 3650
rect 282490 3560 282580 3650
rect 285490 3560 285580 3650
rect 288490 3560 288580 3650
rect 291490 3560 291580 3650
rect 294490 3560 294580 3650
rect 297490 3560 297580 3650
rect -470 2470 -380 2540
rect -470 -530 -380 -460
rect -470 -3530 -380 -3460
rect -470 -6530 -380 -6460
rect -470 -9530 -380 -9460
rect -470 -12530 -380 -12460
rect -470 -15530 -380 -15460
rect -470 -18530 -380 -18460
rect -470 -21530 -380 -21460
rect -470 -24530 -380 -24460
rect -470 -27530 -380 -27460
rect -470 -30530 -380 -30460
rect -470 -33530 -380 -33460
rect -470 -36530 -380 -36460
rect -470 -39530 -380 -39460
rect -470 -42530 -380 -42460
rect -470 -45530 -380 -45460
rect -470 -48530 -380 -48460
rect -470 -51530 -380 -51460
rect -470 -54530 -380 -54460
rect -470 -57530 -380 -57460
rect -470 -60530 -380 -60460
rect -470 -63530 -380 -63460
rect -470 -66530 -380 -66460
rect -470 -69530 -380 -69460
rect -470 -72530 -380 -72460
rect -470 -75530 -380 -75460
rect -470 -78530 -380 -78460
rect -470 -81530 -380 -81460
rect -470 -84530 -380 -84460
rect -470 -87530 -380 -87460
rect -470 -90530 -380 -90460
rect -470 -93530 -380 -93460
rect -470 -96530 -380 -96460
rect -470 -99530 -380 -99460
rect -470 -102530 -380 -102460
rect -470 -105530 -380 -105460
rect -470 -108530 -380 -108460
rect -470 -111530 -380 -111460
rect -470 -114530 -380 -114460
rect -470 -117530 -380 -117460
rect -470 -120530 -380 -120460
rect -470 -123530 -380 -123460
rect -470 -126530 -380 -126460
rect -470 -129530 -380 -129460
rect -470 -132530 -380 -132460
rect -470 -135530 -380 -135460
rect -470 -138530 -380 -138460
rect -470 -141530 -380 -141460
rect -470 -144530 -380 -144460
rect -470 -147530 -380 -147460
rect -470 -150530 -380 -150460
rect -470 -153530 -380 -153460
rect -470 -156530 -380 -156460
rect -470 -159530 -380 -159460
rect -470 -162530 -380 -162460
rect -470 -165530 -380 -165460
rect -470 -168530 -380 -168460
rect -470 -171530 -380 -171460
rect -470 -174530 -380 -174460
rect -470 -177530 -380 -177460
rect -470 -180530 -380 -180460
rect -470 -183530 -380 -183460
rect -470 -186530 -380 -186460
rect -470 -189530 -380 -189460
rect -470 -192530 -380 -192460
rect -470 -195530 -380 -195460
rect -470 -198530 -380 -198460
rect -470 -201530 -380 -201460
rect -470 -204530 -380 -204460
rect -470 -207530 -380 -207460
rect -470 -210530 -380 -210460
rect -470 -213530 -380 -213460
rect -470 -216530 -380 -216460
rect -470 -219530 -380 -219460
rect -470 -222530 -380 -222460
rect -470 -225530 -380 -225460
rect -470 -228530 -380 -228460
rect -470 -231530 -380 -231460
rect -470 -234530 -380 -234460
rect -470 -237530 -380 -237460
rect -470 -240530 -380 -240460
rect -470 -243530 -380 -243460
rect -470 -246530 -380 -246460
rect -470 -249530 -380 -249460
rect -470 -252530 -380 -252460
rect -470 -255530 -380 -255460
rect -470 -258530 -380 -258460
rect -470 -261530 -380 -261460
rect -470 -264530 -380 -264460
rect -470 -267530 -380 -267460
rect -470 -270530 -380 -270460
rect -470 -273530 -380 -273460
rect -470 -276530 -380 -276460
rect -470 -279530 -380 -279460
rect -470 -282530 -380 -282460
rect -470 -285530 -380 -285460
rect -470 -288530 -380 -288460
rect -470 -291530 -380 -291460
rect -470 -294530 -380 -294460
rect 560 -297180 2760 -297080
rect 3560 -297180 5760 -297080
rect 6560 -297180 8760 -297080
rect 9560 -297180 11760 -297080
rect 12560 -297180 14760 -297080
rect 15560 -297180 17760 -297080
rect 18560 -297180 20760 -297080
rect 21560 -297180 23760 -297080
rect 24560 -297180 26760 -297080
rect 27560 -297180 29760 -297080
rect 30560 -297180 32760 -297080
rect 33560 -297180 35760 -297080
rect 36560 -297180 38760 -297080
rect 39560 -297180 41760 -297080
rect 42560 -297180 44760 -297080
rect 45560 -297180 47760 -297080
rect 48560 -297180 50760 -297080
rect 51560 -297180 53760 -297080
rect 54560 -297180 56760 -297080
rect 57560 -297180 59760 -297080
rect 60560 -297180 62760 -297080
rect 63560 -297180 65760 -297080
rect 66560 -297180 68760 -297080
rect 69560 -297180 71760 -297080
rect 72560 -297180 74760 -297080
rect 75560 -297180 77760 -297080
rect 78560 -297180 80760 -297080
rect 81560 -297180 83760 -297080
rect 84560 -297180 86760 -297080
rect 87560 -297180 89760 -297080
rect 90560 -297180 92760 -297080
rect 93560 -297180 95760 -297080
rect 96560 -297180 98760 -297080
rect 99560 -297180 101760 -297080
rect 102560 -297180 104760 -297080
rect 105560 -297180 107760 -297080
rect 108560 -297180 110760 -297080
rect 111560 -297180 113760 -297080
rect 114560 -297180 116760 -297080
rect 117560 -297180 119760 -297080
rect 120560 -297180 122760 -297080
rect 123560 -297180 125760 -297080
rect 126560 -297180 128760 -297080
rect 129560 -297180 131760 -297080
rect 132560 -297180 134760 -297080
rect 135560 -297180 137760 -297080
rect 138560 -297180 140760 -297080
rect 141560 -297180 143760 -297080
rect 144560 -297180 146760 -297080
rect 147560 -297180 149760 -297080
rect 150560 -297180 152760 -297080
rect 153560 -297180 155760 -297080
rect 156560 -297180 158760 -297080
rect 159560 -297180 161760 -297080
rect 162560 -297180 164760 -297080
rect 165560 -297180 167760 -297080
rect 168560 -297180 170760 -297080
rect 171560 -297180 173760 -297080
rect 174560 -297180 176760 -297080
rect 177560 -297180 179760 -297080
rect 180560 -297180 182760 -297080
rect 183560 -297180 185760 -297080
rect 186560 -297180 188760 -297080
rect 189560 -297180 191760 -297080
rect 192560 -297180 194760 -297080
rect 195560 -297180 197760 -297080
rect 198560 -297180 200760 -297080
rect 201560 -297180 203760 -297080
rect 204560 -297180 206760 -297080
rect 207560 -297180 209760 -297080
rect 210560 -297180 212760 -297080
rect 213560 -297180 215760 -297080
rect 216560 -297180 218760 -297080
rect 219560 -297180 221760 -297080
rect 222560 -297180 224760 -297080
rect 225560 -297180 227760 -297080
rect 228560 -297180 230760 -297080
rect 231560 -297180 233760 -297080
rect 234560 -297180 236760 -297080
rect 237560 -297180 239760 -297080
rect 240560 -297180 242760 -297080
rect 243560 -297180 245760 -297080
rect 246560 -297180 248760 -297080
rect 249560 -297180 251760 -297080
rect 252560 -297180 254760 -297080
rect 255560 -297180 257760 -297080
rect 258560 -297180 260760 -297080
rect 261560 -297180 263760 -297080
rect 264560 -297180 266760 -297080
rect 267560 -297180 269760 -297080
rect 270560 -297180 272760 -297080
rect 273560 -297180 275760 -297080
rect 276560 -297180 278760 -297080
rect 279560 -297180 281760 -297080
rect 282560 -297180 284760 -297080
rect 285560 -297180 287760 -297080
rect 288560 -297180 290760 -297080
rect 291560 -297180 293760 -297080
rect 294560 -297180 296760 -297080
rect 297560 -297180 299760 -297080
rect 240 -297700 420 -297500
rect 3240 -297700 3420 -297500
rect 6240 -297700 6420 -297500
rect 9240 -297700 9420 -297500
rect 12240 -297700 12420 -297500
rect 15240 -297700 15420 -297500
rect 18240 -297700 18420 -297500
rect 21240 -297700 21420 -297500
rect 24240 -297700 24420 -297500
rect 27240 -297700 27420 -297500
rect 30240 -297700 30420 -297500
rect 33240 -297700 33420 -297500
rect 36240 -297700 36420 -297500
rect 39240 -297700 39420 -297500
rect 42240 -297700 42420 -297500
rect 45240 -297700 45420 -297500
rect 48240 -297700 48420 -297500
rect 51240 -297700 51420 -297500
rect 54240 -297700 54420 -297500
rect 57240 -297700 57420 -297500
rect 60240 -297700 60420 -297500
rect 63240 -297700 63420 -297500
rect 66240 -297700 66420 -297500
rect 69240 -297700 69420 -297500
rect 72240 -297700 72420 -297500
rect 75240 -297700 75420 -297500
rect 78240 -297700 78420 -297500
rect 81240 -297700 81420 -297500
rect 84240 -297700 84420 -297500
rect 87240 -297700 87420 -297500
rect 90240 -297700 90420 -297500
rect 93240 -297700 93420 -297500
rect 96240 -297700 96420 -297500
rect 99240 -297700 99420 -297500
rect 102240 -297700 102420 -297500
rect 105240 -297700 105420 -297500
rect 108240 -297700 108420 -297500
rect 111240 -297700 111420 -297500
rect 114240 -297700 114420 -297500
rect 117240 -297700 117420 -297500
rect 120240 -297700 120420 -297500
rect 123240 -297700 123420 -297500
rect 126240 -297700 126420 -297500
rect 129240 -297700 129420 -297500
rect 132240 -297700 132420 -297500
rect 135240 -297700 135420 -297500
rect 138240 -297700 138420 -297500
rect 141240 -297700 141420 -297500
rect 144240 -297700 144420 -297500
rect 147240 -297700 147420 -297500
rect 150240 -297700 150420 -297500
rect 153240 -297700 153420 -297500
rect 156240 -297700 156420 -297500
rect 159240 -297700 159420 -297500
rect 162240 -297700 162420 -297500
rect 165240 -297700 165420 -297500
rect 168240 -297700 168420 -297500
rect 171240 -297700 171420 -297500
rect 174240 -297700 174420 -297500
rect 177240 -297700 177420 -297500
rect 180240 -297700 180420 -297500
rect 183240 -297700 183420 -297500
rect 186240 -297700 186420 -297500
rect 189240 -297700 189420 -297500
rect 192240 -297700 192420 -297500
rect 195240 -297700 195420 -297500
rect 198240 -297700 198420 -297500
rect 201240 -297700 201420 -297500
rect 204240 -297700 204420 -297500
rect 207240 -297700 207420 -297500
rect 210240 -297700 210420 -297500
rect 213240 -297700 213420 -297500
rect 216240 -297700 216420 -297500
rect 219240 -297700 219420 -297500
rect 222240 -297700 222420 -297500
rect 225240 -297700 225420 -297500
rect 228240 -297700 228420 -297500
rect 231240 -297700 231420 -297500
rect 234240 -297700 234420 -297500
rect 237240 -297700 237420 -297500
rect 240240 -297700 240420 -297500
rect 243240 -297700 243420 -297500
rect 246240 -297700 246420 -297500
rect 249240 -297700 249420 -297500
rect 252240 -297700 252420 -297500
rect 255240 -297700 255420 -297500
rect 258240 -297700 258420 -297500
rect 261240 -297700 261420 -297500
rect 264240 -297700 264420 -297500
rect 267240 -297700 267420 -297500
rect 270240 -297700 270420 -297500
rect 273240 -297700 273420 -297500
rect 276240 -297700 276420 -297500
rect 279240 -297700 279420 -297500
rect 282240 -297700 282420 -297500
rect 285240 -297700 285420 -297500
rect 288240 -297700 288420 -297500
rect 291240 -297700 291420 -297500
rect 294240 -297700 294420 -297500
rect 297240 -297700 297420 -297500
<< metal4 >>
rect -3000 3650 299200 3660
rect -3000 3560 490 3650
rect 580 3560 3490 3650
rect 3580 3560 6490 3650
rect 6580 3560 9490 3650
rect 9580 3560 12490 3650
rect 12580 3560 15490 3650
rect 15580 3560 18490 3650
rect 18580 3560 21490 3650
rect 21580 3560 24490 3650
rect 24580 3560 27490 3650
rect 27580 3560 30490 3650
rect 30580 3560 33490 3650
rect 33580 3560 36490 3650
rect 36580 3560 39490 3650
rect 39580 3560 42490 3650
rect 42580 3560 45490 3650
rect 45580 3560 48490 3650
rect 48580 3560 51490 3650
rect 51580 3560 54490 3650
rect 54580 3560 57490 3650
rect 57580 3560 60490 3650
rect 60580 3560 63490 3650
rect 63580 3560 66490 3650
rect 66580 3560 69490 3650
rect 69580 3560 72490 3650
rect 72580 3560 75490 3650
rect 75580 3560 78490 3650
rect 78580 3560 81490 3650
rect 81580 3560 84490 3650
rect 84580 3560 87490 3650
rect 87580 3560 90490 3650
rect 90580 3560 93490 3650
rect 93580 3560 96490 3650
rect 96580 3560 99490 3650
rect 99580 3560 102490 3650
rect 102580 3560 105490 3650
rect 105580 3560 108490 3650
rect 108580 3560 111490 3650
rect 111580 3560 114490 3650
rect 114580 3560 117490 3650
rect 117580 3560 120490 3650
rect 120580 3560 123490 3650
rect 123580 3560 126490 3650
rect 126580 3560 129490 3650
rect 129580 3560 132490 3650
rect 132580 3560 135490 3650
rect 135580 3560 138490 3650
rect 138580 3560 141490 3650
rect 141580 3560 144490 3650
rect 144580 3560 147490 3650
rect 147580 3560 150490 3650
rect 150580 3560 153490 3650
rect 153580 3560 156490 3650
rect 156580 3560 159490 3650
rect 159580 3560 162490 3650
rect 162580 3560 165490 3650
rect 165580 3560 168490 3650
rect 168580 3560 171490 3650
rect 171580 3560 174490 3650
rect 174580 3560 177490 3650
rect 177580 3560 180490 3650
rect 180580 3560 183490 3650
rect 183580 3560 186490 3650
rect 186580 3560 189490 3650
rect 189580 3560 192490 3650
rect 192580 3560 195490 3650
rect 195580 3560 198490 3650
rect 198580 3560 201490 3650
rect 201580 3560 204490 3650
rect 204580 3560 207490 3650
rect 207580 3560 210490 3650
rect 210580 3560 213490 3650
rect 213580 3560 216490 3650
rect 216580 3560 219490 3650
rect 219580 3560 222490 3650
rect 222580 3560 225490 3650
rect 225580 3560 228490 3650
rect 228580 3560 231490 3650
rect 231580 3560 234490 3650
rect 234580 3560 237490 3650
rect 237580 3560 240490 3650
rect 240580 3560 243490 3650
rect 243580 3560 246490 3650
rect 246580 3560 249490 3650
rect 249580 3560 252490 3650
rect 252580 3560 255490 3650
rect 255580 3560 258490 3650
rect 258580 3560 261490 3650
rect 261580 3560 264490 3650
rect 264580 3560 267490 3650
rect 267580 3560 270490 3650
rect 270580 3560 273490 3650
rect 273580 3560 276490 3650
rect 276580 3560 279490 3650
rect 279580 3560 282490 3650
rect 282580 3560 285490 3650
rect 285580 3560 288490 3650
rect 288580 3560 291490 3650
rect 291580 3560 294490 3650
rect 294580 3560 297490 3650
rect 297580 3560 299200 3650
rect -3000 3550 299200 3560
rect -480 2540 -370 2600
rect -480 2470 -470 2540
rect -380 2470 -370 2540
rect -480 -460 -370 2470
rect -480 -530 -470 -460
rect -380 -530 -370 -460
rect -480 -3460 -370 -530
rect -480 -3530 -470 -3460
rect -380 -3530 -370 -3460
rect -480 -6460 -370 -3530
rect -480 -6530 -470 -6460
rect -380 -6530 -370 -6460
rect -480 -9460 -370 -6530
rect -480 -9530 -470 -9460
rect -380 -9530 -370 -9460
rect -480 -12460 -370 -9530
rect -480 -12530 -470 -12460
rect -380 -12530 -370 -12460
rect -480 -15460 -370 -12530
rect -480 -15530 -470 -15460
rect -380 -15530 -370 -15460
rect -480 -18460 -370 -15530
rect -480 -18530 -470 -18460
rect -380 -18530 -370 -18460
rect -480 -21460 -370 -18530
rect -480 -21530 -470 -21460
rect -380 -21530 -370 -21460
rect -480 -24460 -370 -21530
rect -480 -24530 -470 -24460
rect -380 -24530 -370 -24460
rect -480 -27460 -370 -24530
rect -480 -27530 -470 -27460
rect -380 -27530 -370 -27460
rect -480 -30460 -370 -27530
rect -480 -30530 -470 -30460
rect -380 -30530 -370 -30460
rect -480 -33460 -370 -30530
rect -480 -33530 -470 -33460
rect -380 -33530 -370 -33460
rect -480 -36460 -370 -33530
rect -480 -36530 -470 -36460
rect -380 -36530 -370 -36460
rect -480 -39460 -370 -36530
rect -480 -39530 -470 -39460
rect -380 -39530 -370 -39460
rect -480 -42460 -370 -39530
rect -480 -42530 -470 -42460
rect -380 -42530 -370 -42460
rect -480 -45460 -370 -42530
rect -480 -45530 -470 -45460
rect -380 -45530 -370 -45460
rect -480 -48460 -370 -45530
rect -480 -48530 -470 -48460
rect -380 -48530 -370 -48460
rect -480 -51460 -370 -48530
rect -480 -51530 -470 -51460
rect -380 -51530 -370 -51460
rect -480 -54460 -370 -51530
rect -480 -54530 -470 -54460
rect -380 -54530 -370 -54460
rect -480 -57460 -370 -54530
rect -480 -57530 -470 -57460
rect -380 -57530 -370 -57460
rect -480 -60460 -370 -57530
rect -480 -60530 -470 -60460
rect -380 -60530 -370 -60460
rect -480 -63460 -370 -60530
rect -480 -63530 -470 -63460
rect -380 -63530 -370 -63460
rect -480 -66460 -370 -63530
rect -480 -66530 -470 -66460
rect -380 -66530 -370 -66460
rect -480 -69460 -370 -66530
rect -480 -69530 -470 -69460
rect -380 -69530 -370 -69460
rect -480 -72460 -370 -69530
rect -480 -72530 -470 -72460
rect -380 -72530 -370 -72460
rect -480 -75460 -370 -72530
rect -480 -75530 -470 -75460
rect -380 -75530 -370 -75460
rect -480 -78460 -370 -75530
rect -480 -78530 -470 -78460
rect -380 -78530 -370 -78460
rect -480 -81460 -370 -78530
rect -480 -81530 -470 -81460
rect -380 -81530 -370 -81460
rect -480 -84460 -370 -81530
rect -480 -84530 -470 -84460
rect -380 -84530 -370 -84460
rect -480 -87460 -370 -84530
rect -480 -87530 -470 -87460
rect -380 -87530 -370 -87460
rect -480 -90460 -370 -87530
rect -480 -90530 -470 -90460
rect -380 -90530 -370 -90460
rect -480 -93460 -370 -90530
rect -480 -93530 -470 -93460
rect -380 -93530 -370 -93460
rect -480 -96460 -370 -93530
rect -480 -96530 -470 -96460
rect -380 -96530 -370 -96460
rect -480 -99460 -370 -96530
rect -480 -99530 -470 -99460
rect -380 -99530 -370 -99460
rect -480 -102460 -370 -99530
rect -480 -102530 -470 -102460
rect -380 -102530 -370 -102460
rect -480 -105460 -370 -102530
rect -480 -105530 -470 -105460
rect -380 -105530 -370 -105460
rect -480 -108460 -370 -105530
rect -480 -108530 -470 -108460
rect -380 -108530 -370 -108460
rect -480 -111460 -370 -108530
rect -480 -111530 -470 -111460
rect -380 -111530 -370 -111460
rect -480 -114460 -370 -111530
rect -480 -114530 -470 -114460
rect -380 -114530 -370 -114460
rect -480 -117460 -370 -114530
rect -480 -117530 -470 -117460
rect -380 -117530 -370 -117460
rect -480 -120460 -370 -117530
rect -480 -120530 -470 -120460
rect -380 -120530 -370 -120460
rect -480 -123460 -370 -120530
rect -480 -123530 -470 -123460
rect -380 -123530 -370 -123460
rect -480 -126460 -370 -123530
rect -480 -126530 -470 -126460
rect -380 -126530 -370 -126460
rect -480 -129460 -370 -126530
rect -480 -129530 -470 -129460
rect -380 -129530 -370 -129460
rect -480 -132460 -370 -129530
rect -480 -132530 -470 -132460
rect -380 -132530 -370 -132460
rect -480 -135460 -370 -132530
rect -480 -135530 -470 -135460
rect -380 -135530 -370 -135460
rect -480 -138460 -370 -135530
rect -480 -138530 -470 -138460
rect -380 -138530 -370 -138460
rect -480 -141460 -370 -138530
rect -480 -141530 -470 -141460
rect -380 -141530 -370 -141460
rect -480 -144460 -370 -141530
rect -480 -144530 -470 -144460
rect -380 -144530 -370 -144460
rect -480 -147460 -370 -144530
rect -480 -147530 -470 -147460
rect -380 -147530 -370 -147460
rect -480 -150460 -370 -147530
rect -480 -150530 -470 -150460
rect -380 -150530 -370 -150460
rect -480 -153460 -370 -150530
rect -480 -153530 -470 -153460
rect -380 -153530 -370 -153460
rect -480 -156460 -370 -153530
rect -480 -156530 -470 -156460
rect -380 -156530 -370 -156460
rect -480 -159460 -370 -156530
rect -480 -159530 -470 -159460
rect -380 -159530 -370 -159460
rect -480 -162460 -370 -159530
rect -480 -162530 -470 -162460
rect -380 -162530 -370 -162460
rect -480 -165460 -370 -162530
rect -480 -165530 -470 -165460
rect -380 -165530 -370 -165460
rect -480 -168460 -370 -165530
rect -480 -168530 -470 -168460
rect -380 -168530 -370 -168460
rect -480 -171460 -370 -168530
rect -480 -171530 -470 -171460
rect -380 -171530 -370 -171460
rect -480 -174460 -370 -171530
rect -480 -174530 -470 -174460
rect -380 -174530 -370 -174460
rect -480 -177460 -370 -174530
rect -480 -177530 -470 -177460
rect -380 -177530 -370 -177460
rect -480 -180460 -370 -177530
rect -480 -180530 -470 -180460
rect -380 -180530 -370 -180460
rect -480 -183460 -370 -180530
rect -480 -183530 -470 -183460
rect -380 -183530 -370 -183460
rect -480 -186460 -370 -183530
rect -480 -186530 -470 -186460
rect -380 -186530 -370 -186460
rect -480 -189460 -370 -186530
rect -480 -189530 -470 -189460
rect -380 -189530 -370 -189460
rect -480 -192460 -370 -189530
rect -480 -192530 -470 -192460
rect -380 -192530 -370 -192460
rect -480 -195460 -370 -192530
rect -480 -195530 -470 -195460
rect -380 -195530 -370 -195460
rect -480 -198460 -370 -195530
rect -480 -198530 -470 -198460
rect -380 -198530 -370 -198460
rect -480 -201460 -370 -198530
rect -480 -201530 -470 -201460
rect -380 -201530 -370 -201460
rect -480 -204460 -370 -201530
rect -480 -204530 -470 -204460
rect -380 -204530 -370 -204460
rect -480 -207460 -370 -204530
rect -480 -207530 -470 -207460
rect -380 -207530 -370 -207460
rect -480 -210460 -370 -207530
rect -480 -210530 -470 -210460
rect -380 -210530 -370 -210460
rect -480 -213460 -370 -210530
rect -480 -213530 -470 -213460
rect -380 -213530 -370 -213460
rect -480 -216460 -370 -213530
rect -480 -216530 -470 -216460
rect -380 -216530 -370 -216460
rect -480 -219460 -370 -216530
rect -480 -219530 -470 -219460
rect -380 -219530 -370 -219460
rect -480 -222460 -370 -219530
rect -480 -222530 -470 -222460
rect -380 -222530 -370 -222460
rect -480 -225460 -370 -222530
rect -480 -225530 -470 -225460
rect -380 -225530 -370 -225460
rect -480 -228460 -370 -225530
rect -480 -228530 -470 -228460
rect -380 -228530 -370 -228460
rect -480 -231460 -370 -228530
rect -480 -231530 -470 -231460
rect -380 -231530 -370 -231460
rect -480 -234460 -370 -231530
rect -480 -234530 -470 -234460
rect -380 -234530 -370 -234460
rect -480 -237460 -370 -234530
rect -480 -237530 -470 -237460
rect -380 -237530 -370 -237460
rect -480 -240460 -370 -237530
rect -480 -240530 -470 -240460
rect -380 -240530 -370 -240460
rect -480 -243460 -370 -240530
rect -480 -243530 -470 -243460
rect -380 -243530 -370 -243460
rect -480 -246460 -370 -243530
rect -480 -246530 -470 -246460
rect -380 -246530 -370 -246460
rect -480 -249460 -370 -246530
rect -480 -249530 -470 -249460
rect -380 -249530 -370 -249460
rect -480 -252460 -370 -249530
rect -480 -252530 -470 -252460
rect -380 -252530 -370 -252460
rect -480 -255460 -370 -252530
rect -480 -255530 -470 -255460
rect -380 -255530 -370 -255460
rect -480 -258460 -370 -255530
rect -480 -258530 -470 -258460
rect -380 -258530 -370 -258460
rect -480 -261460 -370 -258530
rect -480 -261530 -470 -261460
rect -380 -261530 -370 -261460
rect -480 -264460 -370 -261530
rect -480 -264530 -470 -264460
rect -380 -264530 -370 -264460
rect -480 -267460 -370 -264530
rect -480 -267530 -470 -267460
rect -380 -267530 -370 -267460
rect -480 -270460 -370 -267530
rect -480 -270530 -470 -270460
rect -380 -270530 -370 -270460
rect -480 -273460 -370 -270530
rect -480 -273530 -470 -273460
rect -380 -273530 -370 -273460
rect -480 -276460 -370 -273530
rect -480 -276530 -470 -276460
rect -380 -276530 -370 -276460
rect -480 -279460 -370 -276530
rect -480 -279530 -470 -279460
rect -380 -279530 -370 -279460
rect -480 -282460 -370 -279530
rect -480 -282530 -470 -282460
rect -380 -282530 -370 -282460
rect -480 -285460 -370 -282530
rect -480 -285530 -470 -285460
rect -380 -285530 -370 -285460
rect -480 -288460 -370 -285530
rect -480 -288530 -470 -288460
rect -380 -288530 -370 -288460
rect -480 -291460 -370 -288530
rect -480 -291530 -470 -291460
rect -380 -291530 -370 -291460
rect -480 -294460 -370 -291530
rect -480 -294530 -470 -294460
rect -380 -294530 -370 -294460
rect -480 -298600 -370 -294530
rect 2630 -297060 2780 -297000
rect 5630 -297060 5780 -297000
rect 8630 -297060 8780 -297000
rect 11630 -297060 11780 -297000
rect 14630 -297060 14780 -297000
rect 17630 -297060 17780 -297000
rect 20630 -297060 20780 -297000
rect 23630 -297060 23780 -297000
rect 26630 -297060 26780 -297000
rect 29630 -297060 29780 -297000
rect 32630 -297060 32780 -297000
rect 35630 -297060 35780 -297000
rect 38630 -297060 38780 -297000
rect 41630 -297060 41780 -297000
rect 44630 -297060 44780 -297000
rect 47630 -297060 47780 -297000
rect 50630 -297060 50780 -297000
rect 53630 -297060 53780 -297000
rect 56630 -297060 56780 -297000
rect 59630 -297060 59780 -297000
rect 62630 -297060 62780 -297000
rect 65630 -297060 65780 -297000
rect 68630 -297060 68780 -297000
rect 71630 -297060 71780 -297000
rect 74630 -297060 74780 -297000
rect 77630 -297060 77780 -297000
rect 80630 -297060 80780 -297000
rect 83630 -297060 83780 -297000
rect 86630 -297060 86780 -297000
rect 89630 -297060 89780 -297000
rect 92630 -297060 92780 -297000
rect 95630 -297060 95780 -297000
rect 98630 -297060 98780 -297000
rect 101630 -297060 101780 -297000
rect 104630 -297060 104780 -297000
rect 107630 -297060 107780 -297000
rect 110630 -297060 110780 -297000
rect 113630 -297060 113780 -297000
rect 116630 -297060 116780 -297000
rect 119630 -297060 119780 -297000
rect 122630 -297060 122780 -297000
rect 125630 -297060 125780 -297000
rect 128630 -297060 128780 -297000
rect 131630 -297060 131780 -297000
rect 134630 -297060 134780 -297000
rect 137630 -297060 137780 -297000
rect 140630 -297060 140780 -297000
rect 143630 -297060 143780 -297000
rect 146630 -297060 146780 -297000
rect 149630 -297060 149780 -297000
rect 152630 -297060 152780 -297000
rect 155630 -297060 155780 -297000
rect 158630 -297060 158780 -297000
rect 161630 -297060 161780 -297000
rect 164630 -297060 164780 -297000
rect 167630 -297060 167780 -297000
rect 170630 -297060 170780 -297000
rect 173630 -297060 173780 -297000
rect 176630 -297060 176780 -297000
rect 179630 -297060 179780 -297000
rect 182630 -297060 182780 -297000
rect 185630 -297060 185780 -297000
rect 188630 -297060 188780 -297000
rect 191630 -297060 191780 -297000
rect 194630 -297060 194780 -297000
rect 197630 -297060 197780 -297000
rect 200630 -297060 200780 -297000
rect 203630 -297060 203780 -297000
rect 206630 -297060 206780 -297000
rect 209630 -297060 209780 -297000
rect 212630 -297060 212780 -297000
rect 215630 -297060 215780 -297000
rect 218630 -297060 218780 -297000
rect 221630 -297060 221780 -297000
rect 224630 -297060 224780 -297000
rect 227630 -297060 227780 -297000
rect 230630 -297060 230780 -297000
rect 233630 -297060 233780 -297000
rect 236630 -297060 236780 -297000
rect 239630 -297060 239780 -297000
rect 242630 -297060 242780 -297000
rect 245630 -297060 245780 -297000
rect 248630 -297060 248780 -297000
rect 251630 -297060 251780 -297000
rect 254630 -297060 254780 -297000
rect 257630 -297060 257780 -297000
rect 260630 -297060 260780 -297000
rect 263630 -297060 263780 -297000
rect 266630 -297060 266780 -297000
rect 269630 -297060 269780 -297000
rect 272630 -297060 272780 -297000
rect 275630 -297060 275780 -297000
rect 278630 -297060 278780 -297000
rect 281630 -297060 281780 -297000
rect 284630 -297060 284780 -297000
rect 287630 -297060 287780 -297000
rect 290630 -297060 290780 -297000
rect 293630 -297060 293780 -297000
rect 296630 -297060 296780 -297000
rect 299630 -297060 299780 -297000
rect 540 -297080 2780 -297060
rect 540 -297180 560 -297080
rect 2760 -297180 2780 -297080
rect 540 -297200 2780 -297180
rect 3540 -297080 5780 -297060
rect 3540 -297180 3560 -297080
rect 5760 -297180 5780 -297080
rect 3540 -297200 5780 -297180
rect 6540 -297080 8780 -297060
rect 6540 -297180 6560 -297080
rect 8760 -297180 8780 -297080
rect 6540 -297200 8780 -297180
rect 9540 -297080 11780 -297060
rect 9540 -297180 9560 -297080
rect 11760 -297180 11780 -297080
rect 9540 -297200 11780 -297180
rect 12540 -297080 14780 -297060
rect 12540 -297180 12560 -297080
rect 14760 -297180 14780 -297080
rect 12540 -297200 14780 -297180
rect 15540 -297080 17780 -297060
rect 15540 -297180 15560 -297080
rect 17760 -297180 17780 -297080
rect 15540 -297200 17780 -297180
rect 18540 -297080 20780 -297060
rect 18540 -297180 18560 -297080
rect 20760 -297180 20780 -297080
rect 18540 -297200 20780 -297180
rect 21540 -297080 23780 -297060
rect 21540 -297180 21560 -297080
rect 23760 -297180 23780 -297080
rect 21540 -297200 23780 -297180
rect 24540 -297080 26780 -297060
rect 24540 -297180 24560 -297080
rect 26760 -297180 26780 -297080
rect 24540 -297200 26780 -297180
rect 27540 -297080 29780 -297060
rect 27540 -297180 27560 -297080
rect 29760 -297180 29780 -297080
rect 27540 -297200 29780 -297180
rect 30540 -297080 32780 -297060
rect 30540 -297180 30560 -297080
rect 32760 -297180 32780 -297080
rect 30540 -297200 32780 -297180
rect 33540 -297080 35780 -297060
rect 33540 -297180 33560 -297080
rect 35760 -297180 35780 -297080
rect 33540 -297200 35780 -297180
rect 36540 -297080 38780 -297060
rect 36540 -297180 36560 -297080
rect 38760 -297180 38780 -297080
rect 36540 -297200 38780 -297180
rect 39540 -297080 41780 -297060
rect 39540 -297180 39560 -297080
rect 41760 -297180 41780 -297080
rect 39540 -297200 41780 -297180
rect 42540 -297080 44780 -297060
rect 42540 -297180 42560 -297080
rect 44760 -297180 44780 -297080
rect 42540 -297200 44780 -297180
rect 45540 -297080 47780 -297060
rect 45540 -297180 45560 -297080
rect 47760 -297180 47780 -297080
rect 45540 -297200 47780 -297180
rect 48540 -297080 50780 -297060
rect 48540 -297180 48560 -297080
rect 50760 -297180 50780 -297080
rect 48540 -297200 50780 -297180
rect 51540 -297080 53780 -297060
rect 51540 -297180 51560 -297080
rect 53760 -297180 53780 -297080
rect 51540 -297200 53780 -297180
rect 54540 -297080 56780 -297060
rect 54540 -297180 54560 -297080
rect 56760 -297180 56780 -297080
rect 54540 -297200 56780 -297180
rect 57540 -297080 59780 -297060
rect 57540 -297180 57560 -297080
rect 59760 -297180 59780 -297080
rect 57540 -297200 59780 -297180
rect 60540 -297080 62780 -297060
rect 60540 -297180 60560 -297080
rect 62760 -297180 62780 -297080
rect 60540 -297200 62780 -297180
rect 63540 -297080 65780 -297060
rect 63540 -297180 63560 -297080
rect 65760 -297180 65780 -297080
rect 63540 -297200 65780 -297180
rect 66540 -297080 68780 -297060
rect 66540 -297180 66560 -297080
rect 68760 -297180 68780 -297080
rect 66540 -297200 68780 -297180
rect 69540 -297080 71780 -297060
rect 69540 -297180 69560 -297080
rect 71760 -297180 71780 -297080
rect 69540 -297200 71780 -297180
rect 72540 -297080 74780 -297060
rect 72540 -297180 72560 -297080
rect 74760 -297180 74780 -297080
rect 72540 -297200 74780 -297180
rect 75540 -297080 77780 -297060
rect 75540 -297180 75560 -297080
rect 77760 -297180 77780 -297080
rect 75540 -297200 77780 -297180
rect 78540 -297080 80780 -297060
rect 78540 -297180 78560 -297080
rect 80760 -297180 80780 -297080
rect 78540 -297200 80780 -297180
rect 81540 -297080 83780 -297060
rect 81540 -297180 81560 -297080
rect 83760 -297180 83780 -297080
rect 81540 -297200 83780 -297180
rect 84540 -297080 86780 -297060
rect 84540 -297180 84560 -297080
rect 86760 -297180 86780 -297080
rect 84540 -297200 86780 -297180
rect 87540 -297080 89780 -297060
rect 87540 -297180 87560 -297080
rect 89760 -297180 89780 -297080
rect 87540 -297200 89780 -297180
rect 90540 -297080 92780 -297060
rect 90540 -297180 90560 -297080
rect 92760 -297180 92780 -297080
rect 90540 -297200 92780 -297180
rect 93540 -297080 95780 -297060
rect 93540 -297180 93560 -297080
rect 95760 -297180 95780 -297080
rect 93540 -297200 95780 -297180
rect 96540 -297080 98780 -297060
rect 96540 -297180 96560 -297080
rect 98760 -297180 98780 -297080
rect 96540 -297200 98780 -297180
rect 99540 -297080 101780 -297060
rect 99540 -297180 99560 -297080
rect 101760 -297180 101780 -297080
rect 99540 -297200 101780 -297180
rect 102540 -297080 104780 -297060
rect 102540 -297180 102560 -297080
rect 104760 -297180 104780 -297080
rect 102540 -297200 104780 -297180
rect 105540 -297080 107780 -297060
rect 105540 -297180 105560 -297080
rect 107760 -297180 107780 -297080
rect 105540 -297200 107780 -297180
rect 108540 -297080 110780 -297060
rect 108540 -297180 108560 -297080
rect 110760 -297180 110780 -297080
rect 108540 -297200 110780 -297180
rect 111540 -297080 113780 -297060
rect 111540 -297180 111560 -297080
rect 113760 -297180 113780 -297080
rect 111540 -297200 113780 -297180
rect 114540 -297080 116780 -297060
rect 114540 -297180 114560 -297080
rect 116760 -297180 116780 -297080
rect 114540 -297200 116780 -297180
rect 117540 -297080 119780 -297060
rect 117540 -297180 117560 -297080
rect 119760 -297180 119780 -297080
rect 117540 -297200 119780 -297180
rect 120540 -297080 122780 -297060
rect 120540 -297180 120560 -297080
rect 122760 -297180 122780 -297080
rect 120540 -297200 122780 -297180
rect 123540 -297080 125780 -297060
rect 123540 -297180 123560 -297080
rect 125760 -297180 125780 -297080
rect 123540 -297200 125780 -297180
rect 126540 -297080 128780 -297060
rect 126540 -297180 126560 -297080
rect 128760 -297180 128780 -297080
rect 126540 -297200 128780 -297180
rect 129540 -297080 131780 -297060
rect 129540 -297180 129560 -297080
rect 131760 -297180 131780 -297080
rect 129540 -297200 131780 -297180
rect 132540 -297080 134780 -297060
rect 132540 -297180 132560 -297080
rect 134760 -297180 134780 -297080
rect 132540 -297200 134780 -297180
rect 135540 -297080 137780 -297060
rect 135540 -297180 135560 -297080
rect 137760 -297180 137780 -297080
rect 135540 -297200 137780 -297180
rect 138540 -297080 140780 -297060
rect 138540 -297180 138560 -297080
rect 140760 -297180 140780 -297080
rect 138540 -297200 140780 -297180
rect 141540 -297080 143780 -297060
rect 141540 -297180 141560 -297080
rect 143760 -297180 143780 -297080
rect 141540 -297200 143780 -297180
rect 144540 -297080 146780 -297060
rect 144540 -297180 144560 -297080
rect 146760 -297180 146780 -297080
rect 144540 -297200 146780 -297180
rect 147540 -297080 149780 -297060
rect 147540 -297180 147560 -297080
rect 149760 -297180 149780 -297080
rect 147540 -297200 149780 -297180
rect 150540 -297080 152780 -297060
rect 150540 -297180 150560 -297080
rect 152760 -297180 152780 -297080
rect 150540 -297200 152780 -297180
rect 153540 -297080 155780 -297060
rect 153540 -297180 153560 -297080
rect 155760 -297180 155780 -297080
rect 153540 -297200 155780 -297180
rect 156540 -297080 158780 -297060
rect 156540 -297180 156560 -297080
rect 158760 -297180 158780 -297080
rect 156540 -297200 158780 -297180
rect 159540 -297080 161780 -297060
rect 159540 -297180 159560 -297080
rect 161760 -297180 161780 -297080
rect 159540 -297200 161780 -297180
rect 162540 -297080 164780 -297060
rect 162540 -297180 162560 -297080
rect 164760 -297180 164780 -297080
rect 162540 -297200 164780 -297180
rect 165540 -297080 167780 -297060
rect 165540 -297180 165560 -297080
rect 167760 -297180 167780 -297080
rect 165540 -297200 167780 -297180
rect 168540 -297080 170780 -297060
rect 168540 -297180 168560 -297080
rect 170760 -297180 170780 -297080
rect 168540 -297200 170780 -297180
rect 171540 -297080 173780 -297060
rect 171540 -297180 171560 -297080
rect 173760 -297180 173780 -297080
rect 171540 -297200 173780 -297180
rect 174540 -297080 176780 -297060
rect 174540 -297180 174560 -297080
rect 176760 -297180 176780 -297080
rect 174540 -297200 176780 -297180
rect 177540 -297080 179780 -297060
rect 177540 -297180 177560 -297080
rect 179760 -297180 179780 -297080
rect 177540 -297200 179780 -297180
rect 180540 -297080 182780 -297060
rect 180540 -297180 180560 -297080
rect 182760 -297180 182780 -297080
rect 180540 -297200 182780 -297180
rect 183540 -297080 185780 -297060
rect 183540 -297180 183560 -297080
rect 185760 -297180 185780 -297080
rect 183540 -297200 185780 -297180
rect 186540 -297080 188780 -297060
rect 186540 -297180 186560 -297080
rect 188760 -297180 188780 -297080
rect 186540 -297200 188780 -297180
rect 189540 -297080 191780 -297060
rect 189540 -297180 189560 -297080
rect 191760 -297180 191780 -297080
rect 189540 -297200 191780 -297180
rect 192540 -297080 194780 -297060
rect 192540 -297180 192560 -297080
rect 194760 -297180 194780 -297080
rect 192540 -297200 194780 -297180
rect 195540 -297080 197780 -297060
rect 195540 -297180 195560 -297080
rect 197760 -297180 197780 -297080
rect 195540 -297200 197780 -297180
rect 198540 -297080 200780 -297060
rect 198540 -297180 198560 -297080
rect 200760 -297180 200780 -297080
rect 198540 -297200 200780 -297180
rect 201540 -297080 203780 -297060
rect 201540 -297180 201560 -297080
rect 203760 -297180 203780 -297080
rect 201540 -297200 203780 -297180
rect 204540 -297080 206780 -297060
rect 204540 -297180 204560 -297080
rect 206760 -297180 206780 -297080
rect 204540 -297200 206780 -297180
rect 207540 -297080 209780 -297060
rect 207540 -297180 207560 -297080
rect 209760 -297180 209780 -297080
rect 207540 -297200 209780 -297180
rect 210540 -297080 212780 -297060
rect 210540 -297180 210560 -297080
rect 212760 -297180 212780 -297080
rect 210540 -297200 212780 -297180
rect 213540 -297080 215780 -297060
rect 213540 -297180 213560 -297080
rect 215760 -297180 215780 -297080
rect 213540 -297200 215780 -297180
rect 216540 -297080 218780 -297060
rect 216540 -297180 216560 -297080
rect 218760 -297180 218780 -297080
rect 216540 -297200 218780 -297180
rect 219540 -297080 221780 -297060
rect 219540 -297180 219560 -297080
rect 221760 -297180 221780 -297080
rect 219540 -297200 221780 -297180
rect 222540 -297080 224780 -297060
rect 222540 -297180 222560 -297080
rect 224760 -297180 224780 -297080
rect 222540 -297200 224780 -297180
rect 225540 -297080 227780 -297060
rect 225540 -297180 225560 -297080
rect 227760 -297180 227780 -297080
rect 225540 -297200 227780 -297180
rect 228540 -297080 230780 -297060
rect 228540 -297180 228560 -297080
rect 230760 -297180 230780 -297080
rect 228540 -297200 230780 -297180
rect 231540 -297080 233780 -297060
rect 231540 -297180 231560 -297080
rect 233760 -297180 233780 -297080
rect 231540 -297200 233780 -297180
rect 234540 -297080 236780 -297060
rect 234540 -297180 234560 -297080
rect 236760 -297180 236780 -297080
rect 234540 -297200 236780 -297180
rect 237540 -297080 239780 -297060
rect 237540 -297180 237560 -297080
rect 239760 -297180 239780 -297080
rect 237540 -297200 239780 -297180
rect 240540 -297080 242780 -297060
rect 240540 -297180 240560 -297080
rect 242760 -297180 242780 -297080
rect 240540 -297200 242780 -297180
rect 243540 -297080 245780 -297060
rect 243540 -297180 243560 -297080
rect 245760 -297180 245780 -297080
rect 243540 -297200 245780 -297180
rect 246540 -297080 248780 -297060
rect 246540 -297180 246560 -297080
rect 248760 -297180 248780 -297080
rect 246540 -297200 248780 -297180
rect 249540 -297080 251780 -297060
rect 249540 -297180 249560 -297080
rect 251760 -297180 251780 -297080
rect 249540 -297200 251780 -297180
rect 252540 -297080 254780 -297060
rect 252540 -297180 252560 -297080
rect 254760 -297180 254780 -297080
rect 252540 -297200 254780 -297180
rect 255540 -297080 257780 -297060
rect 255540 -297180 255560 -297080
rect 257760 -297180 257780 -297080
rect 255540 -297200 257780 -297180
rect 258540 -297080 260780 -297060
rect 258540 -297180 258560 -297080
rect 260760 -297180 260780 -297080
rect 258540 -297200 260780 -297180
rect 261540 -297080 263780 -297060
rect 261540 -297180 261560 -297080
rect 263760 -297180 263780 -297080
rect 261540 -297200 263780 -297180
rect 264540 -297080 266780 -297060
rect 264540 -297180 264560 -297080
rect 266760 -297180 266780 -297080
rect 264540 -297200 266780 -297180
rect 267540 -297080 269780 -297060
rect 267540 -297180 267560 -297080
rect 269760 -297180 269780 -297080
rect 267540 -297200 269780 -297180
rect 270540 -297080 272780 -297060
rect 270540 -297180 270560 -297080
rect 272760 -297180 272780 -297080
rect 270540 -297200 272780 -297180
rect 273540 -297080 275780 -297060
rect 273540 -297180 273560 -297080
rect 275760 -297180 275780 -297080
rect 273540 -297200 275780 -297180
rect 276540 -297080 278780 -297060
rect 276540 -297180 276560 -297080
rect 278760 -297180 278780 -297080
rect 276540 -297200 278780 -297180
rect 279540 -297080 281780 -297060
rect 279540 -297180 279560 -297080
rect 281760 -297180 281780 -297080
rect 279540 -297200 281780 -297180
rect 282540 -297080 284780 -297060
rect 282540 -297180 282560 -297080
rect 284760 -297180 284780 -297080
rect 282540 -297200 284780 -297180
rect 285540 -297080 287780 -297060
rect 285540 -297180 285560 -297080
rect 287760 -297180 287780 -297080
rect 285540 -297200 287780 -297180
rect 288540 -297080 290780 -297060
rect 288540 -297180 288560 -297080
rect 290760 -297180 290780 -297080
rect 288540 -297200 290780 -297180
rect 291540 -297080 293780 -297060
rect 291540 -297180 291560 -297080
rect 293760 -297180 293780 -297080
rect 291540 -297200 293780 -297180
rect 294540 -297080 296780 -297060
rect 294540 -297180 294560 -297080
rect 296760 -297180 296780 -297080
rect 294540 -297200 296780 -297180
rect 297540 -297080 299780 -297060
rect 297540 -297180 297560 -297080
rect 299760 -297180 299780 -297080
rect 297540 -297200 299780 -297180
rect 220 -297500 440 -297490
rect 220 -297700 240 -297500
rect 420 -297700 440 -297500
rect 220 -298100 440 -297700
rect 3220 -297500 3440 -297490
rect 3220 -297700 3240 -297500
rect 3420 -297700 3440 -297500
rect 3220 -298100 3440 -297700
rect 6220 -297500 6440 -297490
rect 6220 -297700 6240 -297500
rect 6420 -297700 6440 -297500
rect 6220 -298100 6440 -297700
rect 9220 -297500 9440 -297490
rect 9220 -297700 9240 -297500
rect 9420 -297700 9440 -297500
rect 9220 -298100 9440 -297700
rect 12220 -297500 12440 -297490
rect 12220 -297700 12240 -297500
rect 12420 -297700 12440 -297500
rect 12220 -298100 12440 -297700
rect 15220 -297500 15440 -297490
rect 15220 -297700 15240 -297500
rect 15420 -297700 15440 -297500
rect 15220 -298100 15440 -297700
rect 18220 -297500 18440 -297490
rect 18220 -297700 18240 -297500
rect 18420 -297700 18440 -297500
rect 18220 -298100 18440 -297700
rect 21220 -297500 21440 -297490
rect 21220 -297700 21240 -297500
rect 21420 -297700 21440 -297500
rect 21220 -298100 21440 -297700
rect 24220 -297500 24440 -297490
rect 24220 -297700 24240 -297500
rect 24420 -297700 24440 -297500
rect 24220 -298100 24440 -297700
rect 27220 -297500 27440 -297490
rect 27220 -297700 27240 -297500
rect 27420 -297700 27440 -297500
rect 27220 -298100 27440 -297700
rect 30220 -297500 30440 -297490
rect 30220 -297700 30240 -297500
rect 30420 -297700 30440 -297500
rect 30220 -298100 30440 -297700
rect 33220 -297500 33440 -297490
rect 33220 -297700 33240 -297500
rect 33420 -297700 33440 -297500
rect 33220 -298100 33440 -297700
rect 36220 -297500 36440 -297490
rect 36220 -297700 36240 -297500
rect 36420 -297700 36440 -297500
rect 36220 -298100 36440 -297700
rect 39220 -297500 39440 -297490
rect 39220 -297700 39240 -297500
rect 39420 -297700 39440 -297500
rect 39220 -298100 39440 -297700
rect 42220 -297500 42440 -297490
rect 42220 -297700 42240 -297500
rect 42420 -297700 42440 -297500
rect 42220 -298100 42440 -297700
rect 45220 -297500 45440 -297490
rect 45220 -297700 45240 -297500
rect 45420 -297700 45440 -297500
rect 45220 -298100 45440 -297700
rect 48220 -297500 48440 -297490
rect 48220 -297700 48240 -297500
rect 48420 -297700 48440 -297500
rect 48220 -298100 48440 -297700
rect 51220 -297500 51440 -297490
rect 51220 -297700 51240 -297500
rect 51420 -297700 51440 -297500
rect 51220 -298100 51440 -297700
rect 54220 -297500 54440 -297490
rect 54220 -297700 54240 -297500
rect 54420 -297700 54440 -297500
rect 54220 -298100 54440 -297700
rect 57220 -297500 57440 -297490
rect 57220 -297700 57240 -297500
rect 57420 -297700 57440 -297500
rect 57220 -298100 57440 -297700
rect 60220 -297500 60440 -297490
rect 60220 -297700 60240 -297500
rect 60420 -297700 60440 -297500
rect 60220 -298100 60440 -297700
rect 63220 -297500 63440 -297490
rect 63220 -297700 63240 -297500
rect 63420 -297700 63440 -297500
rect 63220 -298100 63440 -297700
rect 66220 -297500 66440 -297490
rect 66220 -297700 66240 -297500
rect 66420 -297700 66440 -297500
rect 66220 -298100 66440 -297700
rect 69220 -297500 69440 -297490
rect 69220 -297700 69240 -297500
rect 69420 -297700 69440 -297500
rect 69220 -298100 69440 -297700
rect 72220 -297500 72440 -297490
rect 72220 -297700 72240 -297500
rect 72420 -297700 72440 -297500
rect 72220 -298100 72440 -297700
rect 75220 -297500 75440 -297490
rect 75220 -297700 75240 -297500
rect 75420 -297700 75440 -297500
rect 75220 -298100 75440 -297700
rect 78220 -297500 78440 -297490
rect 78220 -297700 78240 -297500
rect 78420 -297700 78440 -297500
rect 78220 -298100 78440 -297700
rect 81220 -297500 81440 -297490
rect 81220 -297700 81240 -297500
rect 81420 -297700 81440 -297500
rect 81220 -298100 81440 -297700
rect 84220 -297500 84440 -297490
rect 84220 -297700 84240 -297500
rect 84420 -297700 84440 -297500
rect 84220 -298100 84440 -297700
rect 87220 -297500 87440 -297490
rect 87220 -297700 87240 -297500
rect 87420 -297700 87440 -297500
rect 87220 -298100 87440 -297700
rect 90220 -297500 90440 -297490
rect 90220 -297700 90240 -297500
rect 90420 -297700 90440 -297500
rect 90220 -298100 90440 -297700
rect 93220 -297500 93440 -297490
rect 93220 -297700 93240 -297500
rect 93420 -297700 93440 -297500
rect 93220 -298100 93440 -297700
rect 96220 -297500 96440 -297490
rect 96220 -297700 96240 -297500
rect 96420 -297700 96440 -297500
rect 96220 -298100 96440 -297700
rect 99220 -297500 99440 -297490
rect 99220 -297700 99240 -297500
rect 99420 -297700 99440 -297500
rect 99220 -298100 99440 -297700
rect 102220 -297500 102440 -297490
rect 102220 -297700 102240 -297500
rect 102420 -297700 102440 -297500
rect 102220 -298100 102440 -297700
rect 105220 -297500 105440 -297490
rect 105220 -297700 105240 -297500
rect 105420 -297700 105440 -297500
rect 105220 -298100 105440 -297700
rect 108220 -297500 108440 -297490
rect 108220 -297700 108240 -297500
rect 108420 -297700 108440 -297500
rect 108220 -298100 108440 -297700
rect 111220 -297500 111440 -297490
rect 111220 -297700 111240 -297500
rect 111420 -297700 111440 -297500
rect 111220 -298100 111440 -297700
rect 114220 -297500 114440 -297490
rect 114220 -297700 114240 -297500
rect 114420 -297700 114440 -297500
rect 114220 -298100 114440 -297700
rect 117220 -297500 117440 -297490
rect 117220 -297700 117240 -297500
rect 117420 -297700 117440 -297500
rect 117220 -298100 117440 -297700
rect 120220 -297500 120440 -297490
rect 120220 -297700 120240 -297500
rect 120420 -297700 120440 -297500
rect 120220 -298100 120440 -297700
rect 123220 -297500 123440 -297490
rect 123220 -297700 123240 -297500
rect 123420 -297700 123440 -297500
rect 123220 -298100 123440 -297700
rect 126220 -297500 126440 -297490
rect 126220 -297700 126240 -297500
rect 126420 -297700 126440 -297500
rect 126220 -298100 126440 -297700
rect 129220 -297500 129440 -297490
rect 129220 -297700 129240 -297500
rect 129420 -297700 129440 -297500
rect 129220 -298100 129440 -297700
rect 132220 -297500 132440 -297490
rect 132220 -297700 132240 -297500
rect 132420 -297700 132440 -297500
rect 132220 -298100 132440 -297700
rect 135220 -297500 135440 -297490
rect 135220 -297700 135240 -297500
rect 135420 -297700 135440 -297500
rect 135220 -298100 135440 -297700
rect 138220 -297500 138440 -297490
rect 138220 -297700 138240 -297500
rect 138420 -297700 138440 -297500
rect 138220 -298100 138440 -297700
rect 141220 -297500 141440 -297490
rect 141220 -297700 141240 -297500
rect 141420 -297700 141440 -297500
rect 141220 -298100 141440 -297700
rect 144220 -297500 144440 -297490
rect 144220 -297700 144240 -297500
rect 144420 -297700 144440 -297500
rect 144220 -298100 144440 -297700
rect 147220 -297500 147440 -297490
rect 147220 -297700 147240 -297500
rect 147420 -297700 147440 -297500
rect 147220 -298100 147440 -297700
rect 150220 -297500 150440 -297490
rect 150220 -297700 150240 -297500
rect 150420 -297700 150440 -297500
rect 150220 -298100 150440 -297700
rect 153220 -297500 153440 -297490
rect 153220 -297700 153240 -297500
rect 153420 -297700 153440 -297500
rect 153220 -298100 153440 -297700
rect 156220 -297500 156440 -297490
rect 156220 -297700 156240 -297500
rect 156420 -297700 156440 -297500
rect 156220 -298100 156440 -297700
rect 159220 -297500 159440 -297490
rect 159220 -297700 159240 -297500
rect 159420 -297700 159440 -297500
rect 159220 -298100 159440 -297700
rect 162220 -297500 162440 -297490
rect 162220 -297700 162240 -297500
rect 162420 -297700 162440 -297500
rect 162220 -298100 162440 -297700
rect 165220 -297500 165440 -297490
rect 165220 -297700 165240 -297500
rect 165420 -297700 165440 -297500
rect 165220 -298100 165440 -297700
rect 168220 -297500 168440 -297490
rect 168220 -297700 168240 -297500
rect 168420 -297700 168440 -297500
rect 168220 -298100 168440 -297700
rect 171220 -297500 171440 -297490
rect 171220 -297700 171240 -297500
rect 171420 -297700 171440 -297500
rect 171220 -298100 171440 -297700
rect 174220 -297500 174440 -297490
rect 174220 -297700 174240 -297500
rect 174420 -297700 174440 -297500
rect 174220 -298100 174440 -297700
rect 177220 -297500 177440 -297490
rect 177220 -297700 177240 -297500
rect 177420 -297700 177440 -297500
rect 177220 -298100 177440 -297700
rect 180220 -297500 180440 -297490
rect 180220 -297700 180240 -297500
rect 180420 -297700 180440 -297500
rect 180220 -298100 180440 -297700
rect 183220 -297500 183440 -297490
rect 183220 -297700 183240 -297500
rect 183420 -297700 183440 -297500
rect 183220 -298100 183440 -297700
rect 186220 -297500 186440 -297490
rect 186220 -297700 186240 -297500
rect 186420 -297700 186440 -297500
rect 186220 -298100 186440 -297700
rect 189220 -297500 189440 -297490
rect 189220 -297700 189240 -297500
rect 189420 -297700 189440 -297500
rect 189220 -298100 189440 -297700
rect 192220 -297500 192440 -297490
rect 192220 -297700 192240 -297500
rect 192420 -297700 192440 -297500
rect 192220 -298100 192440 -297700
rect 195220 -297500 195440 -297490
rect 195220 -297700 195240 -297500
rect 195420 -297700 195440 -297500
rect 195220 -298100 195440 -297700
rect 198220 -297500 198440 -297490
rect 198220 -297700 198240 -297500
rect 198420 -297700 198440 -297500
rect 198220 -298100 198440 -297700
rect 201220 -297500 201440 -297490
rect 201220 -297700 201240 -297500
rect 201420 -297700 201440 -297500
rect 201220 -298100 201440 -297700
rect 204220 -297500 204440 -297490
rect 204220 -297700 204240 -297500
rect 204420 -297700 204440 -297500
rect 204220 -298100 204440 -297700
rect 207220 -297500 207440 -297490
rect 207220 -297700 207240 -297500
rect 207420 -297700 207440 -297500
rect 207220 -298100 207440 -297700
rect 210220 -297500 210440 -297490
rect 210220 -297700 210240 -297500
rect 210420 -297700 210440 -297500
rect 210220 -298100 210440 -297700
rect 213220 -297500 213440 -297490
rect 213220 -297700 213240 -297500
rect 213420 -297700 213440 -297500
rect 213220 -298100 213440 -297700
rect 216220 -297500 216440 -297490
rect 216220 -297700 216240 -297500
rect 216420 -297700 216440 -297500
rect 216220 -298100 216440 -297700
rect 219220 -297500 219440 -297490
rect 219220 -297700 219240 -297500
rect 219420 -297700 219440 -297500
rect 219220 -298100 219440 -297700
rect 222220 -297500 222440 -297490
rect 222220 -297700 222240 -297500
rect 222420 -297700 222440 -297500
rect 222220 -298100 222440 -297700
rect 225220 -297500 225440 -297490
rect 225220 -297700 225240 -297500
rect 225420 -297700 225440 -297500
rect 225220 -298100 225440 -297700
rect 228220 -297500 228440 -297490
rect 228220 -297700 228240 -297500
rect 228420 -297700 228440 -297500
rect 228220 -298100 228440 -297700
rect 231220 -297500 231440 -297490
rect 231220 -297700 231240 -297500
rect 231420 -297700 231440 -297500
rect 231220 -298100 231440 -297700
rect 234220 -297500 234440 -297490
rect 234220 -297700 234240 -297500
rect 234420 -297700 234440 -297500
rect 234220 -298100 234440 -297700
rect 237220 -297500 237440 -297490
rect 237220 -297700 237240 -297500
rect 237420 -297700 237440 -297500
rect 237220 -298100 237440 -297700
rect 240220 -297500 240440 -297490
rect 240220 -297700 240240 -297500
rect 240420 -297700 240440 -297500
rect 240220 -298100 240440 -297700
rect 243220 -297500 243440 -297490
rect 243220 -297700 243240 -297500
rect 243420 -297700 243440 -297500
rect 243220 -298100 243440 -297700
rect 246220 -297500 246440 -297490
rect 246220 -297700 246240 -297500
rect 246420 -297700 246440 -297500
rect 246220 -298100 246440 -297700
rect 249220 -297500 249440 -297490
rect 249220 -297700 249240 -297500
rect 249420 -297700 249440 -297500
rect 249220 -298100 249440 -297700
rect 252220 -297500 252440 -297490
rect 252220 -297700 252240 -297500
rect 252420 -297700 252440 -297500
rect 252220 -298100 252440 -297700
rect 255220 -297500 255440 -297490
rect 255220 -297700 255240 -297500
rect 255420 -297700 255440 -297500
rect 255220 -298100 255440 -297700
rect 258220 -297500 258440 -297490
rect 258220 -297700 258240 -297500
rect 258420 -297700 258440 -297500
rect 258220 -298100 258440 -297700
rect 261220 -297500 261440 -297490
rect 261220 -297700 261240 -297500
rect 261420 -297700 261440 -297500
rect 261220 -298100 261440 -297700
rect 264220 -297500 264440 -297490
rect 264220 -297700 264240 -297500
rect 264420 -297700 264440 -297500
rect 264220 -298100 264440 -297700
rect 267220 -297500 267440 -297490
rect 267220 -297700 267240 -297500
rect 267420 -297700 267440 -297500
rect 267220 -298100 267440 -297700
rect 270220 -297500 270440 -297490
rect 270220 -297700 270240 -297500
rect 270420 -297700 270440 -297500
rect 270220 -298100 270440 -297700
rect 273220 -297500 273440 -297490
rect 273220 -297700 273240 -297500
rect 273420 -297700 273440 -297500
rect 273220 -298100 273440 -297700
rect 276220 -297500 276440 -297490
rect 276220 -297700 276240 -297500
rect 276420 -297700 276440 -297500
rect 276220 -298100 276440 -297700
rect 279220 -297500 279440 -297490
rect 279220 -297700 279240 -297500
rect 279420 -297700 279440 -297500
rect 279220 -298100 279440 -297700
rect 282220 -297500 282440 -297490
rect 282220 -297700 282240 -297500
rect 282420 -297700 282440 -297500
rect 282220 -298100 282440 -297700
rect 285220 -297500 285440 -297490
rect 285220 -297700 285240 -297500
rect 285420 -297700 285440 -297500
rect 285220 -298100 285440 -297700
rect 288220 -297500 288440 -297490
rect 288220 -297700 288240 -297500
rect 288420 -297700 288440 -297500
rect 288220 -298100 288440 -297700
rect 291220 -297500 291440 -297490
rect 291220 -297700 291240 -297500
rect 291420 -297700 291440 -297500
rect 291220 -298100 291440 -297700
rect 294220 -297500 294440 -297490
rect 294220 -297700 294240 -297500
rect 294420 -297700 294440 -297500
rect 294220 -298100 294440 -297700
rect 297220 -297500 297440 -297490
rect 297220 -297700 297240 -297500
rect 297420 -297700 297440 -297500
rect 297220 -298100 297440 -297700
<< metal5 >>
rect -2000 2840 0 3160
use pixel  pixel_9801
timestamp 1654712443
transform 1 0 -800 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9800
timestamp 1654712443
transform 1 0 -3800 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9901
timestamp 1654712443
transform 1 0 -800 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9900
timestamp 1654712443
transform 1 0 -3800 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9802
timestamp 1654712443
transform 1 0 2200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9902
timestamp 1654712443
transform 1 0 2200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9803
timestamp 1654712443
transform 1 0 5200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9903
timestamp 1654712443
transform 1 0 5200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9804
timestamp 1654712443
transform 1 0 8200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9904
timestamp 1654712443
transform 1 0 8200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9805
timestamp 1654712443
transform 1 0 11200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9905
timestamp 1654712443
transform 1 0 11200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9806
timestamp 1654712443
transform 1 0 14200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9906
timestamp 1654712443
transform 1 0 14200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9807
timestamp 1654712443
transform 1 0 17200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9907
timestamp 1654712443
transform 1 0 17200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9808
timestamp 1654712443
transform 1 0 20200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9908
timestamp 1654712443
transform 1 0 20200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9809
timestamp 1654712443
transform 1 0 23200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9909
timestamp 1654712443
transform 1 0 23200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9811
timestamp 1654712443
transform 1 0 29200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9810
timestamp 1654712443
transform 1 0 26200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9911
timestamp 1654712443
transform 1 0 29200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9910
timestamp 1654712443
transform 1 0 26200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9812
timestamp 1654712443
transform 1 0 32200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9912
timestamp 1654712443
transform 1 0 32200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9813
timestamp 1654712443
transform 1 0 35200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9913
timestamp 1654712443
transform 1 0 35200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9814
timestamp 1654712443
transform 1 0 38200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9914
timestamp 1654712443
transform 1 0 38200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9815
timestamp 1654712443
transform 1 0 41200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9915
timestamp 1654712443
transform 1 0 41200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9816
timestamp 1654712443
transform 1 0 44200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9916
timestamp 1654712443
transform 1 0 44200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9817
timestamp 1654712443
transform 1 0 47200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9917
timestamp 1654712443
transform 1 0 47200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9818
timestamp 1654712443
transform 1 0 50200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9918
timestamp 1654712443
transform 1 0 50200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9819
timestamp 1654712443
transform 1 0 53200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9919
timestamp 1654712443
transform 1 0 53200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9821
timestamp 1654712443
transform 1 0 59200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9820
timestamp 1654712443
transform 1 0 56200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9921
timestamp 1654712443
transform 1 0 59200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9920
timestamp 1654712443
transform 1 0 56200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9822
timestamp 1654712443
transform 1 0 62200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9922
timestamp 1654712443
transform 1 0 62200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9823
timestamp 1654712443
transform 1 0 65200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9923
timestamp 1654712443
transform 1 0 65200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9824
timestamp 1654712443
transform 1 0 68200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9924
timestamp 1654712443
transform 1 0 68200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9825
timestamp 1654712443
transform 1 0 71200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9925
timestamp 1654712443
transform 1 0 71200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9826
timestamp 1654712443
transform 1 0 74200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9926
timestamp 1654712443
transform 1 0 74200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9827
timestamp 1654712443
transform 1 0 77200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9927
timestamp 1654712443
transform 1 0 77200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9828
timestamp 1654712443
transform 1 0 80200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9928
timestamp 1654712443
transform 1 0 80200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9829
timestamp 1654712443
transform 1 0 83200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9929
timestamp 1654712443
transform 1 0 83200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9830
timestamp 1654712443
transform 1 0 86200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9930
timestamp 1654712443
transform 1 0 86200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9831
timestamp 1654712443
transform 1 0 89200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9832
timestamp 1654712443
transform 1 0 92200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9931
timestamp 1654712443
transform 1 0 89200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9932
timestamp 1654712443
transform 1 0 92200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9833
timestamp 1654712443
transform 1 0 95200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9933
timestamp 1654712443
transform 1 0 95200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9834
timestamp 1654712443
transform 1 0 98200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9934
timestamp 1654712443
transform 1 0 98200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9835
timestamp 1654712443
transform 1 0 101200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9935
timestamp 1654712443
transform 1 0 101200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9836
timestamp 1654712443
transform 1 0 104200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9936
timestamp 1654712443
transform 1 0 104200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9837
timestamp 1654712443
transform 1 0 107200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9937
timestamp 1654712443
transform 1 0 107200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9838
timestamp 1654712443
transform 1 0 110200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9938
timestamp 1654712443
transform 1 0 110200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9839
timestamp 1654712443
transform 1 0 113200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9939
timestamp 1654712443
transform 1 0 113200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9840
timestamp 1654712443
transform 1 0 116200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9940
timestamp 1654712443
transform 1 0 116200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9841
timestamp 1654712443
transform 1 0 119200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9842
timestamp 1654712443
transform 1 0 122200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9941
timestamp 1654712443
transform 1 0 119200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9942
timestamp 1654712443
transform 1 0 122200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9843
timestamp 1654712443
transform 1 0 125200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9943
timestamp 1654712443
transform 1 0 125200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9844
timestamp 1654712443
transform 1 0 128200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9944
timestamp 1654712443
transform 1 0 128200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9845
timestamp 1654712443
transform 1 0 131200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9945
timestamp 1654712443
transform 1 0 131200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9846
timestamp 1654712443
transform 1 0 134200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9946
timestamp 1654712443
transform 1 0 134200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9847
timestamp 1654712443
transform 1 0 137200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9947
timestamp 1654712443
transform 1 0 137200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9848
timestamp 1654712443
transform 1 0 140200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9948
timestamp 1654712443
transform 1 0 140200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9849
timestamp 1654712443
transform 1 0 143200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9949
timestamp 1654712443
transform 1 0 143200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9850
timestamp 1654712443
transform 1 0 146200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9950
timestamp 1654712443
transform 1 0 146200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9851
timestamp 1654712443
transform 1 0 149200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9852
timestamp 1654712443
transform 1 0 152200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9951
timestamp 1654712443
transform 1 0 149200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9952
timestamp 1654712443
transform 1 0 152200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9853
timestamp 1654712443
transform 1 0 155200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9953
timestamp 1654712443
transform 1 0 155200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9854
timestamp 1654712443
transform 1 0 158200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9954
timestamp 1654712443
transform 1 0 158200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9855
timestamp 1654712443
transform 1 0 161200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9955
timestamp 1654712443
transform 1 0 161200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9856
timestamp 1654712443
transform 1 0 164200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9956
timestamp 1654712443
transform 1 0 164200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9857
timestamp 1654712443
transform 1 0 167200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9957
timestamp 1654712443
transform 1 0 167200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9858
timestamp 1654712443
transform 1 0 170200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9958
timestamp 1654712443
transform 1 0 170200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9859
timestamp 1654712443
transform 1 0 173200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9959
timestamp 1654712443
transform 1 0 173200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9860
timestamp 1654712443
transform 1 0 176200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9960
timestamp 1654712443
transform 1 0 176200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9861
timestamp 1654712443
transform 1 0 179200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9961
timestamp 1654712443
transform 1 0 179200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9863
timestamp 1654712443
transform 1 0 185200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9862
timestamp 1654712443
transform 1 0 182200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9963
timestamp 1654712443
transform 1 0 185200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9962
timestamp 1654712443
transform 1 0 182200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9864
timestamp 1654712443
transform 1 0 188200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9964
timestamp 1654712443
transform 1 0 188200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9865
timestamp 1654712443
transform 1 0 191200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9965
timestamp 1654712443
transform 1 0 191200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9866
timestamp 1654712443
transform 1 0 194200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9966
timestamp 1654712443
transform 1 0 194200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9867
timestamp 1654712443
transform 1 0 197200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9967
timestamp 1654712443
transform 1 0 197200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9868
timestamp 1654712443
transform 1 0 200200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9968
timestamp 1654712443
transform 1 0 200200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9869
timestamp 1654712443
transform 1 0 203200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9969
timestamp 1654712443
transform 1 0 203200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9870
timestamp 1654712443
transform 1 0 206200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9970
timestamp 1654712443
transform 1 0 206200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9871
timestamp 1654712443
transform 1 0 209200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9971
timestamp 1654712443
transform 1 0 209200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9873
timestamp 1654712443
transform 1 0 215200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9872
timestamp 1654712443
transform 1 0 212200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9973
timestamp 1654712443
transform 1 0 215200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9972
timestamp 1654712443
transform 1 0 212200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9874
timestamp 1654712443
transform 1 0 218200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9974
timestamp 1654712443
transform 1 0 218200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9875
timestamp 1654712443
transform 1 0 221200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9975
timestamp 1654712443
transform 1 0 221200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9876
timestamp 1654712443
transform 1 0 224200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9976
timestamp 1654712443
transform 1 0 224200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9877
timestamp 1654712443
transform 1 0 227200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9977
timestamp 1654712443
transform 1 0 227200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9878
timestamp 1654712443
transform 1 0 230200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9978
timestamp 1654712443
transform 1 0 230200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9879
timestamp 1654712443
transform 1 0 233200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9979
timestamp 1654712443
transform 1 0 233200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9880
timestamp 1654712443
transform 1 0 236200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9980
timestamp 1654712443
transform 1 0 236200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9881
timestamp 1654712443
transform 1 0 239200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9981
timestamp 1654712443
transform 1 0 239200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9883
timestamp 1654712443
transform 1 0 245200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9882
timestamp 1654712443
transform 1 0 242200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9983
timestamp 1654712443
transform 1 0 245200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9982
timestamp 1654712443
transform 1 0 242200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9884
timestamp 1654712443
transform 1 0 248200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9984
timestamp 1654712443
transform 1 0 248200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9885
timestamp 1654712443
transform 1 0 251200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9985
timestamp 1654712443
transform 1 0 251200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9886
timestamp 1654712443
transform 1 0 254200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9986
timestamp 1654712443
transform 1 0 254200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9887
timestamp 1654712443
transform 1 0 257200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9987
timestamp 1654712443
transform 1 0 257200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9888
timestamp 1654712443
transform 1 0 260200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9988
timestamp 1654712443
transform 1 0 260200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9889
timestamp 1654712443
transform 1 0 263200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9989
timestamp 1654712443
transform 1 0 263200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9890
timestamp 1654712443
transform 1 0 266200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9990
timestamp 1654712443
transform 1 0 266200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9891
timestamp 1654712443
transform 1 0 269200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9991
timestamp 1654712443
transform 1 0 269200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9892
timestamp 1654712443
transform 1 0 272200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9992
timestamp 1654712443
transform 1 0 272200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9893
timestamp 1654712443
transform 1 0 275200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9894
timestamp 1654712443
transform 1 0 278200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9993
timestamp 1654712443
transform 1 0 275200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9994
timestamp 1654712443
transform 1 0 278200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9895
timestamp 1654712443
transform 1 0 281200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9995
timestamp 1654712443
transform 1 0 281200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9896
timestamp 1654712443
transform 1 0 284200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9996
timestamp 1654712443
transform 1 0 284200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9897
timestamp 1654712443
transform 1 0 287200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9997
timestamp 1654712443
transform 1 0 287200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9898
timestamp 1654712443
transform 1 0 290200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9998
timestamp 1654712443
transform 1 0 290200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9899
timestamp 1654712443
transform 1 0 293200 0 1 -291300
box 3640 -2860 6960 460
use pixel  pixel_9999
timestamp 1654712443
transform 1 0 293200 0 1 -294300
box 3640 -2860 6960 460
use pixel  pixel_9701
timestamp 1654712443
transform 1 0 -800 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9700
timestamp 1654712443
transform 1 0 -3800 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9702
timestamp 1654712443
transform 1 0 2200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9703
timestamp 1654712443
transform 1 0 5200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9704
timestamp 1654712443
transform 1 0 8200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9705
timestamp 1654712443
transform 1 0 11200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9706
timestamp 1654712443
transform 1 0 14200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9707
timestamp 1654712443
transform 1 0 17200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9708
timestamp 1654712443
transform 1 0 20200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9709
timestamp 1654712443
transform 1 0 23200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9711
timestamp 1654712443
transform 1 0 29200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9710
timestamp 1654712443
transform 1 0 26200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9712
timestamp 1654712443
transform 1 0 32200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9713
timestamp 1654712443
transform 1 0 35200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9714
timestamp 1654712443
transform 1 0 38200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9715
timestamp 1654712443
transform 1 0 41200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9716
timestamp 1654712443
transform 1 0 44200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9717
timestamp 1654712443
transform 1 0 47200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9718
timestamp 1654712443
transform 1 0 50200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9719
timestamp 1654712443
transform 1 0 53200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9721
timestamp 1654712443
transform 1 0 59200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9720
timestamp 1654712443
transform 1 0 56200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9722
timestamp 1654712443
transform 1 0 62200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9723
timestamp 1654712443
transform 1 0 65200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9724
timestamp 1654712443
transform 1 0 68200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9725
timestamp 1654712443
transform 1 0 71200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9726
timestamp 1654712443
transform 1 0 74200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9727
timestamp 1654712443
transform 1 0 77200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9728
timestamp 1654712443
transform 1 0 80200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9729
timestamp 1654712443
transform 1 0 83200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9730
timestamp 1654712443
transform 1 0 86200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9731
timestamp 1654712443
transform 1 0 89200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9732
timestamp 1654712443
transform 1 0 92200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9733
timestamp 1654712443
transform 1 0 95200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9734
timestamp 1654712443
transform 1 0 98200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9735
timestamp 1654712443
transform 1 0 101200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9736
timestamp 1654712443
transform 1 0 104200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9737
timestamp 1654712443
transform 1 0 107200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9738
timestamp 1654712443
transform 1 0 110200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9739
timestamp 1654712443
transform 1 0 113200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9740
timestamp 1654712443
transform 1 0 116200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9741
timestamp 1654712443
transform 1 0 119200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9742
timestamp 1654712443
transform 1 0 122200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9743
timestamp 1654712443
transform 1 0 125200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9744
timestamp 1654712443
transform 1 0 128200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9745
timestamp 1654712443
transform 1 0 131200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9746
timestamp 1654712443
transform 1 0 134200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9747
timestamp 1654712443
transform 1 0 137200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9748
timestamp 1654712443
transform 1 0 140200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9749
timestamp 1654712443
transform 1 0 143200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9750
timestamp 1654712443
transform 1 0 146200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9751
timestamp 1654712443
transform 1 0 149200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9752
timestamp 1654712443
transform 1 0 152200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9753
timestamp 1654712443
transform 1 0 155200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9754
timestamp 1654712443
transform 1 0 158200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9755
timestamp 1654712443
transform 1 0 161200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9756
timestamp 1654712443
transform 1 0 164200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9757
timestamp 1654712443
transform 1 0 167200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9758
timestamp 1654712443
transform 1 0 170200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9759
timestamp 1654712443
transform 1 0 173200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9760
timestamp 1654712443
transform 1 0 176200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9761
timestamp 1654712443
transform 1 0 179200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9763
timestamp 1654712443
transform 1 0 185200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9762
timestamp 1654712443
transform 1 0 182200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9764
timestamp 1654712443
transform 1 0 188200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9765
timestamp 1654712443
transform 1 0 191200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9766
timestamp 1654712443
transform 1 0 194200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9767
timestamp 1654712443
transform 1 0 197200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9768
timestamp 1654712443
transform 1 0 200200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9769
timestamp 1654712443
transform 1 0 203200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9770
timestamp 1654712443
transform 1 0 206200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9771
timestamp 1654712443
transform 1 0 209200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9773
timestamp 1654712443
transform 1 0 215200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9772
timestamp 1654712443
transform 1 0 212200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9774
timestamp 1654712443
transform 1 0 218200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9775
timestamp 1654712443
transform 1 0 221200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9776
timestamp 1654712443
transform 1 0 224200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9777
timestamp 1654712443
transform 1 0 227200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9778
timestamp 1654712443
transform 1 0 230200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9779
timestamp 1654712443
transform 1 0 233200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9780
timestamp 1654712443
transform 1 0 236200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9781
timestamp 1654712443
transform 1 0 239200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9783
timestamp 1654712443
transform 1 0 245200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9782
timestamp 1654712443
transform 1 0 242200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9784
timestamp 1654712443
transform 1 0 248200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9785
timestamp 1654712443
transform 1 0 251200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9786
timestamp 1654712443
transform 1 0 254200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9787
timestamp 1654712443
transform 1 0 257200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9788
timestamp 1654712443
transform 1 0 260200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9789
timestamp 1654712443
transform 1 0 263200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9790
timestamp 1654712443
transform 1 0 266200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9791
timestamp 1654712443
transform 1 0 269200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9792
timestamp 1654712443
transform 1 0 272200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9793
timestamp 1654712443
transform 1 0 275200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9794
timestamp 1654712443
transform 1 0 278200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9795
timestamp 1654712443
transform 1 0 281200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9796
timestamp 1654712443
transform 1 0 284200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9797
timestamp 1654712443
transform 1 0 287200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9798
timestamp 1654712443
transform 1 0 290200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9799
timestamp 1654712443
transform 1 0 293200 0 1 -288300
box 3640 -2860 6960 460
use pixel  pixel_9601
timestamp 1654712443
transform 1 0 -800 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9600
timestamp 1654712443
transform 1 0 -3800 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9602
timestamp 1654712443
transform 1 0 2200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9603
timestamp 1654712443
transform 1 0 5200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9604
timestamp 1654712443
transform 1 0 8200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9605
timestamp 1654712443
transform 1 0 11200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9606
timestamp 1654712443
transform 1 0 14200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9607
timestamp 1654712443
transform 1 0 17200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9608
timestamp 1654712443
transform 1 0 20200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9609
timestamp 1654712443
transform 1 0 23200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9611
timestamp 1654712443
transform 1 0 29200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9610
timestamp 1654712443
transform 1 0 26200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9612
timestamp 1654712443
transform 1 0 32200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9613
timestamp 1654712443
transform 1 0 35200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9614
timestamp 1654712443
transform 1 0 38200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9615
timestamp 1654712443
transform 1 0 41200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9616
timestamp 1654712443
transform 1 0 44200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9617
timestamp 1654712443
transform 1 0 47200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9618
timestamp 1654712443
transform 1 0 50200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9619
timestamp 1654712443
transform 1 0 53200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9621
timestamp 1654712443
transform 1 0 59200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9620
timestamp 1654712443
transform 1 0 56200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9622
timestamp 1654712443
transform 1 0 62200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9623
timestamp 1654712443
transform 1 0 65200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9624
timestamp 1654712443
transform 1 0 68200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9625
timestamp 1654712443
transform 1 0 71200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9626
timestamp 1654712443
transform 1 0 74200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9627
timestamp 1654712443
transform 1 0 77200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9628
timestamp 1654712443
transform 1 0 80200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9629
timestamp 1654712443
transform 1 0 83200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9630
timestamp 1654712443
transform 1 0 86200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9631
timestamp 1654712443
transform 1 0 89200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9632
timestamp 1654712443
transform 1 0 92200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9633
timestamp 1654712443
transform 1 0 95200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9634
timestamp 1654712443
transform 1 0 98200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9635
timestamp 1654712443
transform 1 0 101200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9636
timestamp 1654712443
transform 1 0 104200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9637
timestamp 1654712443
transform 1 0 107200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9638
timestamp 1654712443
transform 1 0 110200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9639
timestamp 1654712443
transform 1 0 113200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9640
timestamp 1654712443
transform 1 0 116200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9641
timestamp 1654712443
transform 1 0 119200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9642
timestamp 1654712443
transform 1 0 122200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9643
timestamp 1654712443
transform 1 0 125200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9644
timestamp 1654712443
transform 1 0 128200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9645
timestamp 1654712443
transform 1 0 131200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9646
timestamp 1654712443
transform 1 0 134200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9647
timestamp 1654712443
transform 1 0 137200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9648
timestamp 1654712443
transform 1 0 140200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9649
timestamp 1654712443
transform 1 0 143200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9650
timestamp 1654712443
transform 1 0 146200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9651
timestamp 1654712443
transform 1 0 149200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9652
timestamp 1654712443
transform 1 0 152200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9653
timestamp 1654712443
transform 1 0 155200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9654
timestamp 1654712443
transform 1 0 158200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9655
timestamp 1654712443
transform 1 0 161200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9656
timestamp 1654712443
transform 1 0 164200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9657
timestamp 1654712443
transform 1 0 167200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9658
timestamp 1654712443
transform 1 0 170200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9659
timestamp 1654712443
transform 1 0 173200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9660
timestamp 1654712443
transform 1 0 176200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9661
timestamp 1654712443
transform 1 0 179200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9663
timestamp 1654712443
transform 1 0 185200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9662
timestamp 1654712443
transform 1 0 182200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9664
timestamp 1654712443
transform 1 0 188200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9665
timestamp 1654712443
transform 1 0 191200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9666
timestamp 1654712443
transform 1 0 194200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9667
timestamp 1654712443
transform 1 0 197200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9668
timestamp 1654712443
transform 1 0 200200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9669
timestamp 1654712443
transform 1 0 203200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9670
timestamp 1654712443
transform 1 0 206200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9671
timestamp 1654712443
transform 1 0 209200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9673
timestamp 1654712443
transform 1 0 215200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9672
timestamp 1654712443
transform 1 0 212200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9674
timestamp 1654712443
transform 1 0 218200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9675
timestamp 1654712443
transform 1 0 221200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9676
timestamp 1654712443
transform 1 0 224200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9677
timestamp 1654712443
transform 1 0 227200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9678
timestamp 1654712443
transform 1 0 230200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9679
timestamp 1654712443
transform 1 0 233200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9680
timestamp 1654712443
transform 1 0 236200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9681
timestamp 1654712443
transform 1 0 239200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9683
timestamp 1654712443
transform 1 0 245200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9682
timestamp 1654712443
transform 1 0 242200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9684
timestamp 1654712443
transform 1 0 248200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9685
timestamp 1654712443
transform 1 0 251200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9686
timestamp 1654712443
transform 1 0 254200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9687
timestamp 1654712443
transform 1 0 257200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9688
timestamp 1654712443
transform 1 0 260200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9689
timestamp 1654712443
transform 1 0 263200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9690
timestamp 1654712443
transform 1 0 266200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9691
timestamp 1654712443
transform 1 0 269200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9692
timestamp 1654712443
transform 1 0 272200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9693
timestamp 1654712443
transform 1 0 275200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9694
timestamp 1654712443
transform 1 0 278200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9695
timestamp 1654712443
transform 1 0 281200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9696
timestamp 1654712443
transform 1 0 284200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9697
timestamp 1654712443
transform 1 0 287200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9698
timestamp 1654712443
transform 1 0 290200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9699
timestamp 1654712443
transform 1 0 293200 0 1 -285300
box 3640 -2860 6960 460
use pixel  pixel_9501
timestamp 1654712443
transform 1 0 -800 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9500
timestamp 1654712443
transform 1 0 -3800 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9502
timestamp 1654712443
transform 1 0 2200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9503
timestamp 1654712443
transform 1 0 5200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9504
timestamp 1654712443
transform 1 0 8200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9505
timestamp 1654712443
transform 1 0 11200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9506
timestamp 1654712443
transform 1 0 14200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9507
timestamp 1654712443
transform 1 0 17200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9508
timestamp 1654712443
transform 1 0 20200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9509
timestamp 1654712443
transform 1 0 23200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9511
timestamp 1654712443
transform 1 0 29200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9510
timestamp 1654712443
transform 1 0 26200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9512
timestamp 1654712443
transform 1 0 32200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9513
timestamp 1654712443
transform 1 0 35200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9514
timestamp 1654712443
transform 1 0 38200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9515
timestamp 1654712443
transform 1 0 41200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9516
timestamp 1654712443
transform 1 0 44200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9517
timestamp 1654712443
transform 1 0 47200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9518
timestamp 1654712443
transform 1 0 50200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9519
timestamp 1654712443
transform 1 0 53200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9521
timestamp 1654712443
transform 1 0 59200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9520
timestamp 1654712443
transform 1 0 56200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9522
timestamp 1654712443
transform 1 0 62200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9523
timestamp 1654712443
transform 1 0 65200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9524
timestamp 1654712443
transform 1 0 68200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9525
timestamp 1654712443
transform 1 0 71200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9526
timestamp 1654712443
transform 1 0 74200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9527
timestamp 1654712443
transform 1 0 77200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9528
timestamp 1654712443
transform 1 0 80200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9529
timestamp 1654712443
transform 1 0 83200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9530
timestamp 1654712443
transform 1 0 86200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9531
timestamp 1654712443
transform 1 0 89200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9532
timestamp 1654712443
transform 1 0 92200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9533
timestamp 1654712443
transform 1 0 95200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9534
timestamp 1654712443
transform 1 0 98200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9535
timestamp 1654712443
transform 1 0 101200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9536
timestamp 1654712443
transform 1 0 104200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9537
timestamp 1654712443
transform 1 0 107200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9538
timestamp 1654712443
transform 1 0 110200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9539
timestamp 1654712443
transform 1 0 113200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9540
timestamp 1654712443
transform 1 0 116200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9541
timestamp 1654712443
transform 1 0 119200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9542
timestamp 1654712443
transform 1 0 122200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9543
timestamp 1654712443
transform 1 0 125200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9544
timestamp 1654712443
transform 1 0 128200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9545
timestamp 1654712443
transform 1 0 131200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9546
timestamp 1654712443
transform 1 0 134200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9547
timestamp 1654712443
transform 1 0 137200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9548
timestamp 1654712443
transform 1 0 140200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9549
timestamp 1654712443
transform 1 0 143200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9550
timestamp 1654712443
transform 1 0 146200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9551
timestamp 1654712443
transform 1 0 149200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9552
timestamp 1654712443
transform 1 0 152200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9553
timestamp 1654712443
transform 1 0 155200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9554
timestamp 1654712443
transform 1 0 158200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9555
timestamp 1654712443
transform 1 0 161200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9556
timestamp 1654712443
transform 1 0 164200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9557
timestamp 1654712443
transform 1 0 167200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9558
timestamp 1654712443
transform 1 0 170200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9559
timestamp 1654712443
transform 1 0 173200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9560
timestamp 1654712443
transform 1 0 176200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9561
timestamp 1654712443
transform 1 0 179200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9563
timestamp 1654712443
transform 1 0 185200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9562
timestamp 1654712443
transform 1 0 182200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9564
timestamp 1654712443
transform 1 0 188200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9565
timestamp 1654712443
transform 1 0 191200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9566
timestamp 1654712443
transform 1 0 194200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9567
timestamp 1654712443
transform 1 0 197200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9568
timestamp 1654712443
transform 1 0 200200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9569
timestamp 1654712443
transform 1 0 203200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9570
timestamp 1654712443
transform 1 0 206200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9571
timestamp 1654712443
transform 1 0 209200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9573
timestamp 1654712443
transform 1 0 215200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9572
timestamp 1654712443
transform 1 0 212200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9574
timestamp 1654712443
transform 1 0 218200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9575
timestamp 1654712443
transform 1 0 221200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9576
timestamp 1654712443
transform 1 0 224200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9577
timestamp 1654712443
transform 1 0 227200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9578
timestamp 1654712443
transform 1 0 230200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9579
timestamp 1654712443
transform 1 0 233200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9580
timestamp 1654712443
transform 1 0 236200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9581
timestamp 1654712443
transform 1 0 239200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9583
timestamp 1654712443
transform 1 0 245200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9582
timestamp 1654712443
transform 1 0 242200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9584
timestamp 1654712443
transform 1 0 248200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9585
timestamp 1654712443
transform 1 0 251200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9586
timestamp 1654712443
transform 1 0 254200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9587
timestamp 1654712443
transform 1 0 257200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9588
timestamp 1654712443
transform 1 0 260200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9589
timestamp 1654712443
transform 1 0 263200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9590
timestamp 1654712443
transform 1 0 266200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9591
timestamp 1654712443
transform 1 0 269200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9592
timestamp 1654712443
transform 1 0 272200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9593
timestamp 1654712443
transform 1 0 275200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9594
timestamp 1654712443
transform 1 0 278200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9595
timestamp 1654712443
transform 1 0 281200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9596
timestamp 1654712443
transform 1 0 284200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9597
timestamp 1654712443
transform 1 0 287200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9598
timestamp 1654712443
transform 1 0 290200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9599
timestamp 1654712443
transform 1 0 293200 0 1 -282300
box 3640 -2860 6960 460
use pixel  pixel_9401
timestamp 1654712443
transform 1 0 -800 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9400
timestamp 1654712443
transform 1 0 -3800 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9402
timestamp 1654712443
transform 1 0 2200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9403
timestamp 1654712443
transform 1 0 5200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9404
timestamp 1654712443
transform 1 0 8200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9405
timestamp 1654712443
transform 1 0 11200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9406
timestamp 1654712443
transform 1 0 14200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9407
timestamp 1654712443
transform 1 0 17200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9408
timestamp 1654712443
transform 1 0 20200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9409
timestamp 1654712443
transform 1 0 23200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9411
timestamp 1654712443
transform 1 0 29200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9410
timestamp 1654712443
transform 1 0 26200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9412
timestamp 1654712443
transform 1 0 32200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9413
timestamp 1654712443
transform 1 0 35200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9414
timestamp 1654712443
transform 1 0 38200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9415
timestamp 1654712443
transform 1 0 41200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9416
timestamp 1654712443
transform 1 0 44200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9417
timestamp 1654712443
transform 1 0 47200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9418
timestamp 1654712443
transform 1 0 50200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9419
timestamp 1654712443
transform 1 0 53200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9421
timestamp 1654712443
transform 1 0 59200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9420
timestamp 1654712443
transform 1 0 56200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9422
timestamp 1654712443
transform 1 0 62200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9423
timestamp 1654712443
transform 1 0 65200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9424
timestamp 1654712443
transform 1 0 68200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9425
timestamp 1654712443
transform 1 0 71200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9426
timestamp 1654712443
transform 1 0 74200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9427
timestamp 1654712443
transform 1 0 77200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9428
timestamp 1654712443
transform 1 0 80200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9429
timestamp 1654712443
transform 1 0 83200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9430
timestamp 1654712443
transform 1 0 86200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9431
timestamp 1654712443
transform 1 0 89200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9432
timestamp 1654712443
transform 1 0 92200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9433
timestamp 1654712443
transform 1 0 95200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9434
timestamp 1654712443
transform 1 0 98200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9435
timestamp 1654712443
transform 1 0 101200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9436
timestamp 1654712443
transform 1 0 104200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9437
timestamp 1654712443
transform 1 0 107200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9438
timestamp 1654712443
transform 1 0 110200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9439
timestamp 1654712443
transform 1 0 113200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9440
timestamp 1654712443
transform 1 0 116200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9441
timestamp 1654712443
transform 1 0 119200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9442
timestamp 1654712443
transform 1 0 122200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9443
timestamp 1654712443
transform 1 0 125200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9444
timestamp 1654712443
transform 1 0 128200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9445
timestamp 1654712443
transform 1 0 131200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9446
timestamp 1654712443
transform 1 0 134200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9447
timestamp 1654712443
transform 1 0 137200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9448
timestamp 1654712443
transform 1 0 140200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9449
timestamp 1654712443
transform 1 0 143200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9450
timestamp 1654712443
transform 1 0 146200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9451
timestamp 1654712443
transform 1 0 149200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9452
timestamp 1654712443
transform 1 0 152200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9453
timestamp 1654712443
transform 1 0 155200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9454
timestamp 1654712443
transform 1 0 158200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9455
timestamp 1654712443
transform 1 0 161200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9456
timestamp 1654712443
transform 1 0 164200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9457
timestamp 1654712443
transform 1 0 167200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9458
timestamp 1654712443
transform 1 0 170200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9459
timestamp 1654712443
transform 1 0 173200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9460
timestamp 1654712443
transform 1 0 176200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9461
timestamp 1654712443
transform 1 0 179200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9463
timestamp 1654712443
transform 1 0 185200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9462
timestamp 1654712443
transform 1 0 182200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9464
timestamp 1654712443
transform 1 0 188200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9465
timestamp 1654712443
transform 1 0 191200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9466
timestamp 1654712443
transform 1 0 194200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9467
timestamp 1654712443
transform 1 0 197200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9468
timestamp 1654712443
transform 1 0 200200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9469
timestamp 1654712443
transform 1 0 203200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9470
timestamp 1654712443
transform 1 0 206200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9471
timestamp 1654712443
transform 1 0 209200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9473
timestamp 1654712443
transform 1 0 215200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9472
timestamp 1654712443
transform 1 0 212200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9474
timestamp 1654712443
transform 1 0 218200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9475
timestamp 1654712443
transform 1 0 221200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9476
timestamp 1654712443
transform 1 0 224200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9477
timestamp 1654712443
transform 1 0 227200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9478
timestamp 1654712443
transform 1 0 230200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9479
timestamp 1654712443
transform 1 0 233200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9480
timestamp 1654712443
transform 1 0 236200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9481
timestamp 1654712443
transform 1 0 239200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9483
timestamp 1654712443
transform 1 0 245200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9482
timestamp 1654712443
transform 1 0 242200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9484
timestamp 1654712443
transform 1 0 248200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9485
timestamp 1654712443
transform 1 0 251200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9486
timestamp 1654712443
transform 1 0 254200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9487
timestamp 1654712443
transform 1 0 257200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9488
timestamp 1654712443
transform 1 0 260200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9489
timestamp 1654712443
transform 1 0 263200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9490
timestamp 1654712443
transform 1 0 266200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9491
timestamp 1654712443
transform 1 0 269200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9492
timestamp 1654712443
transform 1 0 272200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9493
timestamp 1654712443
transform 1 0 275200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9494
timestamp 1654712443
transform 1 0 278200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9495
timestamp 1654712443
transform 1 0 281200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9496
timestamp 1654712443
transform 1 0 284200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9497
timestamp 1654712443
transform 1 0 287200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9498
timestamp 1654712443
transform 1 0 290200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9499
timestamp 1654712443
transform 1 0 293200 0 1 -279300
box 3640 -2860 6960 460
use pixel  pixel_9301
timestamp 1654712443
transform 1 0 -800 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9300
timestamp 1654712443
transform 1 0 -3800 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9302
timestamp 1654712443
transform 1 0 2200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9303
timestamp 1654712443
transform 1 0 5200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9304
timestamp 1654712443
transform 1 0 8200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9305
timestamp 1654712443
transform 1 0 11200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9306
timestamp 1654712443
transform 1 0 14200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9307
timestamp 1654712443
transform 1 0 17200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9308
timestamp 1654712443
transform 1 0 20200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9309
timestamp 1654712443
transform 1 0 23200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9311
timestamp 1654712443
transform 1 0 29200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9310
timestamp 1654712443
transform 1 0 26200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9312
timestamp 1654712443
transform 1 0 32200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9313
timestamp 1654712443
transform 1 0 35200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9314
timestamp 1654712443
transform 1 0 38200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9315
timestamp 1654712443
transform 1 0 41200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9316
timestamp 1654712443
transform 1 0 44200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9317
timestamp 1654712443
transform 1 0 47200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9318
timestamp 1654712443
transform 1 0 50200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9319
timestamp 1654712443
transform 1 0 53200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9321
timestamp 1654712443
transform 1 0 59200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9320
timestamp 1654712443
transform 1 0 56200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9322
timestamp 1654712443
transform 1 0 62200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9323
timestamp 1654712443
transform 1 0 65200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9324
timestamp 1654712443
transform 1 0 68200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9325
timestamp 1654712443
transform 1 0 71200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9326
timestamp 1654712443
transform 1 0 74200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9327
timestamp 1654712443
transform 1 0 77200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9328
timestamp 1654712443
transform 1 0 80200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9329
timestamp 1654712443
transform 1 0 83200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9330
timestamp 1654712443
transform 1 0 86200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9331
timestamp 1654712443
transform 1 0 89200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9332
timestamp 1654712443
transform 1 0 92200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9333
timestamp 1654712443
transform 1 0 95200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9334
timestamp 1654712443
transform 1 0 98200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9335
timestamp 1654712443
transform 1 0 101200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9336
timestamp 1654712443
transform 1 0 104200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9337
timestamp 1654712443
transform 1 0 107200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9338
timestamp 1654712443
transform 1 0 110200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9339
timestamp 1654712443
transform 1 0 113200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9340
timestamp 1654712443
transform 1 0 116200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9341
timestamp 1654712443
transform 1 0 119200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9342
timestamp 1654712443
transform 1 0 122200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9343
timestamp 1654712443
transform 1 0 125200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9344
timestamp 1654712443
transform 1 0 128200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9345
timestamp 1654712443
transform 1 0 131200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9346
timestamp 1654712443
transform 1 0 134200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9347
timestamp 1654712443
transform 1 0 137200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9348
timestamp 1654712443
transform 1 0 140200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9349
timestamp 1654712443
transform 1 0 143200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9350
timestamp 1654712443
transform 1 0 146200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9351
timestamp 1654712443
transform 1 0 149200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9352
timestamp 1654712443
transform 1 0 152200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9353
timestamp 1654712443
transform 1 0 155200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9354
timestamp 1654712443
transform 1 0 158200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9355
timestamp 1654712443
transform 1 0 161200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9356
timestamp 1654712443
transform 1 0 164200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9357
timestamp 1654712443
transform 1 0 167200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9358
timestamp 1654712443
transform 1 0 170200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9359
timestamp 1654712443
transform 1 0 173200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9360
timestamp 1654712443
transform 1 0 176200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9361
timestamp 1654712443
transform 1 0 179200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9363
timestamp 1654712443
transform 1 0 185200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9362
timestamp 1654712443
transform 1 0 182200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9364
timestamp 1654712443
transform 1 0 188200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9365
timestamp 1654712443
transform 1 0 191200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9366
timestamp 1654712443
transform 1 0 194200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9367
timestamp 1654712443
transform 1 0 197200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9368
timestamp 1654712443
transform 1 0 200200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9369
timestamp 1654712443
transform 1 0 203200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9370
timestamp 1654712443
transform 1 0 206200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9371
timestamp 1654712443
transform 1 0 209200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9373
timestamp 1654712443
transform 1 0 215200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9372
timestamp 1654712443
transform 1 0 212200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9374
timestamp 1654712443
transform 1 0 218200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9375
timestamp 1654712443
transform 1 0 221200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9376
timestamp 1654712443
transform 1 0 224200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9377
timestamp 1654712443
transform 1 0 227200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9378
timestamp 1654712443
transform 1 0 230200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9379
timestamp 1654712443
transform 1 0 233200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9380
timestamp 1654712443
transform 1 0 236200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9381
timestamp 1654712443
transform 1 0 239200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9383
timestamp 1654712443
transform 1 0 245200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9382
timestamp 1654712443
transform 1 0 242200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9384
timestamp 1654712443
transform 1 0 248200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9385
timestamp 1654712443
transform 1 0 251200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9386
timestamp 1654712443
transform 1 0 254200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9387
timestamp 1654712443
transform 1 0 257200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9388
timestamp 1654712443
transform 1 0 260200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9389
timestamp 1654712443
transform 1 0 263200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9390
timestamp 1654712443
transform 1 0 266200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9391
timestamp 1654712443
transform 1 0 269200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9392
timestamp 1654712443
transform 1 0 272200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9393
timestamp 1654712443
transform 1 0 275200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9394
timestamp 1654712443
transform 1 0 278200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9395
timestamp 1654712443
transform 1 0 281200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9396
timestamp 1654712443
transform 1 0 284200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9397
timestamp 1654712443
transform 1 0 287200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9398
timestamp 1654712443
transform 1 0 290200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9399
timestamp 1654712443
transform 1 0 293200 0 1 -276300
box 3640 -2860 6960 460
use pixel  pixel_9201
timestamp 1654712443
transform 1 0 -800 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9200
timestamp 1654712443
transform 1 0 -3800 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9202
timestamp 1654712443
transform 1 0 2200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9203
timestamp 1654712443
transform 1 0 5200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9204
timestamp 1654712443
transform 1 0 8200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9205
timestamp 1654712443
transform 1 0 11200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9206
timestamp 1654712443
transform 1 0 14200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9207
timestamp 1654712443
transform 1 0 17200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9208
timestamp 1654712443
transform 1 0 20200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9209
timestamp 1654712443
transform 1 0 23200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9211
timestamp 1654712443
transform 1 0 29200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9210
timestamp 1654712443
transform 1 0 26200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9212
timestamp 1654712443
transform 1 0 32200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9213
timestamp 1654712443
transform 1 0 35200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9214
timestamp 1654712443
transform 1 0 38200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9215
timestamp 1654712443
transform 1 0 41200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9216
timestamp 1654712443
transform 1 0 44200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9217
timestamp 1654712443
transform 1 0 47200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9218
timestamp 1654712443
transform 1 0 50200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9219
timestamp 1654712443
transform 1 0 53200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9221
timestamp 1654712443
transform 1 0 59200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9220
timestamp 1654712443
transform 1 0 56200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9222
timestamp 1654712443
transform 1 0 62200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9223
timestamp 1654712443
transform 1 0 65200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9224
timestamp 1654712443
transform 1 0 68200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9225
timestamp 1654712443
transform 1 0 71200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9226
timestamp 1654712443
transform 1 0 74200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9227
timestamp 1654712443
transform 1 0 77200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9228
timestamp 1654712443
transform 1 0 80200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9229
timestamp 1654712443
transform 1 0 83200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9230
timestamp 1654712443
transform 1 0 86200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9231
timestamp 1654712443
transform 1 0 89200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9232
timestamp 1654712443
transform 1 0 92200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9233
timestamp 1654712443
transform 1 0 95200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9234
timestamp 1654712443
transform 1 0 98200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9235
timestamp 1654712443
transform 1 0 101200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9236
timestamp 1654712443
transform 1 0 104200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9237
timestamp 1654712443
transform 1 0 107200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9238
timestamp 1654712443
transform 1 0 110200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9239
timestamp 1654712443
transform 1 0 113200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9240
timestamp 1654712443
transform 1 0 116200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9241
timestamp 1654712443
transform 1 0 119200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9242
timestamp 1654712443
transform 1 0 122200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9243
timestamp 1654712443
transform 1 0 125200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9244
timestamp 1654712443
transform 1 0 128200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9245
timestamp 1654712443
transform 1 0 131200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9246
timestamp 1654712443
transform 1 0 134200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9247
timestamp 1654712443
transform 1 0 137200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9248
timestamp 1654712443
transform 1 0 140200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9249
timestamp 1654712443
transform 1 0 143200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9250
timestamp 1654712443
transform 1 0 146200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9251
timestamp 1654712443
transform 1 0 149200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9252
timestamp 1654712443
transform 1 0 152200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9253
timestamp 1654712443
transform 1 0 155200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9254
timestamp 1654712443
transform 1 0 158200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9255
timestamp 1654712443
transform 1 0 161200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9256
timestamp 1654712443
transform 1 0 164200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9257
timestamp 1654712443
transform 1 0 167200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9258
timestamp 1654712443
transform 1 0 170200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9259
timestamp 1654712443
transform 1 0 173200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9260
timestamp 1654712443
transform 1 0 176200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9261
timestamp 1654712443
transform 1 0 179200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9263
timestamp 1654712443
transform 1 0 185200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9262
timestamp 1654712443
transform 1 0 182200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9264
timestamp 1654712443
transform 1 0 188200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9265
timestamp 1654712443
transform 1 0 191200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9266
timestamp 1654712443
transform 1 0 194200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9267
timestamp 1654712443
transform 1 0 197200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9268
timestamp 1654712443
transform 1 0 200200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9269
timestamp 1654712443
transform 1 0 203200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9270
timestamp 1654712443
transform 1 0 206200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9271
timestamp 1654712443
transform 1 0 209200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9273
timestamp 1654712443
transform 1 0 215200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9272
timestamp 1654712443
transform 1 0 212200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9274
timestamp 1654712443
transform 1 0 218200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9275
timestamp 1654712443
transform 1 0 221200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9276
timestamp 1654712443
transform 1 0 224200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9277
timestamp 1654712443
transform 1 0 227200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9278
timestamp 1654712443
transform 1 0 230200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9279
timestamp 1654712443
transform 1 0 233200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9280
timestamp 1654712443
transform 1 0 236200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9281
timestamp 1654712443
transform 1 0 239200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9283
timestamp 1654712443
transform 1 0 245200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9282
timestamp 1654712443
transform 1 0 242200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9284
timestamp 1654712443
transform 1 0 248200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9285
timestamp 1654712443
transform 1 0 251200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9286
timestamp 1654712443
transform 1 0 254200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9287
timestamp 1654712443
transform 1 0 257200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9288
timestamp 1654712443
transform 1 0 260200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9289
timestamp 1654712443
transform 1 0 263200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9290
timestamp 1654712443
transform 1 0 266200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9291
timestamp 1654712443
transform 1 0 269200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9292
timestamp 1654712443
transform 1 0 272200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9293
timestamp 1654712443
transform 1 0 275200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9294
timestamp 1654712443
transform 1 0 278200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9295
timestamp 1654712443
transform 1 0 281200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9296
timestamp 1654712443
transform 1 0 284200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9297
timestamp 1654712443
transform 1 0 287200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9298
timestamp 1654712443
transform 1 0 290200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9299
timestamp 1654712443
transform 1 0 293200 0 1 -273300
box 3640 -2860 6960 460
use pixel  pixel_9101
timestamp 1654712443
transform 1 0 -800 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9100
timestamp 1654712443
transform 1 0 -3800 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9102
timestamp 1654712443
transform 1 0 2200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9103
timestamp 1654712443
transform 1 0 5200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9104
timestamp 1654712443
transform 1 0 8200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9105
timestamp 1654712443
transform 1 0 11200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9106
timestamp 1654712443
transform 1 0 14200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9107
timestamp 1654712443
transform 1 0 17200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9108
timestamp 1654712443
transform 1 0 20200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9109
timestamp 1654712443
transform 1 0 23200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9111
timestamp 1654712443
transform 1 0 29200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9110
timestamp 1654712443
transform 1 0 26200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9112
timestamp 1654712443
transform 1 0 32200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9113
timestamp 1654712443
transform 1 0 35200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9114
timestamp 1654712443
transform 1 0 38200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9115
timestamp 1654712443
transform 1 0 41200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9116
timestamp 1654712443
transform 1 0 44200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9117
timestamp 1654712443
transform 1 0 47200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9118
timestamp 1654712443
transform 1 0 50200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9119
timestamp 1654712443
transform 1 0 53200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9121
timestamp 1654712443
transform 1 0 59200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9120
timestamp 1654712443
transform 1 0 56200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9122
timestamp 1654712443
transform 1 0 62200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9123
timestamp 1654712443
transform 1 0 65200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9124
timestamp 1654712443
transform 1 0 68200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9125
timestamp 1654712443
transform 1 0 71200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9126
timestamp 1654712443
transform 1 0 74200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9127
timestamp 1654712443
transform 1 0 77200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9128
timestamp 1654712443
transform 1 0 80200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9129
timestamp 1654712443
transform 1 0 83200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9130
timestamp 1654712443
transform 1 0 86200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9131
timestamp 1654712443
transform 1 0 89200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9132
timestamp 1654712443
transform 1 0 92200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9133
timestamp 1654712443
transform 1 0 95200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9134
timestamp 1654712443
transform 1 0 98200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9135
timestamp 1654712443
transform 1 0 101200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9136
timestamp 1654712443
transform 1 0 104200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9137
timestamp 1654712443
transform 1 0 107200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9138
timestamp 1654712443
transform 1 0 110200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9139
timestamp 1654712443
transform 1 0 113200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9140
timestamp 1654712443
transform 1 0 116200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9141
timestamp 1654712443
transform 1 0 119200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9142
timestamp 1654712443
transform 1 0 122200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9143
timestamp 1654712443
transform 1 0 125200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9144
timestamp 1654712443
transform 1 0 128200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9145
timestamp 1654712443
transform 1 0 131200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9146
timestamp 1654712443
transform 1 0 134200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9147
timestamp 1654712443
transform 1 0 137200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9148
timestamp 1654712443
transform 1 0 140200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9149
timestamp 1654712443
transform 1 0 143200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9150
timestamp 1654712443
transform 1 0 146200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9151
timestamp 1654712443
transform 1 0 149200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9152
timestamp 1654712443
transform 1 0 152200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9153
timestamp 1654712443
transform 1 0 155200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9154
timestamp 1654712443
transform 1 0 158200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9155
timestamp 1654712443
transform 1 0 161200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9156
timestamp 1654712443
transform 1 0 164200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9157
timestamp 1654712443
transform 1 0 167200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9158
timestamp 1654712443
transform 1 0 170200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9159
timestamp 1654712443
transform 1 0 173200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9160
timestamp 1654712443
transform 1 0 176200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9161
timestamp 1654712443
transform 1 0 179200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9163
timestamp 1654712443
transform 1 0 185200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9162
timestamp 1654712443
transform 1 0 182200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9164
timestamp 1654712443
transform 1 0 188200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9165
timestamp 1654712443
transform 1 0 191200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9166
timestamp 1654712443
transform 1 0 194200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9167
timestamp 1654712443
transform 1 0 197200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9168
timestamp 1654712443
transform 1 0 200200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9169
timestamp 1654712443
transform 1 0 203200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9170
timestamp 1654712443
transform 1 0 206200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9171
timestamp 1654712443
transform 1 0 209200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9173
timestamp 1654712443
transform 1 0 215200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9172
timestamp 1654712443
transform 1 0 212200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9174
timestamp 1654712443
transform 1 0 218200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9175
timestamp 1654712443
transform 1 0 221200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9176
timestamp 1654712443
transform 1 0 224200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9177
timestamp 1654712443
transform 1 0 227200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9178
timestamp 1654712443
transform 1 0 230200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9179
timestamp 1654712443
transform 1 0 233200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9180
timestamp 1654712443
transform 1 0 236200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9181
timestamp 1654712443
transform 1 0 239200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9183
timestamp 1654712443
transform 1 0 245200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9182
timestamp 1654712443
transform 1 0 242200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9184
timestamp 1654712443
transform 1 0 248200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9185
timestamp 1654712443
transform 1 0 251200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9186
timestamp 1654712443
transform 1 0 254200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9187
timestamp 1654712443
transform 1 0 257200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9188
timestamp 1654712443
transform 1 0 260200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9189
timestamp 1654712443
transform 1 0 263200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9190
timestamp 1654712443
transform 1 0 266200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9191
timestamp 1654712443
transform 1 0 269200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9192
timestamp 1654712443
transform 1 0 272200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9193
timestamp 1654712443
transform 1 0 275200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9194
timestamp 1654712443
transform 1 0 278200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9195
timestamp 1654712443
transform 1 0 281200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9196
timestamp 1654712443
transform 1 0 284200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9197
timestamp 1654712443
transform 1 0 287200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9198
timestamp 1654712443
transform 1 0 290200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9199
timestamp 1654712443
transform 1 0 293200 0 1 -270300
box 3640 -2860 6960 460
use pixel  pixel_9001
timestamp 1654712443
transform 1 0 -800 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9000
timestamp 1654712443
transform 1 0 -3800 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9002
timestamp 1654712443
transform 1 0 2200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9003
timestamp 1654712443
transform 1 0 5200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9004
timestamp 1654712443
transform 1 0 8200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9005
timestamp 1654712443
transform 1 0 11200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9006
timestamp 1654712443
transform 1 0 14200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9007
timestamp 1654712443
transform 1 0 17200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9008
timestamp 1654712443
transform 1 0 20200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9009
timestamp 1654712443
transform 1 0 23200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9011
timestamp 1654712443
transform 1 0 29200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9010
timestamp 1654712443
transform 1 0 26200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9012
timestamp 1654712443
transform 1 0 32200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9013
timestamp 1654712443
transform 1 0 35200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9014
timestamp 1654712443
transform 1 0 38200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9015
timestamp 1654712443
transform 1 0 41200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9016
timestamp 1654712443
transform 1 0 44200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9017
timestamp 1654712443
transform 1 0 47200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9018
timestamp 1654712443
transform 1 0 50200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9019
timestamp 1654712443
transform 1 0 53200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9021
timestamp 1654712443
transform 1 0 59200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9020
timestamp 1654712443
transform 1 0 56200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9022
timestamp 1654712443
transform 1 0 62200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9023
timestamp 1654712443
transform 1 0 65200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9024
timestamp 1654712443
transform 1 0 68200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9025
timestamp 1654712443
transform 1 0 71200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9026
timestamp 1654712443
transform 1 0 74200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9027
timestamp 1654712443
transform 1 0 77200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9028
timestamp 1654712443
transform 1 0 80200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9029
timestamp 1654712443
transform 1 0 83200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9030
timestamp 1654712443
transform 1 0 86200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9031
timestamp 1654712443
transform 1 0 89200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9032
timestamp 1654712443
transform 1 0 92200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9033
timestamp 1654712443
transform 1 0 95200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9034
timestamp 1654712443
transform 1 0 98200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9035
timestamp 1654712443
transform 1 0 101200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9036
timestamp 1654712443
transform 1 0 104200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9037
timestamp 1654712443
transform 1 0 107200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9038
timestamp 1654712443
transform 1 0 110200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9039
timestamp 1654712443
transform 1 0 113200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9040
timestamp 1654712443
transform 1 0 116200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9041
timestamp 1654712443
transform 1 0 119200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9042
timestamp 1654712443
transform 1 0 122200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9043
timestamp 1654712443
transform 1 0 125200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9044
timestamp 1654712443
transform 1 0 128200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9045
timestamp 1654712443
transform 1 0 131200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9046
timestamp 1654712443
transform 1 0 134200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9047
timestamp 1654712443
transform 1 0 137200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9048
timestamp 1654712443
transform 1 0 140200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9049
timestamp 1654712443
transform 1 0 143200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9050
timestamp 1654712443
transform 1 0 146200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9051
timestamp 1654712443
transform 1 0 149200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9052
timestamp 1654712443
transform 1 0 152200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9053
timestamp 1654712443
transform 1 0 155200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9054
timestamp 1654712443
transform 1 0 158200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9055
timestamp 1654712443
transform 1 0 161200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9056
timestamp 1654712443
transform 1 0 164200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9057
timestamp 1654712443
transform 1 0 167200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9058
timestamp 1654712443
transform 1 0 170200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9059
timestamp 1654712443
transform 1 0 173200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9060
timestamp 1654712443
transform 1 0 176200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9061
timestamp 1654712443
transform 1 0 179200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9063
timestamp 1654712443
transform 1 0 185200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9062
timestamp 1654712443
transform 1 0 182200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9064
timestamp 1654712443
transform 1 0 188200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9065
timestamp 1654712443
transform 1 0 191200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9066
timestamp 1654712443
transform 1 0 194200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9067
timestamp 1654712443
transform 1 0 197200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9068
timestamp 1654712443
transform 1 0 200200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9069
timestamp 1654712443
transform 1 0 203200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9070
timestamp 1654712443
transform 1 0 206200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9071
timestamp 1654712443
transform 1 0 209200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9073
timestamp 1654712443
transform 1 0 215200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9072
timestamp 1654712443
transform 1 0 212200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9074
timestamp 1654712443
transform 1 0 218200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9075
timestamp 1654712443
transform 1 0 221200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9076
timestamp 1654712443
transform 1 0 224200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9077
timestamp 1654712443
transform 1 0 227200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9078
timestamp 1654712443
transform 1 0 230200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9079
timestamp 1654712443
transform 1 0 233200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9080
timestamp 1654712443
transform 1 0 236200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9081
timestamp 1654712443
transform 1 0 239200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9083
timestamp 1654712443
transform 1 0 245200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9082
timestamp 1654712443
transform 1 0 242200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9084
timestamp 1654712443
transform 1 0 248200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9085
timestamp 1654712443
transform 1 0 251200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9086
timestamp 1654712443
transform 1 0 254200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9087
timestamp 1654712443
transform 1 0 257200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9088
timestamp 1654712443
transform 1 0 260200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9089
timestamp 1654712443
transform 1 0 263200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9090
timestamp 1654712443
transform 1 0 266200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9091
timestamp 1654712443
transform 1 0 269200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9092
timestamp 1654712443
transform 1 0 272200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9094
timestamp 1654712443
transform 1 0 278200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9093
timestamp 1654712443
transform 1 0 275200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9095
timestamp 1654712443
transform 1 0 281200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9096
timestamp 1654712443
transform 1 0 284200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9097
timestamp 1654712443
transform 1 0 287200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9098
timestamp 1654712443
transform 1 0 290200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_9099
timestamp 1654712443
transform 1 0 293200 0 1 -267300
box 3640 -2860 6960 460
use pixel  pixel_8801
timestamp 1654712443
transform 1 0 -800 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8800
timestamp 1654712443
transform 1 0 -3800 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8901
timestamp 1654712443
transform 1 0 -800 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8900
timestamp 1654712443
transform 1 0 -3800 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8802
timestamp 1654712443
transform 1 0 2200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8902
timestamp 1654712443
transform 1 0 2200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8803
timestamp 1654712443
transform 1 0 5200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8903
timestamp 1654712443
transform 1 0 5200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8804
timestamp 1654712443
transform 1 0 8200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8904
timestamp 1654712443
transform 1 0 8200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8805
timestamp 1654712443
transform 1 0 11200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8905
timestamp 1654712443
transform 1 0 11200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8806
timestamp 1654712443
transform 1 0 14200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8906
timestamp 1654712443
transform 1 0 14200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8807
timestamp 1654712443
transform 1 0 17200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8907
timestamp 1654712443
transform 1 0 17200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8808
timestamp 1654712443
transform 1 0 20200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8908
timestamp 1654712443
transform 1 0 20200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8809
timestamp 1654712443
transform 1 0 23200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8909
timestamp 1654712443
transform 1 0 23200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8811
timestamp 1654712443
transform 1 0 29200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8810
timestamp 1654712443
transform 1 0 26200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8911
timestamp 1654712443
transform 1 0 29200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8910
timestamp 1654712443
transform 1 0 26200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8812
timestamp 1654712443
transform 1 0 32200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8912
timestamp 1654712443
transform 1 0 32200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8813
timestamp 1654712443
transform 1 0 35200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8913
timestamp 1654712443
transform 1 0 35200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8814
timestamp 1654712443
transform 1 0 38200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8914
timestamp 1654712443
transform 1 0 38200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8815
timestamp 1654712443
transform 1 0 41200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8915
timestamp 1654712443
transform 1 0 41200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8816
timestamp 1654712443
transform 1 0 44200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8916
timestamp 1654712443
transform 1 0 44200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8817
timestamp 1654712443
transform 1 0 47200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8917
timestamp 1654712443
transform 1 0 47200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8818
timestamp 1654712443
transform 1 0 50200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8918
timestamp 1654712443
transform 1 0 50200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8819
timestamp 1654712443
transform 1 0 53200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8919
timestamp 1654712443
transform 1 0 53200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8821
timestamp 1654712443
transform 1 0 59200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8820
timestamp 1654712443
transform 1 0 56200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8921
timestamp 1654712443
transform 1 0 59200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8920
timestamp 1654712443
transform 1 0 56200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8822
timestamp 1654712443
transform 1 0 62200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8922
timestamp 1654712443
transform 1 0 62200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8823
timestamp 1654712443
transform 1 0 65200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8923
timestamp 1654712443
transform 1 0 65200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8824
timestamp 1654712443
transform 1 0 68200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8924
timestamp 1654712443
transform 1 0 68200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8825
timestamp 1654712443
transform 1 0 71200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8925
timestamp 1654712443
transform 1 0 71200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8826
timestamp 1654712443
transform 1 0 74200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8926
timestamp 1654712443
transform 1 0 74200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8827
timestamp 1654712443
transform 1 0 77200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8927
timestamp 1654712443
transform 1 0 77200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8828
timestamp 1654712443
transform 1 0 80200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8928
timestamp 1654712443
transform 1 0 80200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8829
timestamp 1654712443
transform 1 0 83200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8929
timestamp 1654712443
transform 1 0 83200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8830
timestamp 1654712443
transform 1 0 86200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8930
timestamp 1654712443
transform 1 0 86200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8831
timestamp 1654712443
transform 1 0 89200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8832
timestamp 1654712443
transform 1 0 92200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8931
timestamp 1654712443
transform 1 0 89200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8932
timestamp 1654712443
transform 1 0 92200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8833
timestamp 1654712443
transform 1 0 95200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8933
timestamp 1654712443
transform 1 0 95200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8834
timestamp 1654712443
transform 1 0 98200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8934
timestamp 1654712443
transform 1 0 98200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8835
timestamp 1654712443
transform 1 0 101200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8935
timestamp 1654712443
transform 1 0 101200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8836
timestamp 1654712443
transform 1 0 104200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8936
timestamp 1654712443
transform 1 0 104200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8837
timestamp 1654712443
transform 1 0 107200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8937
timestamp 1654712443
transform 1 0 107200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8838
timestamp 1654712443
transform 1 0 110200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8938
timestamp 1654712443
transform 1 0 110200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8839
timestamp 1654712443
transform 1 0 113200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8939
timestamp 1654712443
transform 1 0 113200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8840
timestamp 1654712443
transform 1 0 116200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8940
timestamp 1654712443
transform 1 0 116200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8841
timestamp 1654712443
transform 1 0 119200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8842
timestamp 1654712443
transform 1 0 122200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8941
timestamp 1654712443
transform 1 0 119200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8942
timestamp 1654712443
transform 1 0 122200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8843
timestamp 1654712443
transform 1 0 125200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8943
timestamp 1654712443
transform 1 0 125200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8844
timestamp 1654712443
transform 1 0 128200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8944
timestamp 1654712443
transform 1 0 128200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8845
timestamp 1654712443
transform 1 0 131200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8945
timestamp 1654712443
transform 1 0 131200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8846
timestamp 1654712443
transform 1 0 134200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8946
timestamp 1654712443
transform 1 0 134200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8847
timestamp 1654712443
transform 1 0 137200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8947
timestamp 1654712443
transform 1 0 137200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8848
timestamp 1654712443
transform 1 0 140200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8948
timestamp 1654712443
transform 1 0 140200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8849
timestamp 1654712443
transform 1 0 143200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8949
timestamp 1654712443
transform 1 0 143200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8850
timestamp 1654712443
transform 1 0 146200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8950
timestamp 1654712443
transform 1 0 146200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8851
timestamp 1654712443
transform 1 0 149200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8852
timestamp 1654712443
transform 1 0 152200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8951
timestamp 1654712443
transform 1 0 149200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8952
timestamp 1654712443
transform 1 0 152200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8853
timestamp 1654712443
transform 1 0 155200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8953
timestamp 1654712443
transform 1 0 155200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8854
timestamp 1654712443
transform 1 0 158200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8954
timestamp 1654712443
transform 1 0 158200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8855
timestamp 1654712443
transform 1 0 161200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8955
timestamp 1654712443
transform 1 0 161200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8856
timestamp 1654712443
transform 1 0 164200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8956
timestamp 1654712443
transform 1 0 164200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8857
timestamp 1654712443
transform 1 0 167200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8957
timestamp 1654712443
transform 1 0 167200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8858
timestamp 1654712443
transform 1 0 170200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8958
timestamp 1654712443
transform 1 0 170200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8859
timestamp 1654712443
transform 1 0 173200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8959
timestamp 1654712443
transform 1 0 173200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8860
timestamp 1654712443
transform 1 0 176200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8960
timestamp 1654712443
transform 1 0 176200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8861
timestamp 1654712443
transform 1 0 179200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8961
timestamp 1654712443
transform 1 0 179200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8863
timestamp 1654712443
transform 1 0 185200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8862
timestamp 1654712443
transform 1 0 182200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8963
timestamp 1654712443
transform 1 0 185200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8962
timestamp 1654712443
transform 1 0 182200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8864
timestamp 1654712443
transform 1 0 188200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8964
timestamp 1654712443
transform 1 0 188200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8865
timestamp 1654712443
transform 1 0 191200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8965
timestamp 1654712443
transform 1 0 191200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8866
timestamp 1654712443
transform 1 0 194200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8966
timestamp 1654712443
transform 1 0 194200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8867
timestamp 1654712443
transform 1 0 197200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8967
timestamp 1654712443
transform 1 0 197200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8868
timestamp 1654712443
transform 1 0 200200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8968
timestamp 1654712443
transform 1 0 200200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8869
timestamp 1654712443
transform 1 0 203200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8969
timestamp 1654712443
transform 1 0 203200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8870
timestamp 1654712443
transform 1 0 206200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8970
timestamp 1654712443
transform 1 0 206200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8871
timestamp 1654712443
transform 1 0 209200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8971
timestamp 1654712443
transform 1 0 209200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8873
timestamp 1654712443
transform 1 0 215200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8872
timestamp 1654712443
transform 1 0 212200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8973
timestamp 1654712443
transform 1 0 215200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8972
timestamp 1654712443
transform 1 0 212200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8874
timestamp 1654712443
transform 1 0 218200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8974
timestamp 1654712443
transform 1 0 218200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8875
timestamp 1654712443
transform 1 0 221200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8975
timestamp 1654712443
transform 1 0 221200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8876
timestamp 1654712443
transform 1 0 224200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8976
timestamp 1654712443
transform 1 0 224200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8877
timestamp 1654712443
transform 1 0 227200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8977
timestamp 1654712443
transform 1 0 227200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8878
timestamp 1654712443
transform 1 0 230200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8978
timestamp 1654712443
transform 1 0 230200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8879
timestamp 1654712443
transform 1 0 233200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8979
timestamp 1654712443
transform 1 0 233200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8880
timestamp 1654712443
transform 1 0 236200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8980
timestamp 1654712443
transform 1 0 236200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8881
timestamp 1654712443
transform 1 0 239200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8981
timestamp 1654712443
transform 1 0 239200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8883
timestamp 1654712443
transform 1 0 245200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8882
timestamp 1654712443
transform 1 0 242200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8983
timestamp 1654712443
transform 1 0 245200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8982
timestamp 1654712443
transform 1 0 242200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8884
timestamp 1654712443
transform 1 0 248200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8984
timestamp 1654712443
transform 1 0 248200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8885
timestamp 1654712443
transform 1 0 251200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8985
timestamp 1654712443
transform 1 0 251200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8886
timestamp 1654712443
transform 1 0 254200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8986
timestamp 1654712443
transform 1 0 254200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8887
timestamp 1654712443
transform 1 0 257200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8987
timestamp 1654712443
transform 1 0 257200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8888
timestamp 1654712443
transform 1 0 260200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8988
timestamp 1654712443
transform 1 0 260200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8889
timestamp 1654712443
transform 1 0 263200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8989
timestamp 1654712443
transform 1 0 263200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8890
timestamp 1654712443
transform 1 0 266200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8990
timestamp 1654712443
transform 1 0 266200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8891
timestamp 1654712443
transform 1 0 269200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8991
timestamp 1654712443
transform 1 0 269200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8892
timestamp 1654712443
transform 1 0 272200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8992
timestamp 1654712443
transform 1 0 272200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8894
timestamp 1654712443
transform 1 0 278200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8893
timestamp 1654712443
transform 1 0 275200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8994
timestamp 1654712443
transform 1 0 278200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8993
timestamp 1654712443
transform 1 0 275200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8895
timestamp 1654712443
transform 1 0 281200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8995
timestamp 1654712443
transform 1 0 281200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8896
timestamp 1654712443
transform 1 0 284200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8996
timestamp 1654712443
transform 1 0 284200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8897
timestamp 1654712443
transform 1 0 287200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8997
timestamp 1654712443
transform 1 0 287200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8898
timestamp 1654712443
transform 1 0 290200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8998
timestamp 1654712443
transform 1 0 290200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8899
timestamp 1654712443
transform 1 0 293200 0 1 -261300
box 3640 -2860 6960 460
use pixel  pixel_8999
timestamp 1654712443
transform 1 0 293200 0 1 -264300
box 3640 -2860 6960 460
use pixel  pixel_8701
timestamp 1654712443
transform 1 0 -800 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8700
timestamp 1654712443
transform 1 0 -3800 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8702
timestamp 1654712443
transform 1 0 2200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8703
timestamp 1654712443
transform 1 0 5200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8704
timestamp 1654712443
transform 1 0 8200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8705
timestamp 1654712443
transform 1 0 11200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8706
timestamp 1654712443
transform 1 0 14200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8707
timestamp 1654712443
transform 1 0 17200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8708
timestamp 1654712443
transform 1 0 20200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8709
timestamp 1654712443
transform 1 0 23200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8711
timestamp 1654712443
transform 1 0 29200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8710
timestamp 1654712443
transform 1 0 26200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8712
timestamp 1654712443
transform 1 0 32200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8713
timestamp 1654712443
transform 1 0 35200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8714
timestamp 1654712443
transform 1 0 38200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8715
timestamp 1654712443
transform 1 0 41200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8716
timestamp 1654712443
transform 1 0 44200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8717
timestamp 1654712443
transform 1 0 47200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8718
timestamp 1654712443
transform 1 0 50200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8719
timestamp 1654712443
transform 1 0 53200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8721
timestamp 1654712443
transform 1 0 59200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8720
timestamp 1654712443
transform 1 0 56200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8722
timestamp 1654712443
transform 1 0 62200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8723
timestamp 1654712443
transform 1 0 65200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8724
timestamp 1654712443
transform 1 0 68200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8725
timestamp 1654712443
transform 1 0 71200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8726
timestamp 1654712443
transform 1 0 74200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8727
timestamp 1654712443
transform 1 0 77200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8728
timestamp 1654712443
transform 1 0 80200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8729
timestamp 1654712443
transform 1 0 83200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8730
timestamp 1654712443
transform 1 0 86200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8731
timestamp 1654712443
transform 1 0 89200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8732
timestamp 1654712443
transform 1 0 92200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8733
timestamp 1654712443
transform 1 0 95200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8734
timestamp 1654712443
transform 1 0 98200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8735
timestamp 1654712443
transform 1 0 101200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8736
timestamp 1654712443
transform 1 0 104200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8737
timestamp 1654712443
transform 1 0 107200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8738
timestamp 1654712443
transform 1 0 110200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8739
timestamp 1654712443
transform 1 0 113200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8740
timestamp 1654712443
transform 1 0 116200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8741
timestamp 1654712443
transform 1 0 119200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8742
timestamp 1654712443
transform 1 0 122200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8743
timestamp 1654712443
transform 1 0 125200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8744
timestamp 1654712443
transform 1 0 128200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8745
timestamp 1654712443
transform 1 0 131200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8746
timestamp 1654712443
transform 1 0 134200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8747
timestamp 1654712443
transform 1 0 137200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8748
timestamp 1654712443
transform 1 0 140200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8749
timestamp 1654712443
transform 1 0 143200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8750
timestamp 1654712443
transform 1 0 146200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8751
timestamp 1654712443
transform 1 0 149200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8752
timestamp 1654712443
transform 1 0 152200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8753
timestamp 1654712443
transform 1 0 155200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8754
timestamp 1654712443
transform 1 0 158200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8755
timestamp 1654712443
transform 1 0 161200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8756
timestamp 1654712443
transform 1 0 164200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8757
timestamp 1654712443
transform 1 0 167200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8758
timestamp 1654712443
transform 1 0 170200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8759
timestamp 1654712443
transform 1 0 173200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8760
timestamp 1654712443
transform 1 0 176200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8761
timestamp 1654712443
transform 1 0 179200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8763
timestamp 1654712443
transform 1 0 185200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8762
timestamp 1654712443
transform 1 0 182200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8764
timestamp 1654712443
transform 1 0 188200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8765
timestamp 1654712443
transform 1 0 191200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8766
timestamp 1654712443
transform 1 0 194200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8767
timestamp 1654712443
transform 1 0 197200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8768
timestamp 1654712443
transform 1 0 200200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8769
timestamp 1654712443
transform 1 0 203200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8770
timestamp 1654712443
transform 1 0 206200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8771
timestamp 1654712443
transform 1 0 209200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8773
timestamp 1654712443
transform 1 0 215200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8772
timestamp 1654712443
transform 1 0 212200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8774
timestamp 1654712443
transform 1 0 218200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8775
timestamp 1654712443
transform 1 0 221200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8776
timestamp 1654712443
transform 1 0 224200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8777
timestamp 1654712443
transform 1 0 227200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8778
timestamp 1654712443
transform 1 0 230200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8779
timestamp 1654712443
transform 1 0 233200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8780
timestamp 1654712443
transform 1 0 236200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8781
timestamp 1654712443
transform 1 0 239200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8783
timestamp 1654712443
transform 1 0 245200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8782
timestamp 1654712443
transform 1 0 242200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8784
timestamp 1654712443
transform 1 0 248200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8785
timestamp 1654712443
transform 1 0 251200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8786
timestamp 1654712443
transform 1 0 254200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8787
timestamp 1654712443
transform 1 0 257200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8788
timestamp 1654712443
transform 1 0 260200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8789
timestamp 1654712443
transform 1 0 263200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8790
timestamp 1654712443
transform 1 0 266200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8791
timestamp 1654712443
transform 1 0 269200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8792
timestamp 1654712443
transform 1 0 272200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8794
timestamp 1654712443
transform 1 0 278200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8793
timestamp 1654712443
transform 1 0 275200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8795
timestamp 1654712443
transform 1 0 281200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8796
timestamp 1654712443
transform 1 0 284200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8797
timestamp 1654712443
transform 1 0 287200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8798
timestamp 1654712443
transform 1 0 290200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8799
timestamp 1654712443
transform 1 0 293200 0 1 -258300
box 3640 -2860 6960 460
use pixel  pixel_8601
timestamp 1654712443
transform 1 0 -800 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8600
timestamp 1654712443
transform 1 0 -3800 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8602
timestamp 1654712443
transform 1 0 2200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8603
timestamp 1654712443
transform 1 0 5200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8604
timestamp 1654712443
transform 1 0 8200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8605
timestamp 1654712443
transform 1 0 11200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8606
timestamp 1654712443
transform 1 0 14200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8607
timestamp 1654712443
transform 1 0 17200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8608
timestamp 1654712443
transform 1 0 20200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8609
timestamp 1654712443
transform 1 0 23200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8611
timestamp 1654712443
transform 1 0 29200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8610
timestamp 1654712443
transform 1 0 26200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8612
timestamp 1654712443
transform 1 0 32200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8613
timestamp 1654712443
transform 1 0 35200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8614
timestamp 1654712443
transform 1 0 38200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8615
timestamp 1654712443
transform 1 0 41200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8616
timestamp 1654712443
transform 1 0 44200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8617
timestamp 1654712443
transform 1 0 47200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8618
timestamp 1654712443
transform 1 0 50200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8619
timestamp 1654712443
transform 1 0 53200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8621
timestamp 1654712443
transform 1 0 59200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8620
timestamp 1654712443
transform 1 0 56200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8622
timestamp 1654712443
transform 1 0 62200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8623
timestamp 1654712443
transform 1 0 65200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8624
timestamp 1654712443
transform 1 0 68200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8625
timestamp 1654712443
transform 1 0 71200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8626
timestamp 1654712443
transform 1 0 74200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8627
timestamp 1654712443
transform 1 0 77200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8628
timestamp 1654712443
transform 1 0 80200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8629
timestamp 1654712443
transform 1 0 83200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8630
timestamp 1654712443
transform 1 0 86200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8631
timestamp 1654712443
transform 1 0 89200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8632
timestamp 1654712443
transform 1 0 92200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8633
timestamp 1654712443
transform 1 0 95200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8634
timestamp 1654712443
transform 1 0 98200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8635
timestamp 1654712443
transform 1 0 101200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8636
timestamp 1654712443
transform 1 0 104200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8637
timestamp 1654712443
transform 1 0 107200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8638
timestamp 1654712443
transform 1 0 110200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8639
timestamp 1654712443
transform 1 0 113200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8640
timestamp 1654712443
transform 1 0 116200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8641
timestamp 1654712443
transform 1 0 119200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8642
timestamp 1654712443
transform 1 0 122200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8643
timestamp 1654712443
transform 1 0 125200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8644
timestamp 1654712443
transform 1 0 128200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8645
timestamp 1654712443
transform 1 0 131200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8646
timestamp 1654712443
transform 1 0 134200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8647
timestamp 1654712443
transform 1 0 137200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8648
timestamp 1654712443
transform 1 0 140200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8649
timestamp 1654712443
transform 1 0 143200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8650
timestamp 1654712443
transform 1 0 146200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8651
timestamp 1654712443
transform 1 0 149200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8652
timestamp 1654712443
transform 1 0 152200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8653
timestamp 1654712443
transform 1 0 155200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8654
timestamp 1654712443
transform 1 0 158200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8655
timestamp 1654712443
transform 1 0 161200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8656
timestamp 1654712443
transform 1 0 164200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8657
timestamp 1654712443
transform 1 0 167200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8658
timestamp 1654712443
transform 1 0 170200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8659
timestamp 1654712443
transform 1 0 173200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8660
timestamp 1654712443
transform 1 0 176200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8661
timestamp 1654712443
transform 1 0 179200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8663
timestamp 1654712443
transform 1 0 185200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8662
timestamp 1654712443
transform 1 0 182200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8664
timestamp 1654712443
transform 1 0 188200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8665
timestamp 1654712443
transform 1 0 191200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8666
timestamp 1654712443
transform 1 0 194200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8667
timestamp 1654712443
transform 1 0 197200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8668
timestamp 1654712443
transform 1 0 200200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8669
timestamp 1654712443
transform 1 0 203200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8670
timestamp 1654712443
transform 1 0 206200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8671
timestamp 1654712443
transform 1 0 209200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8673
timestamp 1654712443
transform 1 0 215200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8672
timestamp 1654712443
transform 1 0 212200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8674
timestamp 1654712443
transform 1 0 218200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8675
timestamp 1654712443
transform 1 0 221200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8676
timestamp 1654712443
transform 1 0 224200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8677
timestamp 1654712443
transform 1 0 227200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8678
timestamp 1654712443
transform 1 0 230200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8679
timestamp 1654712443
transform 1 0 233200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8680
timestamp 1654712443
transform 1 0 236200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8681
timestamp 1654712443
transform 1 0 239200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8683
timestamp 1654712443
transform 1 0 245200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8682
timestamp 1654712443
transform 1 0 242200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8684
timestamp 1654712443
transform 1 0 248200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8685
timestamp 1654712443
transform 1 0 251200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8686
timestamp 1654712443
transform 1 0 254200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8687
timestamp 1654712443
transform 1 0 257200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8688
timestamp 1654712443
transform 1 0 260200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8689
timestamp 1654712443
transform 1 0 263200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8690
timestamp 1654712443
transform 1 0 266200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8691
timestamp 1654712443
transform 1 0 269200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8692
timestamp 1654712443
transform 1 0 272200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8694
timestamp 1654712443
transform 1 0 278200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8693
timestamp 1654712443
transform 1 0 275200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8695
timestamp 1654712443
transform 1 0 281200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8696
timestamp 1654712443
transform 1 0 284200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8697
timestamp 1654712443
transform 1 0 287200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8698
timestamp 1654712443
transform 1 0 290200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8699
timestamp 1654712443
transform 1 0 293200 0 1 -255300
box 3640 -2860 6960 460
use pixel  pixel_8501
timestamp 1654712443
transform 1 0 -800 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8500
timestamp 1654712443
transform 1 0 -3800 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8502
timestamp 1654712443
transform 1 0 2200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8503
timestamp 1654712443
transform 1 0 5200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8504
timestamp 1654712443
transform 1 0 8200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8505
timestamp 1654712443
transform 1 0 11200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8506
timestamp 1654712443
transform 1 0 14200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8507
timestamp 1654712443
transform 1 0 17200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8508
timestamp 1654712443
transform 1 0 20200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8509
timestamp 1654712443
transform 1 0 23200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8511
timestamp 1654712443
transform 1 0 29200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8510
timestamp 1654712443
transform 1 0 26200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8512
timestamp 1654712443
transform 1 0 32200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8513
timestamp 1654712443
transform 1 0 35200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8514
timestamp 1654712443
transform 1 0 38200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8515
timestamp 1654712443
transform 1 0 41200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8516
timestamp 1654712443
transform 1 0 44200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8517
timestamp 1654712443
transform 1 0 47200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8518
timestamp 1654712443
transform 1 0 50200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8519
timestamp 1654712443
transform 1 0 53200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8521
timestamp 1654712443
transform 1 0 59200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8520
timestamp 1654712443
transform 1 0 56200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8522
timestamp 1654712443
transform 1 0 62200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8523
timestamp 1654712443
transform 1 0 65200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8524
timestamp 1654712443
transform 1 0 68200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8525
timestamp 1654712443
transform 1 0 71200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8526
timestamp 1654712443
transform 1 0 74200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8527
timestamp 1654712443
transform 1 0 77200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8528
timestamp 1654712443
transform 1 0 80200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8529
timestamp 1654712443
transform 1 0 83200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8530
timestamp 1654712443
transform 1 0 86200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8531
timestamp 1654712443
transform 1 0 89200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8532
timestamp 1654712443
transform 1 0 92200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8533
timestamp 1654712443
transform 1 0 95200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8534
timestamp 1654712443
transform 1 0 98200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8535
timestamp 1654712443
transform 1 0 101200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8536
timestamp 1654712443
transform 1 0 104200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8537
timestamp 1654712443
transform 1 0 107200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8538
timestamp 1654712443
transform 1 0 110200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8539
timestamp 1654712443
transform 1 0 113200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8540
timestamp 1654712443
transform 1 0 116200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8541
timestamp 1654712443
transform 1 0 119200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8542
timestamp 1654712443
transform 1 0 122200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8543
timestamp 1654712443
transform 1 0 125200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8544
timestamp 1654712443
transform 1 0 128200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8545
timestamp 1654712443
transform 1 0 131200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8546
timestamp 1654712443
transform 1 0 134200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8547
timestamp 1654712443
transform 1 0 137200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8548
timestamp 1654712443
transform 1 0 140200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8549
timestamp 1654712443
transform 1 0 143200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8550
timestamp 1654712443
transform 1 0 146200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8551
timestamp 1654712443
transform 1 0 149200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8552
timestamp 1654712443
transform 1 0 152200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8553
timestamp 1654712443
transform 1 0 155200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8554
timestamp 1654712443
transform 1 0 158200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8555
timestamp 1654712443
transform 1 0 161200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8556
timestamp 1654712443
transform 1 0 164200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8557
timestamp 1654712443
transform 1 0 167200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8558
timestamp 1654712443
transform 1 0 170200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8559
timestamp 1654712443
transform 1 0 173200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8560
timestamp 1654712443
transform 1 0 176200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8561
timestamp 1654712443
transform 1 0 179200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8563
timestamp 1654712443
transform 1 0 185200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8562
timestamp 1654712443
transform 1 0 182200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8564
timestamp 1654712443
transform 1 0 188200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8565
timestamp 1654712443
transform 1 0 191200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8566
timestamp 1654712443
transform 1 0 194200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8567
timestamp 1654712443
transform 1 0 197200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8568
timestamp 1654712443
transform 1 0 200200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8569
timestamp 1654712443
transform 1 0 203200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8570
timestamp 1654712443
transform 1 0 206200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8571
timestamp 1654712443
transform 1 0 209200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8573
timestamp 1654712443
transform 1 0 215200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8572
timestamp 1654712443
transform 1 0 212200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8574
timestamp 1654712443
transform 1 0 218200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8575
timestamp 1654712443
transform 1 0 221200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8576
timestamp 1654712443
transform 1 0 224200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8577
timestamp 1654712443
transform 1 0 227200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8578
timestamp 1654712443
transform 1 0 230200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8579
timestamp 1654712443
transform 1 0 233200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8580
timestamp 1654712443
transform 1 0 236200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8581
timestamp 1654712443
transform 1 0 239200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8583
timestamp 1654712443
transform 1 0 245200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8582
timestamp 1654712443
transform 1 0 242200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8584
timestamp 1654712443
transform 1 0 248200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8585
timestamp 1654712443
transform 1 0 251200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8586
timestamp 1654712443
transform 1 0 254200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8587
timestamp 1654712443
transform 1 0 257200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8588
timestamp 1654712443
transform 1 0 260200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8589
timestamp 1654712443
transform 1 0 263200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8590
timestamp 1654712443
transform 1 0 266200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8591
timestamp 1654712443
transform 1 0 269200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8592
timestamp 1654712443
transform 1 0 272200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8594
timestamp 1654712443
transform 1 0 278200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8593
timestamp 1654712443
transform 1 0 275200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8595
timestamp 1654712443
transform 1 0 281200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8596
timestamp 1654712443
transform 1 0 284200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8597
timestamp 1654712443
transform 1 0 287200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8598
timestamp 1654712443
transform 1 0 290200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8599
timestamp 1654712443
transform 1 0 293200 0 1 -252300
box 3640 -2860 6960 460
use pixel  pixel_8401
timestamp 1654712443
transform 1 0 -800 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8400
timestamp 1654712443
transform 1 0 -3800 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8402
timestamp 1654712443
transform 1 0 2200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8403
timestamp 1654712443
transform 1 0 5200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8404
timestamp 1654712443
transform 1 0 8200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8405
timestamp 1654712443
transform 1 0 11200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8406
timestamp 1654712443
transform 1 0 14200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8407
timestamp 1654712443
transform 1 0 17200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8408
timestamp 1654712443
transform 1 0 20200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8409
timestamp 1654712443
transform 1 0 23200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8411
timestamp 1654712443
transform 1 0 29200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8410
timestamp 1654712443
transform 1 0 26200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8412
timestamp 1654712443
transform 1 0 32200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8413
timestamp 1654712443
transform 1 0 35200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8414
timestamp 1654712443
transform 1 0 38200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8415
timestamp 1654712443
transform 1 0 41200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8416
timestamp 1654712443
transform 1 0 44200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8417
timestamp 1654712443
transform 1 0 47200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8418
timestamp 1654712443
transform 1 0 50200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8419
timestamp 1654712443
transform 1 0 53200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8421
timestamp 1654712443
transform 1 0 59200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8420
timestamp 1654712443
transform 1 0 56200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8422
timestamp 1654712443
transform 1 0 62200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8423
timestamp 1654712443
transform 1 0 65200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8424
timestamp 1654712443
transform 1 0 68200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8425
timestamp 1654712443
transform 1 0 71200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8426
timestamp 1654712443
transform 1 0 74200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8427
timestamp 1654712443
transform 1 0 77200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8428
timestamp 1654712443
transform 1 0 80200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8429
timestamp 1654712443
transform 1 0 83200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8430
timestamp 1654712443
transform 1 0 86200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8431
timestamp 1654712443
transform 1 0 89200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8432
timestamp 1654712443
transform 1 0 92200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8433
timestamp 1654712443
transform 1 0 95200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8434
timestamp 1654712443
transform 1 0 98200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8435
timestamp 1654712443
transform 1 0 101200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8436
timestamp 1654712443
transform 1 0 104200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8437
timestamp 1654712443
transform 1 0 107200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8438
timestamp 1654712443
transform 1 0 110200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8439
timestamp 1654712443
transform 1 0 113200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8440
timestamp 1654712443
transform 1 0 116200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8441
timestamp 1654712443
transform 1 0 119200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8442
timestamp 1654712443
transform 1 0 122200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8443
timestamp 1654712443
transform 1 0 125200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8444
timestamp 1654712443
transform 1 0 128200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8445
timestamp 1654712443
transform 1 0 131200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8446
timestamp 1654712443
transform 1 0 134200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8447
timestamp 1654712443
transform 1 0 137200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8448
timestamp 1654712443
transform 1 0 140200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8449
timestamp 1654712443
transform 1 0 143200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8450
timestamp 1654712443
transform 1 0 146200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8451
timestamp 1654712443
transform 1 0 149200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8452
timestamp 1654712443
transform 1 0 152200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8453
timestamp 1654712443
transform 1 0 155200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8454
timestamp 1654712443
transform 1 0 158200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8455
timestamp 1654712443
transform 1 0 161200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8456
timestamp 1654712443
transform 1 0 164200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8457
timestamp 1654712443
transform 1 0 167200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8458
timestamp 1654712443
transform 1 0 170200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8459
timestamp 1654712443
transform 1 0 173200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8460
timestamp 1654712443
transform 1 0 176200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8461
timestamp 1654712443
transform 1 0 179200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8463
timestamp 1654712443
transform 1 0 185200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8462
timestamp 1654712443
transform 1 0 182200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8464
timestamp 1654712443
transform 1 0 188200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8465
timestamp 1654712443
transform 1 0 191200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8466
timestamp 1654712443
transform 1 0 194200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8467
timestamp 1654712443
transform 1 0 197200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8468
timestamp 1654712443
transform 1 0 200200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8469
timestamp 1654712443
transform 1 0 203200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8470
timestamp 1654712443
transform 1 0 206200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8471
timestamp 1654712443
transform 1 0 209200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8473
timestamp 1654712443
transform 1 0 215200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8472
timestamp 1654712443
transform 1 0 212200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8474
timestamp 1654712443
transform 1 0 218200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8475
timestamp 1654712443
transform 1 0 221200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8476
timestamp 1654712443
transform 1 0 224200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8477
timestamp 1654712443
transform 1 0 227200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8478
timestamp 1654712443
transform 1 0 230200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8479
timestamp 1654712443
transform 1 0 233200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8480
timestamp 1654712443
transform 1 0 236200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8481
timestamp 1654712443
transform 1 0 239200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8483
timestamp 1654712443
transform 1 0 245200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8482
timestamp 1654712443
transform 1 0 242200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8484
timestamp 1654712443
transform 1 0 248200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8485
timestamp 1654712443
transform 1 0 251200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8486
timestamp 1654712443
transform 1 0 254200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8487
timestamp 1654712443
transform 1 0 257200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8488
timestamp 1654712443
transform 1 0 260200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8489
timestamp 1654712443
transform 1 0 263200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8490
timestamp 1654712443
transform 1 0 266200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8491
timestamp 1654712443
transform 1 0 269200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8492
timestamp 1654712443
transform 1 0 272200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8494
timestamp 1654712443
transform 1 0 278200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8493
timestamp 1654712443
transform 1 0 275200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8495
timestamp 1654712443
transform 1 0 281200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8496
timestamp 1654712443
transform 1 0 284200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8497
timestamp 1654712443
transform 1 0 287200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8498
timestamp 1654712443
transform 1 0 290200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8499
timestamp 1654712443
transform 1 0 293200 0 1 -249300
box 3640 -2860 6960 460
use pixel  pixel_8301
timestamp 1654712443
transform 1 0 -800 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8300
timestamp 1654712443
transform 1 0 -3800 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8302
timestamp 1654712443
transform 1 0 2200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8303
timestamp 1654712443
transform 1 0 5200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8304
timestamp 1654712443
transform 1 0 8200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8305
timestamp 1654712443
transform 1 0 11200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8306
timestamp 1654712443
transform 1 0 14200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8307
timestamp 1654712443
transform 1 0 17200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8308
timestamp 1654712443
transform 1 0 20200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8309
timestamp 1654712443
transform 1 0 23200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8311
timestamp 1654712443
transform 1 0 29200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8310
timestamp 1654712443
transform 1 0 26200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8312
timestamp 1654712443
transform 1 0 32200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8313
timestamp 1654712443
transform 1 0 35200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8314
timestamp 1654712443
transform 1 0 38200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8315
timestamp 1654712443
transform 1 0 41200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8316
timestamp 1654712443
transform 1 0 44200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8317
timestamp 1654712443
transform 1 0 47200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8318
timestamp 1654712443
transform 1 0 50200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8319
timestamp 1654712443
transform 1 0 53200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8321
timestamp 1654712443
transform 1 0 59200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8320
timestamp 1654712443
transform 1 0 56200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8322
timestamp 1654712443
transform 1 0 62200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8323
timestamp 1654712443
transform 1 0 65200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8324
timestamp 1654712443
transform 1 0 68200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8325
timestamp 1654712443
transform 1 0 71200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8326
timestamp 1654712443
transform 1 0 74200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8327
timestamp 1654712443
transform 1 0 77200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8328
timestamp 1654712443
transform 1 0 80200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8329
timestamp 1654712443
transform 1 0 83200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8330
timestamp 1654712443
transform 1 0 86200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8331
timestamp 1654712443
transform 1 0 89200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8332
timestamp 1654712443
transform 1 0 92200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8333
timestamp 1654712443
transform 1 0 95200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8334
timestamp 1654712443
transform 1 0 98200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8335
timestamp 1654712443
transform 1 0 101200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8336
timestamp 1654712443
transform 1 0 104200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8337
timestamp 1654712443
transform 1 0 107200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8338
timestamp 1654712443
transform 1 0 110200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8339
timestamp 1654712443
transform 1 0 113200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8340
timestamp 1654712443
transform 1 0 116200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8341
timestamp 1654712443
transform 1 0 119200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8342
timestamp 1654712443
transform 1 0 122200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8343
timestamp 1654712443
transform 1 0 125200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8344
timestamp 1654712443
transform 1 0 128200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8345
timestamp 1654712443
transform 1 0 131200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8346
timestamp 1654712443
transform 1 0 134200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8347
timestamp 1654712443
transform 1 0 137200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8348
timestamp 1654712443
transform 1 0 140200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8349
timestamp 1654712443
transform 1 0 143200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8350
timestamp 1654712443
transform 1 0 146200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8351
timestamp 1654712443
transform 1 0 149200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8352
timestamp 1654712443
transform 1 0 152200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8353
timestamp 1654712443
transform 1 0 155200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8354
timestamp 1654712443
transform 1 0 158200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8355
timestamp 1654712443
transform 1 0 161200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8356
timestamp 1654712443
transform 1 0 164200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8357
timestamp 1654712443
transform 1 0 167200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8358
timestamp 1654712443
transform 1 0 170200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8359
timestamp 1654712443
transform 1 0 173200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8360
timestamp 1654712443
transform 1 0 176200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8361
timestamp 1654712443
transform 1 0 179200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8363
timestamp 1654712443
transform 1 0 185200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8362
timestamp 1654712443
transform 1 0 182200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8364
timestamp 1654712443
transform 1 0 188200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8365
timestamp 1654712443
transform 1 0 191200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8366
timestamp 1654712443
transform 1 0 194200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8367
timestamp 1654712443
transform 1 0 197200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8368
timestamp 1654712443
transform 1 0 200200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8369
timestamp 1654712443
transform 1 0 203200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8370
timestamp 1654712443
transform 1 0 206200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8371
timestamp 1654712443
transform 1 0 209200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8373
timestamp 1654712443
transform 1 0 215200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8372
timestamp 1654712443
transform 1 0 212200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8374
timestamp 1654712443
transform 1 0 218200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8375
timestamp 1654712443
transform 1 0 221200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8376
timestamp 1654712443
transform 1 0 224200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8377
timestamp 1654712443
transform 1 0 227200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8378
timestamp 1654712443
transform 1 0 230200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8379
timestamp 1654712443
transform 1 0 233200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8380
timestamp 1654712443
transform 1 0 236200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8381
timestamp 1654712443
transform 1 0 239200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8383
timestamp 1654712443
transform 1 0 245200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8382
timestamp 1654712443
transform 1 0 242200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8384
timestamp 1654712443
transform 1 0 248200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8385
timestamp 1654712443
transform 1 0 251200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8386
timestamp 1654712443
transform 1 0 254200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8387
timestamp 1654712443
transform 1 0 257200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8388
timestamp 1654712443
transform 1 0 260200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8389
timestamp 1654712443
transform 1 0 263200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8390
timestamp 1654712443
transform 1 0 266200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8391
timestamp 1654712443
transform 1 0 269200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8392
timestamp 1654712443
transform 1 0 272200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8394
timestamp 1654712443
transform 1 0 278200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8393
timestamp 1654712443
transform 1 0 275200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8395
timestamp 1654712443
transform 1 0 281200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8396
timestamp 1654712443
transform 1 0 284200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8397
timestamp 1654712443
transform 1 0 287200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8398
timestamp 1654712443
transform 1 0 290200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8399
timestamp 1654712443
transform 1 0 293200 0 1 -246300
box 3640 -2860 6960 460
use pixel  pixel_8201
timestamp 1654712443
transform 1 0 -800 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8200
timestamp 1654712443
transform 1 0 -3800 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8202
timestamp 1654712443
transform 1 0 2200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8203
timestamp 1654712443
transform 1 0 5200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8204
timestamp 1654712443
transform 1 0 8200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8205
timestamp 1654712443
transform 1 0 11200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8206
timestamp 1654712443
transform 1 0 14200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8207
timestamp 1654712443
transform 1 0 17200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8208
timestamp 1654712443
transform 1 0 20200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8209
timestamp 1654712443
transform 1 0 23200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8211
timestamp 1654712443
transform 1 0 29200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8210
timestamp 1654712443
transform 1 0 26200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8212
timestamp 1654712443
transform 1 0 32200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8213
timestamp 1654712443
transform 1 0 35200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8214
timestamp 1654712443
transform 1 0 38200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8215
timestamp 1654712443
transform 1 0 41200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8216
timestamp 1654712443
transform 1 0 44200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8217
timestamp 1654712443
transform 1 0 47200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8218
timestamp 1654712443
transform 1 0 50200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8219
timestamp 1654712443
transform 1 0 53200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8221
timestamp 1654712443
transform 1 0 59200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8220
timestamp 1654712443
transform 1 0 56200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8222
timestamp 1654712443
transform 1 0 62200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8223
timestamp 1654712443
transform 1 0 65200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8224
timestamp 1654712443
transform 1 0 68200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8225
timestamp 1654712443
transform 1 0 71200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8226
timestamp 1654712443
transform 1 0 74200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8227
timestamp 1654712443
transform 1 0 77200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8228
timestamp 1654712443
transform 1 0 80200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8229
timestamp 1654712443
transform 1 0 83200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8230
timestamp 1654712443
transform 1 0 86200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8231
timestamp 1654712443
transform 1 0 89200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8232
timestamp 1654712443
transform 1 0 92200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8233
timestamp 1654712443
transform 1 0 95200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8234
timestamp 1654712443
transform 1 0 98200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8235
timestamp 1654712443
transform 1 0 101200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8236
timestamp 1654712443
transform 1 0 104200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8237
timestamp 1654712443
transform 1 0 107200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8238
timestamp 1654712443
transform 1 0 110200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8239
timestamp 1654712443
transform 1 0 113200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8240
timestamp 1654712443
transform 1 0 116200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8241
timestamp 1654712443
transform 1 0 119200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8242
timestamp 1654712443
transform 1 0 122200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8243
timestamp 1654712443
transform 1 0 125200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8244
timestamp 1654712443
transform 1 0 128200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8245
timestamp 1654712443
transform 1 0 131200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8246
timestamp 1654712443
transform 1 0 134200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8247
timestamp 1654712443
transform 1 0 137200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8248
timestamp 1654712443
transform 1 0 140200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8249
timestamp 1654712443
transform 1 0 143200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8250
timestamp 1654712443
transform 1 0 146200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8251
timestamp 1654712443
transform 1 0 149200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8252
timestamp 1654712443
transform 1 0 152200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8253
timestamp 1654712443
transform 1 0 155200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8254
timestamp 1654712443
transform 1 0 158200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8255
timestamp 1654712443
transform 1 0 161200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8256
timestamp 1654712443
transform 1 0 164200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8257
timestamp 1654712443
transform 1 0 167200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8258
timestamp 1654712443
transform 1 0 170200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8259
timestamp 1654712443
transform 1 0 173200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8260
timestamp 1654712443
transform 1 0 176200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8261
timestamp 1654712443
transform 1 0 179200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8263
timestamp 1654712443
transform 1 0 185200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8262
timestamp 1654712443
transform 1 0 182200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8264
timestamp 1654712443
transform 1 0 188200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8265
timestamp 1654712443
transform 1 0 191200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8266
timestamp 1654712443
transform 1 0 194200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8267
timestamp 1654712443
transform 1 0 197200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8268
timestamp 1654712443
transform 1 0 200200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8269
timestamp 1654712443
transform 1 0 203200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8270
timestamp 1654712443
transform 1 0 206200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8271
timestamp 1654712443
transform 1 0 209200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8273
timestamp 1654712443
transform 1 0 215200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8272
timestamp 1654712443
transform 1 0 212200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8274
timestamp 1654712443
transform 1 0 218200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8275
timestamp 1654712443
transform 1 0 221200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8276
timestamp 1654712443
transform 1 0 224200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8277
timestamp 1654712443
transform 1 0 227200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8278
timestamp 1654712443
transform 1 0 230200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8279
timestamp 1654712443
transform 1 0 233200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8280
timestamp 1654712443
transform 1 0 236200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8281
timestamp 1654712443
transform 1 0 239200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8283
timestamp 1654712443
transform 1 0 245200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8282
timestamp 1654712443
transform 1 0 242200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8284
timestamp 1654712443
transform 1 0 248200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8285
timestamp 1654712443
transform 1 0 251200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8286
timestamp 1654712443
transform 1 0 254200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8287
timestamp 1654712443
transform 1 0 257200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8288
timestamp 1654712443
transform 1 0 260200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8289
timestamp 1654712443
transform 1 0 263200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8290
timestamp 1654712443
transform 1 0 266200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8291
timestamp 1654712443
transform 1 0 269200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8292
timestamp 1654712443
transform 1 0 272200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8294
timestamp 1654712443
transform 1 0 278200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8293
timestamp 1654712443
transform 1 0 275200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8295
timestamp 1654712443
transform 1 0 281200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8296
timestamp 1654712443
transform 1 0 284200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8297
timestamp 1654712443
transform 1 0 287200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8298
timestamp 1654712443
transform 1 0 290200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8299
timestamp 1654712443
transform 1 0 293200 0 1 -243300
box 3640 -2860 6960 460
use pixel  pixel_8101
timestamp 1654712443
transform 1 0 -800 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8100
timestamp 1654712443
transform 1 0 -3800 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8102
timestamp 1654712443
transform 1 0 2200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8103
timestamp 1654712443
transform 1 0 5200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8104
timestamp 1654712443
transform 1 0 8200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8105
timestamp 1654712443
transform 1 0 11200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8106
timestamp 1654712443
transform 1 0 14200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8107
timestamp 1654712443
transform 1 0 17200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8108
timestamp 1654712443
transform 1 0 20200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8109
timestamp 1654712443
transform 1 0 23200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8111
timestamp 1654712443
transform 1 0 29200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8110
timestamp 1654712443
transform 1 0 26200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8112
timestamp 1654712443
transform 1 0 32200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8113
timestamp 1654712443
transform 1 0 35200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8114
timestamp 1654712443
transform 1 0 38200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8115
timestamp 1654712443
transform 1 0 41200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8116
timestamp 1654712443
transform 1 0 44200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8117
timestamp 1654712443
transform 1 0 47200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8118
timestamp 1654712443
transform 1 0 50200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8119
timestamp 1654712443
transform 1 0 53200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8121
timestamp 1654712443
transform 1 0 59200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8120
timestamp 1654712443
transform 1 0 56200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8122
timestamp 1654712443
transform 1 0 62200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8123
timestamp 1654712443
transform 1 0 65200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8124
timestamp 1654712443
transform 1 0 68200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8125
timestamp 1654712443
transform 1 0 71200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8126
timestamp 1654712443
transform 1 0 74200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8127
timestamp 1654712443
transform 1 0 77200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8128
timestamp 1654712443
transform 1 0 80200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8129
timestamp 1654712443
transform 1 0 83200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8130
timestamp 1654712443
transform 1 0 86200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8131
timestamp 1654712443
transform 1 0 89200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8132
timestamp 1654712443
transform 1 0 92200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8133
timestamp 1654712443
transform 1 0 95200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8134
timestamp 1654712443
transform 1 0 98200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8135
timestamp 1654712443
transform 1 0 101200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8136
timestamp 1654712443
transform 1 0 104200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8137
timestamp 1654712443
transform 1 0 107200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8138
timestamp 1654712443
transform 1 0 110200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8139
timestamp 1654712443
transform 1 0 113200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8140
timestamp 1654712443
transform 1 0 116200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8141
timestamp 1654712443
transform 1 0 119200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8142
timestamp 1654712443
transform 1 0 122200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8143
timestamp 1654712443
transform 1 0 125200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8144
timestamp 1654712443
transform 1 0 128200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8145
timestamp 1654712443
transform 1 0 131200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8146
timestamp 1654712443
transform 1 0 134200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8147
timestamp 1654712443
transform 1 0 137200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8148
timestamp 1654712443
transform 1 0 140200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8149
timestamp 1654712443
transform 1 0 143200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8150
timestamp 1654712443
transform 1 0 146200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8151
timestamp 1654712443
transform 1 0 149200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8152
timestamp 1654712443
transform 1 0 152200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8153
timestamp 1654712443
transform 1 0 155200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8154
timestamp 1654712443
transform 1 0 158200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8155
timestamp 1654712443
transform 1 0 161200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8156
timestamp 1654712443
transform 1 0 164200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8157
timestamp 1654712443
transform 1 0 167200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8158
timestamp 1654712443
transform 1 0 170200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8159
timestamp 1654712443
transform 1 0 173200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8160
timestamp 1654712443
transform 1 0 176200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8161
timestamp 1654712443
transform 1 0 179200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8163
timestamp 1654712443
transform 1 0 185200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8162
timestamp 1654712443
transform 1 0 182200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8164
timestamp 1654712443
transform 1 0 188200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8165
timestamp 1654712443
transform 1 0 191200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8166
timestamp 1654712443
transform 1 0 194200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8167
timestamp 1654712443
transform 1 0 197200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8168
timestamp 1654712443
transform 1 0 200200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8169
timestamp 1654712443
transform 1 0 203200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8170
timestamp 1654712443
transform 1 0 206200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8171
timestamp 1654712443
transform 1 0 209200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8173
timestamp 1654712443
transform 1 0 215200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8172
timestamp 1654712443
transform 1 0 212200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8174
timestamp 1654712443
transform 1 0 218200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8175
timestamp 1654712443
transform 1 0 221200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8176
timestamp 1654712443
transform 1 0 224200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8177
timestamp 1654712443
transform 1 0 227200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8178
timestamp 1654712443
transform 1 0 230200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8179
timestamp 1654712443
transform 1 0 233200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8180
timestamp 1654712443
transform 1 0 236200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8181
timestamp 1654712443
transform 1 0 239200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8183
timestamp 1654712443
transform 1 0 245200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8182
timestamp 1654712443
transform 1 0 242200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8184
timestamp 1654712443
transform 1 0 248200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8185
timestamp 1654712443
transform 1 0 251200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8186
timestamp 1654712443
transform 1 0 254200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8187
timestamp 1654712443
transform 1 0 257200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8188
timestamp 1654712443
transform 1 0 260200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8189
timestamp 1654712443
transform 1 0 263200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8190
timestamp 1654712443
transform 1 0 266200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8191
timestamp 1654712443
transform 1 0 269200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8192
timestamp 1654712443
transform 1 0 272200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8194
timestamp 1654712443
transform 1 0 278200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8193
timestamp 1654712443
transform 1 0 275200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8195
timestamp 1654712443
transform 1 0 281200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8196
timestamp 1654712443
transform 1 0 284200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8197
timestamp 1654712443
transform 1 0 287200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8198
timestamp 1654712443
transform 1 0 290200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8199
timestamp 1654712443
transform 1 0 293200 0 1 -240300
box 3640 -2860 6960 460
use pixel  pixel_8001
timestamp 1654712443
transform 1 0 -800 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8000
timestamp 1654712443
transform 1 0 -3800 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8002
timestamp 1654712443
transform 1 0 2200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8003
timestamp 1654712443
transform 1 0 5200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8004
timestamp 1654712443
transform 1 0 8200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8005
timestamp 1654712443
transform 1 0 11200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8006
timestamp 1654712443
transform 1 0 14200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8007
timestamp 1654712443
transform 1 0 17200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8008
timestamp 1654712443
transform 1 0 20200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8009
timestamp 1654712443
transform 1 0 23200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8011
timestamp 1654712443
transform 1 0 29200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8010
timestamp 1654712443
transform 1 0 26200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8012
timestamp 1654712443
transform 1 0 32200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8013
timestamp 1654712443
transform 1 0 35200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8014
timestamp 1654712443
transform 1 0 38200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8015
timestamp 1654712443
transform 1 0 41200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8016
timestamp 1654712443
transform 1 0 44200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8017
timestamp 1654712443
transform 1 0 47200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8018
timestamp 1654712443
transform 1 0 50200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8019
timestamp 1654712443
transform 1 0 53200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8021
timestamp 1654712443
transform 1 0 59200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8020
timestamp 1654712443
transform 1 0 56200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8022
timestamp 1654712443
transform 1 0 62200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8023
timestamp 1654712443
transform 1 0 65200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8024
timestamp 1654712443
transform 1 0 68200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8025
timestamp 1654712443
transform 1 0 71200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8026
timestamp 1654712443
transform 1 0 74200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8027
timestamp 1654712443
transform 1 0 77200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8028
timestamp 1654712443
transform 1 0 80200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8029
timestamp 1654712443
transform 1 0 83200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8030
timestamp 1654712443
transform 1 0 86200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8031
timestamp 1654712443
transform 1 0 89200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8032
timestamp 1654712443
transform 1 0 92200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8033
timestamp 1654712443
transform 1 0 95200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8034
timestamp 1654712443
transform 1 0 98200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8035
timestamp 1654712443
transform 1 0 101200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8036
timestamp 1654712443
transform 1 0 104200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8037
timestamp 1654712443
transform 1 0 107200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8038
timestamp 1654712443
transform 1 0 110200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8039
timestamp 1654712443
transform 1 0 113200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8040
timestamp 1654712443
transform 1 0 116200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8041
timestamp 1654712443
transform 1 0 119200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8042
timestamp 1654712443
transform 1 0 122200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8043
timestamp 1654712443
transform 1 0 125200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8044
timestamp 1654712443
transform 1 0 128200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8045
timestamp 1654712443
transform 1 0 131200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8046
timestamp 1654712443
transform 1 0 134200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8047
timestamp 1654712443
transform 1 0 137200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8048
timestamp 1654712443
transform 1 0 140200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8049
timestamp 1654712443
transform 1 0 143200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8050
timestamp 1654712443
transform 1 0 146200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8051
timestamp 1654712443
transform 1 0 149200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8052
timestamp 1654712443
transform 1 0 152200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8053
timestamp 1654712443
transform 1 0 155200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8054
timestamp 1654712443
transform 1 0 158200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8055
timestamp 1654712443
transform 1 0 161200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8056
timestamp 1654712443
transform 1 0 164200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8057
timestamp 1654712443
transform 1 0 167200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8058
timestamp 1654712443
transform 1 0 170200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8059
timestamp 1654712443
transform 1 0 173200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8060
timestamp 1654712443
transform 1 0 176200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8061
timestamp 1654712443
transform 1 0 179200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8063
timestamp 1654712443
transform 1 0 185200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8062
timestamp 1654712443
transform 1 0 182200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8064
timestamp 1654712443
transform 1 0 188200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8065
timestamp 1654712443
transform 1 0 191200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8066
timestamp 1654712443
transform 1 0 194200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8067
timestamp 1654712443
transform 1 0 197200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8068
timestamp 1654712443
transform 1 0 200200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8069
timestamp 1654712443
transform 1 0 203200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8070
timestamp 1654712443
transform 1 0 206200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8071
timestamp 1654712443
transform 1 0 209200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8073
timestamp 1654712443
transform 1 0 215200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8072
timestamp 1654712443
transform 1 0 212200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8074
timestamp 1654712443
transform 1 0 218200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8075
timestamp 1654712443
transform 1 0 221200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8076
timestamp 1654712443
transform 1 0 224200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8077
timestamp 1654712443
transform 1 0 227200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8078
timestamp 1654712443
transform 1 0 230200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8079
timestamp 1654712443
transform 1 0 233200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8080
timestamp 1654712443
transform 1 0 236200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8081
timestamp 1654712443
transform 1 0 239200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8083
timestamp 1654712443
transform 1 0 245200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8082
timestamp 1654712443
transform 1 0 242200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8084
timestamp 1654712443
transform 1 0 248200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8085
timestamp 1654712443
transform 1 0 251200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8086
timestamp 1654712443
transform 1 0 254200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8087
timestamp 1654712443
transform 1 0 257200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8088
timestamp 1654712443
transform 1 0 260200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8089
timestamp 1654712443
transform 1 0 263200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8090
timestamp 1654712443
transform 1 0 266200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8091
timestamp 1654712443
transform 1 0 269200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8092
timestamp 1654712443
transform 1 0 272200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8094
timestamp 1654712443
transform 1 0 278200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8093
timestamp 1654712443
transform 1 0 275200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8095
timestamp 1654712443
transform 1 0 281200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8096
timestamp 1654712443
transform 1 0 284200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8097
timestamp 1654712443
transform 1 0 287200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8098
timestamp 1654712443
transform 1 0 290200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_8099
timestamp 1654712443
transform 1 0 293200 0 1 -237300
box 3640 -2860 6960 460
use pixel  pixel_7801
timestamp 1654712443
transform 1 0 -800 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7800
timestamp 1654712443
transform 1 0 -3800 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7901
timestamp 1654712443
transform 1 0 -800 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7900
timestamp 1654712443
transform 1 0 -3800 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7802
timestamp 1654712443
transform 1 0 2200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7902
timestamp 1654712443
transform 1 0 2200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7803
timestamp 1654712443
transform 1 0 5200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7903
timestamp 1654712443
transform 1 0 5200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7804
timestamp 1654712443
transform 1 0 8200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7904
timestamp 1654712443
transform 1 0 8200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7805
timestamp 1654712443
transform 1 0 11200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7905
timestamp 1654712443
transform 1 0 11200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7806
timestamp 1654712443
transform 1 0 14200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7906
timestamp 1654712443
transform 1 0 14200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7807
timestamp 1654712443
transform 1 0 17200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7907
timestamp 1654712443
transform 1 0 17200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7808
timestamp 1654712443
transform 1 0 20200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7908
timestamp 1654712443
transform 1 0 20200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7809
timestamp 1654712443
transform 1 0 23200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7909
timestamp 1654712443
transform 1 0 23200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7811
timestamp 1654712443
transform 1 0 29200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7810
timestamp 1654712443
transform 1 0 26200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7911
timestamp 1654712443
transform 1 0 29200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7910
timestamp 1654712443
transform 1 0 26200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7812
timestamp 1654712443
transform 1 0 32200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7912
timestamp 1654712443
transform 1 0 32200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7813
timestamp 1654712443
transform 1 0 35200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7913
timestamp 1654712443
transform 1 0 35200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7814
timestamp 1654712443
transform 1 0 38200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7914
timestamp 1654712443
transform 1 0 38200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7815
timestamp 1654712443
transform 1 0 41200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7915
timestamp 1654712443
transform 1 0 41200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7816
timestamp 1654712443
transform 1 0 44200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7916
timestamp 1654712443
transform 1 0 44200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7817
timestamp 1654712443
transform 1 0 47200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7917
timestamp 1654712443
transform 1 0 47200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7818
timestamp 1654712443
transform 1 0 50200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7918
timestamp 1654712443
transform 1 0 50200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7819
timestamp 1654712443
transform 1 0 53200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7919
timestamp 1654712443
transform 1 0 53200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7821
timestamp 1654712443
transform 1 0 59200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7820
timestamp 1654712443
transform 1 0 56200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7921
timestamp 1654712443
transform 1 0 59200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7920
timestamp 1654712443
transform 1 0 56200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7822
timestamp 1654712443
transform 1 0 62200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7922
timestamp 1654712443
transform 1 0 62200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7823
timestamp 1654712443
transform 1 0 65200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7923
timestamp 1654712443
transform 1 0 65200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7824
timestamp 1654712443
transform 1 0 68200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7924
timestamp 1654712443
transform 1 0 68200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7825
timestamp 1654712443
transform 1 0 71200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7925
timestamp 1654712443
transform 1 0 71200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7826
timestamp 1654712443
transform 1 0 74200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7926
timestamp 1654712443
transform 1 0 74200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7827
timestamp 1654712443
transform 1 0 77200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7927
timestamp 1654712443
transform 1 0 77200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7828
timestamp 1654712443
transform 1 0 80200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7928
timestamp 1654712443
transform 1 0 80200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7829
timestamp 1654712443
transform 1 0 83200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7929
timestamp 1654712443
transform 1 0 83200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7830
timestamp 1654712443
transform 1 0 86200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7930
timestamp 1654712443
transform 1 0 86200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7831
timestamp 1654712443
transform 1 0 89200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7832
timestamp 1654712443
transform 1 0 92200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7931
timestamp 1654712443
transform 1 0 89200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7932
timestamp 1654712443
transform 1 0 92200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7833
timestamp 1654712443
transform 1 0 95200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7933
timestamp 1654712443
transform 1 0 95200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7834
timestamp 1654712443
transform 1 0 98200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7934
timestamp 1654712443
transform 1 0 98200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7835
timestamp 1654712443
transform 1 0 101200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7935
timestamp 1654712443
transform 1 0 101200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7836
timestamp 1654712443
transform 1 0 104200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7936
timestamp 1654712443
transform 1 0 104200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7837
timestamp 1654712443
transform 1 0 107200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7937
timestamp 1654712443
transform 1 0 107200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7838
timestamp 1654712443
transform 1 0 110200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7938
timestamp 1654712443
transform 1 0 110200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7839
timestamp 1654712443
transform 1 0 113200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7939
timestamp 1654712443
transform 1 0 113200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7840
timestamp 1654712443
transform 1 0 116200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7940
timestamp 1654712443
transform 1 0 116200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7841
timestamp 1654712443
transform 1 0 119200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7842
timestamp 1654712443
transform 1 0 122200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7941
timestamp 1654712443
transform 1 0 119200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7942
timestamp 1654712443
transform 1 0 122200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7843
timestamp 1654712443
transform 1 0 125200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7943
timestamp 1654712443
transform 1 0 125200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7844
timestamp 1654712443
transform 1 0 128200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7944
timestamp 1654712443
transform 1 0 128200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7845
timestamp 1654712443
transform 1 0 131200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7945
timestamp 1654712443
transform 1 0 131200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7846
timestamp 1654712443
transform 1 0 134200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7946
timestamp 1654712443
transform 1 0 134200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7847
timestamp 1654712443
transform 1 0 137200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7947
timestamp 1654712443
transform 1 0 137200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7848
timestamp 1654712443
transform 1 0 140200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7948
timestamp 1654712443
transform 1 0 140200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7849
timestamp 1654712443
transform 1 0 143200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7949
timestamp 1654712443
transform 1 0 143200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7850
timestamp 1654712443
transform 1 0 146200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7950
timestamp 1654712443
transform 1 0 146200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7851
timestamp 1654712443
transform 1 0 149200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7852
timestamp 1654712443
transform 1 0 152200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7951
timestamp 1654712443
transform 1 0 149200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7952
timestamp 1654712443
transform 1 0 152200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7853
timestamp 1654712443
transform 1 0 155200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7953
timestamp 1654712443
transform 1 0 155200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7854
timestamp 1654712443
transform 1 0 158200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7954
timestamp 1654712443
transform 1 0 158200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7855
timestamp 1654712443
transform 1 0 161200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7955
timestamp 1654712443
transform 1 0 161200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7856
timestamp 1654712443
transform 1 0 164200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7956
timestamp 1654712443
transform 1 0 164200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7857
timestamp 1654712443
transform 1 0 167200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7957
timestamp 1654712443
transform 1 0 167200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7858
timestamp 1654712443
transform 1 0 170200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7958
timestamp 1654712443
transform 1 0 170200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7859
timestamp 1654712443
transform 1 0 173200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7959
timestamp 1654712443
transform 1 0 173200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7860
timestamp 1654712443
transform 1 0 176200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7960
timestamp 1654712443
transform 1 0 176200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7861
timestamp 1654712443
transform 1 0 179200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7961
timestamp 1654712443
transform 1 0 179200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7863
timestamp 1654712443
transform 1 0 185200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7862
timestamp 1654712443
transform 1 0 182200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7963
timestamp 1654712443
transform 1 0 185200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7962
timestamp 1654712443
transform 1 0 182200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7864
timestamp 1654712443
transform 1 0 188200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7964
timestamp 1654712443
transform 1 0 188200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7865
timestamp 1654712443
transform 1 0 191200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7965
timestamp 1654712443
transform 1 0 191200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7866
timestamp 1654712443
transform 1 0 194200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7966
timestamp 1654712443
transform 1 0 194200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7867
timestamp 1654712443
transform 1 0 197200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7967
timestamp 1654712443
transform 1 0 197200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7868
timestamp 1654712443
transform 1 0 200200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7968
timestamp 1654712443
transform 1 0 200200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7869
timestamp 1654712443
transform 1 0 203200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7969
timestamp 1654712443
transform 1 0 203200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7870
timestamp 1654712443
transform 1 0 206200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7970
timestamp 1654712443
transform 1 0 206200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7871
timestamp 1654712443
transform 1 0 209200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7971
timestamp 1654712443
transform 1 0 209200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7873
timestamp 1654712443
transform 1 0 215200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7872
timestamp 1654712443
transform 1 0 212200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7973
timestamp 1654712443
transform 1 0 215200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7972
timestamp 1654712443
transform 1 0 212200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7874
timestamp 1654712443
transform 1 0 218200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7974
timestamp 1654712443
transform 1 0 218200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7875
timestamp 1654712443
transform 1 0 221200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7975
timestamp 1654712443
transform 1 0 221200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7876
timestamp 1654712443
transform 1 0 224200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7976
timestamp 1654712443
transform 1 0 224200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7877
timestamp 1654712443
transform 1 0 227200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7977
timestamp 1654712443
transform 1 0 227200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7878
timestamp 1654712443
transform 1 0 230200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7978
timestamp 1654712443
transform 1 0 230200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7879
timestamp 1654712443
transform 1 0 233200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7979
timestamp 1654712443
transform 1 0 233200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7880
timestamp 1654712443
transform 1 0 236200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7980
timestamp 1654712443
transform 1 0 236200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7881
timestamp 1654712443
transform 1 0 239200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7981
timestamp 1654712443
transform 1 0 239200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7883
timestamp 1654712443
transform 1 0 245200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7882
timestamp 1654712443
transform 1 0 242200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7983
timestamp 1654712443
transform 1 0 245200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7982
timestamp 1654712443
transform 1 0 242200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7884
timestamp 1654712443
transform 1 0 248200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7984
timestamp 1654712443
transform 1 0 248200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7885
timestamp 1654712443
transform 1 0 251200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7985
timestamp 1654712443
transform 1 0 251200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7886
timestamp 1654712443
transform 1 0 254200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7986
timestamp 1654712443
transform 1 0 254200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7887
timestamp 1654712443
transform 1 0 257200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7987
timestamp 1654712443
transform 1 0 257200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7888
timestamp 1654712443
transform 1 0 260200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7988
timestamp 1654712443
transform 1 0 260200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7889
timestamp 1654712443
transform 1 0 263200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7989
timestamp 1654712443
transform 1 0 263200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7890
timestamp 1654712443
transform 1 0 266200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7990
timestamp 1654712443
transform 1 0 266200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7891
timestamp 1654712443
transform 1 0 269200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7991
timestamp 1654712443
transform 1 0 269200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7892
timestamp 1654712443
transform 1 0 272200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7992
timestamp 1654712443
transform 1 0 272200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7894
timestamp 1654712443
transform 1 0 278200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7893
timestamp 1654712443
transform 1 0 275200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7994
timestamp 1654712443
transform 1 0 278200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7993
timestamp 1654712443
transform 1 0 275200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7895
timestamp 1654712443
transform 1 0 281200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7995
timestamp 1654712443
transform 1 0 281200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7896
timestamp 1654712443
transform 1 0 284200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7996
timestamp 1654712443
transform 1 0 284200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7897
timestamp 1654712443
transform 1 0 287200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7997
timestamp 1654712443
transform 1 0 287200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7898
timestamp 1654712443
transform 1 0 290200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7998
timestamp 1654712443
transform 1 0 290200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7899
timestamp 1654712443
transform 1 0 293200 0 1 -231300
box 3640 -2860 6960 460
use pixel  pixel_7999
timestamp 1654712443
transform 1 0 293200 0 1 -234300
box 3640 -2860 6960 460
use pixel  pixel_7701
timestamp 1654712443
transform 1 0 -800 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7700
timestamp 1654712443
transform 1 0 -3800 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7702
timestamp 1654712443
transform 1 0 2200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7703
timestamp 1654712443
transform 1 0 5200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7704
timestamp 1654712443
transform 1 0 8200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7705
timestamp 1654712443
transform 1 0 11200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7706
timestamp 1654712443
transform 1 0 14200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7707
timestamp 1654712443
transform 1 0 17200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7708
timestamp 1654712443
transform 1 0 20200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7709
timestamp 1654712443
transform 1 0 23200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7711
timestamp 1654712443
transform 1 0 29200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7710
timestamp 1654712443
transform 1 0 26200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7712
timestamp 1654712443
transform 1 0 32200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7713
timestamp 1654712443
transform 1 0 35200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7714
timestamp 1654712443
transform 1 0 38200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7715
timestamp 1654712443
transform 1 0 41200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7716
timestamp 1654712443
transform 1 0 44200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7717
timestamp 1654712443
transform 1 0 47200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7718
timestamp 1654712443
transform 1 0 50200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7719
timestamp 1654712443
transform 1 0 53200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7721
timestamp 1654712443
transform 1 0 59200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7720
timestamp 1654712443
transform 1 0 56200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7722
timestamp 1654712443
transform 1 0 62200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7723
timestamp 1654712443
transform 1 0 65200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7724
timestamp 1654712443
transform 1 0 68200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7725
timestamp 1654712443
transform 1 0 71200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7726
timestamp 1654712443
transform 1 0 74200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7727
timestamp 1654712443
transform 1 0 77200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7728
timestamp 1654712443
transform 1 0 80200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7729
timestamp 1654712443
transform 1 0 83200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7730
timestamp 1654712443
transform 1 0 86200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7731
timestamp 1654712443
transform 1 0 89200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7732
timestamp 1654712443
transform 1 0 92200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7733
timestamp 1654712443
transform 1 0 95200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7734
timestamp 1654712443
transform 1 0 98200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7735
timestamp 1654712443
transform 1 0 101200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7736
timestamp 1654712443
transform 1 0 104200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7737
timestamp 1654712443
transform 1 0 107200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7738
timestamp 1654712443
transform 1 0 110200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7739
timestamp 1654712443
transform 1 0 113200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7740
timestamp 1654712443
transform 1 0 116200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7741
timestamp 1654712443
transform 1 0 119200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7742
timestamp 1654712443
transform 1 0 122200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7743
timestamp 1654712443
transform 1 0 125200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7744
timestamp 1654712443
transform 1 0 128200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7745
timestamp 1654712443
transform 1 0 131200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7746
timestamp 1654712443
transform 1 0 134200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7747
timestamp 1654712443
transform 1 0 137200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7748
timestamp 1654712443
transform 1 0 140200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7749
timestamp 1654712443
transform 1 0 143200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7750
timestamp 1654712443
transform 1 0 146200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7751
timestamp 1654712443
transform 1 0 149200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7752
timestamp 1654712443
transform 1 0 152200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7753
timestamp 1654712443
transform 1 0 155200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7754
timestamp 1654712443
transform 1 0 158200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7755
timestamp 1654712443
transform 1 0 161200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7756
timestamp 1654712443
transform 1 0 164200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7757
timestamp 1654712443
transform 1 0 167200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7758
timestamp 1654712443
transform 1 0 170200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7759
timestamp 1654712443
transform 1 0 173200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7760
timestamp 1654712443
transform 1 0 176200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7761
timestamp 1654712443
transform 1 0 179200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7763
timestamp 1654712443
transform 1 0 185200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7762
timestamp 1654712443
transform 1 0 182200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7764
timestamp 1654712443
transform 1 0 188200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7765
timestamp 1654712443
transform 1 0 191200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7766
timestamp 1654712443
transform 1 0 194200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7767
timestamp 1654712443
transform 1 0 197200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7768
timestamp 1654712443
transform 1 0 200200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7769
timestamp 1654712443
transform 1 0 203200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7770
timestamp 1654712443
transform 1 0 206200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7771
timestamp 1654712443
transform 1 0 209200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7773
timestamp 1654712443
transform 1 0 215200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7772
timestamp 1654712443
transform 1 0 212200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7774
timestamp 1654712443
transform 1 0 218200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7775
timestamp 1654712443
transform 1 0 221200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7776
timestamp 1654712443
transform 1 0 224200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7777
timestamp 1654712443
transform 1 0 227200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7778
timestamp 1654712443
transform 1 0 230200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7779
timestamp 1654712443
transform 1 0 233200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7780
timestamp 1654712443
transform 1 0 236200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7781
timestamp 1654712443
transform 1 0 239200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7783
timestamp 1654712443
transform 1 0 245200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7782
timestamp 1654712443
transform 1 0 242200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7784
timestamp 1654712443
transform 1 0 248200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7785
timestamp 1654712443
transform 1 0 251200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7786
timestamp 1654712443
transform 1 0 254200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7787
timestamp 1654712443
transform 1 0 257200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7788
timestamp 1654712443
transform 1 0 260200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7789
timestamp 1654712443
transform 1 0 263200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7790
timestamp 1654712443
transform 1 0 266200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7791
timestamp 1654712443
transform 1 0 269200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7792
timestamp 1654712443
transform 1 0 272200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7794
timestamp 1654712443
transform 1 0 278200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7793
timestamp 1654712443
transform 1 0 275200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7795
timestamp 1654712443
transform 1 0 281200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7796
timestamp 1654712443
transform 1 0 284200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7797
timestamp 1654712443
transform 1 0 287200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7798
timestamp 1654712443
transform 1 0 290200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7799
timestamp 1654712443
transform 1 0 293200 0 1 -228300
box 3640 -2860 6960 460
use pixel  pixel_7601
timestamp 1654712443
transform 1 0 -800 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7600
timestamp 1654712443
transform 1 0 -3800 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7602
timestamp 1654712443
transform 1 0 2200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7603
timestamp 1654712443
transform 1 0 5200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7604
timestamp 1654712443
transform 1 0 8200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7605
timestamp 1654712443
transform 1 0 11200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7606
timestamp 1654712443
transform 1 0 14200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7607
timestamp 1654712443
transform 1 0 17200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7608
timestamp 1654712443
transform 1 0 20200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7609
timestamp 1654712443
transform 1 0 23200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7611
timestamp 1654712443
transform 1 0 29200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7610
timestamp 1654712443
transform 1 0 26200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7612
timestamp 1654712443
transform 1 0 32200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7613
timestamp 1654712443
transform 1 0 35200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7614
timestamp 1654712443
transform 1 0 38200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7615
timestamp 1654712443
transform 1 0 41200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7616
timestamp 1654712443
transform 1 0 44200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7617
timestamp 1654712443
transform 1 0 47200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7618
timestamp 1654712443
transform 1 0 50200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7619
timestamp 1654712443
transform 1 0 53200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7621
timestamp 1654712443
transform 1 0 59200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7620
timestamp 1654712443
transform 1 0 56200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7622
timestamp 1654712443
transform 1 0 62200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7623
timestamp 1654712443
transform 1 0 65200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7624
timestamp 1654712443
transform 1 0 68200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7625
timestamp 1654712443
transform 1 0 71200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7626
timestamp 1654712443
transform 1 0 74200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7627
timestamp 1654712443
transform 1 0 77200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7628
timestamp 1654712443
transform 1 0 80200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7629
timestamp 1654712443
transform 1 0 83200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7630
timestamp 1654712443
transform 1 0 86200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7631
timestamp 1654712443
transform 1 0 89200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7632
timestamp 1654712443
transform 1 0 92200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7633
timestamp 1654712443
transform 1 0 95200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7634
timestamp 1654712443
transform 1 0 98200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7635
timestamp 1654712443
transform 1 0 101200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7636
timestamp 1654712443
transform 1 0 104200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7637
timestamp 1654712443
transform 1 0 107200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7638
timestamp 1654712443
transform 1 0 110200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7639
timestamp 1654712443
transform 1 0 113200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7640
timestamp 1654712443
transform 1 0 116200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7641
timestamp 1654712443
transform 1 0 119200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7642
timestamp 1654712443
transform 1 0 122200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7643
timestamp 1654712443
transform 1 0 125200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7644
timestamp 1654712443
transform 1 0 128200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7645
timestamp 1654712443
transform 1 0 131200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7646
timestamp 1654712443
transform 1 0 134200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7647
timestamp 1654712443
transform 1 0 137200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7648
timestamp 1654712443
transform 1 0 140200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7649
timestamp 1654712443
transform 1 0 143200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7650
timestamp 1654712443
transform 1 0 146200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7651
timestamp 1654712443
transform 1 0 149200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7652
timestamp 1654712443
transform 1 0 152200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7653
timestamp 1654712443
transform 1 0 155200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7654
timestamp 1654712443
transform 1 0 158200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7655
timestamp 1654712443
transform 1 0 161200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7656
timestamp 1654712443
transform 1 0 164200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7657
timestamp 1654712443
transform 1 0 167200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7658
timestamp 1654712443
transform 1 0 170200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7659
timestamp 1654712443
transform 1 0 173200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7660
timestamp 1654712443
transform 1 0 176200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7661
timestamp 1654712443
transform 1 0 179200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7663
timestamp 1654712443
transform 1 0 185200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7662
timestamp 1654712443
transform 1 0 182200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7664
timestamp 1654712443
transform 1 0 188200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7665
timestamp 1654712443
transform 1 0 191200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7666
timestamp 1654712443
transform 1 0 194200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7667
timestamp 1654712443
transform 1 0 197200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7668
timestamp 1654712443
transform 1 0 200200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7669
timestamp 1654712443
transform 1 0 203200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7670
timestamp 1654712443
transform 1 0 206200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7671
timestamp 1654712443
transform 1 0 209200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7673
timestamp 1654712443
transform 1 0 215200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7672
timestamp 1654712443
transform 1 0 212200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7674
timestamp 1654712443
transform 1 0 218200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7675
timestamp 1654712443
transform 1 0 221200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7676
timestamp 1654712443
transform 1 0 224200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7677
timestamp 1654712443
transform 1 0 227200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7678
timestamp 1654712443
transform 1 0 230200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7679
timestamp 1654712443
transform 1 0 233200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7680
timestamp 1654712443
transform 1 0 236200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7681
timestamp 1654712443
transform 1 0 239200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7683
timestamp 1654712443
transform 1 0 245200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7682
timestamp 1654712443
transform 1 0 242200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7684
timestamp 1654712443
transform 1 0 248200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7685
timestamp 1654712443
transform 1 0 251200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7686
timestamp 1654712443
transform 1 0 254200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7687
timestamp 1654712443
transform 1 0 257200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7688
timestamp 1654712443
transform 1 0 260200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7689
timestamp 1654712443
transform 1 0 263200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7690
timestamp 1654712443
transform 1 0 266200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7691
timestamp 1654712443
transform 1 0 269200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7692
timestamp 1654712443
transform 1 0 272200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7694
timestamp 1654712443
transform 1 0 278200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7693
timestamp 1654712443
transform 1 0 275200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7695
timestamp 1654712443
transform 1 0 281200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7696
timestamp 1654712443
transform 1 0 284200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7697
timestamp 1654712443
transform 1 0 287200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7698
timestamp 1654712443
transform 1 0 290200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7699
timestamp 1654712443
transform 1 0 293200 0 1 -225300
box 3640 -2860 6960 460
use pixel  pixel_7501
timestamp 1654712443
transform 1 0 -800 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7500
timestamp 1654712443
transform 1 0 -3800 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7502
timestamp 1654712443
transform 1 0 2200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7503
timestamp 1654712443
transform 1 0 5200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7504
timestamp 1654712443
transform 1 0 8200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7505
timestamp 1654712443
transform 1 0 11200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7506
timestamp 1654712443
transform 1 0 14200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7507
timestamp 1654712443
transform 1 0 17200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7508
timestamp 1654712443
transform 1 0 20200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7509
timestamp 1654712443
transform 1 0 23200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7511
timestamp 1654712443
transform 1 0 29200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7510
timestamp 1654712443
transform 1 0 26200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7512
timestamp 1654712443
transform 1 0 32200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7513
timestamp 1654712443
transform 1 0 35200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7514
timestamp 1654712443
transform 1 0 38200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7515
timestamp 1654712443
transform 1 0 41200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7516
timestamp 1654712443
transform 1 0 44200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7517
timestamp 1654712443
transform 1 0 47200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7518
timestamp 1654712443
transform 1 0 50200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7519
timestamp 1654712443
transform 1 0 53200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7521
timestamp 1654712443
transform 1 0 59200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7520
timestamp 1654712443
transform 1 0 56200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7522
timestamp 1654712443
transform 1 0 62200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7523
timestamp 1654712443
transform 1 0 65200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7524
timestamp 1654712443
transform 1 0 68200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7525
timestamp 1654712443
transform 1 0 71200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7526
timestamp 1654712443
transform 1 0 74200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7527
timestamp 1654712443
transform 1 0 77200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7528
timestamp 1654712443
transform 1 0 80200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7529
timestamp 1654712443
transform 1 0 83200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7530
timestamp 1654712443
transform 1 0 86200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7531
timestamp 1654712443
transform 1 0 89200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7532
timestamp 1654712443
transform 1 0 92200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7533
timestamp 1654712443
transform 1 0 95200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7534
timestamp 1654712443
transform 1 0 98200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7535
timestamp 1654712443
transform 1 0 101200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7536
timestamp 1654712443
transform 1 0 104200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7537
timestamp 1654712443
transform 1 0 107200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7538
timestamp 1654712443
transform 1 0 110200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7539
timestamp 1654712443
transform 1 0 113200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7540
timestamp 1654712443
transform 1 0 116200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7541
timestamp 1654712443
transform 1 0 119200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7542
timestamp 1654712443
transform 1 0 122200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7543
timestamp 1654712443
transform 1 0 125200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7544
timestamp 1654712443
transform 1 0 128200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7545
timestamp 1654712443
transform 1 0 131200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7546
timestamp 1654712443
transform 1 0 134200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7547
timestamp 1654712443
transform 1 0 137200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7548
timestamp 1654712443
transform 1 0 140200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7549
timestamp 1654712443
transform 1 0 143200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7550
timestamp 1654712443
transform 1 0 146200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7551
timestamp 1654712443
transform 1 0 149200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7552
timestamp 1654712443
transform 1 0 152200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7553
timestamp 1654712443
transform 1 0 155200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7554
timestamp 1654712443
transform 1 0 158200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7555
timestamp 1654712443
transform 1 0 161200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7556
timestamp 1654712443
transform 1 0 164200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7557
timestamp 1654712443
transform 1 0 167200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7558
timestamp 1654712443
transform 1 0 170200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7559
timestamp 1654712443
transform 1 0 173200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7560
timestamp 1654712443
transform 1 0 176200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7561
timestamp 1654712443
transform 1 0 179200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7563
timestamp 1654712443
transform 1 0 185200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7562
timestamp 1654712443
transform 1 0 182200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7564
timestamp 1654712443
transform 1 0 188200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7565
timestamp 1654712443
transform 1 0 191200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7566
timestamp 1654712443
transform 1 0 194200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7567
timestamp 1654712443
transform 1 0 197200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7568
timestamp 1654712443
transform 1 0 200200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7569
timestamp 1654712443
transform 1 0 203200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7570
timestamp 1654712443
transform 1 0 206200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7571
timestamp 1654712443
transform 1 0 209200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7573
timestamp 1654712443
transform 1 0 215200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7572
timestamp 1654712443
transform 1 0 212200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7574
timestamp 1654712443
transform 1 0 218200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7575
timestamp 1654712443
transform 1 0 221200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7576
timestamp 1654712443
transform 1 0 224200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7577
timestamp 1654712443
transform 1 0 227200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7578
timestamp 1654712443
transform 1 0 230200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7579
timestamp 1654712443
transform 1 0 233200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7580
timestamp 1654712443
transform 1 0 236200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7581
timestamp 1654712443
transform 1 0 239200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7583
timestamp 1654712443
transform 1 0 245200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7582
timestamp 1654712443
transform 1 0 242200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7584
timestamp 1654712443
transform 1 0 248200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7585
timestamp 1654712443
transform 1 0 251200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7586
timestamp 1654712443
transform 1 0 254200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7587
timestamp 1654712443
transform 1 0 257200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7588
timestamp 1654712443
transform 1 0 260200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7589
timestamp 1654712443
transform 1 0 263200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7590
timestamp 1654712443
transform 1 0 266200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7591
timestamp 1654712443
transform 1 0 269200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7592
timestamp 1654712443
transform 1 0 272200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7594
timestamp 1654712443
transform 1 0 278200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7593
timestamp 1654712443
transform 1 0 275200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7595
timestamp 1654712443
transform 1 0 281200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7596
timestamp 1654712443
transform 1 0 284200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7597
timestamp 1654712443
transform 1 0 287200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7598
timestamp 1654712443
transform 1 0 290200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7599
timestamp 1654712443
transform 1 0 293200 0 1 -222300
box 3640 -2860 6960 460
use pixel  pixel_7401
timestamp 1654712443
transform 1 0 -800 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7400
timestamp 1654712443
transform 1 0 -3800 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7402
timestamp 1654712443
transform 1 0 2200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7403
timestamp 1654712443
transform 1 0 5200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7404
timestamp 1654712443
transform 1 0 8200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7405
timestamp 1654712443
transform 1 0 11200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7406
timestamp 1654712443
transform 1 0 14200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7407
timestamp 1654712443
transform 1 0 17200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7408
timestamp 1654712443
transform 1 0 20200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7409
timestamp 1654712443
transform 1 0 23200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7411
timestamp 1654712443
transform 1 0 29200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7410
timestamp 1654712443
transform 1 0 26200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7412
timestamp 1654712443
transform 1 0 32200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7413
timestamp 1654712443
transform 1 0 35200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7414
timestamp 1654712443
transform 1 0 38200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7415
timestamp 1654712443
transform 1 0 41200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7416
timestamp 1654712443
transform 1 0 44200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7417
timestamp 1654712443
transform 1 0 47200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7418
timestamp 1654712443
transform 1 0 50200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7419
timestamp 1654712443
transform 1 0 53200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7421
timestamp 1654712443
transform 1 0 59200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7420
timestamp 1654712443
transform 1 0 56200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7422
timestamp 1654712443
transform 1 0 62200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7423
timestamp 1654712443
transform 1 0 65200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7424
timestamp 1654712443
transform 1 0 68200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7425
timestamp 1654712443
transform 1 0 71200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7426
timestamp 1654712443
transform 1 0 74200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7427
timestamp 1654712443
transform 1 0 77200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7428
timestamp 1654712443
transform 1 0 80200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7429
timestamp 1654712443
transform 1 0 83200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7430
timestamp 1654712443
transform 1 0 86200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7431
timestamp 1654712443
transform 1 0 89200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7432
timestamp 1654712443
transform 1 0 92200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7433
timestamp 1654712443
transform 1 0 95200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7434
timestamp 1654712443
transform 1 0 98200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7435
timestamp 1654712443
transform 1 0 101200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7436
timestamp 1654712443
transform 1 0 104200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7437
timestamp 1654712443
transform 1 0 107200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7438
timestamp 1654712443
transform 1 0 110200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7439
timestamp 1654712443
transform 1 0 113200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7440
timestamp 1654712443
transform 1 0 116200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7441
timestamp 1654712443
transform 1 0 119200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7442
timestamp 1654712443
transform 1 0 122200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7443
timestamp 1654712443
transform 1 0 125200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7444
timestamp 1654712443
transform 1 0 128200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7445
timestamp 1654712443
transform 1 0 131200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7446
timestamp 1654712443
transform 1 0 134200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7447
timestamp 1654712443
transform 1 0 137200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7448
timestamp 1654712443
transform 1 0 140200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7449
timestamp 1654712443
transform 1 0 143200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7450
timestamp 1654712443
transform 1 0 146200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7451
timestamp 1654712443
transform 1 0 149200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7452
timestamp 1654712443
transform 1 0 152200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7453
timestamp 1654712443
transform 1 0 155200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7454
timestamp 1654712443
transform 1 0 158200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7455
timestamp 1654712443
transform 1 0 161200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7456
timestamp 1654712443
transform 1 0 164200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7457
timestamp 1654712443
transform 1 0 167200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7458
timestamp 1654712443
transform 1 0 170200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7459
timestamp 1654712443
transform 1 0 173200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7460
timestamp 1654712443
transform 1 0 176200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7461
timestamp 1654712443
transform 1 0 179200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7463
timestamp 1654712443
transform 1 0 185200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7462
timestamp 1654712443
transform 1 0 182200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7464
timestamp 1654712443
transform 1 0 188200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7465
timestamp 1654712443
transform 1 0 191200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7466
timestamp 1654712443
transform 1 0 194200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7467
timestamp 1654712443
transform 1 0 197200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7468
timestamp 1654712443
transform 1 0 200200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7469
timestamp 1654712443
transform 1 0 203200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7470
timestamp 1654712443
transform 1 0 206200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7471
timestamp 1654712443
transform 1 0 209200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7473
timestamp 1654712443
transform 1 0 215200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7472
timestamp 1654712443
transform 1 0 212200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7474
timestamp 1654712443
transform 1 0 218200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7475
timestamp 1654712443
transform 1 0 221200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7476
timestamp 1654712443
transform 1 0 224200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7477
timestamp 1654712443
transform 1 0 227200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7478
timestamp 1654712443
transform 1 0 230200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7479
timestamp 1654712443
transform 1 0 233200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7480
timestamp 1654712443
transform 1 0 236200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7481
timestamp 1654712443
transform 1 0 239200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7483
timestamp 1654712443
transform 1 0 245200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7482
timestamp 1654712443
transform 1 0 242200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7484
timestamp 1654712443
transform 1 0 248200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7485
timestamp 1654712443
transform 1 0 251200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7486
timestamp 1654712443
transform 1 0 254200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7487
timestamp 1654712443
transform 1 0 257200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7488
timestamp 1654712443
transform 1 0 260200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7489
timestamp 1654712443
transform 1 0 263200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7490
timestamp 1654712443
transform 1 0 266200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7491
timestamp 1654712443
transform 1 0 269200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7492
timestamp 1654712443
transform 1 0 272200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7494
timestamp 1654712443
transform 1 0 278200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7493
timestamp 1654712443
transform 1 0 275200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7495
timestamp 1654712443
transform 1 0 281200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7496
timestamp 1654712443
transform 1 0 284200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7497
timestamp 1654712443
transform 1 0 287200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7498
timestamp 1654712443
transform 1 0 290200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7499
timestamp 1654712443
transform 1 0 293200 0 1 -219300
box 3640 -2860 6960 460
use pixel  pixel_7301
timestamp 1654712443
transform 1 0 -800 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7300
timestamp 1654712443
transform 1 0 -3800 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7302
timestamp 1654712443
transform 1 0 2200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7303
timestamp 1654712443
transform 1 0 5200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7304
timestamp 1654712443
transform 1 0 8200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7305
timestamp 1654712443
transform 1 0 11200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7306
timestamp 1654712443
transform 1 0 14200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7307
timestamp 1654712443
transform 1 0 17200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7308
timestamp 1654712443
transform 1 0 20200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7309
timestamp 1654712443
transform 1 0 23200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7311
timestamp 1654712443
transform 1 0 29200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7310
timestamp 1654712443
transform 1 0 26200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7312
timestamp 1654712443
transform 1 0 32200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7313
timestamp 1654712443
transform 1 0 35200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7314
timestamp 1654712443
transform 1 0 38200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7315
timestamp 1654712443
transform 1 0 41200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7316
timestamp 1654712443
transform 1 0 44200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7317
timestamp 1654712443
transform 1 0 47200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7318
timestamp 1654712443
transform 1 0 50200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7319
timestamp 1654712443
transform 1 0 53200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7321
timestamp 1654712443
transform 1 0 59200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7320
timestamp 1654712443
transform 1 0 56200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7322
timestamp 1654712443
transform 1 0 62200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7323
timestamp 1654712443
transform 1 0 65200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7324
timestamp 1654712443
transform 1 0 68200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7325
timestamp 1654712443
transform 1 0 71200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7326
timestamp 1654712443
transform 1 0 74200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7327
timestamp 1654712443
transform 1 0 77200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7328
timestamp 1654712443
transform 1 0 80200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7329
timestamp 1654712443
transform 1 0 83200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7330
timestamp 1654712443
transform 1 0 86200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7331
timestamp 1654712443
transform 1 0 89200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7332
timestamp 1654712443
transform 1 0 92200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7333
timestamp 1654712443
transform 1 0 95200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7334
timestamp 1654712443
transform 1 0 98200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7335
timestamp 1654712443
transform 1 0 101200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7336
timestamp 1654712443
transform 1 0 104200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7337
timestamp 1654712443
transform 1 0 107200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7338
timestamp 1654712443
transform 1 0 110200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7339
timestamp 1654712443
transform 1 0 113200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7340
timestamp 1654712443
transform 1 0 116200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7341
timestamp 1654712443
transform 1 0 119200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7342
timestamp 1654712443
transform 1 0 122200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7343
timestamp 1654712443
transform 1 0 125200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7344
timestamp 1654712443
transform 1 0 128200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7345
timestamp 1654712443
transform 1 0 131200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7346
timestamp 1654712443
transform 1 0 134200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7347
timestamp 1654712443
transform 1 0 137200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7348
timestamp 1654712443
transform 1 0 140200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7349
timestamp 1654712443
transform 1 0 143200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7350
timestamp 1654712443
transform 1 0 146200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7351
timestamp 1654712443
transform 1 0 149200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7352
timestamp 1654712443
transform 1 0 152200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7353
timestamp 1654712443
transform 1 0 155200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7354
timestamp 1654712443
transform 1 0 158200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7355
timestamp 1654712443
transform 1 0 161200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7356
timestamp 1654712443
transform 1 0 164200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7357
timestamp 1654712443
transform 1 0 167200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7358
timestamp 1654712443
transform 1 0 170200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7359
timestamp 1654712443
transform 1 0 173200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7360
timestamp 1654712443
transform 1 0 176200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7361
timestamp 1654712443
transform 1 0 179200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7363
timestamp 1654712443
transform 1 0 185200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7362
timestamp 1654712443
transform 1 0 182200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7364
timestamp 1654712443
transform 1 0 188200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7365
timestamp 1654712443
transform 1 0 191200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7366
timestamp 1654712443
transform 1 0 194200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7367
timestamp 1654712443
transform 1 0 197200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7368
timestamp 1654712443
transform 1 0 200200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7369
timestamp 1654712443
transform 1 0 203200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7370
timestamp 1654712443
transform 1 0 206200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7371
timestamp 1654712443
transform 1 0 209200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7373
timestamp 1654712443
transform 1 0 215200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7372
timestamp 1654712443
transform 1 0 212200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7374
timestamp 1654712443
transform 1 0 218200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7375
timestamp 1654712443
transform 1 0 221200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7376
timestamp 1654712443
transform 1 0 224200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7377
timestamp 1654712443
transform 1 0 227200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7378
timestamp 1654712443
transform 1 0 230200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7379
timestamp 1654712443
transform 1 0 233200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7380
timestamp 1654712443
transform 1 0 236200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7381
timestamp 1654712443
transform 1 0 239200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7383
timestamp 1654712443
transform 1 0 245200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7382
timestamp 1654712443
transform 1 0 242200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7384
timestamp 1654712443
transform 1 0 248200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7385
timestamp 1654712443
transform 1 0 251200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7386
timestamp 1654712443
transform 1 0 254200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7387
timestamp 1654712443
transform 1 0 257200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7388
timestamp 1654712443
transform 1 0 260200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7389
timestamp 1654712443
transform 1 0 263200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7390
timestamp 1654712443
transform 1 0 266200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7391
timestamp 1654712443
transform 1 0 269200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7392
timestamp 1654712443
transform 1 0 272200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7394
timestamp 1654712443
transform 1 0 278200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7393
timestamp 1654712443
transform 1 0 275200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7395
timestamp 1654712443
transform 1 0 281200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7396
timestamp 1654712443
transform 1 0 284200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7397
timestamp 1654712443
transform 1 0 287200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7398
timestamp 1654712443
transform 1 0 290200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7399
timestamp 1654712443
transform 1 0 293200 0 1 -216300
box 3640 -2860 6960 460
use pixel  pixel_7201
timestamp 1654712443
transform 1 0 -800 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7200
timestamp 1654712443
transform 1 0 -3800 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7202
timestamp 1654712443
transform 1 0 2200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7203
timestamp 1654712443
transform 1 0 5200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7204
timestamp 1654712443
transform 1 0 8200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7205
timestamp 1654712443
transform 1 0 11200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7206
timestamp 1654712443
transform 1 0 14200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7207
timestamp 1654712443
transform 1 0 17200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7208
timestamp 1654712443
transform 1 0 20200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7209
timestamp 1654712443
transform 1 0 23200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7211
timestamp 1654712443
transform 1 0 29200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7210
timestamp 1654712443
transform 1 0 26200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7212
timestamp 1654712443
transform 1 0 32200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7213
timestamp 1654712443
transform 1 0 35200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7214
timestamp 1654712443
transform 1 0 38200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7215
timestamp 1654712443
transform 1 0 41200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7216
timestamp 1654712443
transform 1 0 44200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7217
timestamp 1654712443
transform 1 0 47200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7218
timestamp 1654712443
transform 1 0 50200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7219
timestamp 1654712443
transform 1 0 53200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7221
timestamp 1654712443
transform 1 0 59200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7220
timestamp 1654712443
transform 1 0 56200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7222
timestamp 1654712443
transform 1 0 62200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7223
timestamp 1654712443
transform 1 0 65200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7224
timestamp 1654712443
transform 1 0 68200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7225
timestamp 1654712443
transform 1 0 71200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7226
timestamp 1654712443
transform 1 0 74200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7227
timestamp 1654712443
transform 1 0 77200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7228
timestamp 1654712443
transform 1 0 80200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7229
timestamp 1654712443
transform 1 0 83200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7230
timestamp 1654712443
transform 1 0 86200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7231
timestamp 1654712443
transform 1 0 89200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7232
timestamp 1654712443
transform 1 0 92200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7233
timestamp 1654712443
transform 1 0 95200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7234
timestamp 1654712443
transform 1 0 98200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7235
timestamp 1654712443
transform 1 0 101200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7236
timestamp 1654712443
transform 1 0 104200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7237
timestamp 1654712443
transform 1 0 107200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7238
timestamp 1654712443
transform 1 0 110200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7239
timestamp 1654712443
transform 1 0 113200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7240
timestamp 1654712443
transform 1 0 116200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7241
timestamp 1654712443
transform 1 0 119200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7242
timestamp 1654712443
transform 1 0 122200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7243
timestamp 1654712443
transform 1 0 125200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7244
timestamp 1654712443
transform 1 0 128200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7245
timestamp 1654712443
transform 1 0 131200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7246
timestamp 1654712443
transform 1 0 134200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7247
timestamp 1654712443
transform 1 0 137200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7248
timestamp 1654712443
transform 1 0 140200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7249
timestamp 1654712443
transform 1 0 143200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7250
timestamp 1654712443
transform 1 0 146200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7251
timestamp 1654712443
transform 1 0 149200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7252
timestamp 1654712443
transform 1 0 152200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7253
timestamp 1654712443
transform 1 0 155200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7254
timestamp 1654712443
transform 1 0 158200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7255
timestamp 1654712443
transform 1 0 161200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7256
timestamp 1654712443
transform 1 0 164200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7257
timestamp 1654712443
transform 1 0 167200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7258
timestamp 1654712443
transform 1 0 170200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7259
timestamp 1654712443
transform 1 0 173200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7260
timestamp 1654712443
transform 1 0 176200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7261
timestamp 1654712443
transform 1 0 179200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7263
timestamp 1654712443
transform 1 0 185200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7262
timestamp 1654712443
transform 1 0 182200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7264
timestamp 1654712443
transform 1 0 188200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7265
timestamp 1654712443
transform 1 0 191200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7266
timestamp 1654712443
transform 1 0 194200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7267
timestamp 1654712443
transform 1 0 197200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7268
timestamp 1654712443
transform 1 0 200200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7269
timestamp 1654712443
transform 1 0 203200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7270
timestamp 1654712443
transform 1 0 206200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7271
timestamp 1654712443
transform 1 0 209200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7273
timestamp 1654712443
transform 1 0 215200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7272
timestamp 1654712443
transform 1 0 212200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7274
timestamp 1654712443
transform 1 0 218200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7275
timestamp 1654712443
transform 1 0 221200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7276
timestamp 1654712443
transform 1 0 224200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7277
timestamp 1654712443
transform 1 0 227200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7278
timestamp 1654712443
transform 1 0 230200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7279
timestamp 1654712443
transform 1 0 233200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7280
timestamp 1654712443
transform 1 0 236200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7281
timestamp 1654712443
transform 1 0 239200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7283
timestamp 1654712443
transform 1 0 245200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7282
timestamp 1654712443
transform 1 0 242200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7284
timestamp 1654712443
transform 1 0 248200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7285
timestamp 1654712443
transform 1 0 251200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7286
timestamp 1654712443
transform 1 0 254200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7287
timestamp 1654712443
transform 1 0 257200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7288
timestamp 1654712443
transform 1 0 260200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7289
timestamp 1654712443
transform 1 0 263200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7290
timestamp 1654712443
transform 1 0 266200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7291
timestamp 1654712443
transform 1 0 269200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7292
timestamp 1654712443
transform 1 0 272200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7294
timestamp 1654712443
transform 1 0 278200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7293
timestamp 1654712443
transform 1 0 275200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7295
timestamp 1654712443
transform 1 0 281200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7296
timestamp 1654712443
transform 1 0 284200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7297
timestamp 1654712443
transform 1 0 287200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7298
timestamp 1654712443
transform 1 0 290200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7299
timestamp 1654712443
transform 1 0 293200 0 1 -213300
box 3640 -2860 6960 460
use pixel  pixel_7101
timestamp 1654712443
transform 1 0 -800 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7100
timestamp 1654712443
transform 1 0 -3800 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7102
timestamp 1654712443
transform 1 0 2200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7103
timestamp 1654712443
transform 1 0 5200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7104
timestamp 1654712443
transform 1 0 8200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7105
timestamp 1654712443
transform 1 0 11200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7106
timestamp 1654712443
transform 1 0 14200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7107
timestamp 1654712443
transform 1 0 17200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7108
timestamp 1654712443
transform 1 0 20200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7109
timestamp 1654712443
transform 1 0 23200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7111
timestamp 1654712443
transform 1 0 29200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7110
timestamp 1654712443
transform 1 0 26200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7112
timestamp 1654712443
transform 1 0 32200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7113
timestamp 1654712443
transform 1 0 35200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7114
timestamp 1654712443
transform 1 0 38200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7115
timestamp 1654712443
transform 1 0 41200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7116
timestamp 1654712443
transform 1 0 44200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7117
timestamp 1654712443
transform 1 0 47200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7118
timestamp 1654712443
transform 1 0 50200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7119
timestamp 1654712443
transform 1 0 53200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7121
timestamp 1654712443
transform 1 0 59200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7120
timestamp 1654712443
transform 1 0 56200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7122
timestamp 1654712443
transform 1 0 62200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7123
timestamp 1654712443
transform 1 0 65200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7124
timestamp 1654712443
transform 1 0 68200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7125
timestamp 1654712443
transform 1 0 71200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7126
timestamp 1654712443
transform 1 0 74200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7127
timestamp 1654712443
transform 1 0 77200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7128
timestamp 1654712443
transform 1 0 80200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7129
timestamp 1654712443
transform 1 0 83200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7130
timestamp 1654712443
transform 1 0 86200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7131
timestamp 1654712443
transform 1 0 89200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7132
timestamp 1654712443
transform 1 0 92200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7133
timestamp 1654712443
transform 1 0 95200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7134
timestamp 1654712443
transform 1 0 98200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7135
timestamp 1654712443
transform 1 0 101200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7136
timestamp 1654712443
transform 1 0 104200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7137
timestamp 1654712443
transform 1 0 107200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7138
timestamp 1654712443
transform 1 0 110200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7139
timestamp 1654712443
transform 1 0 113200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7140
timestamp 1654712443
transform 1 0 116200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7141
timestamp 1654712443
transform 1 0 119200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7142
timestamp 1654712443
transform 1 0 122200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7143
timestamp 1654712443
transform 1 0 125200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7144
timestamp 1654712443
transform 1 0 128200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7145
timestamp 1654712443
transform 1 0 131200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7146
timestamp 1654712443
transform 1 0 134200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7147
timestamp 1654712443
transform 1 0 137200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7148
timestamp 1654712443
transform 1 0 140200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7149
timestamp 1654712443
transform 1 0 143200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7150
timestamp 1654712443
transform 1 0 146200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7151
timestamp 1654712443
transform 1 0 149200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7152
timestamp 1654712443
transform 1 0 152200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7153
timestamp 1654712443
transform 1 0 155200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7154
timestamp 1654712443
transform 1 0 158200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7155
timestamp 1654712443
transform 1 0 161200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7156
timestamp 1654712443
transform 1 0 164200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7157
timestamp 1654712443
transform 1 0 167200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7158
timestamp 1654712443
transform 1 0 170200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7159
timestamp 1654712443
transform 1 0 173200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7160
timestamp 1654712443
transform 1 0 176200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7161
timestamp 1654712443
transform 1 0 179200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7163
timestamp 1654712443
transform 1 0 185200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7162
timestamp 1654712443
transform 1 0 182200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7164
timestamp 1654712443
transform 1 0 188200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7165
timestamp 1654712443
transform 1 0 191200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7166
timestamp 1654712443
transform 1 0 194200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7167
timestamp 1654712443
transform 1 0 197200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7168
timestamp 1654712443
transform 1 0 200200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7169
timestamp 1654712443
transform 1 0 203200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7170
timestamp 1654712443
transform 1 0 206200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7171
timestamp 1654712443
transform 1 0 209200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7173
timestamp 1654712443
transform 1 0 215200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7172
timestamp 1654712443
transform 1 0 212200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7174
timestamp 1654712443
transform 1 0 218200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7175
timestamp 1654712443
transform 1 0 221200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7176
timestamp 1654712443
transform 1 0 224200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7177
timestamp 1654712443
transform 1 0 227200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7178
timestamp 1654712443
transform 1 0 230200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7179
timestamp 1654712443
transform 1 0 233200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7180
timestamp 1654712443
transform 1 0 236200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7181
timestamp 1654712443
transform 1 0 239200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7183
timestamp 1654712443
transform 1 0 245200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7182
timestamp 1654712443
transform 1 0 242200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7184
timestamp 1654712443
transform 1 0 248200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7185
timestamp 1654712443
transform 1 0 251200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7186
timestamp 1654712443
transform 1 0 254200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7187
timestamp 1654712443
transform 1 0 257200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7188
timestamp 1654712443
transform 1 0 260200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7189
timestamp 1654712443
transform 1 0 263200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7190
timestamp 1654712443
transform 1 0 266200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7191
timestamp 1654712443
transform 1 0 269200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7192
timestamp 1654712443
transform 1 0 272200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7194
timestamp 1654712443
transform 1 0 278200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7193
timestamp 1654712443
transform 1 0 275200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7195
timestamp 1654712443
transform 1 0 281200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7196
timestamp 1654712443
transform 1 0 284200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7197
timestamp 1654712443
transform 1 0 287200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7198
timestamp 1654712443
transform 1 0 290200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7199
timestamp 1654712443
transform 1 0 293200 0 1 -210300
box 3640 -2860 6960 460
use pixel  pixel_7001
timestamp 1654712443
transform 1 0 -800 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7000
timestamp 1654712443
transform 1 0 -3800 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7002
timestamp 1654712443
transform 1 0 2200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7003
timestamp 1654712443
transform 1 0 5200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7004
timestamp 1654712443
transform 1 0 8200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7005
timestamp 1654712443
transform 1 0 11200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7006
timestamp 1654712443
transform 1 0 14200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7007
timestamp 1654712443
transform 1 0 17200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7008
timestamp 1654712443
transform 1 0 20200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7009
timestamp 1654712443
transform 1 0 23200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7011
timestamp 1654712443
transform 1 0 29200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7010
timestamp 1654712443
transform 1 0 26200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7012
timestamp 1654712443
transform 1 0 32200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7013
timestamp 1654712443
transform 1 0 35200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7014
timestamp 1654712443
transform 1 0 38200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7015
timestamp 1654712443
transform 1 0 41200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7016
timestamp 1654712443
transform 1 0 44200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7017
timestamp 1654712443
transform 1 0 47200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7018
timestamp 1654712443
transform 1 0 50200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7019
timestamp 1654712443
transform 1 0 53200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7021
timestamp 1654712443
transform 1 0 59200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7020
timestamp 1654712443
transform 1 0 56200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7022
timestamp 1654712443
transform 1 0 62200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7023
timestamp 1654712443
transform 1 0 65200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7024
timestamp 1654712443
transform 1 0 68200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7025
timestamp 1654712443
transform 1 0 71200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7026
timestamp 1654712443
transform 1 0 74200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7027
timestamp 1654712443
transform 1 0 77200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7028
timestamp 1654712443
transform 1 0 80200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7029
timestamp 1654712443
transform 1 0 83200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7030
timestamp 1654712443
transform 1 0 86200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7031
timestamp 1654712443
transform 1 0 89200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7032
timestamp 1654712443
transform 1 0 92200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7033
timestamp 1654712443
transform 1 0 95200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7034
timestamp 1654712443
transform 1 0 98200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7035
timestamp 1654712443
transform 1 0 101200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7036
timestamp 1654712443
transform 1 0 104200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7037
timestamp 1654712443
transform 1 0 107200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7038
timestamp 1654712443
transform 1 0 110200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7039
timestamp 1654712443
transform 1 0 113200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7040
timestamp 1654712443
transform 1 0 116200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7041
timestamp 1654712443
transform 1 0 119200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7042
timestamp 1654712443
transform 1 0 122200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7043
timestamp 1654712443
transform 1 0 125200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7044
timestamp 1654712443
transform 1 0 128200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7045
timestamp 1654712443
transform 1 0 131200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7046
timestamp 1654712443
transform 1 0 134200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7047
timestamp 1654712443
transform 1 0 137200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7048
timestamp 1654712443
transform 1 0 140200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7049
timestamp 1654712443
transform 1 0 143200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7050
timestamp 1654712443
transform 1 0 146200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7051
timestamp 1654712443
transform 1 0 149200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7052
timestamp 1654712443
transform 1 0 152200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7053
timestamp 1654712443
transform 1 0 155200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7054
timestamp 1654712443
transform 1 0 158200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7055
timestamp 1654712443
transform 1 0 161200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7056
timestamp 1654712443
transform 1 0 164200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7057
timestamp 1654712443
transform 1 0 167200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7058
timestamp 1654712443
transform 1 0 170200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7059
timestamp 1654712443
transform 1 0 173200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7060
timestamp 1654712443
transform 1 0 176200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7061
timestamp 1654712443
transform 1 0 179200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7063
timestamp 1654712443
transform 1 0 185200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7062
timestamp 1654712443
transform 1 0 182200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7064
timestamp 1654712443
transform 1 0 188200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7065
timestamp 1654712443
transform 1 0 191200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7066
timestamp 1654712443
transform 1 0 194200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7067
timestamp 1654712443
transform 1 0 197200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7068
timestamp 1654712443
transform 1 0 200200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7069
timestamp 1654712443
transform 1 0 203200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7070
timestamp 1654712443
transform 1 0 206200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7071
timestamp 1654712443
transform 1 0 209200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7073
timestamp 1654712443
transform 1 0 215200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7072
timestamp 1654712443
transform 1 0 212200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7074
timestamp 1654712443
transform 1 0 218200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7075
timestamp 1654712443
transform 1 0 221200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7076
timestamp 1654712443
transform 1 0 224200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7077
timestamp 1654712443
transform 1 0 227200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7078
timestamp 1654712443
transform 1 0 230200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7079
timestamp 1654712443
transform 1 0 233200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7080
timestamp 1654712443
transform 1 0 236200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7081
timestamp 1654712443
transform 1 0 239200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7083
timestamp 1654712443
transform 1 0 245200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7082
timestamp 1654712443
transform 1 0 242200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7084
timestamp 1654712443
transform 1 0 248200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7085
timestamp 1654712443
transform 1 0 251200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7086
timestamp 1654712443
transform 1 0 254200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7087
timestamp 1654712443
transform 1 0 257200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7088
timestamp 1654712443
transform 1 0 260200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7089
timestamp 1654712443
transform 1 0 263200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7090
timestamp 1654712443
transform 1 0 266200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7091
timestamp 1654712443
transform 1 0 269200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7092
timestamp 1654712443
transform 1 0 272200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7094
timestamp 1654712443
transform 1 0 278200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7093
timestamp 1654712443
transform 1 0 275200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7095
timestamp 1654712443
transform 1 0 281200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7096
timestamp 1654712443
transform 1 0 284200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7097
timestamp 1654712443
transform 1 0 287200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7098
timestamp 1654712443
transform 1 0 290200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_7099
timestamp 1654712443
transform 1 0 293200 0 1 -207300
box 3640 -2860 6960 460
use pixel  pixel_6901
timestamp 1654712443
transform 1 0 -800 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6900
timestamp 1654712443
transform 1 0 -3800 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6902
timestamp 1654712443
transform 1 0 2200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6903
timestamp 1654712443
transform 1 0 5200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6904
timestamp 1654712443
transform 1 0 8200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6905
timestamp 1654712443
transform 1 0 11200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6906
timestamp 1654712443
transform 1 0 14200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6907
timestamp 1654712443
transform 1 0 17200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6908
timestamp 1654712443
transform 1 0 20200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6909
timestamp 1654712443
transform 1 0 23200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6911
timestamp 1654712443
transform 1 0 29200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6910
timestamp 1654712443
transform 1 0 26200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6912
timestamp 1654712443
transform 1 0 32200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6913
timestamp 1654712443
transform 1 0 35200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6914
timestamp 1654712443
transform 1 0 38200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6915
timestamp 1654712443
transform 1 0 41200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6916
timestamp 1654712443
transform 1 0 44200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6917
timestamp 1654712443
transform 1 0 47200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6918
timestamp 1654712443
transform 1 0 50200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6919
timestamp 1654712443
transform 1 0 53200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6921
timestamp 1654712443
transform 1 0 59200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6920
timestamp 1654712443
transform 1 0 56200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6922
timestamp 1654712443
transform 1 0 62200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6923
timestamp 1654712443
transform 1 0 65200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6924
timestamp 1654712443
transform 1 0 68200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6925
timestamp 1654712443
transform 1 0 71200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6926
timestamp 1654712443
transform 1 0 74200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6927
timestamp 1654712443
transform 1 0 77200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6928
timestamp 1654712443
transform 1 0 80200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6929
timestamp 1654712443
transform 1 0 83200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6930
timestamp 1654712443
transform 1 0 86200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6931
timestamp 1654712443
transform 1 0 89200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6932
timestamp 1654712443
transform 1 0 92200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6933
timestamp 1654712443
transform 1 0 95200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6934
timestamp 1654712443
transform 1 0 98200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6935
timestamp 1654712443
transform 1 0 101200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6936
timestamp 1654712443
transform 1 0 104200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6937
timestamp 1654712443
transform 1 0 107200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6938
timestamp 1654712443
transform 1 0 110200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6939
timestamp 1654712443
transform 1 0 113200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6940
timestamp 1654712443
transform 1 0 116200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6941
timestamp 1654712443
transform 1 0 119200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6942
timestamp 1654712443
transform 1 0 122200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6943
timestamp 1654712443
transform 1 0 125200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6944
timestamp 1654712443
transform 1 0 128200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6945
timestamp 1654712443
transform 1 0 131200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6946
timestamp 1654712443
transform 1 0 134200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6947
timestamp 1654712443
transform 1 0 137200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6948
timestamp 1654712443
transform 1 0 140200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6949
timestamp 1654712443
transform 1 0 143200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6950
timestamp 1654712443
transform 1 0 146200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6951
timestamp 1654712443
transform 1 0 149200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6952
timestamp 1654712443
transform 1 0 152200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6953
timestamp 1654712443
transform 1 0 155200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6954
timestamp 1654712443
transform 1 0 158200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6955
timestamp 1654712443
transform 1 0 161200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6956
timestamp 1654712443
transform 1 0 164200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6957
timestamp 1654712443
transform 1 0 167200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6958
timestamp 1654712443
transform 1 0 170200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6959
timestamp 1654712443
transform 1 0 173200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6960
timestamp 1654712443
transform 1 0 176200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6961
timestamp 1654712443
transform 1 0 179200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6963
timestamp 1654712443
transform 1 0 185200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6962
timestamp 1654712443
transform 1 0 182200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6964
timestamp 1654712443
transform 1 0 188200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6965
timestamp 1654712443
transform 1 0 191200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6966
timestamp 1654712443
transform 1 0 194200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6967
timestamp 1654712443
transform 1 0 197200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6968
timestamp 1654712443
transform 1 0 200200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6969
timestamp 1654712443
transform 1 0 203200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6970
timestamp 1654712443
transform 1 0 206200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6971
timestamp 1654712443
transform 1 0 209200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6973
timestamp 1654712443
transform 1 0 215200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6972
timestamp 1654712443
transform 1 0 212200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6974
timestamp 1654712443
transform 1 0 218200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6975
timestamp 1654712443
transform 1 0 221200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6976
timestamp 1654712443
transform 1 0 224200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6977
timestamp 1654712443
transform 1 0 227200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6978
timestamp 1654712443
transform 1 0 230200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6979
timestamp 1654712443
transform 1 0 233200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6980
timestamp 1654712443
transform 1 0 236200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6981
timestamp 1654712443
transform 1 0 239200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6983
timestamp 1654712443
transform 1 0 245200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6982
timestamp 1654712443
transform 1 0 242200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6984
timestamp 1654712443
transform 1 0 248200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6985
timestamp 1654712443
transform 1 0 251200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6986
timestamp 1654712443
transform 1 0 254200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6987
timestamp 1654712443
transform 1 0 257200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6988
timestamp 1654712443
transform 1 0 260200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6989
timestamp 1654712443
transform 1 0 263200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6990
timestamp 1654712443
transform 1 0 266200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6991
timestamp 1654712443
transform 1 0 269200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6992
timestamp 1654712443
transform 1 0 272200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6994
timestamp 1654712443
transform 1 0 278200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6993
timestamp 1654712443
transform 1 0 275200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6995
timestamp 1654712443
transform 1 0 281200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6996
timestamp 1654712443
transform 1 0 284200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6997
timestamp 1654712443
transform 1 0 287200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6998
timestamp 1654712443
transform 1 0 290200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6999
timestamp 1654712443
transform 1 0 293200 0 1 -204300
box 3640 -2860 6960 460
use pixel  pixel_6701
timestamp 1654712443
transform 1 0 -800 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6801
timestamp 1654712443
transform 1 0 -800 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6700
timestamp 1654712443
transform 1 0 -3800 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6800
timestamp 1654712443
transform 1 0 -3800 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6702
timestamp 1654712443
transform 1 0 2200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6802
timestamp 1654712443
transform 1 0 2200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6703
timestamp 1654712443
transform 1 0 5200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6803
timestamp 1654712443
transform 1 0 5200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6704
timestamp 1654712443
transform 1 0 8200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6804
timestamp 1654712443
transform 1 0 8200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6705
timestamp 1654712443
transform 1 0 11200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6805
timestamp 1654712443
transform 1 0 11200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6706
timestamp 1654712443
transform 1 0 14200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6806
timestamp 1654712443
transform 1 0 14200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6707
timestamp 1654712443
transform 1 0 17200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6807
timestamp 1654712443
transform 1 0 17200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6708
timestamp 1654712443
transform 1 0 20200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6808
timestamp 1654712443
transform 1 0 20200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6709
timestamp 1654712443
transform 1 0 23200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6809
timestamp 1654712443
transform 1 0 23200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6711
timestamp 1654712443
transform 1 0 29200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6811
timestamp 1654712443
transform 1 0 29200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6710
timestamp 1654712443
transform 1 0 26200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6810
timestamp 1654712443
transform 1 0 26200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6712
timestamp 1654712443
transform 1 0 32200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6812
timestamp 1654712443
transform 1 0 32200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6713
timestamp 1654712443
transform 1 0 35200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6813
timestamp 1654712443
transform 1 0 35200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6714
timestamp 1654712443
transform 1 0 38200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6814
timestamp 1654712443
transform 1 0 38200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6715
timestamp 1654712443
transform 1 0 41200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6815
timestamp 1654712443
transform 1 0 41200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6716
timestamp 1654712443
transform 1 0 44200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6816
timestamp 1654712443
transform 1 0 44200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6717
timestamp 1654712443
transform 1 0 47200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6817
timestamp 1654712443
transform 1 0 47200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6718
timestamp 1654712443
transform 1 0 50200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6818
timestamp 1654712443
transform 1 0 50200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6719
timestamp 1654712443
transform 1 0 53200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6819
timestamp 1654712443
transform 1 0 53200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6721
timestamp 1654712443
transform 1 0 59200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6821
timestamp 1654712443
transform 1 0 59200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6720
timestamp 1654712443
transform 1 0 56200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6820
timestamp 1654712443
transform 1 0 56200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6722
timestamp 1654712443
transform 1 0 62200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6822
timestamp 1654712443
transform 1 0 62200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6723
timestamp 1654712443
transform 1 0 65200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6823
timestamp 1654712443
transform 1 0 65200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6724
timestamp 1654712443
transform 1 0 68200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6824
timestamp 1654712443
transform 1 0 68200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6725
timestamp 1654712443
transform 1 0 71200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6825
timestamp 1654712443
transform 1 0 71200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6726
timestamp 1654712443
transform 1 0 74200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6826
timestamp 1654712443
transform 1 0 74200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6727
timestamp 1654712443
transform 1 0 77200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6827
timestamp 1654712443
transform 1 0 77200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6728
timestamp 1654712443
transform 1 0 80200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6828
timestamp 1654712443
transform 1 0 80200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6729
timestamp 1654712443
transform 1 0 83200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6829
timestamp 1654712443
transform 1 0 83200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6730
timestamp 1654712443
transform 1 0 86200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6830
timestamp 1654712443
transform 1 0 86200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6731
timestamp 1654712443
transform 1 0 89200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6732
timestamp 1654712443
transform 1 0 92200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6831
timestamp 1654712443
transform 1 0 89200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6832
timestamp 1654712443
transform 1 0 92200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6733
timestamp 1654712443
transform 1 0 95200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6833
timestamp 1654712443
transform 1 0 95200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6734
timestamp 1654712443
transform 1 0 98200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6834
timestamp 1654712443
transform 1 0 98200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6735
timestamp 1654712443
transform 1 0 101200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6835
timestamp 1654712443
transform 1 0 101200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6736
timestamp 1654712443
transform 1 0 104200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6836
timestamp 1654712443
transform 1 0 104200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6737
timestamp 1654712443
transform 1 0 107200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6837
timestamp 1654712443
transform 1 0 107200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6738
timestamp 1654712443
transform 1 0 110200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6838
timestamp 1654712443
transform 1 0 110200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6739
timestamp 1654712443
transform 1 0 113200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6839
timestamp 1654712443
transform 1 0 113200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6740
timestamp 1654712443
transform 1 0 116200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6840
timestamp 1654712443
transform 1 0 116200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6741
timestamp 1654712443
transform 1 0 119200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6742
timestamp 1654712443
transform 1 0 122200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6841
timestamp 1654712443
transform 1 0 119200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6842
timestamp 1654712443
transform 1 0 122200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6743
timestamp 1654712443
transform 1 0 125200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6843
timestamp 1654712443
transform 1 0 125200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6744
timestamp 1654712443
transform 1 0 128200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6844
timestamp 1654712443
transform 1 0 128200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6745
timestamp 1654712443
transform 1 0 131200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6845
timestamp 1654712443
transform 1 0 131200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6746
timestamp 1654712443
transform 1 0 134200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6846
timestamp 1654712443
transform 1 0 134200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6747
timestamp 1654712443
transform 1 0 137200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6847
timestamp 1654712443
transform 1 0 137200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6748
timestamp 1654712443
transform 1 0 140200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6848
timestamp 1654712443
transform 1 0 140200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6749
timestamp 1654712443
transform 1 0 143200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6849
timestamp 1654712443
transform 1 0 143200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6750
timestamp 1654712443
transform 1 0 146200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6850
timestamp 1654712443
transform 1 0 146200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6751
timestamp 1654712443
transform 1 0 149200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6752
timestamp 1654712443
transform 1 0 152200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6851
timestamp 1654712443
transform 1 0 149200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6852
timestamp 1654712443
transform 1 0 152200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6753
timestamp 1654712443
transform 1 0 155200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6853
timestamp 1654712443
transform 1 0 155200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6754
timestamp 1654712443
transform 1 0 158200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6854
timestamp 1654712443
transform 1 0 158200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6755
timestamp 1654712443
transform 1 0 161200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6855
timestamp 1654712443
transform 1 0 161200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6756
timestamp 1654712443
transform 1 0 164200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6856
timestamp 1654712443
transform 1 0 164200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6757
timestamp 1654712443
transform 1 0 167200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6857
timestamp 1654712443
transform 1 0 167200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6758
timestamp 1654712443
transform 1 0 170200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6858
timestamp 1654712443
transform 1 0 170200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6759
timestamp 1654712443
transform 1 0 173200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6859
timestamp 1654712443
transform 1 0 173200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6760
timestamp 1654712443
transform 1 0 176200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6860
timestamp 1654712443
transform 1 0 176200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6761
timestamp 1654712443
transform 1 0 179200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6861
timestamp 1654712443
transform 1 0 179200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6763
timestamp 1654712443
transform 1 0 185200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6863
timestamp 1654712443
transform 1 0 185200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6762
timestamp 1654712443
transform 1 0 182200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6862
timestamp 1654712443
transform 1 0 182200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6764
timestamp 1654712443
transform 1 0 188200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6864
timestamp 1654712443
transform 1 0 188200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6765
timestamp 1654712443
transform 1 0 191200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6865
timestamp 1654712443
transform 1 0 191200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6766
timestamp 1654712443
transform 1 0 194200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6866
timestamp 1654712443
transform 1 0 194200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6767
timestamp 1654712443
transform 1 0 197200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6867
timestamp 1654712443
transform 1 0 197200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6768
timestamp 1654712443
transform 1 0 200200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6868
timestamp 1654712443
transform 1 0 200200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6769
timestamp 1654712443
transform 1 0 203200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6869
timestamp 1654712443
transform 1 0 203200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6770
timestamp 1654712443
transform 1 0 206200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6870
timestamp 1654712443
transform 1 0 206200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6771
timestamp 1654712443
transform 1 0 209200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6871
timestamp 1654712443
transform 1 0 209200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6773
timestamp 1654712443
transform 1 0 215200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6873
timestamp 1654712443
transform 1 0 215200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6772
timestamp 1654712443
transform 1 0 212200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6872
timestamp 1654712443
transform 1 0 212200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6774
timestamp 1654712443
transform 1 0 218200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6874
timestamp 1654712443
transform 1 0 218200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6775
timestamp 1654712443
transform 1 0 221200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6875
timestamp 1654712443
transform 1 0 221200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6776
timestamp 1654712443
transform 1 0 224200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6876
timestamp 1654712443
transform 1 0 224200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6777
timestamp 1654712443
transform 1 0 227200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6877
timestamp 1654712443
transform 1 0 227200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6778
timestamp 1654712443
transform 1 0 230200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6878
timestamp 1654712443
transform 1 0 230200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6779
timestamp 1654712443
transform 1 0 233200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6879
timestamp 1654712443
transform 1 0 233200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6780
timestamp 1654712443
transform 1 0 236200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6880
timestamp 1654712443
transform 1 0 236200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6781
timestamp 1654712443
transform 1 0 239200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6881
timestamp 1654712443
transform 1 0 239200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6783
timestamp 1654712443
transform 1 0 245200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6883
timestamp 1654712443
transform 1 0 245200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6782
timestamp 1654712443
transform 1 0 242200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6882
timestamp 1654712443
transform 1 0 242200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6784
timestamp 1654712443
transform 1 0 248200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6884
timestamp 1654712443
transform 1 0 248200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6785
timestamp 1654712443
transform 1 0 251200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6885
timestamp 1654712443
transform 1 0 251200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6786
timestamp 1654712443
transform 1 0 254200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6886
timestamp 1654712443
transform 1 0 254200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6787
timestamp 1654712443
transform 1 0 257200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6887
timestamp 1654712443
transform 1 0 257200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6788
timestamp 1654712443
transform 1 0 260200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6888
timestamp 1654712443
transform 1 0 260200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6789
timestamp 1654712443
transform 1 0 263200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6889
timestamp 1654712443
transform 1 0 263200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6790
timestamp 1654712443
transform 1 0 266200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6890
timestamp 1654712443
transform 1 0 266200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6791
timestamp 1654712443
transform 1 0 269200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6891
timestamp 1654712443
transform 1 0 269200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6792
timestamp 1654712443
transform 1 0 272200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6892
timestamp 1654712443
transform 1 0 272200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6794
timestamp 1654712443
transform 1 0 278200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6894
timestamp 1654712443
transform 1 0 278200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6793
timestamp 1654712443
transform 1 0 275200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6893
timestamp 1654712443
transform 1 0 275200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6795
timestamp 1654712443
transform 1 0 281200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6895
timestamp 1654712443
transform 1 0 281200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6796
timestamp 1654712443
transform 1 0 284200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6896
timestamp 1654712443
transform 1 0 284200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6797
timestamp 1654712443
transform 1 0 287200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6897
timestamp 1654712443
transform 1 0 287200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6798
timestamp 1654712443
transform 1 0 290200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6898
timestamp 1654712443
transform 1 0 290200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6799
timestamp 1654712443
transform 1 0 293200 0 1 -198300
box 3640 -2860 6960 460
use pixel  pixel_6899
timestamp 1654712443
transform 1 0 293200 0 1 -201300
box 3640 -2860 6960 460
use pixel  pixel_6601
timestamp 1654712443
transform 1 0 -800 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6600
timestamp 1654712443
transform 1 0 -3800 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6602
timestamp 1654712443
transform 1 0 2200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6603
timestamp 1654712443
transform 1 0 5200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6604
timestamp 1654712443
transform 1 0 8200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6605
timestamp 1654712443
transform 1 0 11200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6606
timestamp 1654712443
transform 1 0 14200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6607
timestamp 1654712443
transform 1 0 17200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6608
timestamp 1654712443
transform 1 0 20200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6609
timestamp 1654712443
transform 1 0 23200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6611
timestamp 1654712443
transform 1 0 29200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6610
timestamp 1654712443
transform 1 0 26200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6612
timestamp 1654712443
transform 1 0 32200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6613
timestamp 1654712443
transform 1 0 35200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6614
timestamp 1654712443
transform 1 0 38200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6615
timestamp 1654712443
transform 1 0 41200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6616
timestamp 1654712443
transform 1 0 44200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6617
timestamp 1654712443
transform 1 0 47200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6618
timestamp 1654712443
transform 1 0 50200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6619
timestamp 1654712443
transform 1 0 53200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6621
timestamp 1654712443
transform 1 0 59200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6620
timestamp 1654712443
transform 1 0 56200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6622
timestamp 1654712443
transform 1 0 62200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6623
timestamp 1654712443
transform 1 0 65200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6624
timestamp 1654712443
transform 1 0 68200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6625
timestamp 1654712443
transform 1 0 71200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6626
timestamp 1654712443
transform 1 0 74200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6627
timestamp 1654712443
transform 1 0 77200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6628
timestamp 1654712443
transform 1 0 80200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6629
timestamp 1654712443
transform 1 0 83200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6630
timestamp 1654712443
transform 1 0 86200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6631
timestamp 1654712443
transform 1 0 89200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6632
timestamp 1654712443
transform 1 0 92200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6633
timestamp 1654712443
transform 1 0 95200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6634
timestamp 1654712443
transform 1 0 98200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6635
timestamp 1654712443
transform 1 0 101200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6636
timestamp 1654712443
transform 1 0 104200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6637
timestamp 1654712443
transform 1 0 107200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6638
timestamp 1654712443
transform 1 0 110200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6639
timestamp 1654712443
transform 1 0 113200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6640
timestamp 1654712443
transform 1 0 116200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6641
timestamp 1654712443
transform 1 0 119200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6642
timestamp 1654712443
transform 1 0 122200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6643
timestamp 1654712443
transform 1 0 125200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6644
timestamp 1654712443
transform 1 0 128200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6645
timestamp 1654712443
transform 1 0 131200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6646
timestamp 1654712443
transform 1 0 134200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6647
timestamp 1654712443
transform 1 0 137200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6648
timestamp 1654712443
transform 1 0 140200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6649
timestamp 1654712443
transform 1 0 143200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6650
timestamp 1654712443
transform 1 0 146200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6651
timestamp 1654712443
transform 1 0 149200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6652
timestamp 1654712443
transform 1 0 152200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6653
timestamp 1654712443
transform 1 0 155200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6654
timestamp 1654712443
transform 1 0 158200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6655
timestamp 1654712443
transform 1 0 161200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6656
timestamp 1654712443
transform 1 0 164200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6657
timestamp 1654712443
transform 1 0 167200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6658
timestamp 1654712443
transform 1 0 170200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6659
timestamp 1654712443
transform 1 0 173200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6660
timestamp 1654712443
transform 1 0 176200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6661
timestamp 1654712443
transform 1 0 179200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6663
timestamp 1654712443
transform 1 0 185200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6662
timestamp 1654712443
transform 1 0 182200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6664
timestamp 1654712443
transform 1 0 188200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6665
timestamp 1654712443
transform 1 0 191200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6666
timestamp 1654712443
transform 1 0 194200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6667
timestamp 1654712443
transform 1 0 197200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6668
timestamp 1654712443
transform 1 0 200200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6669
timestamp 1654712443
transform 1 0 203200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6670
timestamp 1654712443
transform 1 0 206200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6671
timestamp 1654712443
transform 1 0 209200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6673
timestamp 1654712443
transform 1 0 215200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6672
timestamp 1654712443
transform 1 0 212200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6674
timestamp 1654712443
transform 1 0 218200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6675
timestamp 1654712443
transform 1 0 221200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6676
timestamp 1654712443
transform 1 0 224200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6677
timestamp 1654712443
transform 1 0 227200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6678
timestamp 1654712443
transform 1 0 230200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6679
timestamp 1654712443
transform 1 0 233200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6680
timestamp 1654712443
transform 1 0 236200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6681
timestamp 1654712443
transform 1 0 239200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6683
timestamp 1654712443
transform 1 0 245200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6682
timestamp 1654712443
transform 1 0 242200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6684
timestamp 1654712443
transform 1 0 248200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6685
timestamp 1654712443
transform 1 0 251200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6686
timestamp 1654712443
transform 1 0 254200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6687
timestamp 1654712443
transform 1 0 257200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6688
timestamp 1654712443
transform 1 0 260200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6689
timestamp 1654712443
transform 1 0 263200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6690
timestamp 1654712443
transform 1 0 266200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6691
timestamp 1654712443
transform 1 0 269200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6692
timestamp 1654712443
transform 1 0 272200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6694
timestamp 1654712443
transform 1 0 278200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6693
timestamp 1654712443
transform 1 0 275200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6695
timestamp 1654712443
transform 1 0 281200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6696
timestamp 1654712443
transform 1 0 284200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6697
timestamp 1654712443
transform 1 0 287200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6698
timestamp 1654712443
transform 1 0 290200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6699
timestamp 1654712443
transform 1 0 293200 0 1 -195300
box 3640 -2860 6960 460
use pixel  pixel_6501
timestamp 1654712443
transform 1 0 -800 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6500
timestamp 1654712443
transform 1 0 -3800 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6502
timestamp 1654712443
transform 1 0 2200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6503
timestamp 1654712443
transform 1 0 5200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6504
timestamp 1654712443
transform 1 0 8200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6505
timestamp 1654712443
transform 1 0 11200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6506
timestamp 1654712443
transform 1 0 14200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6507
timestamp 1654712443
transform 1 0 17200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6508
timestamp 1654712443
transform 1 0 20200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6509
timestamp 1654712443
transform 1 0 23200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6511
timestamp 1654712443
transform 1 0 29200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6510
timestamp 1654712443
transform 1 0 26200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6512
timestamp 1654712443
transform 1 0 32200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6513
timestamp 1654712443
transform 1 0 35200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6514
timestamp 1654712443
transform 1 0 38200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6515
timestamp 1654712443
transform 1 0 41200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6516
timestamp 1654712443
transform 1 0 44200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6517
timestamp 1654712443
transform 1 0 47200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6518
timestamp 1654712443
transform 1 0 50200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6519
timestamp 1654712443
transform 1 0 53200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6521
timestamp 1654712443
transform 1 0 59200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6520
timestamp 1654712443
transform 1 0 56200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6522
timestamp 1654712443
transform 1 0 62200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6523
timestamp 1654712443
transform 1 0 65200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6524
timestamp 1654712443
transform 1 0 68200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6525
timestamp 1654712443
transform 1 0 71200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6526
timestamp 1654712443
transform 1 0 74200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6527
timestamp 1654712443
transform 1 0 77200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6528
timestamp 1654712443
transform 1 0 80200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6529
timestamp 1654712443
transform 1 0 83200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6530
timestamp 1654712443
transform 1 0 86200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6531
timestamp 1654712443
transform 1 0 89200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6532
timestamp 1654712443
transform 1 0 92200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6533
timestamp 1654712443
transform 1 0 95200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6534
timestamp 1654712443
transform 1 0 98200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6535
timestamp 1654712443
transform 1 0 101200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6536
timestamp 1654712443
transform 1 0 104200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6537
timestamp 1654712443
transform 1 0 107200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6538
timestamp 1654712443
transform 1 0 110200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6539
timestamp 1654712443
transform 1 0 113200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6540
timestamp 1654712443
transform 1 0 116200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6541
timestamp 1654712443
transform 1 0 119200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6542
timestamp 1654712443
transform 1 0 122200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6543
timestamp 1654712443
transform 1 0 125200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6544
timestamp 1654712443
transform 1 0 128200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6545
timestamp 1654712443
transform 1 0 131200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6546
timestamp 1654712443
transform 1 0 134200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6547
timestamp 1654712443
transform 1 0 137200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6548
timestamp 1654712443
transform 1 0 140200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6549
timestamp 1654712443
transform 1 0 143200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6550
timestamp 1654712443
transform 1 0 146200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6551
timestamp 1654712443
transform 1 0 149200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6552
timestamp 1654712443
transform 1 0 152200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6553
timestamp 1654712443
transform 1 0 155200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6554
timestamp 1654712443
transform 1 0 158200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6555
timestamp 1654712443
transform 1 0 161200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6556
timestamp 1654712443
transform 1 0 164200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6557
timestamp 1654712443
transform 1 0 167200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6558
timestamp 1654712443
transform 1 0 170200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6559
timestamp 1654712443
transform 1 0 173200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6560
timestamp 1654712443
transform 1 0 176200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6561
timestamp 1654712443
transform 1 0 179200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6563
timestamp 1654712443
transform 1 0 185200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6562
timestamp 1654712443
transform 1 0 182200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6564
timestamp 1654712443
transform 1 0 188200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6565
timestamp 1654712443
transform 1 0 191200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6566
timestamp 1654712443
transform 1 0 194200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6567
timestamp 1654712443
transform 1 0 197200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6568
timestamp 1654712443
transform 1 0 200200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6569
timestamp 1654712443
transform 1 0 203200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6570
timestamp 1654712443
transform 1 0 206200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6571
timestamp 1654712443
transform 1 0 209200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6573
timestamp 1654712443
transform 1 0 215200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6572
timestamp 1654712443
transform 1 0 212200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6574
timestamp 1654712443
transform 1 0 218200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6575
timestamp 1654712443
transform 1 0 221200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6576
timestamp 1654712443
transform 1 0 224200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6577
timestamp 1654712443
transform 1 0 227200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6578
timestamp 1654712443
transform 1 0 230200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6579
timestamp 1654712443
transform 1 0 233200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6580
timestamp 1654712443
transform 1 0 236200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6581
timestamp 1654712443
transform 1 0 239200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6583
timestamp 1654712443
transform 1 0 245200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6582
timestamp 1654712443
transform 1 0 242200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6584
timestamp 1654712443
transform 1 0 248200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6585
timestamp 1654712443
transform 1 0 251200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6586
timestamp 1654712443
transform 1 0 254200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6587
timestamp 1654712443
transform 1 0 257200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6588
timestamp 1654712443
transform 1 0 260200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6589
timestamp 1654712443
transform 1 0 263200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6590
timestamp 1654712443
transform 1 0 266200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6591
timestamp 1654712443
transform 1 0 269200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6592
timestamp 1654712443
transform 1 0 272200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6594
timestamp 1654712443
transform 1 0 278200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6593
timestamp 1654712443
transform 1 0 275200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6595
timestamp 1654712443
transform 1 0 281200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6596
timestamp 1654712443
transform 1 0 284200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6597
timestamp 1654712443
transform 1 0 287200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6598
timestamp 1654712443
transform 1 0 290200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6599
timestamp 1654712443
transform 1 0 293200 0 1 -192300
box 3640 -2860 6960 460
use pixel  pixel_6401
timestamp 1654712443
transform 1 0 -800 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6400
timestamp 1654712443
transform 1 0 -3800 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6402
timestamp 1654712443
transform 1 0 2200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6403
timestamp 1654712443
transform 1 0 5200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6404
timestamp 1654712443
transform 1 0 8200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6405
timestamp 1654712443
transform 1 0 11200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6406
timestamp 1654712443
transform 1 0 14200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6407
timestamp 1654712443
transform 1 0 17200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6408
timestamp 1654712443
transform 1 0 20200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6409
timestamp 1654712443
transform 1 0 23200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6411
timestamp 1654712443
transform 1 0 29200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6410
timestamp 1654712443
transform 1 0 26200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6412
timestamp 1654712443
transform 1 0 32200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6413
timestamp 1654712443
transform 1 0 35200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6414
timestamp 1654712443
transform 1 0 38200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6415
timestamp 1654712443
transform 1 0 41200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6416
timestamp 1654712443
transform 1 0 44200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6417
timestamp 1654712443
transform 1 0 47200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6418
timestamp 1654712443
transform 1 0 50200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6419
timestamp 1654712443
transform 1 0 53200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6421
timestamp 1654712443
transform 1 0 59200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6420
timestamp 1654712443
transform 1 0 56200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6422
timestamp 1654712443
transform 1 0 62200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6423
timestamp 1654712443
transform 1 0 65200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6424
timestamp 1654712443
transform 1 0 68200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6425
timestamp 1654712443
transform 1 0 71200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6426
timestamp 1654712443
transform 1 0 74200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6427
timestamp 1654712443
transform 1 0 77200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6428
timestamp 1654712443
transform 1 0 80200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6429
timestamp 1654712443
transform 1 0 83200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6430
timestamp 1654712443
transform 1 0 86200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6431
timestamp 1654712443
transform 1 0 89200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6432
timestamp 1654712443
transform 1 0 92200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6433
timestamp 1654712443
transform 1 0 95200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6434
timestamp 1654712443
transform 1 0 98200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6435
timestamp 1654712443
transform 1 0 101200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6436
timestamp 1654712443
transform 1 0 104200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6437
timestamp 1654712443
transform 1 0 107200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6438
timestamp 1654712443
transform 1 0 110200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6439
timestamp 1654712443
transform 1 0 113200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6440
timestamp 1654712443
transform 1 0 116200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6441
timestamp 1654712443
transform 1 0 119200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6442
timestamp 1654712443
transform 1 0 122200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6443
timestamp 1654712443
transform 1 0 125200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6444
timestamp 1654712443
transform 1 0 128200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6445
timestamp 1654712443
transform 1 0 131200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6446
timestamp 1654712443
transform 1 0 134200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6447
timestamp 1654712443
transform 1 0 137200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6448
timestamp 1654712443
transform 1 0 140200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6449
timestamp 1654712443
transform 1 0 143200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6450
timestamp 1654712443
transform 1 0 146200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6451
timestamp 1654712443
transform 1 0 149200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6452
timestamp 1654712443
transform 1 0 152200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6453
timestamp 1654712443
transform 1 0 155200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6454
timestamp 1654712443
transform 1 0 158200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6455
timestamp 1654712443
transform 1 0 161200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6456
timestamp 1654712443
transform 1 0 164200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6457
timestamp 1654712443
transform 1 0 167200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6458
timestamp 1654712443
transform 1 0 170200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6459
timestamp 1654712443
transform 1 0 173200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6460
timestamp 1654712443
transform 1 0 176200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6461
timestamp 1654712443
transform 1 0 179200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6463
timestamp 1654712443
transform 1 0 185200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6462
timestamp 1654712443
transform 1 0 182200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6464
timestamp 1654712443
transform 1 0 188200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6465
timestamp 1654712443
transform 1 0 191200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6466
timestamp 1654712443
transform 1 0 194200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6467
timestamp 1654712443
transform 1 0 197200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6468
timestamp 1654712443
transform 1 0 200200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6469
timestamp 1654712443
transform 1 0 203200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6470
timestamp 1654712443
transform 1 0 206200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6471
timestamp 1654712443
transform 1 0 209200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6473
timestamp 1654712443
transform 1 0 215200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6472
timestamp 1654712443
transform 1 0 212200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6474
timestamp 1654712443
transform 1 0 218200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6475
timestamp 1654712443
transform 1 0 221200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6476
timestamp 1654712443
transform 1 0 224200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6477
timestamp 1654712443
transform 1 0 227200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6478
timestamp 1654712443
transform 1 0 230200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6479
timestamp 1654712443
transform 1 0 233200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6480
timestamp 1654712443
transform 1 0 236200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6481
timestamp 1654712443
transform 1 0 239200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6483
timestamp 1654712443
transform 1 0 245200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6482
timestamp 1654712443
transform 1 0 242200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6484
timestamp 1654712443
transform 1 0 248200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6485
timestamp 1654712443
transform 1 0 251200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6486
timestamp 1654712443
transform 1 0 254200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6487
timestamp 1654712443
transform 1 0 257200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6488
timestamp 1654712443
transform 1 0 260200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6489
timestamp 1654712443
transform 1 0 263200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6490
timestamp 1654712443
transform 1 0 266200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6491
timestamp 1654712443
transform 1 0 269200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6492
timestamp 1654712443
transform 1 0 272200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6494
timestamp 1654712443
transform 1 0 278200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6493
timestamp 1654712443
transform 1 0 275200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6495
timestamp 1654712443
transform 1 0 281200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6496
timestamp 1654712443
transform 1 0 284200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6497
timestamp 1654712443
transform 1 0 287200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6498
timestamp 1654712443
transform 1 0 290200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6499
timestamp 1654712443
transform 1 0 293200 0 1 -189300
box 3640 -2860 6960 460
use pixel  pixel_6301
timestamp 1654712443
transform 1 0 -800 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6300
timestamp 1654712443
transform 1 0 -3800 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6302
timestamp 1654712443
transform 1 0 2200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6303
timestamp 1654712443
transform 1 0 5200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6304
timestamp 1654712443
transform 1 0 8200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6305
timestamp 1654712443
transform 1 0 11200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6306
timestamp 1654712443
transform 1 0 14200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6307
timestamp 1654712443
transform 1 0 17200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6308
timestamp 1654712443
transform 1 0 20200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6309
timestamp 1654712443
transform 1 0 23200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6311
timestamp 1654712443
transform 1 0 29200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6310
timestamp 1654712443
transform 1 0 26200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6312
timestamp 1654712443
transform 1 0 32200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6313
timestamp 1654712443
transform 1 0 35200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6314
timestamp 1654712443
transform 1 0 38200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6315
timestamp 1654712443
transform 1 0 41200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6316
timestamp 1654712443
transform 1 0 44200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6317
timestamp 1654712443
transform 1 0 47200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6318
timestamp 1654712443
transform 1 0 50200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6319
timestamp 1654712443
transform 1 0 53200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6321
timestamp 1654712443
transform 1 0 59200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6320
timestamp 1654712443
transform 1 0 56200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6322
timestamp 1654712443
transform 1 0 62200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6323
timestamp 1654712443
transform 1 0 65200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6324
timestamp 1654712443
transform 1 0 68200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6325
timestamp 1654712443
transform 1 0 71200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6326
timestamp 1654712443
transform 1 0 74200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6327
timestamp 1654712443
transform 1 0 77200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6328
timestamp 1654712443
transform 1 0 80200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6329
timestamp 1654712443
transform 1 0 83200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6330
timestamp 1654712443
transform 1 0 86200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6331
timestamp 1654712443
transform 1 0 89200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6332
timestamp 1654712443
transform 1 0 92200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6333
timestamp 1654712443
transform 1 0 95200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6334
timestamp 1654712443
transform 1 0 98200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6335
timestamp 1654712443
transform 1 0 101200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6336
timestamp 1654712443
transform 1 0 104200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6337
timestamp 1654712443
transform 1 0 107200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6338
timestamp 1654712443
transform 1 0 110200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6339
timestamp 1654712443
transform 1 0 113200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6340
timestamp 1654712443
transform 1 0 116200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6341
timestamp 1654712443
transform 1 0 119200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6342
timestamp 1654712443
transform 1 0 122200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6343
timestamp 1654712443
transform 1 0 125200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6344
timestamp 1654712443
transform 1 0 128200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6345
timestamp 1654712443
transform 1 0 131200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6346
timestamp 1654712443
transform 1 0 134200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6347
timestamp 1654712443
transform 1 0 137200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6348
timestamp 1654712443
transform 1 0 140200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6349
timestamp 1654712443
transform 1 0 143200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6350
timestamp 1654712443
transform 1 0 146200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6351
timestamp 1654712443
transform 1 0 149200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6352
timestamp 1654712443
transform 1 0 152200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6353
timestamp 1654712443
transform 1 0 155200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6354
timestamp 1654712443
transform 1 0 158200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6355
timestamp 1654712443
transform 1 0 161200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6356
timestamp 1654712443
transform 1 0 164200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6357
timestamp 1654712443
transform 1 0 167200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6358
timestamp 1654712443
transform 1 0 170200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6359
timestamp 1654712443
transform 1 0 173200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6360
timestamp 1654712443
transform 1 0 176200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6361
timestamp 1654712443
transform 1 0 179200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6363
timestamp 1654712443
transform 1 0 185200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6362
timestamp 1654712443
transform 1 0 182200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6364
timestamp 1654712443
transform 1 0 188200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6365
timestamp 1654712443
transform 1 0 191200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6366
timestamp 1654712443
transform 1 0 194200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6367
timestamp 1654712443
transform 1 0 197200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6368
timestamp 1654712443
transform 1 0 200200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6369
timestamp 1654712443
transform 1 0 203200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6370
timestamp 1654712443
transform 1 0 206200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6371
timestamp 1654712443
transform 1 0 209200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6373
timestamp 1654712443
transform 1 0 215200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6372
timestamp 1654712443
transform 1 0 212200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6374
timestamp 1654712443
transform 1 0 218200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6375
timestamp 1654712443
transform 1 0 221200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6376
timestamp 1654712443
transform 1 0 224200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6377
timestamp 1654712443
transform 1 0 227200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6378
timestamp 1654712443
transform 1 0 230200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6379
timestamp 1654712443
transform 1 0 233200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6380
timestamp 1654712443
transform 1 0 236200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6381
timestamp 1654712443
transform 1 0 239200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6383
timestamp 1654712443
transform 1 0 245200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6382
timestamp 1654712443
transform 1 0 242200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6384
timestamp 1654712443
transform 1 0 248200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6385
timestamp 1654712443
transform 1 0 251200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6386
timestamp 1654712443
transform 1 0 254200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6387
timestamp 1654712443
transform 1 0 257200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6388
timestamp 1654712443
transform 1 0 260200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6389
timestamp 1654712443
transform 1 0 263200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6390
timestamp 1654712443
transform 1 0 266200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6391
timestamp 1654712443
transform 1 0 269200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6392
timestamp 1654712443
transform 1 0 272200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6394
timestamp 1654712443
transform 1 0 278200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6393
timestamp 1654712443
transform 1 0 275200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6395
timestamp 1654712443
transform 1 0 281200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6396
timestamp 1654712443
transform 1 0 284200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6397
timestamp 1654712443
transform 1 0 287200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6398
timestamp 1654712443
transform 1 0 290200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6399
timestamp 1654712443
transform 1 0 293200 0 1 -186300
box 3640 -2860 6960 460
use pixel  pixel_6201
timestamp 1654712443
transform 1 0 -800 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6200
timestamp 1654712443
transform 1 0 -3800 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6202
timestamp 1654712443
transform 1 0 2200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6203
timestamp 1654712443
transform 1 0 5200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6204
timestamp 1654712443
transform 1 0 8200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6205
timestamp 1654712443
transform 1 0 11200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6206
timestamp 1654712443
transform 1 0 14200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6207
timestamp 1654712443
transform 1 0 17200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6208
timestamp 1654712443
transform 1 0 20200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6209
timestamp 1654712443
transform 1 0 23200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6211
timestamp 1654712443
transform 1 0 29200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6210
timestamp 1654712443
transform 1 0 26200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6212
timestamp 1654712443
transform 1 0 32200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6213
timestamp 1654712443
transform 1 0 35200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6214
timestamp 1654712443
transform 1 0 38200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6215
timestamp 1654712443
transform 1 0 41200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6216
timestamp 1654712443
transform 1 0 44200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6217
timestamp 1654712443
transform 1 0 47200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6218
timestamp 1654712443
transform 1 0 50200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6219
timestamp 1654712443
transform 1 0 53200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6221
timestamp 1654712443
transform 1 0 59200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6220
timestamp 1654712443
transform 1 0 56200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6222
timestamp 1654712443
transform 1 0 62200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6223
timestamp 1654712443
transform 1 0 65200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6224
timestamp 1654712443
transform 1 0 68200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6225
timestamp 1654712443
transform 1 0 71200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6226
timestamp 1654712443
transform 1 0 74200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6227
timestamp 1654712443
transform 1 0 77200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6228
timestamp 1654712443
transform 1 0 80200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6229
timestamp 1654712443
transform 1 0 83200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6230
timestamp 1654712443
transform 1 0 86200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6231
timestamp 1654712443
transform 1 0 89200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6232
timestamp 1654712443
transform 1 0 92200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6233
timestamp 1654712443
transform 1 0 95200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6234
timestamp 1654712443
transform 1 0 98200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6235
timestamp 1654712443
transform 1 0 101200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6236
timestamp 1654712443
transform 1 0 104200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6237
timestamp 1654712443
transform 1 0 107200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6238
timestamp 1654712443
transform 1 0 110200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6239
timestamp 1654712443
transform 1 0 113200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6240
timestamp 1654712443
transform 1 0 116200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6241
timestamp 1654712443
transform 1 0 119200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6242
timestamp 1654712443
transform 1 0 122200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6243
timestamp 1654712443
transform 1 0 125200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6244
timestamp 1654712443
transform 1 0 128200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6245
timestamp 1654712443
transform 1 0 131200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6246
timestamp 1654712443
transform 1 0 134200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6247
timestamp 1654712443
transform 1 0 137200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6248
timestamp 1654712443
transform 1 0 140200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6249
timestamp 1654712443
transform 1 0 143200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6250
timestamp 1654712443
transform 1 0 146200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6251
timestamp 1654712443
transform 1 0 149200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6252
timestamp 1654712443
transform 1 0 152200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6253
timestamp 1654712443
transform 1 0 155200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6254
timestamp 1654712443
transform 1 0 158200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6255
timestamp 1654712443
transform 1 0 161200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6256
timestamp 1654712443
transform 1 0 164200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6257
timestamp 1654712443
transform 1 0 167200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6258
timestamp 1654712443
transform 1 0 170200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6259
timestamp 1654712443
transform 1 0 173200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6260
timestamp 1654712443
transform 1 0 176200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6261
timestamp 1654712443
transform 1 0 179200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6263
timestamp 1654712443
transform 1 0 185200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6262
timestamp 1654712443
transform 1 0 182200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6264
timestamp 1654712443
transform 1 0 188200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6265
timestamp 1654712443
transform 1 0 191200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6266
timestamp 1654712443
transform 1 0 194200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6267
timestamp 1654712443
transform 1 0 197200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6268
timestamp 1654712443
transform 1 0 200200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6269
timestamp 1654712443
transform 1 0 203200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6270
timestamp 1654712443
transform 1 0 206200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6271
timestamp 1654712443
transform 1 0 209200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6273
timestamp 1654712443
transform 1 0 215200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6272
timestamp 1654712443
transform 1 0 212200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6274
timestamp 1654712443
transform 1 0 218200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6275
timestamp 1654712443
transform 1 0 221200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6276
timestamp 1654712443
transform 1 0 224200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6277
timestamp 1654712443
transform 1 0 227200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6278
timestamp 1654712443
transform 1 0 230200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6279
timestamp 1654712443
transform 1 0 233200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6280
timestamp 1654712443
transform 1 0 236200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6281
timestamp 1654712443
transform 1 0 239200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6283
timestamp 1654712443
transform 1 0 245200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6282
timestamp 1654712443
transform 1 0 242200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6284
timestamp 1654712443
transform 1 0 248200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6285
timestamp 1654712443
transform 1 0 251200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6286
timestamp 1654712443
transform 1 0 254200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6287
timestamp 1654712443
transform 1 0 257200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6288
timestamp 1654712443
transform 1 0 260200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6289
timestamp 1654712443
transform 1 0 263200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6290
timestamp 1654712443
transform 1 0 266200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6291
timestamp 1654712443
transform 1 0 269200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6292
timestamp 1654712443
transform 1 0 272200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6294
timestamp 1654712443
transform 1 0 278200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6293
timestamp 1654712443
transform 1 0 275200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6295
timestamp 1654712443
transform 1 0 281200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6296
timestamp 1654712443
transform 1 0 284200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6297
timestamp 1654712443
transform 1 0 287200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6298
timestamp 1654712443
transform 1 0 290200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6299
timestamp 1654712443
transform 1 0 293200 0 1 -183300
box 3640 -2860 6960 460
use pixel  pixel_6101
timestamp 1654712443
transform 1 0 -800 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6100
timestamp 1654712443
transform 1 0 -3800 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6102
timestamp 1654712443
transform 1 0 2200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6103
timestamp 1654712443
transform 1 0 5200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6104
timestamp 1654712443
transform 1 0 8200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6105
timestamp 1654712443
transform 1 0 11200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6106
timestamp 1654712443
transform 1 0 14200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6107
timestamp 1654712443
transform 1 0 17200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6108
timestamp 1654712443
transform 1 0 20200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6109
timestamp 1654712443
transform 1 0 23200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6111
timestamp 1654712443
transform 1 0 29200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6110
timestamp 1654712443
transform 1 0 26200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6112
timestamp 1654712443
transform 1 0 32200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6113
timestamp 1654712443
transform 1 0 35200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6114
timestamp 1654712443
transform 1 0 38200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6115
timestamp 1654712443
transform 1 0 41200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6116
timestamp 1654712443
transform 1 0 44200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6117
timestamp 1654712443
transform 1 0 47200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6118
timestamp 1654712443
transform 1 0 50200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6119
timestamp 1654712443
transform 1 0 53200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6121
timestamp 1654712443
transform 1 0 59200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6120
timestamp 1654712443
transform 1 0 56200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6122
timestamp 1654712443
transform 1 0 62200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6123
timestamp 1654712443
transform 1 0 65200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6124
timestamp 1654712443
transform 1 0 68200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6125
timestamp 1654712443
transform 1 0 71200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6126
timestamp 1654712443
transform 1 0 74200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6127
timestamp 1654712443
transform 1 0 77200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6128
timestamp 1654712443
transform 1 0 80200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6129
timestamp 1654712443
transform 1 0 83200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6130
timestamp 1654712443
transform 1 0 86200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6131
timestamp 1654712443
transform 1 0 89200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6132
timestamp 1654712443
transform 1 0 92200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6133
timestamp 1654712443
transform 1 0 95200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6134
timestamp 1654712443
transform 1 0 98200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6135
timestamp 1654712443
transform 1 0 101200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6136
timestamp 1654712443
transform 1 0 104200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6137
timestamp 1654712443
transform 1 0 107200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6138
timestamp 1654712443
transform 1 0 110200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6139
timestamp 1654712443
transform 1 0 113200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6140
timestamp 1654712443
transform 1 0 116200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6141
timestamp 1654712443
transform 1 0 119200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6142
timestamp 1654712443
transform 1 0 122200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6143
timestamp 1654712443
transform 1 0 125200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6144
timestamp 1654712443
transform 1 0 128200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6145
timestamp 1654712443
transform 1 0 131200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6146
timestamp 1654712443
transform 1 0 134200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6147
timestamp 1654712443
transform 1 0 137200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6148
timestamp 1654712443
transform 1 0 140200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6149
timestamp 1654712443
transform 1 0 143200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6150
timestamp 1654712443
transform 1 0 146200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6151
timestamp 1654712443
transform 1 0 149200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6152
timestamp 1654712443
transform 1 0 152200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6153
timestamp 1654712443
transform 1 0 155200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6154
timestamp 1654712443
transform 1 0 158200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6155
timestamp 1654712443
transform 1 0 161200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6156
timestamp 1654712443
transform 1 0 164200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6157
timestamp 1654712443
transform 1 0 167200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6158
timestamp 1654712443
transform 1 0 170200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6159
timestamp 1654712443
transform 1 0 173200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6160
timestamp 1654712443
transform 1 0 176200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6161
timestamp 1654712443
transform 1 0 179200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6163
timestamp 1654712443
transform 1 0 185200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6162
timestamp 1654712443
transform 1 0 182200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6164
timestamp 1654712443
transform 1 0 188200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6165
timestamp 1654712443
transform 1 0 191200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6166
timestamp 1654712443
transform 1 0 194200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6167
timestamp 1654712443
transform 1 0 197200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6168
timestamp 1654712443
transform 1 0 200200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6169
timestamp 1654712443
transform 1 0 203200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6170
timestamp 1654712443
transform 1 0 206200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6171
timestamp 1654712443
transform 1 0 209200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6173
timestamp 1654712443
transform 1 0 215200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6172
timestamp 1654712443
transform 1 0 212200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6174
timestamp 1654712443
transform 1 0 218200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6175
timestamp 1654712443
transform 1 0 221200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6176
timestamp 1654712443
transform 1 0 224200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6177
timestamp 1654712443
transform 1 0 227200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6178
timestamp 1654712443
transform 1 0 230200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6179
timestamp 1654712443
transform 1 0 233200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6180
timestamp 1654712443
transform 1 0 236200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6181
timestamp 1654712443
transform 1 0 239200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6183
timestamp 1654712443
transform 1 0 245200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6182
timestamp 1654712443
transform 1 0 242200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6184
timestamp 1654712443
transform 1 0 248200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6185
timestamp 1654712443
transform 1 0 251200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6186
timestamp 1654712443
transform 1 0 254200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6187
timestamp 1654712443
transform 1 0 257200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6188
timestamp 1654712443
transform 1 0 260200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6189
timestamp 1654712443
transform 1 0 263200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6190
timestamp 1654712443
transform 1 0 266200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6191
timestamp 1654712443
transform 1 0 269200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6192
timestamp 1654712443
transform 1 0 272200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6194
timestamp 1654712443
transform 1 0 278200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6193
timestamp 1654712443
transform 1 0 275200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6195
timestamp 1654712443
transform 1 0 281200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6196
timestamp 1654712443
transform 1 0 284200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6197
timestamp 1654712443
transform 1 0 287200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6198
timestamp 1654712443
transform 1 0 290200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6199
timestamp 1654712443
transform 1 0 293200 0 1 -180300
box 3640 -2860 6960 460
use pixel  pixel_6001
timestamp 1654712443
transform 1 0 -800 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6000
timestamp 1654712443
transform 1 0 -3800 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6002
timestamp 1654712443
transform 1 0 2200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6003
timestamp 1654712443
transform 1 0 5200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6004
timestamp 1654712443
transform 1 0 8200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6005
timestamp 1654712443
transform 1 0 11200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6006
timestamp 1654712443
transform 1 0 14200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6007
timestamp 1654712443
transform 1 0 17200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6008
timestamp 1654712443
transform 1 0 20200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6009
timestamp 1654712443
transform 1 0 23200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6011
timestamp 1654712443
transform 1 0 29200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6010
timestamp 1654712443
transform 1 0 26200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6012
timestamp 1654712443
transform 1 0 32200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6013
timestamp 1654712443
transform 1 0 35200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6014
timestamp 1654712443
transform 1 0 38200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6015
timestamp 1654712443
transform 1 0 41200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6016
timestamp 1654712443
transform 1 0 44200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6017
timestamp 1654712443
transform 1 0 47200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6018
timestamp 1654712443
transform 1 0 50200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6019
timestamp 1654712443
transform 1 0 53200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6021
timestamp 1654712443
transform 1 0 59200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6020
timestamp 1654712443
transform 1 0 56200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6022
timestamp 1654712443
transform 1 0 62200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6023
timestamp 1654712443
transform 1 0 65200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6024
timestamp 1654712443
transform 1 0 68200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6025
timestamp 1654712443
transform 1 0 71200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6026
timestamp 1654712443
transform 1 0 74200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6027
timestamp 1654712443
transform 1 0 77200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6028
timestamp 1654712443
transform 1 0 80200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6029
timestamp 1654712443
transform 1 0 83200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6030
timestamp 1654712443
transform 1 0 86200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6031
timestamp 1654712443
transform 1 0 89200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6032
timestamp 1654712443
transform 1 0 92200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6033
timestamp 1654712443
transform 1 0 95200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6034
timestamp 1654712443
transform 1 0 98200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6035
timestamp 1654712443
transform 1 0 101200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6036
timestamp 1654712443
transform 1 0 104200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6037
timestamp 1654712443
transform 1 0 107200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6038
timestamp 1654712443
transform 1 0 110200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6039
timestamp 1654712443
transform 1 0 113200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6040
timestamp 1654712443
transform 1 0 116200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6041
timestamp 1654712443
transform 1 0 119200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6042
timestamp 1654712443
transform 1 0 122200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6043
timestamp 1654712443
transform 1 0 125200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6044
timestamp 1654712443
transform 1 0 128200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6045
timestamp 1654712443
transform 1 0 131200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6046
timestamp 1654712443
transform 1 0 134200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6047
timestamp 1654712443
transform 1 0 137200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6048
timestamp 1654712443
transform 1 0 140200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6049
timestamp 1654712443
transform 1 0 143200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6050
timestamp 1654712443
transform 1 0 146200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6051
timestamp 1654712443
transform 1 0 149200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6052
timestamp 1654712443
transform 1 0 152200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6053
timestamp 1654712443
transform 1 0 155200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6054
timestamp 1654712443
transform 1 0 158200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6055
timestamp 1654712443
transform 1 0 161200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6056
timestamp 1654712443
transform 1 0 164200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6057
timestamp 1654712443
transform 1 0 167200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6058
timestamp 1654712443
transform 1 0 170200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6059
timestamp 1654712443
transform 1 0 173200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6060
timestamp 1654712443
transform 1 0 176200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6061
timestamp 1654712443
transform 1 0 179200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6063
timestamp 1654712443
transform 1 0 185200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6062
timestamp 1654712443
transform 1 0 182200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6064
timestamp 1654712443
transform 1 0 188200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6065
timestamp 1654712443
transform 1 0 191200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6066
timestamp 1654712443
transform 1 0 194200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6067
timestamp 1654712443
transform 1 0 197200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6068
timestamp 1654712443
transform 1 0 200200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6069
timestamp 1654712443
transform 1 0 203200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6070
timestamp 1654712443
transform 1 0 206200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6071
timestamp 1654712443
transform 1 0 209200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6073
timestamp 1654712443
transform 1 0 215200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6072
timestamp 1654712443
transform 1 0 212200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6074
timestamp 1654712443
transform 1 0 218200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6075
timestamp 1654712443
transform 1 0 221200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6076
timestamp 1654712443
transform 1 0 224200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6077
timestamp 1654712443
transform 1 0 227200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6078
timestamp 1654712443
transform 1 0 230200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6079
timestamp 1654712443
transform 1 0 233200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6080
timestamp 1654712443
transform 1 0 236200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6081
timestamp 1654712443
transform 1 0 239200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6083
timestamp 1654712443
transform 1 0 245200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6082
timestamp 1654712443
transform 1 0 242200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6084
timestamp 1654712443
transform 1 0 248200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6085
timestamp 1654712443
transform 1 0 251200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6086
timestamp 1654712443
transform 1 0 254200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6087
timestamp 1654712443
transform 1 0 257200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6088
timestamp 1654712443
transform 1 0 260200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6089
timestamp 1654712443
transform 1 0 263200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6090
timestamp 1654712443
transform 1 0 266200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6091
timestamp 1654712443
transform 1 0 269200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6092
timestamp 1654712443
transform 1 0 272200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6094
timestamp 1654712443
transform 1 0 278200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6093
timestamp 1654712443
transform 1 0 275200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6095
timestamp 1654712443
transform 1 0 281200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6096
timestamp 1654712443
transform 1 0 284200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6097
timestamp 1654712443
transform 1 0 287200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6098
timestamp 1654712443
transform 1 0 290200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_6099
timestamp 1654712443
transform 1 0 293200 0 1 -177300
box 3640 -2860 6960 460
use pixel  pixel_5901
timestamp 1654712443
transform 1 0 -800 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5900
timestamp 1654712443
transform 1 0 -3800 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5902
timestamp 1654712443
transform 1 0 2200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5903
timestamp 1654712443
transform 1 0 5200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5904
timestamp 1654712443
transform 1 0 8200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5905
timestamp 1654712443
transform 1 0 11200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5906
timestamp 1654712443
transform 1 0 14200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5907
timestamp 1654712443
transform 1 0 17200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5908
timestamp 1654712443
transform 1 0 20200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5909
timestamp 1654712443
transform 1 0 23200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5911
timestamp 1654712443
transform 1 0 29200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5910
timestamp 1654712443
transform 1 0 26200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5912
timestamp 1654712443
transform 1 0 32200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5913
timestamp 1654712443
transform 1 0 35200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5914
timestamp 1654712443
transform 1 0 38200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5915
timestamp 1654712443
transform 1 0 41200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5916
timestamp 1654712443
transform 1 0 44200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5917
timestamp 1654712443
transform 1 0 47200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5918
timestamp 1654712443
transform 1 0 50200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5919
timestamp 1654712443
transform 1 0 53200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5921
timestamp 1654712443
transform 1 0 59200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5920
timestamp 1654712443
transform 1 0 56200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5922
timestamp 1654712443
transform 1 0 62200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5923
timestamp 1654712443
transform 1 0 65200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5924
timestamp 1654712443
transform 1 0 68200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5925
timestamp 1654712443
transform 1 0 71200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5926
timestamp 1654712443
transform 1 0 74200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5927
timestamp 1654712443
transform 1 0 77200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5928
timestamp 1654712443
transform 1 0 80200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5929
timestamp 1654712443
transform 1 0 83200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5930
timestamp 1654712443
transform 1 0 86200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5931
timestamp 1654712443
transform 1 0 89200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5932
timestamp 1654712443
transform 1 0 92200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5933
timestamp 1654712443
transform 1 0 95200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5934
timestamp 1654712443
transform 1 0 98200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5935
timestamp 1654712443
transform 1 0 101200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5936
timestamp 1654712443
transform 1 0 104200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5937
timestamp 1654712443
transform 1 0 107200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5938
timestamp 1654712443
transform 1 0 110200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5939
timestamp 1654712443
transform 1 0 113200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5940
timestamp 1654712443
transform 1 0 116200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5942
timestamp 1654712443
transform 1 0 122200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5941
timestamp 1654712443
transform 1 0 119200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5943
timestamp 1654712443
transform 1 0 125200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5944
timestamp 1654712443
transform 1 0 128200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5945
timestamp 1654712443
transform 1 0 131200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5946
timestamp 1654712443
transform 1 0 134200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5947
timestamp 1654712443
transform 1 0 137200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5948
timestamp 1654712443
transform 1 0 140200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5949
timestamp 1654712443
transform 1 0 143200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5950
timestamp 1654712443
transform 1 0 146200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5952
timestamp 1654712443
transform 1 0 152200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5951
timestamp 1654712443
transform 1 0 149200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5953
timestamp 1654712443
transform 1 0 155200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5954
timestamp 1654712443
transform 1 0 158200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5955
timestamp 1654712443
transform 1 0 161200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5956
timestamp 1654712443
transform 1 0 164200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5957
timestamp 1654712443
transform 1 0 167200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5958
timestamp 1654712443
transform 1 0 170200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5959
timestamp 1654712443
transform 1 0 173200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5960
timestamp 1654712443
transform 1 0 176200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5961
timestamp 1654712443
transform 1 0 179200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5963
timestamp 1654712443
transform 1 0 185200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5962
timestamp 1654712443
transform 1 0 182200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5964
timestamp 1654712443
transform 1 0 188200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5965
timestamp 1654712443
transform 1 0 191200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5966
timestamp 1654712443
transform 1 0 194200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5967
timestamp 1654712443
transform 1 0 197200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5968
timestamp 1654712443
transform 1 0 200200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5969
timestamp 1654712443
transform 1 0 203200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5970
timestamp 1654712443
transform 1 0 206200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5971
timestamp 1654712443
transform 1 0 209200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5973
timestamp 1654712443
transform 1 0 215200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5972
timestamp 1654712443
transform 1 0 212200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5974
timestamp 1654712443
transform 1 0 218200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5975
timestamp 1654712443
transform 1 0 221200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5976
timestamp 1654712443
transform 1 0 224200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5977
timestamp 1654712443
transform 1 0 227200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5978
timestamp 1654712443
transform 1 0 230200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5979
timestamp 1654712443
transform 1 0 233200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5980
timestamp 1654712443
transform 1 0 236200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5981
timestamp 1654712443
transform 1 0 239200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5983
timestamp 1654712443
transform 1 0 245200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5982
timestamp 1654712443
transform 1 0 242200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5984
timestamp 1654712443
transform 1 0 248200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5985
timestamp 1654712443
transform 1 0 251200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5986
timestamp 1654712443
transform 1 0 254200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5987
timestamp 1654712443
transform 1 0 257200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5988
timestamp 1654712443
transform 1 0 260200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5989
timestamp 1654712443
transform 1 0 263200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5990
timestamp 1654712443
transform 1 0 266200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5991
timestamp 1654712443
transform 1 0 269200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5992
timestamp 1654712443
transform 1 0 272200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5994
timestamp 1654712443
transform 1 0 278200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5993
timestamp 1654712443
transform 1 0 275200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5995
timestamp 1654712443
transform 1 0 281200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5996
timestamp 1654712443
transform 1 0 284200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5997
timestamp 1654712443
transform 1 0 287200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5998
timestamp 1654712443
transform 1 0 290200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5999
timestamp 1654712443
transform 1 0 293200 0 1 -174300
box 3640 -2860 6960 460
use pixel  pixel_5701
timestamp 1654712443
transform 1 0 -800 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5801
timestamp 1654712443
transform 1 0 -800 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5700
timestamp 1654712443
transform 1 0 -3800 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5800
timestamp 1654712443
transform 1 0 -3800 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5702
timestamp 1654712443
transform 1 0 2200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5802
timestamp 1654712443
transform 1 0 2200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5703
timestamp 1654712443
transform 1 0 5200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5803
timestamp 1654712443
transform 1 0 5200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5704
timestamp 1654712443
transform 1 0 8200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5804
timestamp 1654712443
transform 1 0 8200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5705
timestamp 1654712443
transform 1 0 11200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5805
timestamp 1654712443
transform 1 0 11200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5706
timestamp 1654712443
transform 1 0 14200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5806
timestamp 1654712443
transform 1 0 14200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5707
timestamp 1654712443
transform 1 0 17200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5807
timestamp 1654712443
transform 1 0 17200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5708
timestamp 1654712443
transform 1 0 20200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5808
timestamp 1654712443
transform 1 0 20200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5709
timestamp 1654712443
transform 1 0 23200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5809
timestamp 1654712443
transform 1 0 23200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5711
timestamp 1654712443
transform 1 0 29200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5811
timestamp 1654712443
transform 1 0 29200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5710
timestamp 1654712443
transform 1 0 26200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5810
timestamp 1654712443
transform 1 0 26200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5712
timestamp 1654712443
transform 1 0 32200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5812
timestamp 1654712443
transform 1 0 32200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5713
timestamp 1654712443
transform 1 0 35200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5813
timestamp 1654712443
transform 1 0 35200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5714
timestamp 1654712443
transform 1 0 38200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5814
timestamp 1654712443
transform 1 0 38200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5715
timestamp 1654712443
transform 1 0 41200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5815
timestamp 1654712443
transform 1 0 41200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5716
timestamp 1654712443
transform 1 0 44200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5816
timestamp 1654712443
transform 1 0 44200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5717
timestamp 1654712443
transform 1 0 47200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5817
timestamp 1654712443
transform 1 0 47200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5718
timestamp 1654712443
transform 1 0 50200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5818
timestamp 1654712443
transform 1 0 50200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5719
timestamp 1654712443
transform 1 0 53200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5819
timestamp 1654712443
transform 1 0 53200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5721
timestamp 1654712443
transform 1 0 59200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5821
timestamp 1654712443
transform 1 0 59200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5720
timestamp 1654712443
transform 1 0 56200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5820
timestamp 1654712443
transform 1 0 56200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5722
timestamp 1654712443
transform 1 0 62200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5822
timestamp 1654712443
transform 1 0 62200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5723
timestamp 1654712443
transform 1 0 65200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5823
timestamp 1654712443
transform 1 0 65200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5724
timestamp 1654712443
transform 1 0 68200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5824
timestamp 1654712443
transform 1 0 68200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5725
timestamp 1654712443
transform 1 0 71200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5825
timestamp 1654712443
transform 1 0 71200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5726
timestamp 1654712443
transform 1 0 74200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5826
timestamp 1654712443
transform 1 0 74200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5727
timestamp 1654712443
transform 1 0 77200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5827
timestamp 1654712443
transform 1 0 77200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5728
timestamp 1654712443
transform 1 0 80200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5828
timestamp 1654712443
transform 1 0 80200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5729
timestamp 1654712443
transform 1 0 83200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5829
timestamp 1654712443
transform 1 0 83200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5730
timestamp 1654712443
transform 1 0 86200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5830
timestamp 1654712443
transform 1 0 86200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5731
timestamp 1654712443
transform 1 0 89200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5732
timestamp 1654712443
transform 1 0 92200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5831
timestamp 1654712443
transform 1 0 89200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5832
timestamp 1654712443
transform 1 0 92200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5733
timestamp 1654712443
transform 1 0 95200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5833
timestamp 1654712443
transform 1 0 95200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5734
timestamp 1654712443
transform 1 0 98200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5834
timestamp 1654712443
transform 1 0 98200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5735
timestamp 1654712443
transform 1 0 101200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5835
timestamp 1654712443
transform 1 0 101200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5736
timestamp 1654712443
transform 1 0 104200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5836
timestamp 1654712443
transform 1 0 104200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5737
timestamp 1654712443
transform 1 0 107200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5837
timestamp 1654712443
transform 1 0 107200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5738
timestamp 1654712443
transform 1 0 110200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5838
timestamp 1654712443
transform 1 0 110200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5739
timestamp 1654712443
transform 1 0 113200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5839
timestamp 1654712443
transform 1 0 113200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5740
timestamp 1654712443
transform 1 0 116200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5840
timestamp 1654712443
transform 1 0 116200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5742
timestamp 1654712443
transform 1 0 122200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5741
timestamp 1654712443
transform 1 0 119200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5842
timestamp 1654712443
transform 1 0 122200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5841
timestamp 1654712443
transform 1 0 119200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5743
timestamp 1654712443
transform 1 0 125200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5843
timestamp 1654712443
transform 1 0 125200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5744
timestamp 1654712443
transform 1 0 128200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5844
timestamp 1654712443
transform 1 0 128200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5745
timestamp 1654712443
transform 1 0 131200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5845
timestamp 1654712443
transform 1 0 131200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5746
timestamp 1654712443
transform 1 0 134200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5846
timestamp 1654712443
transform 1 0 134200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5747
timestamp 1654712443
transform 1 0 137200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5847
timestamp 1654712443
transform 1 0 137200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5748
timestamp 1654712443
transform 1 0 140200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5848
timestamp 1654712443
transform 1 0 140200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5749
timestamp 1654712443
transform 1 0 143200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5849
timestamp 1654712443
transform 1 0 143200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5750
timestamp 1654712443
transform 1 0 146200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5850
timestamp 1654712443
transform 1 0 146200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5752
timestamp 1654712443
transform 1 0 152200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5751
timestamp 1654712443
transform 1 0 149200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5852
timestamp 1654712443
transform 1 0 152200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5851
timestamp 1654712443
transform 1 0 149200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5753
timestamp 1654712443
transform 1 0 155200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5853
timestamp 1654712443
transform 1 0 155200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5754
timestamp 1654712443
transform 1 0 158200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5854
timestamp 1654712443
transform 1 0 158200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5755
timestamp 1654712443
transform 1 0 161200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5855
timestamp 1654712443
transform 1 0 161200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5756
timestamp 1654712443
transform 1 0 164200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5856
timestamp 1654712443
transform 1 0 164200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5757
timestamp 1654712443
transform 1 0 167200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5857
timestamp 1654712443
transform 1 0 167200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5758
timestamp 1654712443
transform 1 0 170200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5858
timestamp 1654712443
transform 1 0 170200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5759
timestamp 1654712443
transform 1 0 173200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5859
timestamp 1654712443
transform 1 0 173200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5760
timestamp 1654712443
transform 1 0 176200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5860
timestamp 1654712443
transform 1 0 176200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5761
timestamp 1654712443
transform 1 0 179200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5861
timestamp 1654712443
transform 1 0 179200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5763
timestamp 1654712443
transform 1 0 185200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5863
timestamp 1654712443
transform 1 0 185200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5762
timestamp 1654712443
transform 1 0 182200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5862
timestamp 1654712443
transform 1 0 182200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5764
timestamp 1654712443
transform 1 0 188200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5864
timestamp 1654712443
transform 1 0 188200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5765
timestamp 1654712443
transform 1 0 191200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5865
timestamp 1654712443
transform 1 0 191200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5766
timestamp 1654712443
transform 1 0 194200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5866
timestamp 1654712443
transform 1 0 194200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5767
timestamp 1654712443
transform 1 0 197200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5867
timestamp 1654712443
transform 1 0 197200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5768
timestamp 1654712443
transform 1 0 200200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5868
timestamp 1654712443
transform 1 0 200200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5769
timestamp 1654712443
transform 1 0 203200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5869
timestamp 1654712443
transform 1 0 203200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5770
timestamp 1654712443
transform 1 0 206200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5870
timestamp 1654712443
transform 1 0 206200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5771
timestamp 1654712443
transform 1 0 209200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5871
timestamp 1654712443
transform 1 0 209200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5773
timestamp 1654712443
transform 1 0 215200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5873
timestamp 1654712443
transform 1 0 215200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5772
timestamp 1654712443
transform 1 0 212200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5872
timestamp 1654712443
transform 1 0 212200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5774
timestamp 1654712443
transform 1 0 218200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5874
timestamp 1654712443
transform 1 0 218200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5775
timestamp 1654712443
transform 1 0 221200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5875
timestamp 1654712443
transform 1 0 221200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5776
timestamp 1654712443
transform 1 0 224200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5876
timestamp 1654712443
transform 1 0 224200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5777
timestamp 1654712443
transform 1 0 227200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5877
timestamp 1654712443
transform 1 0 227200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5778
timestamp 1654712443
transform 1 0 230200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5878
timestamp 1654712443
transform 1 0 230200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5779
timestamp 1654712443
transform 1 0 233200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5879
timestamp 1654712443
transform 1 0 233200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5780
timestamp 1654712443
transform 1 0 236200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5880
timestamp 1654712443
transform 1 0 236200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5781
timestamp 1654712443
transform 1 0 239200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5881
timestamp 1654712443
transform 1 0 239200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5783
timestamp 1654712443
transform 1 0 245200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5883
timestamp 1654712443
transform 1 0 245200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5782
timestamp 1654712443
transform 1 0 242200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5882
timestamp 1654712443
transform 1 0 242200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5784
timestamp 1654712443
transform 1 0 248200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5884
timestamp 1654712443
transform 1 0 248200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5785
timestamp 1654712443
transform 1 0 251200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5885
timestamp 1654712443
transform 1 0 251200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5786
timestamp 1654712443
transform 1 0 254200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5886
timestamp 1654712443
transform 1 0 254200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5787
timestamp 1654712443
transform 1 0 257200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5887
timestamp 1654712443
transform 1 0 257200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5788
timestamp 1654712443
transform 1 0 260200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5888
timestamp 1654712443
transform 1 0 260200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5789
timestamp 1654712443
transform 1 0 263200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5889
timestamp 1654712443
transform 1 0 263200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5790
timestamp 1654712443
transform 1 0 266200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5890
timestamp 1654712443
transform 1 0 266200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5791
timestamp 1654712443
transform 1 0 269200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5891
timestamp 1654712443
transform 1 0 269200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5792
timestamp 1654712443
transform 1 0 272200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5892
timestamp 1654712443
transform 1 0 272200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5794
timestamp 1654712443
transform 1 0 278200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5894
timestamp 1654712443
transform 1 0 278200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5793
timestamp 1654712443
transform 1 0 275200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5893
timestamp 1654712443
transform 1 0 275200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5795
timestamp 1654712443
transform 1 0 281200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5895
timestamp 1654712443
transform 1 0 281200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5796
timestamp 1654712443
transform 1 0 284200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5896
timestamp 1654712443
transform 1 0 284200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5797
timestamp 1654712443
transform 1 0 287200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5897
timestamp 1654712443
transform 1 0 287200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5798
timestamp 1654712443
transform 1 0 290200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5898
timestamp 1654712443
transform 1 0 290200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5799
timestamp 1654712443
transform 1 0 293200 0 1 -168300
box 3640 -2860 6960 460
use pixel  pixel_5899
timestamp 1654712443
transform 1 0 293200 0 1 -171300
box 3640 -2860 6960 460
use pixel  pixel_5601
timestamp 1654712443
transform 1 0 -800 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5600
timestamp 1654712443
transform 1 0 -3800 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5602
timestamp 1654712443
transform 1 0 2200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5603
timestamp 1654712443
transform 1 0 5200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5604
timestamp 1654712443
transform 1 0 8200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5605
timestamp 1654712443
transform 1 0 11200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5606
timestamp 1654712443
transform 1 0 14200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5607
timestamp 1654712443
transform 1 0 17200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5608
timestamp 1654712443
transform 1 0 20200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5609
timestamp 1654712443
transform 1 0 23200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5611
timestamp 1654712443
transform 1 0 29200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5610
timestamp 1654712443
transform 1 0 26200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5612
timestamp 1654712443
transform 1 0 32200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5613
timestamp 1654712443
transform 1 0 35200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5614
timestamp 1654712443
transform 1 0 38200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5615
timestamp 1654712443
transform 1 0 41200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5616
timestamp 1654712443
transform 1 0 44200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5617
timestamp 1654712443
transform 1 0 47200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5618
timestamp 1654712443
transform 1 0 50200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5619
timestamp 1654712443
transform 1 0 53200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5621
timestamp 1654712443
transform 1 0 59200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5620
timestamp 1654712443
transform 1 0 56200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5622
timestamp 1654712443
transform 1 0 62200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5623
timestamp 1654712443
transform 1 0 65200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5624
timestamp 1654712443
transform 1 0 68200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5625
timestamp 1654712443
transform 1 0 71200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5626
timestamp 1654712443
transform 1 0 74200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5627
timestamp 1654712443
transform 1 0 77200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5628
timestamp 1654712443
transform 1 0 80200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5629
timestamp 1654712443
transform 1 0 83200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5630
timestamp 1654712443
transform 1 0 86200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5631
timestamp 1654712443
transform 1 0 89200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5632
timestamp 1654712443
transform 1 0 92200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5633
timestamp 1654712443
transform 1 0 95200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5634
timestamp 1654712443
transform 1 0 98200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5635
timestamp 1654712443
transform 1 0 101200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5636
timestamp 1654712443
transform 1 0 104200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5637
timestamp 1654712443
transform 1 0 107200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5638
timestamp 1654712443
transform 1 0 110200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5639
timestamp 1654712443
transform 1 0 113200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5640
timestamp 1654712443
transform 1 0 116200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5642
timestamp 1654712443
transform 1 0 122200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5641
timestamp 1654712443
transform 1 0 119200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5643
timestamp 1654712443
transform 1 0 125200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5644
timestamp 1654712443
transform 1 0 128200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5645
timestamp 1654712443
transform 1 0 131200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5646
timestamp 1654712443
transform 1 0 134200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5647
timestamp 1654712443
transform 1 0 137200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5648
timestamp 1654712443
transform 1 0 140200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5649
timestamp 1654712443
transform 1 0 143200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5650
timestamp 1654712443
transform 1 0 146200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5652
timestamp 1654712443
transform 1 0 152200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5651
timestamp 1654712443
transform 1 0 149200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5653
timestamp 1654712443
transform 1 0 155200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5654
timestamp 1654712443
transform 1 0 158200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5655
timestamp 1654712443
transform 1 0 161200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5656
timestamp 1654712443
transform 1 0 164200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5657
timestamp 1654712443
transform 1 0 167200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5658
timestamp 1654712443
transform 1 0 170200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5659
timestamp 1654712443
transform 1 0 173200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5660
timestamp 1654712443
transform 1 0 176200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5661
timestamp 1654712443
transform 1 0 179200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5663
timestamp 1654712443
transform 1 0 185200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5662
timestamp 1654712443
transform 1 0 182200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5664
timestamp 1654712443
transform 1 0 188200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5665
timestamp 1654712443
transform 1 0 191200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5666
timestamp 1654712443
transform 1 0 194200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5667
timestamp 1654712443
transform 1 0 197200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5668
timestamp 1654712443
transform 1 0 200200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5669
timestamp 1654712443
transform 1 0 203200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5670
timestamp 1654712443
transform 1 0 206200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5671
timestamp 1654712443
transform 1 0 209200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5673
timestamp 1654712443
transform 1 0 215200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5672
timestamp 1654712443
transform 1 0 212200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5674
timestamp 1654712443
transform 1 0 218200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5675
timestamp 1654712443
transform 1 0 221200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5676
timestamp 1654712443
transform 1 0 224200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5677
timestamp 1654712443
transform 1 0 227200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5678
timestamp 1654712443
transform 1 0 230200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5679
timestamp 1654712443
transform 1 0 233200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5680
timestamp 1654712443
transform 1 0 236200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5681
timestamp 1654712443
transform 1 0 239200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5683
timestamp 1654712443
transform 1 0 245200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5682
timestamp 1654712443
transform 1 0 242200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5684
timestamp 1654712443
transform 1 0 248200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5685
timestamp 1654712443
transform 1 0 251200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5686
timestamp 1654712443
transform 1 0 254200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5687
timestamp 1654712443
transform 1 0 257200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5688
timestamp 1654712443
transform 1 0 260200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5689
timestamp 1654712443
transform 1 0 263200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5690
timestamp 1654712443
transform 1 0 266200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5691
timestamp 1654712443
transform 1 0 269200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5692
timestamp 1654712443
transform 1 0 272200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5694
timestamp 1654712443
transform 1 0 278200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5693
timestamp 1654712443
transform 1 0 275200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5695
timestamp 1654712443
transform 1 0 281200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5696
timestamp 1654712443
transform 1 0 284200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5697
timestamp 1654712443
transform 1 0 287200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5698
timestamp 1654712443
transform 1 0 290200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5699
timestamp 1654712443
transform 1 0 293200 0 1 -165300
box 3640 -2860 6960 460
use pixel  pixel_5501
timestamp 1654712443
transform 1 0 -800 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5500
timestamp 1654712443
transform 1 0 -3800 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5502
timestamp 1654712443
transform 1 0 2200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5503
timestamp 1654712443
transform 1 0 5200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5504
timestamp 1654712443
transform 1 0 8200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5505
timestamp 1654712443
transform 1 0 11200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5506
timestamp 1654712443
transform 1 0 14200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5507
timestamp 1654712443
transform 1 0 17200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5508
timestamp 1654712443
transform 1 0 20200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5509
timestamp 1654712443
transform 1 0 23200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5511
timestamp 1654712443
transform 1 0 29200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5510
timestamp 1654712443
transform 1 0 26200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5512
timestamp 1654712443
transform 1 0 32200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5513
timestamp 1654712443
transform 1 0 35200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5514
timestamp 1654712443
transform 1 0 38200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5515
timestamp 1654712443
transform 1 0 41200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5516
timestamp 1654712443
transform 1 0 44200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5517
timestamp 1654712443
transform 1 0 47200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5518
timestamp 1654712443
transform 1 0 50200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5519
timestamp 1654712443
transform 1 0 53200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5521
timestamp 1654712443
transform 1 0 59200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5520
timestamp 1654712443
transform 1 0 56200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5522
timestamp 1654712443
transform 1 0 62200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5523
timestamp 1654712443
transform 1 0 65200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5524
timestamp 1654712443
transform 1 0 68200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5525
timestamp 1654712443
transform 1 0 71200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5526
timestamp 1654712443
transform 1 0 74200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5527
timestamp 1654712443
transform 1 0 77200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5528
timestamp 1654712443
transform 1 0 80200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5529
timestamp 1654712443
transform 1 0 83200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5530
timestamp 1654712443
transform 1 0 86200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5531
timestamp 1654712443
transform 1 0 89200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5532
timestamp 1654712443
transform 1 0 92200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5533
timestamp 1654712443
transform 1 0 95200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5534
timestamp 1654712443
transform 1 0 98200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5535
timestamp 1654712443
transform 1 0 101200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5536
timestamp 1654712443
transform 1 0 104200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5537
timestamp 1654712443
transform 1 0 107200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5538
timestamp 1654712443
transform 1 0 110200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5539
timestamp 1654712443
transform 1 0 113200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5540
timestamp 1654712443
transform 1 0 116200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5542
timestamp 1654712443
transform 1 0 122200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5541
timestamp 1654712443
transform 1 0 119200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5543
timestamp 1654712443
transform 1 0 125200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5544
timestamp 1654712443
transform 1 0 128200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5545
timestamp 1654712443
transform 1 0 131200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5546
timestamp 1654712443
transform 1 0 134200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5547
timestamp 1654712443
transform 1 0 137200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5548
timestamp 1654712443
transform 1 0 140200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5549
timestamp 1654712443
transform 1 0 143200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5550
timestamp 1654712443
transform 1 0 146200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5552
timestamp 1654712443
transform 1 0 152200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5551
timestamp 1654712443
transform 1 0 149200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5553
timestamp 1654712443
transform 1 0 155200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5554
timestamp 1654712443
transform 1 0 158200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5555
timestamp 1654712443
transform 1 0 161200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5556
timestamp 1654712443
transform 1 0 164200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5557
timestamp 1654712443
transform 1 0 167200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5558
timestamp 1654712443
transform 1 0 170200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5559
timestamp 1654712443
transform 1 0 173200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5560
timestamp 1654712443
transform 1 0 176200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5561
timestamp 1654712443
transform 1 0 179200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5563
timestamp 1654712443
transform 1 0 185200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5562
timestamp 1654712443
transform 1 0 182200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5564
timestamp 1654712443
transform 1 0 188200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5565
timestamp 1654712443
transform 1 0 191200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5566
timestamp 1654712443
transform 1 0 194200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5567
timestamp 1654712443
transform 1 0 197200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5568
timestamp 1654712443
transform 1 0 200200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5569
timestamp 1654712443
transform 1 0 203200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5570
timestamp 1654712443
transform 1 0 206200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5571
timestamp 1654712443
transform 1 0 209200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5573
timestamp 1654712443
transform 1 0 215200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5572
timestamp 1654712443
transform 1 0 212200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5574
timestamp 1654712443
transform 1 0 218200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5575
timestamp 1654712443
transform 1 0 221200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5576
timestamp 1654712443
transform 1 0 224200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5577
timestamp 1654712443
transform 1 0 227200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5578
timestamp 1654712443
transform 1 0 230200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5579
timestamp 1654712443
transform 1 0 233200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5580
timestamp 1654712443
transform 1 0 236200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5581
timestamp 1654712443
transform 1 0 239200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5583
timestamp 1654712443
transform 1 0 245200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5582
timestamp 1654712443
transform 1 0 242200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5584
timestamp 1654712443
transform 1 0 248200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5585
timestamp 1654712443
transform 1 0 251200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5586
timestamp 1654712443
transform 1 0 254200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5587
timestamp 1654712443
transform 1 0 257200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5588
timestamp 1654712443
transform 1 0 260200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5589
timestamp 1654712443
transform 1 0 263200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5590
timestamp 1654712443
transform 1 0 266200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5591
timestamp 1654712443
transform 1 0 269200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5592
timestamp 1654712443
transform 1 0 272200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5594
timestamp 1654712443
transform 1 0 278200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5593
timestamp 1654712443
transform 1 0 275200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5595
timestamp 1654712443
transform 1 0 281200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5596
timestamp 1654712443
transform 1 0 284200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5597
timestamp 1654712443
transform 1 0 287200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5598
timestamp 1654712443
transform 1 0 290200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5599
timestamp 1654712443
transform 1 0 293200 0 1 -162300
box 3640 -2860 6960 460
use pixel  pixel_5401
timestamp 1654712443
transform 1 0 -800 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5400
timestamp 1654712443
transform 1 0 -3800 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5402
timestamp 1654712443
transform 1 0 2200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5403
timestamp 1654712443
transform 1 0 5200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5404
timestamp 1654712443
transform 1 0 8200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5405
timestamp 1654712443
transform 1 0 11200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5406
timestamp 1654712443
transform 1 0 14200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5407
timestamp 1654712443
transform 1 0 17200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5408
timestamp 1654712443
transform 1 0 20200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5409
timestamp 1654712443
transform 1 0 23200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5411
timestamp 1654712443
transform 1 0 29200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5410
timestamp 1654712443
transform 1 0 26200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5412
timestamp 1654712443
transform 1 0 32200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5413
timestamp 1654712443
transform 1 0 35200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5414
timestamp 1654712443
transform 1 0 38200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5415
timestamp 1654712443
transform 1 0 41200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5416
timestamp 1654712443
transform 1 0 44200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5417
timestamp 1654712443
transform 1 0 47200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5418
timestamp 1654712443
transform 1 0 50200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5419
timestamp 1654712443
transform 1 0 53200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5421
timestamp 1654712443
transform 1 0 59200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5420
timestamp 1654712443
transform 1 0 56200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5422
timestamp 1654712443
transform 1 0 62200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5423
timestamp 1654712443
transform 1 0 65200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5424
timestamp 1654712443
transform 1 0 68200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5425
timestamp 1654712443
transform 1 0 71200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5426
timestamp 1654712443
transform 1 0 74200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5427
timestamp 1654712443
transform 1 0 77200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5428
timestamp 1654712443
transform 1 0 80200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5429
timestamp 1654712443
transform 1 0 83200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5430
timestamp 1654712443
transform 1 0 86200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5431
timestamp 1654712443
transform 1 0 89200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5432
timestamp 1654712443
transform 1 0 92200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5433
timestamp 1654712443
transform 1 0 95200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5434
timestamp 1654712443
transform 1 0 98200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5435
timestamp 1654712443
transform 1 0 101200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5436
timestamp 1654712443
transform 1 0 104200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5437
timestamp 1654712443
transform 1 0 107200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5438
timestamp 1654712443
transform 1 0 110200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5439
timestamp 1654712443
transform 1 0 113200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5440
timestamp 1654712443
transform 1 0 116200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5442
timestamp 1654712443
transform 1 0 122200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5441
timestamp 1654712443
transform 1 0 119200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5443
timestamp 1654712443
transform 1 0 125200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5444
timestamp 1654712443
transform 1 0 128200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5445
timestamp 1654712443
transform 1 0 131200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5446
timestamp 1654712443
transform 1 0 134200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5447
timestamp 1654712443
transform 1 0 137200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5448
timestamp 1654712443
transform 1 0 140200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5449
timestamp 1654712443
transform 1 0 143200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5450
timestamp 1654712443
transform 1 0 146200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5452
timestamp 1654712443
transform 1 0 152200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5451
timestamp 1654712443
transform 1 0 149200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5453
timestamp 1654712443
transform 1 0 155200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5454
timestamp 1654712443
transform 1 0 158200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5455
timestamp 1654712443
transform 1 0 161200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5456
timestamp 1654712443
transform 1 0 164200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5457
timestamp 1654712443
transform 1 0 167200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5458
timestamp 1654712443
transform 1 0 170200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5459
timestamp 1654712443
transform 1 0 173200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5460
timestamp 1654712443
transform 1 0 176200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5461
timestamp 1654712443
transform 1 0 179200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5463
timestamp 1654712443
transform 1 0 185200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5462
timestamp 1654712443
transform 1 0 182200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5464
timestamp 1654712443
transform 1 0 188200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5465
timestamp 1654712443
transform 1 0 191200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5466
timestamp 1654712443
transform 1 0 194200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5467
timestamp 1654712443
transform 1 0 197200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5468
timestamp 1654712443
transform 1 0 200200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5469
timestamp 1654712443
transform 1 0 203200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5470
timestamp 1654712443
transform 1 0 206200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5471
timestamp 1654712443
transform 1 0 209200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5473
timestamp 1654712443
transform 1 0 215200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5472
timestamp 1654712443
transform 1 0 212200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5474
timestamp 1654712443
transform 1 0 218200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5475
timestamp 1654712443
transform 1 0 221200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5476
timestamp 1654712443
transform 1 0 224200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5477
timestamp 1654712443
transform 1 0 227200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5478
timestamp 1654712443
transform 1 0 230200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5479
timestamp 1654712443
transform 1 0 233200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5480
timestamp 1654712443
transform 1 0 236200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5481
timestamp 1654712443
transform 1 0 239200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5483
timestamp 1654712443
transform 1 0 245200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5482
timestamp 1654712443
transform 1 0 242200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5484
timestamp 1654712443
transform 1 0 248200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5485
timestamp 1654712443
transform 1 0 251200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5486
timestamp 1654712443
transform 1 0 254200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5487
timestamp 1654712443
transform 1 0 257200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5488
timestamp 1654712443
transform 1 0 260200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5489
timestamp 1654712443
transform 1 0 263200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5490
timestamp 1654712443
transform 1 0 266200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5491
timestamp 1654712443
transform 1 0 269200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5492
timestamp 1654712443
transform 1 0 272200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5494
timestamp 1654712443
transform 1 0 278200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5493
timestamp 1654712443
transform 1 0 275200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5495
timestamp 1654712443
transform 1 0 281200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5496
timestamp 1654712443
transform 1 0 284200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5497
timestamp 1654712443
transform 1 0 287200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5498
timestamp 1654712443
transform 1 0 290200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5499
timestamp 1654712443
transform 1 0 293200 0 1 -159300
box 3640 -2860 6960 460
use pixel  pixel_5301
timestamp 1654712443
transform 1 0 -800 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5300
timestamp 1654712443
transform 1 0 -3800 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5302
timestamp 1654712443
transform 1 0 2200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5303
timestamp 1654712443
transform 1 0 5200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5304
timestamp 1654712443
transform 1 0 8200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5305
timestamp 1654712443
transform 1 0 11200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5306
timestamp 1654712443
transform 1 0 14200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5307
timestamp 1654712443
transform 1 0 17200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5308
timestamp 1654712443
transform 1 0 20200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5309
timestamp 1654712443
transform 1 0 23200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5311
timestamp 1654712443
transform 1 0 29200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5310
timestamp 1654712443
transform 1 0 26200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5312
timestamp 1654712443
transform 1 0 32200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5313
timestamp 1654712443
transform 1 0 35200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5314
timestamp 1654712443
transform 1 0 38200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5315
timestamp 1654712443
transform 1 0 41200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5316
timestamp 1654712443
transform 1 0 44200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5317
timestamp 1654712443
transform 1 0 47200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5318
timestamp 1654712443
transform 1 0 50200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5319
timestamp 1654712443
transform 1 0 53200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5321
timestamp 1654712443
transform 1 0 59200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5320
timestamp 1654712443
transform 1 0 56200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5322
timestamp 1654712443
transform 1 0 62200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5323
timestamp 1654712443
transform 1 0 65200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5324
timestamp 1654712443
transform 1 0 68200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5325
timestamp 1654712443
transform 1 0 71200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5326
timestamp 1654712443
transform 1 0 74200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5327
timestamp 1654712443
transform 1 0 77200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5328
timestamp 1654712443
transform 1 0 80200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5329
timestamp 1654712443
transform 1 0 83200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5330
timestamp 1654712443
transform 1 0 86200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5331
timestamp 1654712443
transform 1 0 89200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5332
timestamp 1654712443
transform 1 0 92200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5333
timestamp 1654712443
transform 1 0 95200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5334
timestamp 1654712443
transform 1 0 98200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5335
timestamp 1654712443
transform 1 0 101200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5336
timestamp 1654712443
transform 1 0 104200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5337
timestamp 1654712443
transform 1 0 107200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5338
timestamp 1654712443
transform 1 0 110200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5339
timestamp 1654712443
transform 1 0 113200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5340
timestamp 1654712443
transform 1 0 116200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5342
timestamp 1654712443
transform 1 0 122200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5341
timestamp 1654712443
transform 1 0 119200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5343
timestamp 1654712443
transform 1 0 125200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5344
timestamp 1654712443
transform 1 0 128200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5345
timestamp 1654712443
transform 1 0 131200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5346
timestamp 1654712443
transform 1 0 134200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5347
timestamp 1654712443
transform 1 0 137200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5348
timestamp 1654712443
transform 1 0 140200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5349
timestamp 1654712443
transform 1 0 143200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5350
timestamp 1654712443
transform 1 0 146200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5352
timestamp 1654712443
transform 1 0 152200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5351
timestamp 1654712443
transform 1 0 149200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5353
timestamp 1654712443
transform 1 0 155200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5354
timestamp 1654712443
transform 1 0 158200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5355
timestamp 1654712443
transform 1 0 161200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5356
timestamp 1654712443
transform 1 0 164200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5357
timestamp 1654712443
transform 1 0 167200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5358
timestamp 1654712443
transform 1 0 170200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5359
timestamp 1654712443
transform 1 0 173200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5360
timestamp 1654712443
transform 1 0 176200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5361
timestamp 1654712443
transform 1 0 179200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5363
timestamp 1654712443
transform 1 0 185200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5362
timestamp 1654712443
transform 1 0 182200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5364
timestamp 1654712443
transform 1 0 188200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5365
timestamp 1654712443
transform 1 0 191200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5366
timestamp 1654712443
transform 1 0 194200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5367
timestamp 1654712443
transform 1 0 197200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5368
timestamp 1654712443
transform 1 0 200200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5369
timestamp 1654712443
transform 1 0 203200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5370
timestamp 1654712443
transform 1 0 206200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5371
timestamp 1654712443
transform 1 0 209200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5373
timestamp 1654712443
transform 1 0 215200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5372
timestamp 1654712443
transform 1 0 212200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5374
timestamp 1654712443
transform 1 0 218200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5375
timestamp 1654712443
transform 1 0 221200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5376
timestamp 1654712443
transform 1 0 224200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5377
timestamp 1654712443
transform 1 0 227200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5378
timestamp 1654712443
transform 1 0 230200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5379
timestamp 1654712443
transform 1 0 233200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5380
timestamp 1654712443
transform 1 0 236200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5381
timestamp 1654712443
transform 1 0 239200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5383
timestamp 1654712443
transform 1 0 245200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5382
timestamp 1654712443
transform 1 0 242200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5384
timestamp 1654712443
transform 1 0 248200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5385
timestamp 1654712443
transform 1 0 251200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5386
timestamp 1654712443
transform 1 0 254200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5387
timestamp 1654712443
transform 1 0 257200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5388
timestamp 1654712443
transform 1 0 260200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5389
timestamp 1654712443
transform 1 0 263200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5390
timestamp 1654712443
transform 1 0 266200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5391
timestamp 1654712443
transform 1 0 269200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5392
timestamp 1654712443
transform 1 0 272200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5394
timestamp 1654712443
transform 1 0 278200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5393
timestamp 1654712443
transform 1 0 275200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5395
timestamp 1654712443
transform 1 0 281200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5396
timestamp 1654712443
transform 1 0 284200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5397
timestamp 1654712443
transform 1 0 287200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5398
timestamp 1654712443
transform 1 0 290200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5399
timestamp 1654712443
transform 1 0 293200 0 1 -156300
box 3640 -2860 6960 460
use pixel  pixel_5201
timestamp 1654712443
transform 1 0 -800 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5200
timestamp 1654712443
transform 1 0 -3800 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5202
timestamp 1654712443
transform 1 0 2200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5203
timestamp 1654712443
transform 1 0 5200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5204
timestamp 1654712443
transform 1 0 8200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5205
timestamp 1654712443
transform 1 0 11200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5206
timestamp 1654712443
transform 1 0 14200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5207
timestamp 1654712443
transform 1 0 17200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5208
timestamp 1654712443
transform 1 0 20200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5209
timestamp 1654712443
transform 1 0 23200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5211
timestamp 1654712443
transform 1 0 29200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5210
timestamp 1654712443
transform 1 0 26200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5212
timestamp 1654712443
transform 1 0 32200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5213
timestamp 1654712443
transform 1 0 35200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5214
timestamp 1654712443
transform 1 0 38200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5215
timestamp 1654712443
transform 1 0 41200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5216
timestamp 1654712443
transform 1 0 44200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5217
timestamp 1654712443
transform 1 0 47200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5218
timestamp 1654712443
transform 1 0 50200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5219
timestamp 1654712443
transform 1 0 53200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5221
timestamp 1654712443
transform 1 0 59200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5220
timestamp 1654712443
transform 1 0 56200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5222
timestamp 1654712443
transform 1 0 62200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5223
timestamp 1654712443
transform 1 0 65200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5224
timestamp 1654712443
transform 1 0 68200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5225
timestamp 1654712443
transform 1 0 71200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5226
timestamp 1654712443
transform 1 0 74200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5227
timestamp 1654712443
transform 1 0 77200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5228
timestamp 1654712443
transform 1 0 80200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5229
timestamp 1654712443
transform 1 0 83200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5230
timestamp 1654712443
transform 1 0 86200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5231
timestamp 1654712443
transform 1 0 89200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5232
timestamp 1654712443
transform 1 0 92200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5233
timestamp 1654712443
transform 1 0 95200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5234
timestamp 1654712443
transform 1 0 98200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5235
timestamp 1654712443
transform 1 0 101200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5236
timestamp 1654712443
transform 1 0 104200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5237
timestamp 1654712443
transform 1 0 107200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5238
timestamp 1654712443
transform 1 0 110200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5239
timestamp 1654712443
transform 1 0 113200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5240
timestamp 1654712443
transform 1 0 116200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5242
timestamp 1654712443
transform 1 0 122200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5241
timestamp 1654712443
transform 1 0 119200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5243
timestamp 1654712443
transform 1 0 125200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5244
timestamp 1654712443
transform 1 0 128200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5245
timestamp 1654712443
transform 1 0 131200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5246
timestamp 1654712443
transform 1 0 134200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5247
timestamp 1654712443
transform 1 0 137200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5248
timestamp 1654712443
transform 1 0 140200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5249
timestamp 1654712443
transform 1 0 143200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5250
timestamp 1654712443
transform 1 0 146200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5252
timestamp 1654712443
transform 1 0 152200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5251
timestamp 1654712443
transform 1 0 149200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5253
timestamp 1654712443
transform 1 0 155200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5254
timestamp 1654712443
transform 1 0 158200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5255
timestamp 1654712443
transform 1 0 161200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5256
timestamp 1654712443
transform 1 0 164200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5257
timestamp 1654712443
transform 1 0 167200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5258
timestamp 1654712443
transform 1 0 170200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5259
timestamp 1654712443
transform 1 0 173200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5260
timestamp 1654712443
transform 1 0 176200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5261
timestamp 1654712443
transform 1 0 179200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5263
timestamp 1654712443
transform 1 0 185200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5262
timestamp 1654712443
transform 1 0 182200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5264
timestamp 1654712443
transform 1 0 188200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5265
timestamp 1654712443
transform 1 0 191200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5266
timestamp 1654712443
transform 1 0 194200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5267
timestamp 1654712443
transform 1 0 197200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5268
timestamp 1654712443
transform 1 0 200200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5269
timestamp 1654712443
transform 1 0 203200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5270
timestamp 1654712443
transform 1 0 206200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5271
timestamp 1654712443
transform 1 0 209200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5273
timestamp 1654712443
transform 1 0 215200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5272
timestamp 1654712443
transform 1 0 212200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5274
timestamp 1654712443
transform 1 0 218200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5275
timestamp 1654712443
transform 1 0 221200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5276
timestamp 1654712443
transform 1 0 224200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5277
timestamp 1654712443
transform 1 0 227200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5278
timestamp 1654712443
transform 1 0 230200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5279
timestamp 1654712443
transform 1 0 233200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5280
timestamp 1654712443
transform 1 0 236200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5281
timestamp 1654712443
transform 1 0 239200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5283
timestamp 1654712443
transform 1 0 245200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5282
timestamp 1654712443
transform 1 0 242200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5284
timestamp 1654712443
transform 1 0 248200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5285
timestamp 1654712443
transform 1 0 251200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5286
timestamp 1654712443
transform 1 0 254200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5287
timestamp 1654712443
transform 1 0 257200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5288
timestamp 1654712443
transform 1 0 260200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5289
timestamp 1654712443
transform 1 0 263200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5290
timestamp 1654712443
transform 1 0 266200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5291
timestamp 1654712443
transform 1 0 269200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5292
timestamp 1654712443
transform 1 0 272200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5294
timestamp 1654712443
transform 1 0 278200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5293
timestamp 1654712443
transform 1 0 275200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5295
timestamp 1654712443
transform 1 0 281200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5296
timestamp 1654712443
transform 1 0 284200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5297
timestamp 1654712443
transform 1 0 287200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5298
timestamp 1654712443
transform 1 0 290200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5299
timestamp 1654712443
transform 1 0 293200 0 1 -153300
box 3640 -2860 6960 460
use pixel  pixel_5101
timestamp 1654712443
transform 1 0 -800 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5100
timestamp 1654712443
transform 1 0 -3800 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5102
timestamp 1654712443
transform 1 0 2200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5103
timestamp 1654712443
transform 1 0 5200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5104
timestamp 1654712443
transform 1 0 8200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5105
timestamp 1654712443
transform 1 0 11200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5106
timestamp 1654712443
transform 1 0 14200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5107
timestamp 1654712443
transform 1 0 17200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5108
timestamp 1654712443
transform 1 0 20200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5109
timestamp 1654712443
transform 1 0 23200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5111
timestamp 1654712443
transform 1 0 29200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5110
timestamp 1654712443
transform 1 0 26200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5112
timestamp 1654712443
transform 1 0 32200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5113
timestamp 1654712443
transform 1 0 35200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5114
timestamp 1654712443
transform 1 0 38200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5115
timestamp 1654712443
transform 1 0 41200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5116
timestamp 1654712443
transform 1 0 44200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5117
timestamp 1654712443
transform 1 0 47200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5118
timestamp 1654712443
transform 1 0 50200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5119
timestamp 1654712443
transform 1 0 53200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5121
timestamp 1654712443
transform 1 0 59200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5120
timestamp 1654712443
transform 1 0 56200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5122
timestamp 1654712443
transform 1 0 62200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5123
timestamp 1654712443
transform 1 0 65200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5124
timestamp 1654712443
transform 1 0 68200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5125
timestamp 1654712443
transform 1 0 71200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5126
timestamp 1654712443
transform 1 0 74200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5127
timestamp 1654712443
transform 1 0 77200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5128
timestamp 1654712443
transform 1 0 80200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5129
timestamp 1654712443
transform 1 0 83200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5130
timestamp 1654712443
transform 1 0 86200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5131
timestamp 1654712443
transform 1 0 89200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5132
timestamp 1654712443
transform 1 0 92200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5133
timestamp 1654712443
transform 1 0 95200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5134
timestamp 1654712443
transform 1 0 98200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5135
timestamp 1654712443
transform 1 0 101200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5136
timestamp 1654712443
transform 1 0 104200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5137
timestamp 1654712443
transform 1 0 107200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5138
timestamp 1654712443
transform 1 0 110200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5139
timestamp 1654712443
transform 1 0 113200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5140
timestamp 1654712443
transform 1 0 116200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5142
timestamp 1654712443
transform 1 0 122200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5141
timestamp 1654712443
transform 1 0 119200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5143
timestamp 1654712443
transform 1 0 125200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5144
timestamp 1654712443
transform 1 0 128200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5145
timestamp 1654712443
transform 1 0 131200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5146
timestamp 1654712443
transform 1 0 134200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5147
timestamp 1654712443
transform 1 0 137200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5148
timestamp 1654712443
transform 1 0 140200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5149
timestamp 1654712443
transform 1 0 143200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5150
timestamp 1654712443
transform 1 0 146200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5152
timestamp 1654712443
transform 1 0 152200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5151
timestamp 1654712443
transform 1 0 149200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5153
timestamp 1654712443
transform 1 0 155200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5154
timestamp 1654712443
transform 1 0 158200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5155
timestamp 1654712443
transform 1 0 161200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5156
timestamp 1654712443
transform 1 0 164200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5157
timestamp 1654712443
transform 1 0 167200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5158
timestamp 1654712443
transform 1 0 170200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5159
timestamp 1654712443
transform 1 0 173200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5160
timestamp 1654712443
transform 1 0 176200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5161
timestamp 1654712443
transform 1 0 179200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5163
timestamp 1654712443
transform 1 0 185200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5162
timestamp 1654712443
transform 1 0 182200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5164
timestamp 1654712443
transform 1 0 188200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5165
timestamp 1654712443
transform 1 0 191200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5166
timestamp 1654712443
transform 1 0 194200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5167
timestamp 1654712443
transform 1 0 197200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5168
timestamp 1654712443
transform 1 0 200200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5169
timestamp 1654712443
transform 1 0 203200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5170
timestamp 1654712443
transform 1 0 206200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5171
timestamp 1654712443
transform 1 0 209200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5173
timestamp 1654712443
transform 1 0 215200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5172
timestamp 1654712443
transform 1 0 212200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5174
timestamp 1654712443
transform 1 0 218200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5175
timestamp 1654712443
transform 1 0 221200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5176
timestamp 1654712443
transform 1 0 224200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5177
timestamp 1654712443
transform 1 0 227200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5178
timestamp 1654712443
transform 1 0 230200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5179
timestamp 1654712443
transform 1 0 233200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5180
timestamp 1654712443
transform 1 0 236200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5181
timestamp 1654712443
transform 1 0 239200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5183
timestamp 1654712443
transform 1 0 245200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5182
timestamp 1654712443
transform 1 0 242200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5184
timestamp 1654712443
transform 1 0 248200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5185
timestamp 1654712443
transform 1 0 251200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5186
timestamp 1654712443
transform 1 0 254200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5187
timestamp 1654712443
transform 1 0 257200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5188
timestamp 1654712443
transform 1 0 260200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5189
timestamp 1654712443
transform 1 0 263200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5190
timestamp 1654712443
transform 1 0 266200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5191
timestamp 1654712443
transform 1 0 269200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5192
timestamp 1654712443
transform 1 0 272200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5194
timestamp 1654712443
transform 1 0 278200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5193
timestamp 1654712443
transform 1 0 275200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5195
timestamp 1654712443
transform 1 0 281200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5196
timestamp 1654712443
transform 1 0 284200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5197
timestamp 1654712443
transform 1 0 287200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5198
timestamp 1654712443
transform 1 0 290200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5199
timestamp 1654712443
transform 1 0 293200 0 1 -150300
box 3640 -2860 6960 460
use pixel  pixel_5001
timestamp 1654712443
transform 1 0 -800 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5000
timestamp 1654712443
transform 1 0 -3800 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5002
timestamp 1654712443
transform 1 0 2200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5003
timestamp 1654712443
transform 1 0 5200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5004
timestamp 1654712443
transform 1 0 8200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5005
timestamp 1654712443
transform 1 0 11200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5006
timestamp 1654712443
transform 1 0 14200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5007
timestamp 1654712443
transform 1 0 17200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5008
timestamp 1654712443
transform 1 0 20200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5009
timestamp 1654712443
transform 1 0 23200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5011
timestamp 1654712443
transform 1 0 29200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5010
timestamp 1654712443
transform 1 0 26200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5012
timestamp 1654712443
transform 1 0 32200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5013
timestamp 1654712443
transform 1 0 35200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5014
timestamp 1654712443
transform 1 0 38200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5015
timestamp 1654712443
transform 1 0 41200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5016
timestamp 1654712443
transform 1 0 44200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5017
timestamp 1654712443
transform 1 0 47200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5018
timestamp 1654712443
transform 1 0 50200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5019
timestamp 1654712443
transform 1 0 53200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5021
timestamp 1654712443
transform 1 0 59200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5020
timestamp 1654712443
transform 1 0 56200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5022
timestamp 1654712443
transform 1 0 62200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5023
timestamp 1654712443
transform 1 0 65200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5024
timestamp 1654712443
transform 1 0 68200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5025
timestamp 1654712443
transform 1 0 71200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5026
timestamp 1654712443
transform 1 0 74200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5027
timestamp 1654712443
transform 1 0 77200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5028
timestamp 1654712443
transform 1 0 80200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5029
timestamp 1654712443
transform 1 0 83200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5030
timestamp 1654712443
transform 1 0 86200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5031
timestamp 1654712443
transform 1 0 89200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5032
timestamp 1654712443
transform 1 0 92200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5033
timestamp 1654712443
transform 1 0 95200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5034
timestamp 1654712443
transform 1 0 98200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5035
timestamp 1654712443
transform 1 0 101200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5036
timestamp 1654712443
transform 1 0 104200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5037
timestamp 1654712443
transform 1 0 107200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5038
timestamp 1654712443
transform 1 0 110200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5039
timestamp 1654712443
transform 1 0 113200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5040
timestamp 1654712443
transform 1 0 116200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5042
timestamp 1654712443
transform 1 0 122200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5041
timestamp 1654712443
transform 1 0 119200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5043
timestamp 1654712443
transform 1 0 125200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5044
timestamp 1654712443
transform 1 0 128200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5045
timestamp 1654712443
transform 1 0 131200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5046
timestamp 1654712443
transform 1 0 134200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5047
timestamp 1654712443
transform 1 0 137200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5048
timestamp 1654712443
transform 1 0 140200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5049
timestamp 1654712443
transform 1 0 143200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5050
timestamp 1654712443
transform 1 0 146200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5052
timestamp 1654712443
transform 1 0 152200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5051
timestamp 1654712443
transform 1 0 149200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5053
timestamp 1654712443
transform 1 0 155200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5054
timestamp 1654712443
transform 1 0 158200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5055
timestamp 1654712443
transform 1 0 161200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5056
timestamp 1654712443
transform 1 0 164200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5057
timestamp 1654712443
transform 1 0 167200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5058
timestamp 1654712443
transform 1 0 170200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5059
timestamp 1654712443
transform 1 0 173200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5060
timestamp 1654712443
transform 1 0 176200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5061
timestamp 1654712443
transform 1 0 179200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5063
timestamp 1654712443
transform 1 0 185200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5062
timestamp 1654712443
transform 1 0 182200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5064
timestamp 1654712443
transform 1 0 188200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5065
timestamp 1654712443
transform 1 0 191200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5066
timestamp 1654712443
transform 1 0 194200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5067
timestamp 1654712443
transform 1 0 197200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5068
timestamp 1654712443
transform 1 0 200200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5069
timestamp 1654712443
transform 1 0 203200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5070
timestamp 1654712443
transform 1 0 206200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5071
timestamp 1654712443
transform 1 0 209200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5073
timestamp 1654712443
transform 1 0 215200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5072
timestamp 1654712443
transform 1 0 212200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5074
timestamp 1654712443
transform 1 0 218200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5075
timestamp 1654712443
transform 1 0 221200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5076
timestamp 1654712443
transform 1 0 224200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5077
timestamp 1654712443
transform 1 0 227200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5078
timestamp 1654712443
transform 1 0 230200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5079
timestamp 1654712443
transform 1 0 233200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5080
timestamp 1654712443
transform 1 0 236200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5081
timestamp 1654712443
transform 1 0 239200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5083
timestamp 1654712443
transform 1 0 245200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5082
timestamp 1654712443
transform 1 0 242200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5084
timestamp 1654712443
transform 1 0 248200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5085
timestamp 1654712443
transform 1 0 251200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5086
timestamp 1654712443
transform 1 0 254200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5087
timestamp 1654712443
transform 1 0 257200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5088
timestamp 1654712443
transform 1 0 260200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5089
timestamp 1654712443
transform 1 0 263200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5090
timestamp 1654712443
transform 1 0 266200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5091
timestamp 1654712443
transform 1 0 269200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5092
timestamp 1654712443
transform 1 0 272200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5094
timestamp 1654712443
transform 1 0 278200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5093
timestamp 1654712443
transform 1 0 275200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5095
timestamp 1654712443
transform 1 0 281200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5096
timestamp 1654712443
transform 1 0 284200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5097
timestamp 1654712443
transform 1 0 287200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5098
timestamp 1654712443
transform 1 0 290200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_5099
timestamp 1654712443
transform 1 0 293200 0 1 -147300
box 3640 -2860 6960 460
use pixel  pixel_4901
timestamp 1654712443
transform 1 0 -800 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4900
timestamp 1654712443
transform 1 0 -3800 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4902
timestamp 1654712443
transform 1 0 2200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4903
timestamp 1654712443
transform 1 0 5200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4904
timestamp 1654712443
transform 1 0 8200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4905
timestamp 1654712443
transform 1 0 11200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4906
timestamp 1654712443
transform 1 0 14200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4907
timestamp 1654712443
transform 1 0 17200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4908
timestamp 1654712443
transform 1 0 20200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4909
timestamp 1654712443
transform 1 0 23200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4911
timestamp 1654712443
transform 1 0 29200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4910
timestamp 1654712443
transform 1 0 26200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4912
timestamp 1654712443
transform 1 0 32200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4913
timestamp 1654712443
transform 1 0 35200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4914
timestamp 1654712443
transform 1 0 38200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4915
timestamp 1654712443
transform 1 0 41200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4916
timestamp 1654712443
transform 1 0 44200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4917
timestamp 1654712443
transform 1 0 47200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4918
timestamp 1654712443
transform 1 0 50200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4919
timestamp 1654712443
transform 1 0 53200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4921
timestamp 1654712443
transform 1 0 59200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4920
timestamp 1654712443
transform 1 0 56200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4922
timestamp 1654712443
transform 1 0 62200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4923
timestamp 1654712443
transform 1 0 65200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4924
timestamp 1654712443
transform 1 0 68200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4925
timestamp 1654712443
transform 1 0 71200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4926
timestamp 1654712443
transform 1 0 74200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4927
timestamp 1654712443
transform 1 0 77200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4928
timestamp 1654712443
transform 1 0 80200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4929
timestamp 1654712443
transform 1 0 83200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4930
timestamp 1654712443
transform 1 0 86200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4931
timestamp 1654712443
transform 1 0 89200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4932
timestamp 1654712443
transform 1 0 92200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4933
timestamp 1654712443
transform 1 0 95200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4934
timestamp 1654712443
transform 1 0 98200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4935
timestamp 1654712443
transform 1 0 101200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4936
timestamp 1654712443
transform 1 0 104200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4937
timestamp 1654712443
transform 1 0 107200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4938
timestamp 1654712443
transform 1 0 110200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4939
timestamp 1654712443
transform 1 0 113200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4940
timestamp 1654712443
transform 1 0 116200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4942
timestamp 1654712443
transform 1 0 122200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4941
timestamp 1654712443
transform 1 0 119200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4943
timestamp 1654712443
transform 1 0 125200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4944
timestamp 1654712443
transform 1 0 128200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4945
timestamp 1654712443
transform 1 0 131200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4946
timestamp 1654712443
transform 1 0 134200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4947
timestamp 1654712443
transform 1 0 137200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4948
timestamp 1654712443
transform 1 0 140200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4949
timestamp 1654712443
transform 1 0 143200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4950
timestamp 1654712443
transform 1 0 146200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4952
timestamp 1654712443
transform 1 0 152200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4951
timestamp 1654712443
transform 1 0 149200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4953
timestamp 1654712443
transform 1 0 155200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4954
timestamp 1654712443
transform 1 0 158200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4955
timestamp 1654712443
transform 1 0 161200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4956
timestamp 1654712443
transform 1 0 164200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4957
timestamp 1654712443
transform 1 0 167200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4958
timestamp 1654712443
transform 1 0 170200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4959
timestamp 1654712443
transform 1 0 173200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4960
timestamp 1654712443
transform 1 0 176200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4961
timestamp 1654712443
transform 1 0 179200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4963
timestamp 1654712443
transform 1 0 185200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4962
timestamp 1654712443
transform 1 0 182200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4964
timestamp 1654712443
transform 1 0 188200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4965
timestamp 1654712443
transform 1 0 191200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4966
timestamp 1654712443
transform 1 0 194200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4967
timestamp 1654712443
transform 1 0 197200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4968
timestamp 1654712443
transform 1 0 200200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4969
timestamp 1654712443
transform 1 0 203200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4970
timestamp 1654712443
transform 1 0 206200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4971
timestamp 1654712443
transform 1 0 209200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4973
timestamp 1654712443
transform 1 0 215200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4972
timestamp 1654712443
transform 1 0 212200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4974
timestamp 1654712443
transform 1 0 218200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4975
timestamp 1654712443
transform 1 0 221200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4976
timestamp 1654712443
transform 1 0 224200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4977
timestamp 1654712443
transform 1 0 227200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4978
timestamp 1654712443
transform 1 0 230200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4979
timestamp 1654712443
transform 1 0 233200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4980
timestamp 1654712443
transform 1 0 236200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4981
timestamp 1654712443
transform 1 0 239200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4983
timestamp 1654712443
transform 1 0 245200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4982
timestamp 1654712443
transform 1 0 242200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4984
timestamp 1654712443
transform 1 0 248200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4985
timestamp 1654712443
transform 1 0 251200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4986
timestamp 1654712443
transform 1 0 254200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4987
timestamp 1654712443
transform 1 0 257200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4988
timestamp 1654712443
transform 1 0 260200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4989
timestamp 1654712443
transform 1 0 263200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4990
timestamp 1654712443
transform 1 0 266200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4991
timestamp 1654712443
transform 1 0 269200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4992
timestamp 1654712443
transform 1 0 272200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4994
timestamp 1654712443
transform 1 0 278200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4993
timestamp 1654712443
transform 1 0 275200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4995
timestamp 1654712443
transform 1 0 281200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4996
timestamp 1654712443
transform 1 0 284200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4997
timestamp 1654712443
transform 1 0 287200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4998
timestamp 1654712443
transform 1 0 290200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4999
timestamp 1654712443
transform 1 0 293200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_4701
timestamp 1654712443
transform 1 0 -800 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4801
timestamp 1654712443
transform 1 0 -800 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4700
timestamp 1654712443
transform 1 0 -3800 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4800
timestamp 1654712443
transform 1 0 -3800 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4702
timestamp 1654712443
transform 1 0 2200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4802
timestamp 1654712443
transform 1 0 2200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4703
timestamp 1654712443
transform 1 0 5200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4803
timestamp 1654712443
transform 1 0 5200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4704
timestamp 1654712443
transform 1 0 8200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4804
timestamp 1654712443
transform 1 0 8200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4705
timestamp 1654712443
transform 1 0 11200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4805
timestamp 1654712443
transform 1 0 11200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4706
timestamp 1654712443
transform 1 0 14200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4806
timestamp 1654712443
transform 1 0 14200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4707
timestamp 1654712443
transform 1 0 17200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4807
timestamp 1654712443
transform 1 0 17200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4708
timestamp 1654712443
transform 1 0 20200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4808
timestamp 1654712443
transform 1 0 20200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4709
timestamp 1654712443
transform 1 0 23200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4809
timestamp 1654712443
transform 1 0 23200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4711
timestamp 1654712443
transform 1 0 29200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4811
timestamp 1654712443
transform 1 0 29200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4710
timestamp 1654712443
transform 1 0 26200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4810
timestamp 1654712443
transform 1 0 26200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4712
timestamp 1654712443
transform 1 0 32200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4812
timestamp 1654712443
transform 1 0 32200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4713
timestamp 1654712443
transform 1 0 35200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4813
timestamp 1654712443
transform 1 0 35200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4714
timestamp 1654712443
transform 1 0 38200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4814
timestamp 1654712443
transform 1 0 38200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4715
timestamp 1654712443
transform 1 0 41200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4815
timestamp 1654712443
transform 1 0 41200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4716
timestamp 1654712443
transform 1 0 44200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4816
timestamp 1654712443
transform 1 0 44200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4717
timestamp 1654712443
transform 1 0 47200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4817
timestamp 1654712443
transform 1 0 47200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4718
timestamp 1654712443
transform 1 0 50200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4818
timestamp 1654712443
transform 1 0 50200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4719
timestamp 1654712443
transform 1 0 53200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4819
timestamp 1654712443
transform 1 0 53200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4721
timestamp 1654712443
transform 1 0 59200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4821
timestamp 1654712443
transform 1 0 59200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4720
timestamp 1654712443
transform 1 0 56200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4820
timestamp 1654712443
transform 1 0 56200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4722
timestamp 1654712443
transform 1 0 62200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4822
timestamp 1654712443
transform 1 0 62200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4723
timestamp 1654712443
transform 1 0 65200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4823
timestamp 1654712443
transform 1 0 65200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4724
timestamp 1654712443
transform 1 0 68200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4824
timestamp 1654712443
transform 1 0 68200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4725
timestamp 1654712443
transform 1 0 71200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4825
timestamp 1654712443
transform 1 0 71200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4726
timestamp 1654712443
transform 1 0 74200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4826
timestamp 1654712443
transform 1 0 74200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4727
timestamp 1654712443
transform 1 0 77200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4827
timestamp 1654712443
transform 1 0 77200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4728
timestamp 1654712443
transform 1 0 80200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4828
timestamp 1654712443
transform 1 0 80200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4729
timestamp 1654712443
transform 1 0 83200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4829
timestamp 1654712443
transform 1 0 83200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4730
timestamp 1654712443
transform 1 0 86200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4830
timestamp 1654712443
transform 1 0 86200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4731
timestamp 1654712443
transform 1 0 89200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4732
timestamp 1654712443
transform 1 0 92200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4831
timestamp 1654712443
transform 1 0 89200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4832
timestamp 1654712443
transform 1 0 92200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4733
timestamp 1654712443
transform 1 0 95200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4833
timestamp 1654712443
transform 1 0 95200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4734
timestamp 1654712443
transform 1 0 98200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4834
timestamp 1654712443
transform 1 0 98200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4735
timestamp 1654712443
transform 1 0 101200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4835
timestamp 1654712443
transform 1 0 101200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4736
timestamp 1654712443
transform 1 0 104200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4836
timestamp 1654712443
transform 1 0 104200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4737
timestamp 1654712443
transform 1 0 107200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4837
timestamp 1654712443
transform 1 0 107200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4738
timestamp 1654712443
transform 1 0 110200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4838
timestamp 1654712443
transform 1 0 110200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4739
timestamp 1654712443
transform 1 0 113200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4839
timestamp 1654712443
transform 1 0 113200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4740
timestamp 1654712443
transform 1 0 116200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4840
timestamp 1654712443
transform 1 0 116200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4742
timestamp 1654712443
transform 1 0 122200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4842
timestamp 1654712443
transform 1 0 122200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4741
timestamp 1654712443
transform 1 0 119200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4841
timestamp 1654712443
transform 1 0 119200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4743
timestamp 1654712443
transform 1 0 125200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4843
timestamp 1654712443
transform 1 0 125200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4744
timestamp 1654712443
transform 1 0 128200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4844
timestamp 1654712443
transform 1 0 128200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4745
timestamp 1654712443
transform 1 0 131200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4845
timestamp 1654712443
transform 1 0 131200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4746
timestamp 1654712443
transform 1 0 134200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4846
timestamp 1654712443
transform 1 0 134200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4747
timestamp 1654712443
transform 1 0 137200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4847
timestamp 1654712443
transform 1 0 137200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4748
timestamp 1654712443
transform 1 0 140200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4848
timestamp 1654712443
transform 1 0 140200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4749
timestamp 1654712443
transform 1 0 143200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4849
timestamp 1654712443
transform 1 0 143200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4750
timestamp 1654712443
transform 1 0 146200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4850
timestamp 1654712443
transform 1 0 146200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4752
timestamp 1654712443
transform 1 0 152200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4852
timestamp 1654712443
transform 1 0 152200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4751
timestamp 1654712443
transform 1 0 149200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4851
timestamp 1654712443
transform 1 0 149200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4753
timestamp 1654712443
transform 1 0 155200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4853
timestamp 1654712443
transform 1 0 155200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4754
timestamp 1654712443
transform 1 0 158200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4854
timestamp 1654712443
transform 1 0 158200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4755
timestamp 1654712443
transform 1 0 161200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4855
timestamp 1654712443
transform 1 0 161200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4756
timestamp 1654712443
transform 1 0 164200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4856
timestamp 1654712443
transform 1 0 164200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4757
timestamp 1654712443
transform 1 0 167200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4857
timestamp 1654712443
transform 1 0 167200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4758
timestamp 1654712443
transform 1 0 170200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4858
timestamp 1654712443
transform 1 0 170200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4759
timestamp 1654712443
transform 1 0 173200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4859
timestamp 1654712443
transform 1 0 173200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4760
timestamp 1654712443
transform 1 0 176200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4860
timestamp 1654712443
transform 1 0 176200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4761
timestamp 1654712443
transform 1 0 179200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4861
timestamp 1654712443
transform 1 0 179200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4763
timestamp 1654712443
transform 1 0 185200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4863
timestamp 1654712443
transform 1 0 185200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4762
timestamp 1654712443
transform 1 0 182200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4862
timestamp 1654712443
transform 1 0 182200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4764
timestamp 1654712443
transform 1 0 188200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4864
timestamp 1654712443
transform 1 0 188200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4765
timestamp 1654712443
transform 1 0 191200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4865
timestamp 1654712443
transform 1 0 191200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4766
timestamp 1654712443
transform 1 0 194200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4866
timestamp 1654712443
transform 1 0 194200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4767
timestamp 1654712443
transform 1 0 197200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4867
timestamp 1654712443
transform 1 0 197200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4768
timestamp 1654712443
transform 1 0 200200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4868
timestamp 1654712443
transform 1 0 200200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4769
timestamp 1654712443
transform 1 0 203200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4869
timestamp 1654712443
transform 1 0 203200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4770
timestamp 1654712443
transform 1 0 206200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4870
timestamp 1654712443
transform 1 0 206200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4771
timestamp 1654712443
transform 1 0 209200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4871
timestamp 1654712443
transform 1 0 209200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4773
timestamp 1654712443
transform 1 0 215200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4873
timestamp 1654712443
transform 1 0 215200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4772
timestamp 1654712443
transform 1 0 212200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4872
timestamp 1654712443
transform 1 0 212200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4774
timestamp 1654712443
transform 1 0 218200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4874
timestamp 1654712443
transform 1 0 218200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4775
timestamp 1654712443
transform 1 0 221200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4875
timestamp 1654712443
transform 1 0 221200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4776
timestamp 1654712443
transform 1 0 224200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4876
timestamp 1654712443
transform 1 0 224200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4777
timestamp 1654712443
transform 1 0 227200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4877
timestamp 1654712443
transform 1 0 227200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4778
timestamp 1654712443
transform 1 0 230200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4878
timestamp 1654712443
transform 1 0 230200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4779
timestamp 1654712443
transform 1 0 233200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4879
timestamp 1654712443
transform 1 0 233200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4780
timestamp 1654712443
transform 1 0 236200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4880
timestamp 1654712443
transform 1 0 236200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4781
timestamp 1654712443
transform 1 0 239200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4881
timestamp 1654712443
transform 1 0 239200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4783
timestamp 1654712443
transform 1 0 245200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4883
timestamp 1654712443
transform 1 0 245200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4782
timestamp 1654712443
transform 1 0 242200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4882
timestamp 1654712443
transform 1 0 242200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4784
timestamp 1654712443
transform 1 0 248200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4884
timestamp 1654712443
transform 1 0 248200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4785
timestamp 1654712443
transform 1 0 251200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4885
timestamp 1654712443
transform 1 0 251200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4786
timestamp 1654712443
transform 1 0 254200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4886
timestamp 1654712443
transform 1 0 254200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4787
timestamp 1654712443
transform 1 0 257200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4887
timestamp 1654712443
transform 1 0 257200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4788
timestamp 1654712443
transform 1 0 260200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4888
timestamp 1654712443
transform 1 0 260200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4789
timestamp 1654712443
transform 1 0 263200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4889
timestamp 1654712443
transform 1 0 263200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4790
timestamp 1654712443
transform 1 0 266200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4890
timestamp 1654712443
transform 1 0 266200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4791
timestamp 1654712443
transform 1 0 269200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4891
timestamp 1654712443
transform 1 0 269200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4792
timestamp 1654712443
transform 1 0 272200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4892
timestamp 1654712443
transform 1 0 272200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4794
timestamp 1654712443
transform 1 0 278200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4894
timestamp 1654712443
transform 1 0 278200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4793
timestamp 1654712443
transform 1 0 275200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4893
timestamp 1654712443
transform 1 0 275200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4795
timestamp 1654712443
transform 1 0 281200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4895
timestamp 1654712443
transform 1 0 281200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4796
timestamp 1654712443
transform 1 0 284200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4896
timestamp 1654712443
transform 1 0 284200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4797
timestamp 1654712443
transform 1 0 287200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4897
timestamp 1654712443
transform 1 0 287200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4798
timestamp 1654712443
transform 1 0 290200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4898
timestamp 1654712443
transform 1 0 290200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4799
timestamp 1654712443
transform 1 0 293200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_4899
timestamp 1654712443
transform 1 0 293200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_4601
timestamp 1654712443
transform 1 0 -800 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4600
timestamp 1654712443
transform 1 0 -3800 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4602
timestamp 1654712443
transform 1 0 2200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4603
timestamp 1654712443
transform 1 0 5200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4604
timestamp 1654712443
transform 1 0 8200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4605
timestamp 1654712443
transform 1 0 11200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4606
timestamp 1654712443
transform 1 0 14200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4607
timestamp 1654712443
transform 1 0 17200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4608
timestamp 1654712443
transform 1 0 20200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4609
timestamp 1654712443
transform 1 0 23200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4611
timestamp 1654712443
transform 1 0 29200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4610
timestamp 1654712443
transform 1 0 26200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4612
timestamp 1654712443
transform 1 0 32200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4613
timestamp 1654712443
transform 1 0 35200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4614
timestamp 1654712443
transform 1 0 38200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4615
timestamp 1654712443
transform 1 0 41200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4616
timestamp 1654712443
transform 1 0 44200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4617
timestamp 1654712443
transform 1 0 47200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4618
timestamp 1654712443
transform 1 0 50200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4619
timestamp 1654712443
transform 1 0 53200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4621
timestamp 1654712443
transform 1 0 59200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4620
timestamp 1654712443
transform 1 0 56200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4622
timestamp 1654712443
transform 1 0 62200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4623
timestamp 1654712443
transform 1 0 65200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4624
timestamp 1654712443
transform 1 0 68200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4625
timestamp 1654712443
transform 1 0 71200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4626
timestamp 1654712443
transform 1 0 74200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4627
timestamp 1654712443
transform 1 0 77200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4628
timestamp 1654712443
transform 1 0 80200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4629
timestamp 1654712443
transform 1 0 83200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4630
timestamp 1654712443
transform 1 0 86200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4631
timestamp 1654712443
transform 1 0 89200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4632
timestamp 1654712443
transform 1 0 92200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4633
timestamp 1654712443
transform 1 0 95200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4634
timestamp 1654712443
transform 1 0 98200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4635
timestamp 1654712443
transform 1 0 101200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4636
timestamp 1654712443
transform 1 0 104200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4637
timestamp 1654712443
transform 1 0 107200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4638
timestamp 1654712443
transform 1 0 110200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4639
timestamp 1654712443
transform 1 0 113200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4640
timestamp 1654712443
transform 1 0 116200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4642
timestamp 1654712443
transform 1 0 122200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4641
timestamp 1654712443
transform 1 0 119200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4643
timestamp 1654712443
transform 1 0 125200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4644
timestamp 1654712443
transform 1 0 128200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4645
timestamp 1654712443
transform 1 0 131200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4646
timestamp 1654712443
transform 1 0 134200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4647
timestamp 1654712443
transform 1 0 137200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4648
timestamp 1654712443
transform 1 0 140200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4649
timestamp 1654712443
transform 1 0 143200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4650
timestamp 1654712443
transform 1 0 146200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4652
timestamp 1654712443
transform 1 0 152200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4651
timestamp 1654712443
transform 1 0 149200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4653
timestamp 1654712443
transform 1 0 155200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4654
timestamp 1654712443
transform 1 0 158200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4655
timestamp 1654712443
transform 1 0 161200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4656
timestamp 1654712443
transform 1 0 164200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4657
timestamp 1654712443
transform 1 0 167200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4658
timestamp 1654712443
transform 1 0 170200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4659
timestamp 1654712443
transform 1 0 173200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4660
timestamp 1654712443
transform 1 0 176200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4661
timestamp 1654712443
transform 1 0 179200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4663
timestamp 1654712443
transform 1 0 185200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4662
timestamp 1654712443
transform 1 0 182200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4664
timestamp 1654712443
transform 1 0 188200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4665
timestamp 1654712443
transform 1 0 191200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4666
timestamp 1654712443
transform 1 0 194200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4667
timestamp 1654712443
transform 1 0 197200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4668
timestamp 1654712443
transform 1 0 200200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4669
timestamp 1654712443
transform 1 0 203200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4670
timestamp 1654712443
transform 1 0 206200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4671
timestamp 1654712443
transform 1 0 209200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4673
timestamp 1654712443
transform 1 0 215200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4672
timestamp 1654712443
transform 1 0 212200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4674
timestamp 1654712443
transform 1 0 218200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4675
timestamp 1654712443
transform 1 0 221200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4676
timestamp 1654712443
transform 1 0 224200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4677
timestamp 1654712443
transform 1 0 227200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4678
timestamp 1654712443
transform 1 0 230200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4679
timestamp 1654712443
transform 1 0 233200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4680
timestamp 1654712443
transform 1 0 236200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4681
timestamp 1654712443
transform 1 0 239200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4683
timestamp 1654712443
transform 1 0 245200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4682
timestamp 1654712443
transform 1 0 242200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4684
timestamp 1654712443
transform 1 0 248200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4685
timestamp 1654712443
transform 1 0 251200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4686
timestamp 1654712443
transform 1 0 254200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4687
timestamp 1654712443
transform 1 0 257200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4688
timestamp 1654712443
transform 1 0 260200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4689
timestamp 1654712443
transform 1 0 263200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4690
timestamp 1654712443
transform 1 0 266200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4691
timestamp 1654712443
transform 1 0 269200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4692
timestamp 1654712443
transform 1 0 272200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4694
timestamp 1654712443
transform 1 0 278200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4693
timestamp 1654712443
transform 1 0 275200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4695
timestamp 1654712443
transform 1 0 281200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4696
timestamp 1654712443
transform 1 0 284200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4697
timestamp 1654712443
transform 1 0 287200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4698
timestamp 1654712443
transform 1 0 290200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4699
timestamp 1654712443
transform 1 0 293200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_4501
timestamp 1654712443
transform 1 0 -800 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4500
timestamp 1654712443
transform 1 0 -3800 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4502
timestamp 1654712443
transform 1 0 2200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4503
timestamp 1654712443
transform 1 0 5200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4504
timestamp 1654712443
transform 1 0 8200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4505
timestamp 1654712443
transform 1 0 11200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4506
timestamp 1654712443
transform 1 0 14200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4507
timestamp 1654712443
transform 1 0 17200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4508
timestamp 1654712443
transform 1 0 20200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4509
timestamp 1654712443
transform 1 0 23200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4511
timestamp 1654712443
transform 1 0 29200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4510
timestamp 1654712443
transform 1 0 26200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4512
timestamp 1654712443
transform 1 0 32200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4513
timestamp 1654712443
transform 1 0 35200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4514
timestamp 1654712443
transform 1 0 38200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4515
timestamp 1654712443
transform 1 0 41200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4516
timestamp 1654712443
transform 1 0 44200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4517
timestamp 1654712443
transform 1 0 47200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4518
timestamp 1654712443
transform 1 0 50200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4519
timestamp 1654712443
transform 1 0 53200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4521
timestamp 1654712443
transform 1 0 59200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4520
timestamp 1654712443
transform 1 0 56200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4522
timestamp 1654712443
transform 1 0 62200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4523
timestamp 1654712443
transform 1 0 65200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4524
timestamp 1654712443
transform 1 0 68200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4525
timestamp 1654712443
transform 1 0 71200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4526
timestamp 1654712443
transform 1 0 74200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4527
timestamp 1654712443
transform 1 0 77200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4528
timestamp 1654712443
transform 1 0 80200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4529
timestamp 1654712443
transform 1 0 83200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4530
timestamp 1654712443
transform 1 0 86200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4531
timestamp 1654712443
transform 1 0 89200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4532
timestamp 1654712443
transform 1 0 92200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4533
timestamp 1654712443
transform 1 0 95200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4534
timestamp 1654712443
transform 1 0 98200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4535
timestamp 1654712443
transform 1 0 101200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4536
timestamp 1654712443
transform 1 0 104200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4537
timestamp 1654712443
transform 1 0 107200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4538
timestamp 1654712443
transform 1 0 110200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4539
timestamp 1654712443
transform 1 0 113200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4540
timestamp 1654712443
transform 1 0 116200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4542
timestamp 1654712443
transform 1 0 122200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4541
timestamp 1654712443
transform 1 0 119200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4543
timestamp 1654712443
transform 1 0 125200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4544
timestamp 1654712443
transform 1 0 128200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4545
timestamp 1654712443
transform 1 0 131200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4546
timestamp 1654712443
transform 1 0 134200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4547
timestamp 1654712443
transform 1 0 137200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4548
timestamp 1654712443
transform 1 0 140200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4549
timestamp 1654712443
transform 1 0 143200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4550
timestamp 1654712443
transform 1 0 146200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4552
timestamp 1654712443
transform 1 0 152200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4551
timestamp 1654712443
transform 1 0 149200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4553
timestamp 1654712443
transform 1 0 155200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4554
timestamp 1654712443
transform 1 0 158200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4555
timestamp 1654712443
transform 1 0 161200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4556
timestamp 1654712443
transform 1 0 164200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4557
timestamp 1654712443
transform 1 0 167200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4558
timestamp 1654712443
transform 1 0 170200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4559
timestamp 1654712443
transform 1 0 173200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4560
timestamp 1654712443
transform 1 0 176200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4561
timestamp 1654712443
transform 1 0 179200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4563
timestamp 1654712443
transform 1 0 185200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4562
timestamp 1654712443
transform 1 0 182200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4564
timestamp 1654712443
transform 1 0 188200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4565
timestamp 1654712443
transform 1 0 191200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4566
timestamp 1654712443
transform 1 0 194200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4567
timestamp 1654712443
transform 1 0 197200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4568
timestamp 1654712443
transform 1 0 200200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4569
timestamp 1654712443
transform 1 0 203200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4570
timestamp 1654712443
transform 1 0 206200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4571
timestamp 1654712443
transform 1 0 209200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4573
timestamp 1654712443
transform 1 0 215200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4572
timestamp 1654712443
transform 1 0 212200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4574
timestamp 1654712443
transform 1 0 218200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4575
timestamp 1654712443
transform 1 0 221200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4576
timestamp 1654712443
transform 1 0 224200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4577
timestamp 1654712443
transform 1 0 227200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4578
timestamp 1654712443
transform 1 0 230200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4579
timestamp 1654712443
transform 1 0 233200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4580
timestamp 1654712443
transform 1 0 236200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4581
timestamp 1654712443
transform 1 0 239200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4583
timestamp 1654712443
transform 1 0 245200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4582
timestamp 1654712443
transform 1 0 242200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4584
timestamp 1654712443
transform 1 0 248200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4585
timestamp 1654712443
transform 1 0 251200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4586
timestamp 1654712443
transform 1 0 254200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4587
timestamp 1654712443
transform 1 0 257200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4588
timestamp 1654712443
transform 1 0 260200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4589
timestamp 1654712443
transform 1 0 263200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4590
timestamp 1654712443
transform 1 0 266200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4591
timestamp 1654712443
transform 1 0 269200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4592
timestamp 1654712443
transform 1 0 272200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4594
timestamp 1654712443
transform 1 0 278200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4593
timestamp 1654712443
transform 1 0 275200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4595
timestamp 1654712443
transform 1 0 281200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4596
timestamp 1654712443
transform 1 0 284200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4597
timestamp 1654712443
transform 1 0 287200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4598
timestamp 1654712443
transform 1 0 290200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4599
timestamp 1654712443
transform 1 0 293200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_4401
timestamp 1654712443
transform 1 0 -800 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4400
timestamp 1654712443
transform 1 0 -3800 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4402
timestamp 1654712443
transform 1 0 2200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4403
timestamp 1654712443
transform 1 0 5200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4404
timestamp 1654712443
transform 1 0 8200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4405
timestamp 1654712443
transform 1 0 11200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4406
timestamp 1654712443
transform 1 0 14200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4407
timestamp 1654712443
transform 1 0 17200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4408
timestamp 1654712443
transform 1 0 20200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4409
timestamp 1654712443
transform 1 0 23200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4411
timestamp 1654712443
transform 1 0 29200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4410
timestamp 1654712443
transform 1 0 26200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4412
timestamp 1654712443
transform 1 0 32200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4413
timestamp 1654712443
transform 1 0 35200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4414
timestamp 1654712443
transform 1 0 38200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4415
timestamp 1654712443
transform 1 0 41200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4416
timestamp 1654712443
transform 1 0 44200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4417
timestamp 1654712443
transform 1 0 47200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4418
timestamp 1654712443
transform 1 0 50200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4419
timestamp 1654712443
transform 1 0 53200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4421
timestamp 1654712443
transform 1 0 59200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4420
timestamp 1654712443
transform 1 0 56200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4422
timestamp 1654712443
transform 1 0 62200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4423
timestamp 1654712443
transform 1 0 65200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4424
timestamp 1654712443
transform 1 0 68200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4425
timestamp 1654712443
transform 1 0 71200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4426
timestamp 1654712443
transform 1 0 74200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4427
timestamp 1654712443
transform 1 0 77200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4428
timestamp 1654712443
transform 1 0 80200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4429
timestamp 1654712443
transform 1 0 83200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4430
timestamp 1654712443
transform 1 0 86200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4431
timestamp 1654712443
transform 1 0 89200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4432
timestamp 1654712443
transform 1 0 92200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4433
timestamp 1654712443
transform 1 0 95200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4434
timestamp 1654712443
transform 1 0 98200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4435
timestamp 1654712443
transform 1 0 101200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4436
timestamp 1654712443
transform 1 0 104200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4437
timestamp 1654712443
transform 1 0 107200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4438
timestamp 1654712443
transform 1 0 110200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4439
timestamp 1654712443
transform 1 0 113200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4440
timestamp 1654712443
transform 1 0 116200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4442
timestamp 1654712443
transform 1 0 122200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4441
timestamp 1654712443
transform 1 0 119200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4443
timestamp 1654712443
transform 1 0 125200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4444
timestamp 1654712443
transform 1 0 128200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4445
timestamp 1654712443
transform 1 0 131200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4446
timestamp 1654712443
transform 1 0 134200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4447
timestamp 1654712443
transform 1 0 137200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4448
timestamp 1654712443
transform 1 0 140200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4449
timestamp 1654712443
transform 1 0 143200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4450
timestamp 1654712443
transform 1 0 146200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4452
timestamp 1654712443
transform 1 0 152200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4451
timestamp 1654712443
transform 1 0 149200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4453
timestamp 1654712443
transform 1 0 155200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4454
timestamp 1654712443
transform 1 0 158200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4455
timestamp 1654712443
transform 1 0 161200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4456
timestamp 1654712443
transform 1 0 164200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4457
timestamp 1654712443
transform 1 0 167200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4458
timestamp 1654712443
transform 1 0 170200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4459
timestamp 1654712443
transform 1 0 173200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4460
timestamp 1654712443
transform 1 0 176200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4461
timestamp 1654712443
transform 1 0 179200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4463
timestamp 1654712443
transform 1 0 185200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4462
timestamp 1654712443
transform 1 0 182200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4464
timestamp 1654712443
transform 1 0 188200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4465
timestamp 1654712443
transform 1 0 191200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4466
timestamp 1654712443
transform 1 0 194200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4467
timestamp 1654712443
transform 1 0 197200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4468
timestamp 1654712443
transform 1 0 200200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4469
timestamp 1654712443
transform 1 0 203200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4470
timestamp 1654712443
transform 1 0 206200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4471
timestamp 1654712443
transform 1 0 209200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4473
timestamp 1654712443
transform 1 0 215200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4472
timestamp 1654712443
transform 1 0 212200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4474
timestamp 1654712443
transform 1 0 218200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4475
timestamp 1654712443
transform 1 0 221200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4476
timestamp 1654712443
transform 1 0 224200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4477
timestamp 1654712443
transform 1 0 227200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4478
timestamp 1654712443
transform 1 0 230200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4479
timestamp 1654712443
transform 1 0 233200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4480
timestamp 1654712443
transform 1 0 236200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4481
timestamp 1654712443
transform 1 0 239200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4483
timestamp 1654712443
transform 1 0 245200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4482
timestamp 1654712443
transform 1 0 242200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4484
timestamp 1654712443
transform 1 0 248200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4485
timestamp 1654712443
transform 1 0 251200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4486
timestamp 1654712443
transform 1 0 254200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4487
timestamp 1654712443
transform 1 0 257200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4488
timestamp 1654712443
transform 1 0 260200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4489
timestamp 1654712443
transform 1 0 263200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4490
timestamp 1654712443
transform 1 0 266200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4491
timestamp 1654712443
transform 1 0 269200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4492
timestamp 1654712443
transform 1 0 272200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4494
timestamp 1654712443
transform 1 0 278200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4493
timestamp 1654712443
transform 1 0 275200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4495
timestamp 1654712443
transform 1 0 281200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4496
timestamp 1654712443
transform 1 0 284200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4497
timestamp 1654712443
transform 1 0 287200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4498
timestamp 1654712443
transform 1 0 290200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4499
timestamp 1654712443
transform 1 0 293200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_4301
timestamp 1654712443
transform 1 0 -800 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4300
timestamp 1654712443
transform 1 0 -3800 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4302
timestamp 1654712443
transform 1 0 2200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4303
timestamp 1654712443
transform 1 0 5200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4304
timestamp 1654712443
transform 1 0 8200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4305
timestamp 1654712443
transform 1 0 11200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4306
timestamp 1654712443
transform 1 0 14200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4307
timestamp 1654712443
transform 1 0 17200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4308
timestamp 1654712443
transform 1 0 20200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4309
timestamp 1654712443
transform 1 0 23200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4311
timestamp 1654712443
transform 1 0 29200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4310
timestamp 1654712443
transform 1 0 26200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4312
timestamp 1654712443
transform 1 0 32200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4313
timestamp 1654712443
transform 1 0 35200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4314
timestamp 1654712443
transform 1 0 38200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4315
timestamp 1654712443
transform 1 0 41200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4316
timestamp 1654712443
transform 1 0 44200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4317
timestamp 1654712443
transform 1 0 47200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4318
timestamp 1654712443
transform 1 0 50200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4319
timestamp 1654712443
transform 1 0 53200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4321
timestamp 1654712443
transform 1 0 59200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4320
timestamp 1654712443
transform 1 0 56200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4322
timestamp 1654712443
transform 1 0 62200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4323
timestamp 1654712443
transform 1 0 65200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4324
timestamp 1654712443
transform 1 0 68200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4325
timestamp 1654712443
transform 1 0 71200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4326
timestamp 1654712443
transform 1 0 74200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4327
timestamp 1654712443
transform 1 0 77200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4328
timestamp 1654712443
transform 1 0 80200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4329
timestamp 1654712443
transform 1 0 83200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4330
timestamp 1654712443
transform 1 0 86200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4331
timestamp 1654712443
transform 1 0 89200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4332
timestamp 1654712443
transform 1 0 92200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4333
timestamp 1654712443
transform 1 0 95200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4334
timestamp 1654712443
transform 1 0 98200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4335
timestamp 1654712443
transform 1 0 101200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4336
timestamp 1654712443
transform 1 0 104200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4337
timestamp 1654712443
transform 1 0 107200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4338
timestamp 1654712443
transform 1 0 110200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4339
timestamp 1654712443
transform 1 0 113200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4340
timestamp 1654712443
transform 1 0 116200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4342
timestamp 1654712443
transform 1 0 122200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4341
timestamp 1654712443
transform 1 0 119200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4343
timestamp 1654712443
transform 1 0 125200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4344
timestamp 1654712443
transform 1 0 128200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4345
timestamp 1654712443
transform 1 0 131200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4346
timestamp 1654712443
transform 1 0 134200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4347
timestamp 1654712443
transform 1 0 137200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4348
timestamp 1654712443
transform 1 0 140200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4349
timestamp 1654712443
transform 1 0 143200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4350
timestamp 1654712443
transform 1 0 146200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4352
timestamp 1654712443
transform 1 0 152200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4351
timestamp 1654712443
transform 1 0 149200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4353
timestamp 1654712443
transform 1 0 155200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4354
timestamp 1654712443
transform 1 0 158200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4355
timestamp 1654712443
transform 1 0 161200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4356
timestamp 1654712443
transform 1 0 164200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4357
timestamp 1654712443
transform 1 0 167200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4358
timestamp 1654712443
transform 1 0 170200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4359
timestamp 1654712443
transform 1 0 173200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4360
timestamp 1654712443
transform 1 0 176200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4361
timestamp 1654712443
transform 1 0 179200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4363
timestamp 1654712443
transform 1 0 185200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4362
timestamp 1654712443
transform 1 0 182200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4364
timestamp 1654712443
transform 1 0 188200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4365
timestamp 1654712443
transform 1 0 191200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4366
timestamp 1654712443
transform 1 0 194200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4367
timestamp 1654712443
transform 1 0 197200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4368
timestamp 1654712443
transform 1 0 200200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4369
timestamp 1654712443
transform 1 0 203200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4370
timestamp 1654712443
transform 1 0 206200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4371
timestamp 1654712443
transform 1 0 209200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4373
timestamp 1654712443
transform 1 0 215200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4372
timestamp 1654712443
transform 1 0 212200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4374
timestamp 1654712443
transform 1 0 218200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4375
timestamp 1654712443
transform 1 0 221200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4376
timestamp 1654712443
transform 1 0 224200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4377
timestamp 1654712443
transform 1 0 227200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4378
timestamp 1654712443
transform 1 0 230200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4379
timestamp 1654712443
transform 1 0 233200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4380
timestamp 1654712443
transform 1 0 236200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4381
timestamp 1654712443
transform 1 0 239200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4383
timestamp 1654712443
transform 1 0 245200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4382
timestamp 1654712443
transform 1 0 242200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4384
timestamp 1654712443
transform 1 0 248200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4385
timestamp 1654712443
transform 1 0 251200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4386
timestamp 1654712443
transform 1 0 254200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4387
timestamp 1654712443
transform 1 0 257200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4388
timestamp 1654712443
transform 1 0 260200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4389
timestamp 1654712443
transform 1 0 263200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4390
timestamp 1654712443
transform 1 0 266200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4391
timestamp 1654712443
transform 1 0 269200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4392
timestamp 1654712443
transform 1 0 272200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4394
timestamp 1654712443
transform 1 0 278200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4393
timestamp 1654712443
transform 1 0 275200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4395
timestamp 1654712443
transform 1 0 281200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4396
timestamp 1654712443
transform 1 0 284200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4397
timestamp 1654712443
transform 1 0 287200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4398
timestamp 1654712443
transform 1 0 290200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4399
timestamp 1654712443
transform 1 0 293200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_4201
timestamp 1654712443
transform 1 0 -800 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4200
timestamp 1654712443
transform 1 0 -3800 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4202
timestamp 1654712443
transform 1 0 2200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4203
timestamp 1654712443
transform 1 0 5200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4204
timestamp 1654712443
transform 1 0 8200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4205
timestamp 1654712443
transform 1 0 11200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4206
timestamp 1654712443
transform 1 0 14200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4207
timestamp 1654712443
transform 1 0 17200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4208
timestamp 1654712443
transform 1 0 20200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4209
timestamp 1654712443
transform 1 0 23200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4211
timestamp 1654712443
transform 1 0 29200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4210
timestamp 1654712443
transform 1 0 26200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4212
timestamp 1654712443
transform 1 0 32200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4213
timestamp 1654712443
transform 1 0 35200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4214
timestamp 1654712443
transform 1 0 38200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4215
timestamp 1654712443
transform 1 0 41200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4216
timestamp 1654712443
transform 1 0 44200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4217
timestamp 1654712443
transform 1 0 47200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4218
timestamp 1654712443
transform 1 0 50200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4219
timestamp 1654712443
transform 1 0 53200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4221
timestamp 1654712443
transform 1 0 59200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4220
timestamp 1654712443
transform 1 0 56200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4222
timestamp 1654712443
transform 1 0 62200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4223
timestamp 1654712443
transform 1 0 65200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4224
timestamp 1654712443
transform 1 0 68200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4225
timestamp 1654712443
transform 1 0 71200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4226
timestamp 1654712443
transform 1 0 74200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4227
timestamp 1654712443
transform 1 0 77200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4228
timestamp 1654712443
transform 1 0 80200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4229
timestamp 1654712443
transform 1 0 83200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4230
timestamp 1654712443
transform 1 0 86200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4231
timestamp 1654712443
transform 1 0 89200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4232
timestamp 1654712443
transform 1 0 92200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4233
timestamp 1654712443
transform 1 0 95200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4234
timestamp 1654712443
transform 1 0 98200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4235
timestamp 1654712443
transform 1 0 101200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4236
timestamp 1654712443
transform 1 0 104200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4237
timestamp 1654712443
transform 1 0 107200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4238
timestamp 1654712443
transform 1 0 110200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4239
timestamp 1654712443
transform 1 0 113200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4240
timestamp 1654712443
transform 1 0 116200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4242
timestamp 1654712443
transform 1 0 122200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4241
timestamp 1654712443
transform 1 0 119200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4243
timestamp 1654712443
transform 1 0 125200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4244
timestamp 1654712443
transform 1 0 128200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4245
timestamp 1654712443
transform 1 0 131200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4246
timestamp 1654712443
transform 1 0 134200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4247
timestamp 1654712443
transform 1 0 137200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4248
timestamp 1654712443
transform 1 0 140200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4249
timestamp 1654712443
transform 1 0 143200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4250
timestamp 1654712443
transform 1 0 146200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4252
timestamp 1654712443
transform 1 0 152200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4251
timestamp 1654712443
transform 1 0 149200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4253
timestamp 1654712443
transform 1 0 155200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4254
timestamp 1654712443
transform 1 0 158200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4255
timestamp 1654712443
transform 1 0 161200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4256
timestamp 1654712443
transform 1 0 164200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4257
timestamp 1654712443
transform 1 0 167200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4258
timestamp 1654712443
transform 1 0 170200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4259
timestamp 1654712443
transform 1 0 173200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4260
timestamp 1654712443
transform 1 0 176200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4261
timestamp 1654712443
transform 1 0 179200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4263
timestamp 1654712443
transform 1 0 185200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4262
timestamp 1654712443
transform 1 0 182200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4264
timestamp 1654712443
transform 1 0 188200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4265
timestamp 1654712443
transform 1 0 191200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4266
timestamp 1654712443
transform 1 0 194200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4267
timestamp 1654712443
transform 1 0 197200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4268
timestamp 1654712443
transform 1 0 200200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4269
timestamp 1654712443
transform 1 0 203200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4270
timestamp 1654712443
transform 1 0 206200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4271
timestamp 1654712443
transform 1 0 209200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4273
timestamp 1654712443
transform 1 0 215200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4272
timestamp 1654712443
transform 1 0 212200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4274
timestamp 1654712443
transform 1 0 218200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4275
timestamp 1654712443
transform 1 0 221200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4276
timestamp 1654712443
transform 1 0 224200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4277
timestamp 1654712443
transform 1 0 227200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4278
timestamp 1654712443
transform 1 0 230200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4279
timestamp 1654712443
transform 1 0 233200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4280
timestamp 1654712443
transform 1 0 236200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4281
timestamp 1654712443
transform 1 0 239200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4283
timestamp 1654712443
transform 1 0 245200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4282
timestamp 1654712443
transform 1 0 242200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4284
timestamp 1654712443
transform 1 0 248200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4285
timestamp 1654712443
transform 1 0 251200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4286
timestamp 1654712443
transform 1 0 254200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4287
timestamp 1654712443
transform 1 0 257200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4288
timestamp 1654712443
transform 1 0 260200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4289
timestamp 1654712443
transform 1 0 263200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4290
timestamp 1654712443
transform 1 0 266200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4291
timestamp 1654712443
transform 1 0 269200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4292
timestamp 1654712443
transform 1 0 272200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4294
timestamp 1654712443
transform 1 0 278200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4293
timestamp 1654712443
transform 1 0 275200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4295
timestamp 1654712443
transform 1 0 281200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4296
timestamp 1654712443
transform 1 0 284200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4297
timestamp 1654712443
transform 1 0 287200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4298
timestamp 1654712443
transform 1 0 290200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4299
timestamp 1654712443
transform 1 0 293200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_4101
timestamp 1654712443
transform 1 0 -800 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4100
timestamp 1654712443
transform 1 0 -3800 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4102
timestamp 1654712443
transform 1 0 2200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4103
timestamp 1654712443
transform 1 0 5200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4104
timestamp 1654712443
transform 1 0 8200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4105
timestamp 1654712443
transform 1 0 11200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4106
timestamp 1654712443
transform 1 0 14200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4107
timestamp 1654712443
transform 1 0 17200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4108
timestamp 1654712443
transform 1 0 20200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4109
timestamp 1654712443
transform 1 0 23200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4111
timestamp 1654712443
transform 1 0 29200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4110
timestamp 1654712443
transform 1 0 26200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4112
timestamp 1654712443
transform 1 0 32200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4113
timestamp 1654712443
transform 1 0 35200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4114
timestamp 1654712443
transform 1 0 38200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4115
timestamp 1654712443
transform 1 0 41200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4116
timestamp 1654712443
transform 1 0 44200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4117
timestamp 1654712443
transform 1 0 47200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4118
timestamp 1654712443
transform 1 0 50200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4119
timestamp 1654712443
transform 1 0 53200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4121
timestamp 1654712443
transform 1 0 59200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4120
timestamp 1654712443
transform 1 0 56200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4122
timestamp 1654712443
transform 1 0 62200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4123
timestamp 1654712443
transform 1 0 65200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4124
timestamp 1654712443
transform 1 0 68200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4125
timestamp 1654712443
transform 1 0 71200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4126
timestamp 1654712443
transform 1 0 74200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4127
timestamp 1654712443
transform 1 0 77200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4128
timestamp 1654712443
transform 1 0 80200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4129
timestamp 1654712443
transform 1 0 83200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4130
timestamp 1654712443
transform 1 0 86200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4131
timestamp 1654712443
transform 1 0 89200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4132
timestamp 1654712443
transform 1 0 92200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4133
timestamp 1654712443
transform 1 0 95200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4134
timestamp 1654712443
transform 1 0 98200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4135
timestamp 1654712443
transform 1 0 101200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4136
timestamp 1654712443
transform 1 0 104200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4137
timestamp 1654712443
transform 1 0 107200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4138
timestamp 1654712443
transform 1 0 110200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4139
timestamp 1654712443
transform 1 0 113200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4140
timestamp 1654712443
transform 1 0 116200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4142
timestamp 1654712443
transform 1 0 122200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4141
timestamp 1654712443
transform 1 0 119200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4143
timestamp 1654712443
transform 1 0 125200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4144
timestamp 1654712443
transform 1 0 128200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4145
timestamp 1654712443
transform 1 0 131200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4146
timestamp 1654712443
transform 1 0 134200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4147
timestamp 1654712443
transform 1 0 137200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4148
timestamp 1654712443
transform 1 0 140200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4149
timestamp 1654712443
transform 1 0 143200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4150
timestamp 1654712443
transform 1 0 146200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4152
timestamp 1654712443
transform 1 0 152200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4151
timestamp 1654712443
transform 1 0 149200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4153
timestamp 1654712443
transform 1 0 155200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4154
timestamp 1654712443
transform 1 0 158200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4155
timestamp 1654712443
transform 1 0 161200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4156
timestamp 1654712443
transform 1 0 164200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4157
timestamp 1654712443
transform 1 0 167200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4158
timestamp 1654712443
transform 1 0 170200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4159
timestamp 1654712443
transform 1 0 173200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4160
timestamp 1654712443
transform 1 0 176200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4161
timestamp 1654712443
transform 1 0 179200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4163
timestamp 1654712443
transform 1 0 185200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4162
timestamp 1654712443
transform 1 0 182200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4164
timestamp 1654712443
transform 1 0 188200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4165
timestamp 1654712443
transform 1 0 191200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4166
timestamp 1654712443
transform 1 0 194200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4167
timestamp 1654712443
transform 1 0 197200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4168
timestamp 1654712443
transform 1 0 200200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4169
timestamp 1654712443
transform 1 0 203200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4170
timestamp 1654712443
transform 1 0 206200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4171
timestamp 1654712443
transform 1 0 209200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4173
timestamp 1654712443
transform 1 0 215200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4172
timestamp 1654712443
transform 1 0 212200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4174
timestamp 1654712443
transform 1 0 218200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4175
timestamp 1654712443
transform 1 0 221200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4176
timestamp 1654712443
transform 1 0 224200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4177
timestamp 1654712443
transform 1 0 227200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4178
timestamp 1654712443
transform 1 0 230200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4179
timestamp 1654712443
transform 1 0 233200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4180
timestamp 1654712443
transform 1 0 236200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4181
timestamp 1654712443
transform 1 0 239200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4183
timestamp 1654712443
transform 1 0 245200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4182
timestamp 1654712443
transform 1 0 242200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4184
timestamp 1654712443
transform 1 0 248200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4185
timestamp 1654712443
transform 1 0 251200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4186
timestamp 1654712443
transform 1 0 254200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4187
timestamp 1654712443
transform 1 0 257200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4188
timestamp 1654712443
transform 1 0 260200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4189
timestamp 1654712443
transform 1 0 263200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4190
timestamp 1654712443
transform 1 0 266200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4191
timestamp 1654712443
transform 1 0 269200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4192
timestamp 1654712443
transform 1 0 272200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4194
timestamp 1654712443
transform 1 0 278200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4193
timestamp 1654712443
transform 1 0 275200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4195
timestamp 1654712443
transform 1 0 281200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4196
timestamp 1654712443
transform 1 0 284200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4197
timestamp 1654712443
transform 1 0 287200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4198
timestamp 1654712443
transform 1 0 290200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4199
timestamp 1654712443
transform 1 0 293200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_4001
timestamp 1654712443
transform 1 0 -800 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4000
timestamp 1654712443
transform 1 0 -3800 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4002
timestamp 1654712443
transform 1 0 2200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4003
timestamp 1654712443
transform 1 0 5200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4004
timestamp 1654712443
transform 1 0 8200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4005
timestamp 1654712443
transform 1 0 11200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4006
timestamp 1654712443
transform 1 0 14200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4007
timestamp 1654712443
transform 1 0 17200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4008
timestamp 1654712443
transform 1 0 20200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4009
timestamp 1654712443
transform 1 0 23200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4011
timestamp 1654712443
transform 1 0 29200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4010
timestamp 1654712443
transform 1 0 26200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4012
timestamp 1654712443
transform 1 0 32200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4013
timestamp 1654712443
transform 1 0 35200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4014
timestamp 1654712443
transform 1 0 38200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4015
timestamp 1654712443
transform 1 0 41200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4016
timestamp 1654712443
transform 1 0 44200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4017
timestamp 1654712443
transform 1 0 47200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4018
timestamp 1654712443
transform 1 0 50200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4019
timestamp 1654712443
transform 1 0 53200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4021
timestamp 1654712443
transform 1 0 59200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4020
timestamp 1654712443
transform 1 0 56200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4022
timestamp 1654712443
transform 1 0 62200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4023
timestamp 1654712443
transform 1 0 65200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4024
timestamp 1654712443
transform 1 0 68200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4025
timestamp 1654712443
transform 1 0 71200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4026
timestamp 1654712443
transform 1 0 74200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4027
timestamp 1654712443
transform 1 0 77200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4028
timestamp 1654712443
transform 1 0 80200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4029
timestamp 1654712443
transform 1 0 83200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4030
timestamp 1654712443
transform 1 0 86200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4031
timestamp 1654712443
transform 1 0 89200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4032
timestamp 1654712443
transform 1 0 92200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4033
timestamp 1654712443
transform 1 0 95200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4034
timestamp 1654712443
transform 1 0 98200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4035
timestamp 1654712443
transform 1 0 101200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4036
timestamp 1654712443
transform 1 0 104200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4037
timestamp 1654712443
transform 1 0 107200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4038
timestamp 1654712443
transform 1 0 110200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4039
timestamp 1654712443
transform 1 0 113200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4040
timestamp 1654712443
transform 1 0 116200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4042
timestamp 1654712443
transform 1 0 122200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4041
timestamp 1654712443
transform 1 0 119200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4043
timestamp 1654712443
transform 1 0 125200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4044
timestamp 1654712443
transform 1 0 128200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4045
timestamp 1654712443
transform 1 0 131200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4046
timestamp 1654712443
transform 1 0 134200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4047
timestamp 1654712443
transform 1 0 137200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4048
timestamp 1654712443
transform 1 0 140200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4049
timestamp 1654712443
transform 1 0 143200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4050
timestamp 1654712443
transform 1 0 146200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4052
timestamp 1654712443
transform 1 0 152200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4051
timestamp 1654712443
transform 1 0 149200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4053
timestamp 1654712443
transform 1 0 155200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4054
timestamp 1654712443
transform 1 0 158200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4055
timestamp 1654712443
transform 1 0 161200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4056
timestamp 1654712443
transform 1 0 164200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4057
timestamp 1654712443
transform 1 0 167200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4058
timestamp 1654712443
transform 1 0 170200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4059
timestamp 1654712443
transform 1 0 173200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4060
timestamp 1654712443
transform 1 0 176200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4061
timestamp 1654712443
transform 1 0 179200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4063
timestamp 1654712443
transform 1 0 185200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4062
timestamp 1654712443
transform 1 0 182200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4064
timestamp 1654712443
transform 1 0 188200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4065
timestamp 1654712443
transform 1 0 191200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4066
timestamp 1654712443
transform 1 0 194200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4067
timestamp 1654712443
transform 1 0 197200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4068
timestamp 1654712443
transform 1 0 200200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4069
timestamp 1654712443
transform 1 0 203200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4070
timestamp 1654712443
transform 1 0 206200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4071
timestamp 1654712443
transform 1 0 209200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4073
timestamp 1654712443
transform 1 0 215200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4072
timestamp 1654712443
transform 1 0 212200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4074
timestamp 1654712443
transform 1 0 218200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4075
timestamp 1654712443
transform 1 0 221200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4076
timestamp 1654712443
transform 1 0 224200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4077
timestamp 1654712443
transform 1 0 227200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4078
timestamp 1654712443
transform 1 0 230200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4079
timestamp 1654712443
transform 1 0 233200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4080
timestamp 1654712443
transform 1 0 236200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4081
timestamp 1654712443
transform 1 0 239200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4083
timestamp 1654712443
transform 1 0 245200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4082
timestamp 1654712443
transform 1 0 242200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4084
timestamp 1654712443
transform 1 0 248200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4085
timestamp 1654712443
transform 1 0 251200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4086
timestamp 1654712443
transform 1 0 254200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4087
timestamp 1654712443
transform 1 0 257200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4088
timestamp 1654712443
transform 1 0 260200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4089
timestamp 1654712443
transform 1 0 263200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4090
timestamp 1654712443
transform 1 0 266200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4091
timestamp 1654712443
transform 1 0 269200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4092
timestamp 1654712443
transform 1 0 272200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4094
timestamp 1654712443
transform 1 0 278200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4093
timestamp 1654712443
transform 1 0 275200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4095
timestamp 1654712443
transform 1 0 281200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4096
timestamp 1654712443
transform 1 0 284200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4097
timestamp 1654712443
transform 1 0 287200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4098
timestamp 1654712443
transform 1 0 290200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_4099
timestamp 1654712443
transform 1 0 293200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_3901
timestamp 1654712443
transform 1 0 -800 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3900
timestamp 1654712443
transform 1 0 -3800 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3902
timestamp 1654712443
transform 1 0 2200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3903
timestamp 1654712443
transform 1 0 5200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3904
timestamp 1654712443
transform 1 0 8200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3905
timestamp 1654712443
transform 1 0 11200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3906
timestamp 1654712443
transform 1 0 14200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3907
timestamp 1654712443
transform 1 0 17200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3908
timestamp 1654712443
transform 1 0 20200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3909
timestamp 1654712443
transform 1 0 23200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3911
timestamp 1654712443
transform 1 0 29200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3910
timestamp 1654712443
transform 1 0 26200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3912
timestamp 1654712443
transform 1 0 32200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3913
timestamp 1654712443
transform 1 0 35200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3914
timestamp 1654712443
transform 1 0 38200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3915
timestamp 1654712443
transform 1 0 41200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3916
timestamp 1654712443
transform 1 0 44200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3917
timestamp 1654712443
transform 1 0 47200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3918
timestamp 1654712443
transform 1 0 50200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3919
timestamp 1654712443
transform 1 0 53200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3921
timestamp 1654712443
transform 1 0 59200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3920
timestamp 1654712443
transform 1 0 56200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3922
timestamp 1654712443
transform 1 0 62200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3923
timestamp 1654712443
transform 1 0 65200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3924
timestamp 1654712443
transform 1 0 68200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3925
timestamp 1654712443
transform 1 0 71200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3926
timestamp 1654712443
transform 1 0 74200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3927
timestamp 1654712443
transform 1 0 77200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3928
timestamp 1654712443
transform 1 0 80200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3929
timestamp 1654712443
transform 1 0 83200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3930
timestamp 1654712443
transform 1 0 86200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3931
timestamp 1654712443
transform 1 0 89200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3932
timestamp 1654712443
transform 1 0 92200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3933
timestamp 1654712443
transform 1 0 95200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3934
timestamp 1654712443
transform 1 0 98200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3935
timestamp 1654712443
transform 1 0 101200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3936
timestamp 1654712443
transform 1 0 104200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3937
timestamp 1654712443
transform 1 0 107200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3938
timestamp 1654712443
transform 1 0 110200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3939
timestamp 1654712443
transform 1 0 113200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3940
timestamp 1654712443
transform 1 0 116200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3942
timestamp 1654712443
transform 1 0 122200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3941
timestamp 1654712443
transform 1 0 119200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3943
timestamp 1654712443
transform 1 0 125200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3944
timestamp 1654712443
transform 1 0 128200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3945
timestamp 1654712443
transform 1 0 131200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3946
timestamp 1654712443
transform 1 0 134200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3947
timestamp 1654712443
transform 1 0 137200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3948
timestamp 1654712443
transform 1 0 140200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3949
timestamp 1654712443
transform 1 0 143200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3950
timestamp 1654712443
transform 1 0 146200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3952
timestamp 1654712443
transform 1 0 152200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3951
timestamp 1654712443
transform 1 0 149200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3953
timestamp 1654712443
transform 1 0 155200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3954
timestamp 1654712443
transform 1 0 158200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3955
timestamp 1654712443
transform 1 0 161200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3956
timestamp 1654712443
transform 1 0 164200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3957
timestamp 1654712443
transform 1 0 167200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3958
timestamp 1654712443
transform 1 0 170200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3959
timestamp 1654712443
transform 1 0 173200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3960
timestamp 1654712443
transform 1 0 176200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3961
timestamp 1654712443
transform 1 0 179200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3963
timestamp 1654712443
transform 1 0 185200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3962
timestamp 1654712443
transform 1 0 182200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3964
timestamp 1654712443
transform 1 0 188200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3965
timestamp 1654712443
transform 1 0 191200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3966
timestamp 1654712443
transform 1 0 194200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3967
timestamp 1654712443
transform 1 0 197200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3968
timestamp 1654712443
transform 1 0 200200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3969
timestamp 1654712443
transform 1 0 203200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3970
timestamp 1654712443
transform 1 0 206200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3971
timestamp 1654712443
transform 1 0 209200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3973
timestamp 1654712443
transform 1 0 215200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3972
timestamp 1654712443
transform 1 0 212200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3974
timestamp 1654712443
transform 1 0 218200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3975
timestamp 1654712443
transform 1 0 221200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3976
timestamp 1654712443
transform 1 0 224200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3977
timestamp 1654712443
transform 1 0 227200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3978
timestamp 1654712443
transform 1 0 230200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3979
timestamp 1654712443
transform 1 0 233200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3980
timestamp 1654712443
transform 1 0 236200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3981
timestamp 1654712443
transform 1 0 239200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3983
timestamp 1654712443
transform 1 0 245200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3982
timestamp 1654712443
transform 1 0 242200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3984
timestamp 1654712443
transform 1 0 248200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3985
timestamp 1654712443
transform 1 0 251200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3986
timestamp 1654712443
transform 1 0 254200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3987
timestamp 1654712443
transform 1 0 257200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3988
timestamp 1654712443
transform 1 0 260200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3989
timestamp 1654712443
transform 1 0 263200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3990
timestamp 1654712443
transform 1 0 266200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3991
timestamp 1654712443
transform 1 0 269200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3992
timestamp 1654712443
transform 1 0 272200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3994
timestamp 1654712443
transform 1 0 278200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3993
timestamp 1654712443
transform 1 0 275200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3995
timestamp 1654712443
transform 1 0 281200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3996
timestamp 1654712443
transform 1 0 284200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3997
timestamp 1654712443
transform 1 0 287200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3998
timestamp 1654712443
transform 1 0 290200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3999
timestamp 1654712443
transform 1 0 293200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_3801
timestamp 1654712443
transform 1 0 -800 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3800
timestamp 1654712443
transform 1 0 -3800 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3802
timestamp 1654712443
transform 1 0 2200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3803
timestamp 1654712443
transform 1 0 5200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3804
timestamp 1654712443
transform 1 0 8200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3805
timestamp 1654712443
transform 1 0 11200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3806
timestamp 1654712443
transform 1 0 14200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3807
timestamp 1654712443
transform 1 0 17200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3808
timestamp 1654712443
transform 1 0 20200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3809
timestamp 1654712443
transform 1 0 23200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3811
timestamp 1654712443
transform 1 0 29200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3810
timestamp 1654712443
transform 1 0 26200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3812
timestamp 1654712443
transform 1 0 32200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3813
timestamp 1654712443
transform 1 0 35200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3814
timestamp 1654712443
transform 1 0 38200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3815
timestamp 1654712443
transform 1 0 41200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3816
timestamp 1654712443
transform 1 0 44200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3817
timestamp 1654712443
transform 1 0 47200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3818
timestamp 1654712443
transform 1 0 50200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3819
timestamp 1654712443
transform 1 0 53200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3821
timestamp 1654712443
transform 1 0 59200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3820
timestamp 1654712443
transform 1 0 56200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3822
timestamp 1654712443
transform 1 0 62200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3823
timestamp 1654712443
transform 1 0 65200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3824
timestamp 1654712443
transform 1 0 68200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3825
timestamp 1654712443
transform 1 0 71200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3826
timestamp 1654712443
transform 1 0 74200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3827
timestamp 1654712443
transform 1 0 77200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3828
timestamp 1654712443
transform 1 0 80200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3829
timestamp 1654712443
transform 1 0 83200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3830
timestamp 1654712443
transform 1 0 86200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3832
timestamp 1654712443
transform 1 0 92200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3831
timestamp 1654712443
transform 1 0 89200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3833
timestamp 1654712443
transform 1 0 95200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3834
timestamp 1654712443
transform 1 0 98200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3835
timestamp 1654712443
transform 1 0 101200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3836
timestamp 1654712443
transform 1 0 104200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3837
timestamp 1654712443
transform 1 0 107200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3838
timestamp 1654712443
transform 1 0 110200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3839
timestamp 1654712443
transform 1 0 113200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3840
timestamp 1654712443
transform 1 0 116200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3842
timestamp 1654712443
transform 1 0 122200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3841
timestamp 1654712443
transform 1 0 119200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3843
timestamp 1654712443
transform 1 0 125200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3844
timestamp 1654712443
transform 1 0 128200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3845
timestamp 1654712443
transform 1 0 131200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3846
timestamp 1654712443
transform 1 0 134200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3847
timestamp 1654712443
transform 1 0 137200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3848
timestamp 1654712443
transform 1 0 140200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3849
timestamp 1654712443
transform 1 0 143200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3850
timestamp 1654712443
transform 1 0 146200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3852
timestamp 1654712443
transform 1 0 152200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3851
timestamp 1654712443
transform 1 0 149200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3853
timestamp 1654712443
transform 1 0 155200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3854
timestamp 1654712443
transform 1 0 158200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3855
timestamp 1654712443
transform 1 0 161200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3856
timestamp 1654712443
transform 1 0 164200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3857
timestamp 1654712443
transform 1 0 167200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3858
timestamp 1654712443
transform 1 0 170200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3859
timestamp 1654712443
transform 1 0 173200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3860
timestamp 1654712443
transform 1 0 176200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3861
timestamp 1654712443
transform 1 0 179200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3863
timestamp 1654712443
transform 1 0 185200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3862
timestamp 1654712443
transform 1 0 182200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3864
timestamp 1654712443
transform 1 0 188200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3865
timestamp 1654712443
transform 1 0 191200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3866
timestamp 1654712443
transform 1 0 194200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3867
timestamp 1654712443
transform 1 0 197200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3868
timestamp 1654712443
transform 1 0 200200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3869
timestamp 1654712443
transform 1 0 203200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3870
timestamp 1654712443
transform 1 0 206200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3871
timestamp 1654712443
transform 1 0 209200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3873
timestamp 1654712443
transform 1 0 215200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3872
timestamp 1654712443
transform 1 0 212200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3874
timestamp 1654712443
transform 1 0 218200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3875
timestamp 1654712443
transform 1 0 221200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3876
timestamp 1654712443
transform 1 0 224200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3877
timestamp 1654712443
transform 1 0 227200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3878
timestamp 1654712443
transform 1 0 230200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3879
timestamp 1654712443
transform 1 0 233200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3880
timestamp 1654712443
transform 1 0 236200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3881
timestamp 1654712443
transform 1 0 239200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3883
timestamp 1654712443
transform 1 0 245200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3882
timestamp 1654712443
transform 1 0 242200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3884
timestamp 1654712443
transform 1 0 248200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3885
timestamp 1654712443
transform 1 0 251200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3886
timestamp 1654712443
transform 1 0 254200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3887
timestamp 1654712443
transform 1 0 257200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3888
timestamp 1654712443
transform 1 0 260200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3889
timestamp 1654712443
transform 1 0 263200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3890
timestamp 1654712443
transform 1 0 266200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3891
timestamp 1654712443
transform 1 0 269200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3892
timestamp 1654712443
transform 1 0 272200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3894
timestamp 1654712443
transform 1 0 278200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3893
timestamp 1654712443
transform 1 0 275200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3895
timestamp 1654712443
transform 1 0 281200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3896
timestamp 1654712443
transform 1 0 284200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3897
timestamp 1654712443
transform 1 0 287200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3898
timestamp 1654712443
transform 1 0 290200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3899
timestamp 1654712443
transform 1 0 293200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_3601
timestamp 1654712443
transform 1 0 -800 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3600
timestamp 1654712443
transform 1 0 -3800 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3701
timestamp 1654712443
transform 1 0 -800 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3700
timestamp 1654712443
transform 1 0 -3800 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3602
timestamp 1654712443
transform 1 0 2200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3702
timestamp 1654712443
transform 1 0 2200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3603
timestamp 1654712443
transform 1 0 5200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3703
timestamp 1654712443
transform 1 0 5200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3604
timestamp 1654712443
transform 1 0 8200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3704
timestamp 1654712443
transform 1 0 8200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3605
timestamp 1654712443
transform 1 0 11200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3705
timestamp 1654712443
transform 1 0 11200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3606
timestamp 1654712443
transform 1 0 14200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3706
timestamp 1654712443
transform 1 0 14200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3607
timestamp 1654712443
transform 1 0 17200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3707
timestamp 1654712443
transform 1 0 17200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3608
timestamp 1654712443
transform 1 0 20200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3708
timestamp 1654712443
transform 1 0 20200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3609
timestamp 1654712443
transform 1 0 23200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3709
timestamp 1654712443
transform 1 0 23200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3611
timestamp 1654712443
transform 1 0 29200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3610
timestamp 1654712443
transform 1 0 26200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3711
timestamp 1654712443
transform 1 0 29200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3710
timestamp 1654712443
transform 1 0 26200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3612
timestamp 1654712443
transform 1 0 32200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3712
timestamp 1654712443
transform 1 0 32200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3613
timestamp 1654712443
transform 1 0 35200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3713
timestamp 1654712443
transform 1 0 35200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3614
timestamp 1654712443
transform 1 0 38200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3714
timestamp 1654712443
transform 1 0 38200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3615
timestamp 1654712443
transform 1 0 41200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3715
timestamp 1654712443
transform 1 0 41200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3616
timestamp 1654712443
transform 1 0 44200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3716
timestamp 1654712443
transform 1 0 44200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3617
timestamp 1654712443
transform 1 0 47200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3717
timestamp 1654712443
transform 1 0 47200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3618
timestamp 1654712443
transform 1 0 50200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3718
timestamp 1654712443
transform 1 0 50200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3619
timestamp 1654712443
transform 1 0 53200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3719
timestamp 1654712443
transform 1 0 53200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3621
timestamp 1654712443
transform 1 0 59200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3620
timestamp 1654712443
transform 1 0 56200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3721
timestamp 1654712443
transform 1 0 59200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3720
timestamp 1654712443
transform 1 0 56200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3622
timestamp 1654712443
transform 1 0 62200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3722
timestamp 1654712443
transform 1 0 62200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3623
timestamp 1654712443
transform 1 0 65200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3723
timestamp 1654712443
transform 1 0 65200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3624
timestamp 1654712443
transform 1 0 68200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3724
timestamp 1654712443
transform 1 0 68200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3625
timestamp 1654712443
transform 1 0 71200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3725
timestamp 1654712443
transform 1 0 71200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3626
timestamp 1654712443
transform 1 0 74200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3726
timestamp 1654712443
transform 1 0 74200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3627
timestamp 1654712443
transform 1 0 77200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3727
timestamp 1654712443
transform 1 0 77200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3628
timestamp 1654712443
transform 1 0 80200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3728
timestamp 1654712443
transform 1 0 80200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3629
timestamp 1654712443
transform 1 0 83200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3729
timestamp 1654712443
transform 1 0 83200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3630
timestamp 1654712443
transform 1 0 86200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3730
timestamp 1654712443
transform 1 0 86200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3632
timestamp 1654712443
transform 1 0 92200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3631
timestamp 1654712443
transform 1 0 89200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3732
timestamp 1654712443
transform 1 0 92200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3731
timestamp 1654712443
transform 1 0 89200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3633
timestamp 1654712443
transform 1 0 95200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3733
timestamp 1654712443
transform 1 0 95200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3634
timestamp 1654712443
transform 1 0 98200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3734
timestamp 1654712443
transform 1 0 98200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3635
timestamp 1654712443
transform 1 0 101200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3735
timestamp 1654712443
transform 1 0 101200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3636
timestamp 1654712443
transform 1 0 104200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3736
timestamp 1654712443
transform 1 0 104200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3637
timestamp 1654712443
transform 1 0 107200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3737
timestamp 1654712443
transform 1 0 107200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3638
timestamp 1654712443
transform 1 0 110200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3738
timestamp 1654712443
transform 1 0 110200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3639
timestamp 1654712443
transform 1 0 113200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3739
timestamp 1654712443
transform 1 0 113200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3640
timestamp 1654712443
transform 1 0 116200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3740
timestamp 1654712443
transform 1 0 116200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3642
timestamp 1654712443
transform 1 0 122200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3641
timestamp 1654712443
transform 1 0 119200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3742
timestamp 1654712443
transform 1 0 122200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3741
timestamp 1654712443
transform 1 0 119200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3643
timestamp 1654712443
transform 1 0 125200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3743
timestamp 1654712443
transform 1 0 125200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3644
timestamp 1654712443
transform 1 0 128200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3744
timestamp 1654712443
transform 1 0 128200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3645
timestamp 1654712443
transform 1 0 131200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3745
timestamp 1654712443
transform 1 0 131200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3646
timestamp 1654712443
transform 1 0 134200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3746
timestamp 1654712443
transform 1 0 134200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3647
timestamp 1654712443
transform 1 0 137200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3747
timestamp 1654712443
transform 1 0 137200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3648
timestamp 1654712443
transform 1 0 140200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3748
timestamp 1654712443
transform 1 0 140200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3649
timestamp 1654712443
transform 1 0 143200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3749
timestamp 1654712443
transform 1 0 143200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3650
timestamp 1654712443
transform 1 0 146200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3750
timestamp 1654712443
transform 1 0 146200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3652
timestamp 1654712443
transform 1 0 152200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3651
timestamp 1654712443
transform 1 0 149200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3752
timestamp 1654712443
transform 1 0 152200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3751
timestamp 1654712443
transform 1 0 149200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3653
timestamp 1654712443
transform 1 0 155200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3753
timestamp 1654712443
transform 1 0 155200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3654
timestamp 1654712443
transform 1 0 158200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3754
timestamp 1654712443
transform 1 0 158200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3655
timestamp 1654712443
transform 1 0 161200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3755
timestamp 1654712443
transform 1 0 161200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3656
timestamp 1654712443
transform 1 0 164200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3756
timestamp 1654712443
transform 1 0 164200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3657
timestamp 1654712443
transform 1 0 167200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3757
timestamp 1654712443
transform 1 0 167200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3658
timestamp 1654712443
transform 1 0 170200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3758
timestamp 1654712443
transform 1 0 170200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3659
timestamp 1654712443
transform 1 0 173200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3759
timestamp 1654712443
transform 1 0 173200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3660
timestamp 1654712443
transform 1 0 176200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3760
timestamp 1654712443
transform 1 0 176200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3661
timestamp 1654712443
transform 1 0 179200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3761
timestamp 1654712443
transform 1 0 179200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3663
timestamp 1654712443
transform 1 0 185200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3662
timestamp 1654712443
transform 1 0 182200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3763
timestamp 1654712443
transform 1 0 185200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3762
timestamp 1654712443
transform 1 0 182200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3664
timestamp 1654712443
transform 1 0 188200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3764
timestamp 1654712443
transform 1 0 188200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3665
timestamp 1654712443
transform 1 0 191200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3765
timestamp 1654712443
transform 1 0 191200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3666
timestamp 1654712443
transform 1 0 194200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3766
timestamp 1654712443
transform 1 0 194200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3667
timestamp 1654712443
transform 1 0 197200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3767
timestamp 1654712443
transform 1 0 197200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3668
timestamp 1654712443
transform 1 0 200200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3768
timestamp 1654712443
transform 1 0 200200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3669
timestamp 1654712443
transform 1 0 203200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3769
timestamp 1654712443
transform 1 0 203200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3670
timestamp 1654712443
transform 1 0 206200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3770
timestamp 1654712443
transform 1 0 206200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3671
timestamp 1654712443
transform 1 0 209200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3771
timestamp 1654712443
transform 1 0 209200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3673
timestamp 1654712443
transform 1 0 215200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3672
timestamp 1654712443
transform 1 0 212200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3773
timestamp 1654712443
transform 1 0 215200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3772
timestamp 1654712443
transform 1 0 212200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3674
timestamp 1654712443
transform 1 0 218200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3774
timestamp 1654712443
transform 1 0 218200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3675
timestamp 1654712443
transform 1 0 221200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3775
timestamp 1654712443
transform 1 0 221200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3676
timestamp 1654712443
transform 1 0 224200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3776
timestamp 1654712443
transform 1 0 224200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3677
timestamp 1654712443
transform 1 0 227200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3777
timestamp 1654712443
transform 1 0 227200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3678
timestamp 1654712443
transform 1 0 230200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3778
timestamp 1654712443
transform 1 0 230200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3679
timestamp 1654712443
transform 1 0 233200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3779
timestamp 1654712443
transform 1 0 233200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3680
timestamp 1654712443
transform 1 0 236200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3780
timestamp 1654712443
transform 1 0 236200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3681
timestamp 1654712443
transform 1 0 239200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3781
timestamp 1654712443
transform 1 0 239200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3683
timestamp 1654712443
transform 1 0 245200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3682
timestamp 1654712443
transform 1 0 242200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3783
timestamp 1654712443
transform 1 0 245200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3782
timestamp 1654712443
transform 1 0 242200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3684
timestamp 1654712443
transform 1 0 248200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3784
timestamp 1654712443
transform 1 0 248200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3685
timestamp 1654712443
transform 1 0 251200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3785
timestamp 1654712443
transform 1 0 251200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3686
timestamp 1654712443
transform 1 0 254200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3786
timestamp 1654712443
transform 1 0 254200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3687
timestamp 1654712443
transform 1 0 257200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3787
timestamp 1654712443
transform 1 0 257200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3688
timestamp 1654712443
transform 1 0 260200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3788
timestamp 1654712443
transform 1 0 260200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3689
timestamp 1654712443
transform 1 0 263200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3789
timestamp 1654712443
transform 1 0 263200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3690
timestamp 1654712443
transform 1 0 266200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3790
timestamp 1654712443
transform 1 0 266200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3691
timestamp 1654712443
transform 1 0 269200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3791
timestamp 1654712443
transform 1 0 269200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3692
timestamp 1654712443
transform 1 0 272200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3792
timestamp 1654712443
transform 1 0 272200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3694
timestamp 1654712443
transform 1 0 278200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3693
timestamp 1654712443
transform 1 0 275200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3794
timestamp 1654712443
transform 1 0 278200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3793
timestamp 1654712443
transform 1 0 275200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3695
timestamp 1654712443
transform 1 0 281200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3795
timestamp 1654712443
transform 1 0 281200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3696
timestamp 1654712443
transform 1 0 284200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3796
timestamp 1654712443
transform 1 0 284200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3697
timestamp 1654712443
transform 1 0 287200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3797
timestamp 1654712443
transform 1 0 287200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3698
timestamp 1654712443
transform 1 0 290200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3798
timestamp 1654712443
transform 1 0 290200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3699
timestamp 1654712443
transform 1 0 293200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_3799
timestamp 1654712443
transform 1 0 293200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_3501
timestamp 1654712443
transform 1 0 -800 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3500
timestamp 1654712443
transform 1 0 -3800 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3502
timestamp 1654712443
transform 1 0 2200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3503
timestamp 1654712443
transform 1 0 5200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3504
timestamp 1654712443
transform 1 0 8200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3505
timestamp 1654712443
transform 1 0 11200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3506
timestamp 1654712443
transform 1 0 14200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3507
timestamp 1654712443
transform 1 0 17200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3508
timestamp 1654712443
transform 1 0 20200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3509
timestamp 1654712443
transform 1 0 23200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3511
timestamp 1654712443
transform 1 0 29200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3510
timestamp 1654712443
transform 1 0 26200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3512
timestamp 1654712443
transform 1 0 32200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3513
timestamp 1654712443
transform 1 0 35200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3514
timestamp 1654712443
transform 1 0 38200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3515
timestamp 1654712443
transform 1 0 41200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3516
timestamp 1654712443
transform 1 0 44200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3517
timestamp 1654712443
transform 1 0 47200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3518
timestamp 1654712443
transform 1 0 50200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3519
timestamp 1654712443
transform 1 0 53200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3521
timestamp 1654712443
transform 1 0 59200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3520
timestamp 1654712443
transform 1 0 56200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3522
timestamp 1654712443
transform 1 0 62200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3523
timestamp 1654712443
transform 1 0 65200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3524
timestamp 1654712443
transform 1 0 68200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3525
timestamp 1654712443
transform 1 0 71200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3526
timestamp 1654712443
transform 1 0 74200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3527
timestamp 1654712443
transform 1 0 77200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3528
timestamp 1654712443
transform 1 0 80200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3529
timestamp 1654712443
transform 1 0 83200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3530
timestamp 1654712443
transform 1 0 86200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3532
timestamp 1654712443
transform 1 0 92200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3531
timestamp 1654712443
transform 1 0 89200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3533
timestamp 1654712443
transform 1 0 95200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3534
timestamp 1654712443
transform 1 0 98200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3535
timestamp 1654712443
transform 1 0 101200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3536
timestamp 1654712443
transform 1 0 104200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3537
timestamp 1654712443
transform 1 0 107200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3538
timestamp 1654712443
transform 1 0 110200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3539
timestamp 1654712443
transform 1 0 113200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3540
timestamp 1654712443
transform 1 0 116200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3542
timestamp 1654712443
transform 1 0 122200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3541
timestamp 1654712443
transform 1 0 119200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3543
timestamp 1654712443
transform 1 0 125200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3544
timestamp 1654712443
transform 1 0 128200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3545
timestamp 1654712443
transform 1 0 131200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3546
timestamp 1654712443
transform 1 0 134200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3547
timestamp 1654712443
transform 1 0 137200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3548
timestamp 1654712443
transform 1 0 140200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3549
timestamp 1654712443
transform 1 0 143200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3550
timestamp 1654712443
transform 1 0 146200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3552
timestamp 1654712443
transform 1 0 152200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3551
timestamp 1654712443
transform 1 0 149200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3553
timestamp 1654712443
transform 1 0 155200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3554
timestamp 1654712443
transform 1 0 158200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3555
timestamp 1654712443
transform 1 0 161200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3556
timestamp 1654712443
transform 1 0 164200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3557
timestamp 1654712443
transform 1 0 167200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3558
timestamp 1654712443
transform 1 0 170200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3559
timestamp 1654712443
transform 1 0 173200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3560
timestamp 1654712443
transform 1 0 176200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3561
timestamp 1654712443
transform 1 0 179200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3563
timestamp 1654712443
transform 1 0 185200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3562
timestamp 1654712443
transform 1 0 182200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3564
timestamp 1654712443
transform 1 0 188200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3565
timestamp 1654712443
transform 1 0 191200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3566
timestamp 1654712443
transform 1 0 194200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3567
timestamp 1654712443
transform 1 0 197200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3568
timestamp 1654712443
transform 1 0 200200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3569
timestamp 1654712443
transform 1 0 203200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3570
timestamp 1654712443
transform 1 0 206200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3571
timestamp 1654712443
transform 1 0 209200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3573
timestamp 1654712443
transform 1 0 215200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3572
timestamp 1654712443
transform 1 0 212200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3574
timestamp 1654712443
transform 1 0 218200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3575
timestamp 1654712443
transform 1 0 221200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3576
timestamp 1654712443
transform 1 0 224200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3577
timestamp 1654712443
transform 1 0 227200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3578
timestamp 1654712443
transform 1 0 230200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3579
timestamp 1654712443
transform 1 0 233200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3580
timestamp 1654712443
transform 1 0 236200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3581
timestamp 1654712443
transform 1 0 239200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3583
timestamp 1654712443
transform 1 0 245200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3582
timestamp 1654712443
transform 1 0 242200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3584
timestamp 1654712443
transform 1 0 248200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3585
timestamp 1654712443
transform 1 0 251200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3586
timestamp 1654712443
transform 1 0 254200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3587
timestamp 1654712443
transform 1 0 257200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3588
timestamp 1654712443
transform 1 0 260200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3589
timestamp 1654712443
transform 1 0 263200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3590
timestamp 1654712443
transform 1 0 266200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3591
timestamp 1654712443
transform 1 0 269200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3592
timestamp 1654712443
transform 1 0 272200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3594
timestamp 1654712443
transform 1 0 278200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3593
timestamp 1654712443
transform 1 0 275200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3595
timestamp 1654712443
transform 1 0 281200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3596
timestamp 1654712443
transform 1 0 284200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3597
timestamp 1654712443
transform 1 0 287200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3598
timestamp 1654712443
transform 1 0 290200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3599
timestamp 1654712443
transform 1 0 293200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_3401
timestamp 1654712443
transform 1 0 -800 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3400
timestamp 1654712443
transform 1 0 -3800 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3402
timestamp 1654712443
transform 1 0 2200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3403
timestamp 1654712443
transform 1 0 5200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3404
timestamp 1654712443
transform 1 0 8200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3405
timestamp 1654712443
transform 1 0 11200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3406
timestamp 1654712443
transform 1 0 14200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3407
timestamp 1654712443
transform 1 0 17200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3408
timestamp 1654712443
transform 1 0 20200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3409
timestamp 1654712443
transform 1 0 23200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3411
timestamp 1654712443
transform 1 0 29200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3410
timestamp 1654712443
transform 1 0 26200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3412
timestamp 1654712443
transform 1 0 32200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3413
timestamp 1654712443
transform 1 0 35200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3414
timestamp 1654712443
transform 1 0 38200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3415
timestamp 1654712443
transform 1 0 41200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3416
timestamp 1654712443
transform 1 0 44200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3417
timestamp 1654712443
transform 1 0 47200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3418
timestamp 1654712443
transform 1 0 50200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3419
timestamp 1654712443
transform 1 0 53200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3421
timestamp 1654712443
transform 1 0 59200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3420
timestamp 1654712443
transform 1 0 56200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3422
timestamp 1654712443
transform 1 0 62200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3423
timestamp 1654712443
transform 1 0 65200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3424
timestamp 1654712443
transform 1 0 68200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3425
timestamp 1654712443
transform 1 0 71200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3426
timestamp 1654712443
transform 1 0 74200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3427
timestamp 1654712443
transform 1 0 77200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3428
timestamp 1654712443
transform 1 0 80200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3429
timestamp 1654712443
transform 1 0 83200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3430
timestamp 1654712443
transform 1 0 86200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3432
timestamp 1654712443
transform 1 0 92200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3431
timestamp 1654712443
transform 1 0 89200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3433
timestamp 1654712443
transform 1 0 95200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3434
timestamp 1654712443
transform 1 0 98200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3435
timestamp 1654712443
transform 1 0 101200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3436
timestamp 1654712443
transform 1 0 104200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3437
timestamp 1654712443
transform 1 0 107200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3438
timestamp 1654712443
transform 1 0 110200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3439
timestamp 1654712443
transform 1 0 113200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3440
timestamp 1654712443
transform 1 0 116200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3442
timestamp 1654712443
transform 1 0 122200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3441
timestamp 1654712443
transform 1 0 119200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3443
timestamp 1654712443
transform 1 0 125200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3444
timestamp 1654712443
transform 1 0 128200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3445
timestamp 1654712443
transform 1 0 131200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3446
timestamp 1654712443
transform 1 0 134200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3447
timestamp 1654712443
transform 1 0 137200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3448
timestamp 1654712443
transform 1 0 140200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3449
timestamp 1654712443
transform 1 0 143200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3450
timestamp 1654712443
transform 1 0 146200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3452
timestamp 1654712443
transform 1 0 152200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3451
timestamp 1654712443
transform 1 0 149200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3453
timestamp 1654712443
transform 1 0 155200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3454
timestamp 1654712443
transform 1 0 158200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3455
timestamp 1654712443
transform 1 0 161200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3456
timestamp 1654712443
transform 1 0 164200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3457
timestamp 1654712443
transform 1 0 167200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3458
timestamp 1654712443
transform 1 0 170200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3459
timestamp 1654712443
transform 1 0 173200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3460
timestamp 1654712443
transform 1 0 176200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3461
timestamp 1654712443
transform 1 0 179200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3463
timestamp 1654712443
transform 1 0 185200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3462
timestamp 1654712443
transform 1 0 182200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3464
timestamp 1654712443
transform 1 0 188200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3465
timestamp 1654712443
transform 1 0 191200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3466
timestamp 1654712443
transform 1 0 194200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3467
timestamp 1654712443
transform 1 0 197200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3468
timestamp 1654712443
transform 1 0 200200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3469
timestamp 1654712443
transform 1 0 203200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3470
timestamp 1654712443
transform 1 0 206200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3471
timestamp 1654712443
transform 1 0 209200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3473
timestamp 1654712443
transform 1 0 215200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3472
timestamp 1654712443
transform 1 0 212200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3474
timestamp 1654712443
transform 1 0 218200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3475
timestamp 1654712443
transform 1 0 221200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3476
timestamp 1654712443
transform 1 0 224200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3477
timestamp 1654712443
transform 1 0 227200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3478
timestamp 1654712443
transform 1 0 230200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3479
timestamp 1654712443
transform 1 0 233200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3480
timestamp 1654712443
transform 1 0 236200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3481
timestamp 1654712443
transform 1 0 239200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3483
timestamp 1654712443
transform 1 0 245200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3482
timestamp 1654712443
transform 1 0 242200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3484
timestamp 1654712443
transform 1 0 248200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3485
timestamp 1654712443
transform 1 0 251200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3486
timestamp 1654712443
transform 1 0 254200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3487
timestamp 1654712443
transform 1 0 257200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3488
timestamp 1654712443
transform 1 0 260200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3489
timestamp 1654712443
transform 1 0 263200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3490
timestamp 1654712443
transform 1 0 266200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3491
timestamp 1654712443
transform 1 0 269200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3492
timestamp 1654712443
transform 1 0 272200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3494
timestamp 1654712443
transform 1 0 278200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3493
timestamp 1654712443
transform 1 0 275200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3495
timestamp 1654712443
transform 1 0 281200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3496
timestamp 1654712443
transform 1 0 284200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3497
timestamp 1654712443
transform 1 0 287200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3498
timestamp 1654712443
transform 1 0 290200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3499
timestamp 1654712443
transform 1 0 293200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_3301
timestamp 1654712443
transform 1 0 -800 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3300
timestamp 1654712443
transform 1 0 -3800 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3302
timestamp 1654712443
transform 1 0 2200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3303
timestamp 1654712443
transform 1 0 5200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3304
timestamp 1654712443
transform 1 0 8200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3305
timestamp 1654712443
transform 1 0 11200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3306
timestamp 1654712443
transform 1 0 14200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3307
timestamp 1654712443
transform 1 0 17200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3308
timestamp 1654712443
transform 1 0 20200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3309
timestamp 1654712443
transform 1 0 23200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3311
timestamp 1654712443
transform 1 0 29200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3310
timestamp 1654712443
transform 1 0 26200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3312
timestamp 1654712443
transform 1 0 32200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3313
timestamp 1654712443
transform 1 0 35200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3314
timestamp 1654712443
transform 1 0 38200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3315
timestamp 1654712443
transform 1 0 41200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3316
timestamp 1654712443
transform 1 0 44200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3317
timestamp 1654712443
transform 1 0 47200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3318
timestamp 1654712443
transform 1 0 50200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3319
timestamp 1654712443
transform 1 0 53200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3321
timestamp 1654712443
transform 1 0 59200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3320
timestamp 1654712443
transform 1 0 56200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3322
timestamp 1654712443
transform 1 0 62200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3323
timestamp 1654712443
transform 1 0 65200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3324
timestamp 1654712443
transform 1 0 68200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3325
timestamp 1654712443
transform 1 0 71200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3326
timestamp 1654712443
transform 1 0 74200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3327
timestamp 1654712443
transform 1 0 77200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3328
timestamp 1654712443
transform 1 0 80200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3329
timestamp 1654712443
transform 1 0 83200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3330
timestamp 1654712443
transform 1 0 86200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3332
timestamp 1654712443
transform 1 0 92200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3331
timestamp 1654712443
transform 1 0 89200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3333
timestamp 1654712443
transform 1 0 95200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3334
timestamp 1654712443
transform 1 0 98200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3335
timestamp 1654712443
transform 1 0 101200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3336
timestamp 1654712443
transform 1 0 104200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3337
timestamp 1654712443
transform 1 0 107200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3338
timestamp 1654712443
transform 1 0 110200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3339
timestamp 1654712443
transform 1 0 113200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3340
timestamp 1654712443
transform 1 0 116200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3342
timestamp 1654712443
transform 1 0 122200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3341
timestamp 1654712443
transform 1 0 119200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3343
timestamp 1654712443
transform 1 0 125200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3344
timestamp 1654712443
transform 1 0 128200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3345
timestamp 1654712443
transform 1 0 131200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3346
timestamp 1654712443
transform 1 0 134200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3347
timestamp 1654712443
transform 1 0 137200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3348
timestamp 1654712443
transform 1 0 140200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3349
timestamp 1654712443
transform 1 0 143200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3350
timestamp 1654712443
transform 1 0 146200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3352
timestamp 1654712443
transform 1 0 152200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3351
timestamp 1654712443
transform 1 0 149200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3353
timestamp 1654712443
transform 1 0 155200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3354
timestamp 1654712443
transform 1 0 158200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3355
timestamp 1654712443
transform 1 0 161200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3356
timestamp 1654712443
transform 1 0 164200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3357
timestamp 1654712443
transform 1 0 167200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3358
timestamp 1654712443
transform 1 0 170200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3359
timestamp 1654712443
transform 1 0 173200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3360
timestamp 1654712443
transform 1 0 176200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3361
timestamp 1654712443
transform 1 0 179200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3363
timestamp 1654712443
transform 1 0 185200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3362
timestamp 1654712443
transform 1 0 182200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3364
timestamp 1654712443
transform 1 0 188200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3365
timestamp 1654712443
transform 1 0 191200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3366
timestamp 1654712443
transform 1 0 194200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3367
timestamp 1654712443
transform 1 0 197200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3368
timestamp 1654712443
transform 1 0 200200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3369
timestamp 1654712443
transform 1 0 203200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3370
timestamp 1654712443
transform 1 0 206200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3371
timestamp 1654712443
transform 1 0 209200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3373
timestamp 1654712443
transform 1 0 215200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3372
timestamp 1654712443
transform 1 0 212200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3374
timestamp 1654712443
transform 1 0 218200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3375
timestamp 1654712443
transform 1 0 221200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3376
timestamp 1654712443
transform 1 0 224200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3377
timestamp 1654712443
transform 1 0 227200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3378
timestamp 1654712443
transform 1 0 230200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3379
timestamp 1654712443
transform 1 0 233200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3380
timestamp 1654712443
transform 1 0 236200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3381
timestamp 1654712443
transform 1 0 239200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3383
timestamp 1654712443
transform 1 0 245200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3382
timestamp 1654712443
transform 1 0 242200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3384
timestamp 1654712443
transform 1 0 248200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3385
timestamp 1654712443
transform 1 0 251200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3386
timestamp 1654712443
transform 1 0 254200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3387
timestamp 1654712443
transform 1 0 257200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3388
timestamp 1654712443
transform 1 0 260200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3389
timestamp 1654712443
transform 1 0 263200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3390
timestamp 1654712443
transform 1 0 266200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3391
timestamp 1654712443
transform 1 0 269200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3392
timestamp 1654712443
transform 1 0 272200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3394
timestamp 1654712443
transform 1 0 278200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3393
timestamp 1654712443
transform 1 0 275200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3395
timestamp 1654712443
transform 1 0 281200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3396
timestamp 1654712443
transform 1 0 284200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3397
timestamp 1654712443
transform 1 0 287200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3398
timestamp 1654712443
transform 1 0 290200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3399
timestamp 1654712443
transform 1 0 293200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_3201
timestamp 1654712443
transform 1 0 -800 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3200
timestamp 1654712443
transform 1 0 -3800 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3202
timestamp 1654712443
transform 1 0 2200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3203
timestamp 1654712443
transform 1 0 5200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3204
timestamp 1654712443
transform 1 0 8200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3205
timestamp 1654712443
transform 1 0 11200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3206
timestamp 1654712443
transform 1 0 14200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3207
timestamp 1654712443
transform 1 0 17200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3208
timestamp 1654712443
transform 1 0 20200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3209
timestamp 1654712443
transform 1 0 23200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3211
timestamp 1654712443
transform 1 0 29200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3210
timestamp 1654712443
transform 1 0 26200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3212
timestamp 1654712443
transform 1 0 32200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3213
timestamp 1654712443
transform 1 0 35200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3214
timestamp 1654712443
transform 1 0 38200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3215
timestamp 1654712443
transform 1 0 41200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3216
timestamp 1654712443
transform 1 0 44200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3217
timestamp 1654712443
transform 1 0 47200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3218
timestamp 1654712443
transform 1 0 50200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3219
timestamp 1654712443
transform 1 0 53200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3221
timestamp 1654712443
transform 1 0 59200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3220
timestamp 1654712443
transform 1 0 56200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3222
timestamp 1654712443
transform 1 0 62200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3223
timestamp 1654712443
transform 1 0 65200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3224
timestamp 1654712443
transform 1 0 68200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3225
timestamp 1654712443
transform 1 0 71200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3226
timestamp 1654712443
transform 1 0 74200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3227
timestamp 1654712443
transform 1 0 77200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3228
timestamp 1654712443
transform 1 0 80200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3229
timestamp 1654712443
transform 1 0 83200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3230
timestamp 1654712443
transform 1 0 86200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3232
timestamp 1654712443
transform 1 0 92200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3231
timestamp 1654712443
transform 1 0 89200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3233
timestamp 1654712443
transform 1 0 95200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3234
timestamp 1654712443
transform 1 0 98200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3235
timestamp 1654712443
transform 1 0 101200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3236
timestamp 1654712443
transform 1 0 104200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3237
timestamp 1654712443
transform 1 0 107200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3238
timestamp 1654712443
transform 1 0 110200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3239
timestamp 1654712443
transform 1 0 113200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3240
timestamp 1654712443
transform 1 0 116200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3242
timestamp 1654712443
transform 1 0 122200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3241
timestamp 1654712443
transform 1 0 119200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3243
timestamp 1654712443
transform 1 0 125200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3244
timestamp 1654712443
transform 1 0 128200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3245
timestamp 1654712443
transform 1 0 131200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3246
timestamp 1654712443
transform 1 0 134200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3247
timestamp 1654712443
transform 1 0 137200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3248
timestamp 1654712443
transform 1 0 140200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3249
timestamp 1654712443
transform 1 0 143200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3250
timestamp 1654712443
transform 1 0 146200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3252
timestamp 1654712443
transform 1 0 152200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3251
timestamp 1654712443
transform 1 0 149200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3253
timestamp 1654712443
transform 1 0 155200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3254
timestamp 1654712443
transform 1 0 158200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3255
timestamp 1654712443
transform 1 0 161200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3256
timestamp 1654712443
transform 1 0 164200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3257
timestamp 1654712443
transform 1 0 167200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3258
timestamp 1654712443
transform 1 0 170200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3259
timestamp 1654712443
transform 1 0 173200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3260
timestamp 1654712443
transform 1 0 176200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3261
timestamp 1654712443
transform 1 0 179200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3263
timestamp 1654712443
transform 1 0 185200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3262
timestamp 1654712443
transform 1 0 182200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3264
timestamp 1654712443
transform 1 0 188200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3265
timestamp 1654712443
transform 1 0 191200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3266
timestamp 1654712443
transform 1 0 194200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3267
timestamp 1654712443
transform 1 0 197200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3268
timestamp 1654712443
transform 1 0 200200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3269
timestamp 1654712443
transform 1 0 203200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3270
timestamp 1654712443
transform 1 0 206200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3271
timestamp 1654712443
transform 1 0 209200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3273
timestamp 1654712443
transform 1 0 215200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3272
timestamp 1654712443
transform 1 0 212200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3274
timestamp 1654712443
transform 1 0 218200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3275
timestamp 1654712443
transform 1 0 221200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3276
timestamp 1654712443
transform 1 0 224200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3277
timestamp 1654712443
transform 1 0 227200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3278
timestamp 1654712443
transform 1 0 230200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3279
timestamp 1654712443
transform 1 0 233200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3280
timestamp 1654712443
transform 1 0 236200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3281
timestamp 1654712443
transform 1 0 239200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3283
timestamp 1654712443
transform 1 0 245200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3282
timestamp 1654712443
transform 1 0 242200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3284
timestamp 1654712443
transform 1 0 248200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3285
timestamp 1654712443
transform 1 0 251200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3286
timestamp 1654712443
transform 1 0 254200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3287
timestamp 1654712443
transform 1 0 257200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3288
timestamp 1654712443
transform 1 0 260200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3289
timestamp 1654712443
transform 1 0 263200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3290
timestamp 1654712443
transform 1 0 266200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3291
timestamp 1654712443
transform 1 0 269200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3292
timestamp 1654712443
transform 1 0 272200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3294
timestamp 1654712443
transform 1 0 278200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3293
timestamp 1654712443
transform 1 0 275200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3295
timestamp 1654712443
transform 1 0 281200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3296
timestamp 1654712443
transform 1 0 284200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3297
timestamp 1654712443
transform 1 0 287200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3298
timestamp 1654712443
transform 1 0 290200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3299
timestamp 1654712443
transform 1 0 293200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_3101
timestamp 1654712443
transform 1 0 -800 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3100
timestamp 1654712443
transform 1 0 -3800 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3102
timestamp 1654712443
transform 1 0 2200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3103
timestamp 1654712443
transform 1 0 5200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3104
timestamp 1654712443
transform 1 0 8200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3105
timestamp 1654712443
transform 1 0 11200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3106
timestamp 1654712443
transform 1 0 14200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3107
timestamp 1654712443
transform 1 0 17200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3108
timestamp 1654712443
transform 1 0 20200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3109
timestamp 1654712443
transform 1 0 23200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3111
timestamp 1654712443
transform 1 0 29200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3110
timestamp 1654712443
transform 1 0 26200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3112
timestamp 1654712443
transform 1 0 32200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3113
timestamp 1654712443
transform 1 0 35200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3114
timestamp 1654712443
transform 1 0 38200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3115
timestamp 1654712443
transform 1 0 41200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3116
timestamp 1654712443
transform 1 0 44200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3117
timestamp 1654712443
transform 1 0 47200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3118
timestamp 1654712443
transform 1 0 50200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3119
timestamp 1654712443
transform 1 0 53200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3121
timestamp 1654712443
transform 1 0 59200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3120
timestamp 1654712443
transform 1 0 56200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3122
timestamp 1654712443
transform 1 0 62200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3123
timestamp 1654712443
transform 1 0 65200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3124
timestamp 1654712443
transform 1 0 68200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3125
timestamp 1654712443
transform 1 0 71200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3126
timestamp 1654712443
transform 1 0 74200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3127
timestamp 1654712443
transform 1 0 77200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3128
timestamp 1654712443
transform 1 0 80200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3129
timestamp 1654712443
transform 1 0 83200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3130
timestamp 1654712443
transform 1 0 86200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3132
timestamp 1654712443
transform 1 0 92200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3131
timestamp 1654712443
transform 1 0 89200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3133
timestamp 1654712443
transform 1 0 95200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3134
timestamp 1654712443
transform 1 0 98200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3135
timestamp 1654712443
transform 1 0 101200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3136
timestamp 1654712443
transform 1 0 104200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3137
timestamp 1654712443
transform 1 0 107200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3138
timestamp 1654712443
transform 1 0 110200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3139
timestamp 1654712443
transform 1 0 113200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3140
timestamp 1654712443
transform 1 0 116200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3142
timestamp 1654712443
transform 1 0 122200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3141
timestamp 1654712443
transform 1 0 119200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3143
timestamp 1654712443
transform 1 0 125200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3144
timestamp 1654712443
transform 1 0 128200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3145
timestamp 1654712443
transform 1 0 131200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3146
timestamp 1654712443
transform 1 0 134200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3147
timestamp 1654712443
transform 1 0 137200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3148
timestamp 1654712443
transform 1 0 140200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3149
timestamp 1654712443
transform 1 0 143200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3150
timestamp 1654712443
transform 1 0 146200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3152
timestamp 1654712443
transform 1 0 152200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3151
timestamp 1654712443
transform 1 0 149200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3153
timestamp 1654712443
transform 1 0 155200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3154
timestamp 1654712443
transform 1 0 158200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3155
timestamp 1654712443
transform 1 0 161200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3156
timestamp 1654712443
transform 1 0 164200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3157
timestamp 1654712443
transform 1 0 167200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3158
timestamp 1654712443
transform 1 0 170200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3159
timestamp 1654712443
transform 1 0 173200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3160
timestamp 1654712443
transform 1 0 176200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3161
timestamp 1654712443
transform 1 0 179200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3163
timestamp 1654712443
transform 1 0 185200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3162
timestamp 1654712443
transform 1 0 182200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3164
timestamp 1654712443
transform 1 0 188200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3165
timestamp 1654712443
transform 1 0 191200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3166
timestamp 1654712443
transform 1 0 194200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3167
timestamp 1654712443
transform 1 0 197200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3168
timestamp 1654712443
transform 1 0 200200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3169
timestamp 1654712443
transform 1 0 203200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3170
timestamp 1654712443
transform 1 0 206200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3171
timestamp 1654712443
transform 1 0 209200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3173
timestamp 1654712443
transform 1 0 215200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3172
timestamp 1654712443
transform 1 0 212200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3174
timestamp 1654712443
transform 1 0 218200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3175
timestamp 1654712443
transform 1 0 221200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3176
timestamp 1654712443
transform 1 0 224200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3177
timestamp 1654712443
transform 1 0 227200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3178
timestamp 1654712443
transform 1 0 230200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3179
timestamp 1654712443
transform 1 0 233200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3180
timestamp 1654712443
transform 1 0 236200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3181
timestamp 1654712443
transform 1 0 239200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3183
timestamp 1654712443
transform 1 0 245200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3182
timestamp 1654712443
transform 1 0 242200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3184
timestamp 1654712443
transform 1 0 248200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3185
timestamp 1654712443
transform 1 0 251200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3186
timestamp 1654712443
transform 1 0 254200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3187
timestamp 1654712443
transform 1 0 257200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3188
timestamp 1654712443
transform 1 0 260200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3189
timestamp 1654712443
transform 1 0 263200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3190
timestamp 1654712443
transform 1 0 266200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3191
timestamp 1654712443
transform 1 0 269200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3192
timestamp 1654712443
transform 1 0 272200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3194
timestamp 1654712443
transform 1 0 278200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3193
timestamp 1654712443
transform 1 0 275200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3195
timestamp 1654712443
transform 1 0 281200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3196
timestamp 1654712443
transform 1 0 284200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3197
timestamp 1654712443
transform 1 0 287200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3198
timestamp 1654712443
transform 1 0 290200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3199
timestamp 1654712443
transform 1 0 293200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_3001
timestamp 1654712443
transform 1 0 -800 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3000
timestamp 1654712443
transform 1 0 -3800 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3002
timestamp 1654712443
transform 1 0 2200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3003
timestamp 1654712443
transform 1 0 5200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3004
timestamp 1654712443
transform 1 0 8200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3005
timestamp 1654712443
transform 1 0 11200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3006
timestamp 1654712443
transform 1 0 14200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3007
timestamp 1654712443
transform 1 0 17200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3008
timestamp 1654712443
transform 1 0 20200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3009
timestamp 1654712443
transform 1 0 23200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3011
timestamp 1654712443
transform 1 0 29200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3010
timestamp 1654712443
transform 1 0 26200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3012
timestamp 1654712443
transform 1 0 32200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3013
timestamp 1654712443
transform 1 0 35200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3014
timestamp 1654712443
transform 1 0 38200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3015
timestamp 1654712443
transform 1 0 41200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3016
timestamp 1654712443
transform 1 0 44200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3017
timestamp 1654712443
transform 1 0 47200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3018
timestamp 1654712443
transform 1 0 50200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3019
timestamp 1654712443
transform 1 0 53200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3021
timestamp 1654712443
transform 1 0 59200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3020
timestamp 1654712443
transform 1 0 56200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3022
timestamp 1654712443
transform 1 0 62200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3023
timestamp 1654712443
transform 1 0 65200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3024
timestamp 1654712443
transform 1 0 68200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3025
timestamp 1654712443
transform 1 0 71200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3026
timestamp 1654712443
transform 1 0 74200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3027
timestamp 1654712443
transform 1 0 77200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3028
timestamp 1654712443
transform 1 0 80200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3029
timestamp 1654712443
transform 1 0 83200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3030
timestamp 1654712443
transform 1 0 86200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3032
timestamp 1654712443
transform 1 0 92200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3031
timestamp 1654712443
transform 1 0 89200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3033
timestamp 1654712443
transform 1 0 95200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3034
timestamp 1654712443
transform 1 0 98200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3035
timestamp 1654712443
transform 1 0 101200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3036
timestamp 1654712443
transform 1 0 104200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3037
timestamp 1654712443
transform 1 0 107200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3038
timestamp 1654712443
transform 1 0 110200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3039
timestamp 1654712443
transform 1 0 113200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3040
timestamp 1654712443
transform 1 0 116200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3042
timestamp 1654712443
transform 1 0 122200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3041
timestamp 1654712443
transform 1 0 119200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3043
timestamp 1654712443
transform 1 0 125200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3044
timestamp 1654712443
transform 1 0 128200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3045
timestamp 1654712443
transform 1 0 131200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3046
timestamp 1654712443
transform 1 0 134200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3047
timestamp 1654712443
transform 1 0 137200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3048
timestamp 1654712443
transform 1 0 140200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3049
timestamp 1654712443
transform 1 0 143200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3050
timestamp 1654712443
transform 1 0 146200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3052
timestamp 1654712443
transform 1 0 152200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3051
timestamp 1654712443
transform 1 0 149200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3053
timestamp 1654712443
transform 1 0 155200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3054
timestamp 1654712443
transform 1 0 158200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3055
timestamp 1654712443
transform 1 0 161200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3056
timestamp 1654712443
transform 1 0 164200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3057
timestamp 1654712443
transform 1 0 167200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3058
timestamp 1654712443
transform 1 0 170200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3059
timestamp 1654712443
transform 1 0 173200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3060
timestamp 1654712443
transform 1 0 176200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3061
timestamp 1654712443
transform 1 0 179200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3063
timestamp 1654712443
transform 1 0 185200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3062
timestamp 1654712443
transform 1 0 182200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3064
timestamp 1654712443
transform 1 0 188200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3065
timestamp 1654712443
transform 1 0 191200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3066
timestamp 1654712443
transform 1 0 194200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3067
timestamp 1654712443
transform 1 0 197200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3068
timestamp 1654712443
transform 1 0 200200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3069
timestamp 1654712443
transform 1 0 203200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3070
timestamp 1654712443
transform 1 0 206200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3071
timestamp 1654712443
transform 1 0 209200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3073
timestamp 1654712443
transform 1 0 215200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3072
timestamp 1654712443
transform 1 0 212200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3074
timestamp 1654712443
transform 1 0 218200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3075
timestamp 1654712443
transform 1 0 221200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3076
timestamp 1654712443
transform 1 0 224200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3077
timestamp 1654712443
transform 1 0 227200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3078
timestamp 1654712443
transform 1 0 230200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3079
timestamp 1654712443
transform 1 0 233200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3080
timestamp 1654712443
transform 1 0 236200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3081
timestamp 1654712443
transform 1 0 239200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3083
timestamp 1654712443
transform 1 0 245200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3082
timestamp 1654712443
transform 1 0 242200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3084
timestamp 1654712443
transform 1 0 248200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3085
timestamp 1654712443
transform 1 0 251200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3086
timestamp 1654712443
transform 1 0 254200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3087
timestamp 1654712443
transform 1 0 257200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3088
timestamp 1654712443
transform 1 0 260200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3089
timestamp 1654712443
transform 1 0 263200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3090
timestamp 1654712443
transform 1 0 266200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3091
timestamp 1654712443
transform 1 0 269200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3092
timestamp 1654712443
transform 1 0 272200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3094
timestamp 1654712443
transform 1 0 278200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3093
timestamp 1654712443
transform 1 0 275200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3095
timestamp 1654712443
transform 1 0 281200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3096
timestamp 1654712443
transform 1 0 284200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3097
timestamp 1654712443
transform 1 0 287200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3098
timestamp 1654712443
transform 1 0 290200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_3099
timestamp 1654712443
transform 1 0 293200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_2901
timestamp 1654712443
transform 1 0 -800 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2900
timestamp 1654712443
transform 1 0 -3800 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2902
timestamp 1654712443
transform 1 0 2200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2903
timestamp 1654712443
transform 1 0 5200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2904
timestamp 1654712443
transform 1 0 8200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2905
timestamp 1654712443
transform 1 0 11200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2906
timestamp 1654712443
transform 1 0 14200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2907
timestamp 1654712443
transform 1 0 17200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2908
timestamp 1654712443
transform 1 0 20200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2909
timestamp 1654712443
transform 1 0 23200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2911
timestamp 1654712443
transform 1 0 29200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2910
timestamp 1654712443
transform 1 0 26200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2912
timestamp 1654712443
transform 1 0 32200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2913
timestamp 1654712443
transform 1 0 35200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2914
timestamp 1654712443
transform 1 0 38200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2915
timestamp 1654712443
transform 1 0 41200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2916
timestamp 1654712443
transform 1 0 44200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2917
timestamp 1654712443
transform 1 0 47200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2918
timestamp 1654712443
transform 1 0 50200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2919
timestamp 1654712443
transform 1 0 53200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2921
timestamp 1654712443
transform 1 0 59200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2920
timestamp 1654712443
transform 1 0 56200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2922
timestamp 1654712443
transform 1 0 62200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2923
timestamp 1654712443
transform 1 0 65200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2924
timestamp 1654712443
transform 1 0 68200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2925
timestamp 1654712443
transform 1 0 71200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2926
timestamp 1654712443
transform 1 0 74200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2927
timestamp 1654712443
transform 1 0 77200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2928
timestamp 1654712443
transform 1 0 80200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2929
timestamp 1654712443
transform 1 0 83200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2930
timestamp 1654712443
transform 1 0 86200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2932
timestamp 1654712443
transform 1 0 92200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2931
timestamp 1654712443
transform 1 0 89200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2933
timestamp 1654712443
transform 1 0 95200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2934
timestamp 1654712443
transform 1 0 98200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2935
timestamp 1654712443
transform 1 0 101200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2936
timestamp 1654712443
transform 1 0 104200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2937
timestamp 1654712443
transform 1 0 107200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2938
timestamp 1654712443
transform 1 0 110200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2939
timestamp 1654712443
transform 1 0 113200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2940
timestamp 1654712443
transform 1 0 116200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2942
timestamp 1654712443
transform 1 0 122200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2941
timestamp 1654712443
transform 1 0 119200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2943
timestamp 1654712443
transform 1 0 125200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2944
timestamp 1654712443
transform 1 0 128200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2945
timestamp 1654712443
transform 1 0 131200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2946
timestamp 1654712443
transform 1 0 134200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2947
timestamp 1654712443
transform 1 0 137200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2948
timestamp 1654712443
transform 1 0 140200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2949
timestamp 1654712443
transform 1 0 143200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2950
timestamp 1654712443
transform 1 0 146200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2952
timestamp 1654712443
transform 1 0 152200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2951
timestamp 1654712443
transform 1 0 149200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2953
timestamp 1654712443
transform 1 0 155200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2954
timestamp 1654712443
transform 1 0 158200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2955
timestamp 1654712443
transform 1 0 161200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2956
timestamp 1654712443
transform 1 0 164200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2957
timestamp 1654712443
transform 1 0 167200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2958
timestamp 1654712443
transform 1 0 170200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2959
timestamp 1654712443
transform 1 0 173200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2960
timestamp 1654712443
transform 1 0 176200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2961
timestamp 1654712443
transform 1 0 179200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2963
timestamp 1654712443
transform 1 0 185200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2962
timestamp 1654712443
transform 1 0 182200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2964
timestamp 1654712443
transform 1 0 188200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2965
timestamp 1654712443
transform 1 0 191200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2966
timestamp 1654712443
transform 1 0 194200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2967
timestamp 1654712443
transform 1 0 197200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2968
timestamp 1654712443
transform 1 0 200200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2969
timestamp 1654712443
transform 1 0 203200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2970
timestamp 1654712443
transform 1 0 206200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2971
timestamp 1654712443
transform 1 0 209200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2973
timestamp 1654712443
transform 1 0 215200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2972
timestamp 1654712443
transform 1 0 212200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2974
timestamp 1654712443
transform 1 0 218200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2975
timestamp 1654712443
transform 1 0 221200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2976
timestamp 1654712443
transform 1 0 224200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2977
timestamp 1654712443
transform 1 0 227200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2978
timestamp 1654712443
transform 1 0 230200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2979
timestamp 1654712443
transform 1 0 233200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2980
timestamp 1654712443
transform 1 0 236200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2981
timestamp 1654712443
transform 1 0 239200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2983
timestamp 1654712443
transform 1 0 245200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2982
timestamp 1654712443
transform 1 0 242200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2984
timestamp 1654712443
transform 1 0 248200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2985
timestamp 1654712443
transform 1 0 251200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2986
timestamp 1654712443
transform 1 0 254200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2987
timestamp 1654712443
transform 1 0 257200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2988
timestamp 1654712443
transform 1 0 260200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2989
timestamp 1654712443
transform 1 0 263200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2990
timestamp 1654712443
transform 1 0 266200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2991
timestamp 1654712443
transform 1 0 269200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2992
timestamp 1654712443
transform 1 0 272200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2994
timestamp 1654712443
transform 1 0 278200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2993
timestamp 1654712443
transform 1 0 275200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2995
timestamp 1654712443
transform 1 0 281200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2996
timestamp 1654712443
transform 1 0 284200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2997
timestamp 1654712443
transform 1 0 287200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2998
timestamp 1654712443
transform 1 0 290200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2999
timestamp 1654712443
transform 1 0 293200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_2801
timestamp 1654712443
transform 1 0 -800 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2800
timestamp 1654712443
transform 1 0 -3800 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2802
timestamp 1654712443
transform 1 0 2200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2803
timestamp 1654712443
transform 1 0 5200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2804
timestamp 1654712443
transform 1 0 8200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2805
timestamp 1654712443
transform 1 0 11200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2806
timestamp 1654712443
transform 1 0 14200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2807
timestamp 1654712443
transform 1 0 17200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2808
timestamp 1654712443
transform 1 0 20200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2809
timestamp 1654712443
transform 1 0 23200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2811
timestamp 1654712443
transform 1 0 29200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2810
timestamp 1654712443
transform 1 0 26200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2812
timestamp 1654712443
transform 1 0 32200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2813
timestamp 1654712443
transform 1 0 35200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2814
timestamp 1654712443
transform 1 0 38200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2815
timestamp 1654712443
transform 1 0 41200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2816
timestamp 1654712443
transform 1 0 44200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2817
timestamp 1654712443
transform 1 0 47200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2818
timestamp 1654712443
transform 1 0 50200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2819
timestamp 1654712443
transform 1 0 53200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2821
timestamp 1654712443
transform 1 0 59200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2820
timestamp 1654712443
transform 1 0 56200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2822
timestamp 1654712443
transform 1 0 62200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2823
timestamp 1654712443
transform 1 0 65200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2824
timestamp 1654712443
transform 1 0 68200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2825
timestamp 1654712443
transform 1 0 71200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2826
timestamp 1654712443
transform 1 0 74200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2827
timestamp 1654712443
transform 1 0 77200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2828
timestamp 1654712443
transform 1 0 80200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2829
timestamp 1654712443
transform 1 0 83200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2830
timestamp 1654712443
transform 1 0 86200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2832
timestamp 1654712443
transform 1 0 92200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2831
timestamp 1654712443
transform 1 0 89200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2833
timestamp 1654712443
transform 1 0 95200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2834
timestamp 1654712443
transform 1 0 98200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2835
timestamp 1654712443
transform 1 0 101200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2836
timestamp 1654712443
transform 1 0 104200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2837
timestamp 1654712443
transform 1 0 107200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2838
timestamp 1654712443
transform 1 0 110200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2839
timestamp 1654712443
transform 1 0 113200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2840
timestamp 1654712443
transform 1 0 116200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2842
timestamp 1654712443
transform 1 0 122200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2841
timestamp 1654712443
transform 1 0 119200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2843
timestamp 1654712443
transform 1 0 125200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2844
timestamp 1654712443
transform 1 0 128200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2845
timestamp 1654712443
transform 1 0 131200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2846
timestamp 1654712443
transform 1 0 134200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2847
timestamp 1654712443
transform 1 0 137200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2848
timestamp 1654712443
transform 1 0 140200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2849
timestamp 1654712443
transform 1 0 143200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2850
timestamp 1654712443
transform 1 0 146200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2852
timestamp 1654712443
transform 1 0 152200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2851
timestamp 1654712443
transform 1 0 149200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2853
timestamp 1654712443
transform 1 0 155200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2854
timestamp 1654712443
transform 1 0 158200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2855
timestamp 1654712443
transform 1 0 161200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2856
timestamp 1654712443
transform 1 0 164200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2857
timestamp 1654712443
transform 1 0 167200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2858
timestamp 1654712443
transform 1 0 170200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2859
timestamp 1654712443
transform 1 0 173200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2860
timestamp 1654712443
transform 1 0 176200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2861
timestamp 1654712443
transform 1 0 179200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2863
timestamp 1654712443
transform 1 0 185200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2862
timestamp 1654712443
transform 1 0 182200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2864
timestamp 1654712443
transform 1 0 188200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2865
timestamp 1654712443
transform 1 0 191200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2866
timestamp 1654712443
transform 1 0 194200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2867
timestamp 1654712443
transform 1 0 197200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2868
timestamp 1654712443
transform 1 0 200200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2869
timestamp 1654712443
transform 1 0 203200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2870
timestamp 1654712443
transform 1 0 206200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2871
timestamp 1654712443
transform 1 0 209200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2873
timestamp 1654712443
transform 1 0 215200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2872
timestamp 1654712443
transform 1 0 212200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2874
timestamp 1654712443
transform 1 0 218200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2875
timestamp 1654712443
transform 1 0 221200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2876
timestamp 1654712443
transform 1 0 224200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2877
timestamp 1654712443
transform 1 0 227200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2878
timestamp 1654712443
transform 1 0 230200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2879
timestamp 1654712443
transform 1 0 233200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2880
timestamp 1654712443
transform 1 0 236200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2881
timestamp 1654712443
transform 1 0 239200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2883
timestamp 1654712443
transform 1 0 245200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2882
timestamp 1654712443
transform 1 0 242200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2884
timestamp 1654712443
transform 1 0 248200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2885
timestamp 1654712443
transform 1 0 251200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2886
timestamp 1654712443
transform 1 0 254200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2887
timestamp 1654712443
transform 1 0 257200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2888
timestamp 1654712443
transform 1 0 260200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2889
timestamp 1654712443
transform 1 0 263200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2890
timestamp 1654712443
transform 1 0 266200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2891
timestamp 1654712443
transform 1 0 269200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2892
timestamp 1654712443
transform 1 0 272200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2894
timestamp 1654712443
transform 1 0 278200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2893
timestamp 1654712443
transform 1 0 275200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2895
timestamp 1654712443
transform 1 0 281200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2896
timestamp 1654712443
transform 1 0 284200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2897
timestamp 1654712443
transform 1 0 287200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2898
timestamp 1654712443
transform 1 0 290200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2899
timestamp 1654712443
transform 1 0 293200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_2601
timestamp 1654712443
transform 1 0 -800 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2600
timestamp 1654712443
transform 1 0 -3800 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2701
timestamp 1654712443
transform 1 0 -800 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2700
timestamp 1654712443
transform 1 0 -3800 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2602
timestamp 1654712443
transform 1 0 2200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2702
timestamp 1654712443
transform 1 0 2200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2603
timestamp 1654712443
transform 1 0 5200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2703
timestamp 1654712443
transform 1 0 5200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2604
timestamp 1654712443
transform 1 0 8200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2704
timestamp 1654712443
transform 1 0 8200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2605
timestamp 1654712443
transform 1 0 11200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2705
timestamp 1654712443
transform 1 0 11200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2606
timestamp 1654712443
transform 1 0 14200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2706
timestamp 1654712443
transform 1 0 14200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2607
timestamp 1654712443
transform 1 0 17200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2707
timestamp 1654712443
transform 1 0 17200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2608
timestamp 1654712443
transform 1 0 20200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2708
timestamp 1654712443
transform 1 0 20200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2609
timestamp 1654712443
transform 1 0 23200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2709
timestamp 1654712443
transform 1 0 23200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2611
timestamp 1654712443
transform 1 0 29200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2610
timestamp 1654712443
transform 1 0 26200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2711
timestamp 1654712443
transform 1 0 29200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2710
timestamp 1654712443
transform 1 0 26200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2612
timestamp 1654712443
transform 1 0 32200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2712
timestamp 1654712443
transform 1 0 32200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2613
timestamp 1654712443
transform 1 0 35200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2713
timestamp 1654712443
transform 1 0 35200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2614
timestamp 1654712443
transform 1 0 38200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2714
timestamp 1654712443
transform 1 0 38200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2615
timestamp 1654712443
transform 1 0 41200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2715
timestamp 1654712443
transform 1 0 41200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2616
timestamp 1654712443
transform 1 0 44200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2716
timestamp 1654712443
transform 1 0 44200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2617
timestamp 1654712443
transform 1 0 47200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2717
timestamp 1654712443
transform 1 0 47200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2618
timestamp 1654712443
transform 1 0 50200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2718
timestamp 1654712443
transform 1 0 50200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2619
timestamp 1654712443
transform 1 0 53200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2719
timestamp 1654712443
transform 1 0 53200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2621
timestamp 1654712443
transform 1 0 59200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2620
timestamp 1654712443
transform 1 0 56200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2721
timestamp 1654712443
transform 1 0 59200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2720
timestamp 1654712443
transform 1 0 56200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2622
timestamp 1654712443
transform 1 0 62200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2722
timestamp 1654712443
transform 1 0 62200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2623
timestamp 1654712443
transform 1 0 65200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2723
timestamp 1654712443
transform 1 0 65200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2624
timestamp 1654712443
transform 1 0 68200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2724
timestamp 1654712443
transform 1 0 68200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2625
timestamp 1654712443
transform 1 0 71200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2725
timestamp 1654712443
transform 1 0 71200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2626
timestamp 1654712443
transform 1 0 74200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2726
timestamp 1654712443
transform 1 0 74200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2627
timestamp 1654712443
transform 1 0 77200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2727
timestamp 1654712443
transform 1 0 77200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2628
timestamp 1654712443
transform 1 0 80200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2728
timestamp 1654712443
transform 1 0 80200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2629
timestamp 1654712443
transform 1 0 83200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2729
timestamp 1654712443
transform 1 0 83200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2630
timestamp 1654712443
transform 1 0 86200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2730
timestamp 1654712443
transform 1 0 86200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2632
timestamp 1654712443
transform 1 0 92200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2631
timestamp 1654712443
transform 1 0 89200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2732
timestamp 1654712443
transform 1 0 92200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2731
timestamp 1654712443
transform 1 0 89200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2633
timestamp 1654712443
transform 1 0 95200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2733
timestamp 1654712443
transform 1 0 95200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2634
timestamp 1654712443
transform 1 0 98200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2734
timestamp 1654712443
transform 1 0 98200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2635
timestamp 1654712443
transform 1 0 101200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2735
timestamp 1654712443
transform 1 0 101200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2636
timestamp 1654712443
transform 1 0 104200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2736
timestamp 1654712443
transform 1 0 104200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2637
timestamp 1654712443
transform 1 0 107200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2737
timestamp 1654712443
transform 1 0 107200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2638
timestamp 1654712443
transform 1 0 110200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2738
timestamp 1654712443
transform 1 0 110200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2639
timestamp 1654712443
transform 1 0 113200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2739
timestamp 1654712443
transform 1 0 113200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2640
timestamp 1654712443
transform 1 0 116200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2740
timestamp 1654712443
transform 1 0 116200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2642
timestamp 1654712443
transform 1 0 122200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2641
timestamp 1654712443
transform 1 0 119200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2742
timestamp 1654712443
transform 1 0 122200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2741
timestamp 1654712443
transform 1 0 119200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2643
timestamp 1654712443
transform 1 0 125200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2743
timestamp 1654712443
transform 1 0 125200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2644
timestamp 1654712443
transform 1 0 128200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2744
timestamp 1654712443
transform 1 0 128200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2645
timestamp 1654712443
transform 1 0 131200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2745
timestamp 1654712443
transform 1 0 131200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2646
timestamp 1654712443
transform 1 0 134200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2746
timestamp 1654712443
transform 1 0 134200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2647
timestamp 1654712443
transform 1 0 137200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2747
timestamp 1654712443
transform 1 0 137200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2648
timestamp 1654712443
transform 1 0 140200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2748
timestamp 1654712443
transform 1 0 140200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2649
timestamp 1654712443
transform 1 0 143200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2749
timestamp 1654712443
transform 1 0 143200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2650
timestamp 1654712443
transform 1 0 146200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2750
timestamp 1654712443
transform 1 0 146200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2652
timestamp 1654712443
transform 1 0 152200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2651
timestamp 1654712443
transform 1 0 149200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2752
timestamp 1654712443
transform 1 0 152200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2751
timestamp 1654712443
transform 1 0 149200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2653
timestamp 1654712443
transform 1 0 155200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2753
timestamp 1654712443
transform 1 0 155200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2654
timestamp 1654712443
transform 1 0 158200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2754
timestamp 1654712443
transform 1 0 158200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2655
timestamp 1654712443
transform 1 0 161200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2755
timestamp 1654712443
transform 1 0 161200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2656
timestamp 1654712443
transform 1 0 164200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2756
timestamp 1654712443
transform 1 0 164200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2657
timestamp 1654712443
transform 1 0 167200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2757
timestamp 1654712443
transform 1 0 167200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2658
timestamp 1654712443
transform 1 0 170200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2758
timestamp 1654712443
transform 1 0 170200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2659
timestamp 1654712443
transform 1 0 173200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2759
timestamp 1654712443
transform 1 0 173200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2660
timestamp 1654712443
transform 1 0 176200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2760
timestamp 1654712443
transform 1 0 176200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2661
timestamp 1654712443
transform 1 0 179200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2761
timestamp 1654712443
transform 1 0 179200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2663
timestamp 1654712443
transform 1 0 185200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2662
timestamp 1654712443
transform 1 0 182200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2763
timestamp 1654712443
transform 1 0 185200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2762
timestamp 1654712443
transform 1 0 182200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2664
timestamp 1654712443
transform 1 0 188200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2764
timestamp 1654712443
transform 1 0 188200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2665
timestamp 1654712443
transform 1 0 191200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2765
timestamp 1654712443
transform 1 0 191200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2666
timestamp 1654712443
transform 1 0 194200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2766
timestamp 1654712443
transform 1 0 194200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2667
timestamp 1654712443
transform 1 0 197200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2767
timestamp 1654712443
transform 1 0 197200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2668
timestamp 1654712443
transform 1 0 200200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2768
timestamp 1654712443
transform 1 0 200200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2669
timestamp 1654712443
transform 1 0 203200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2769
timestamp 1654712443
transform 1 0 203200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2670
timestamp 1654712443
transform 1 0 206200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2770
timestamp 1654712443
transform 1 0 206200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2671
timestamp 1654712443
transform 1 0 209200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2771
timestamp 1654712443
transform 1 0 209200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2673
timestamp 1654712443
transform 1 0 215200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2672
timestamp 1654712443
transform 1 0 212200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2773
timestamp 1654712443
transform 1 0 215200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2772
timestamp 1654712443
transform 1 0 212200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2674
timestamp 1654712443
transform 1 0 218200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2774
timestamp 1654712443
transform 1 0 218200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2675
timestamp 1654712443
transform 1 0 221200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2775
timestamp 1654712443
transform 1 0 221200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2676
timestamp 1654712443
transform 1 0 224200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2776
timestamp 1654712443
transform 1 0 224200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2677
timestamp 1654712443
transform 1 0 227200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2777
timestamp 1654712443
transform 1 0 227200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2678
timestamp 1654712443
transform 1 0 230200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2778
timestamp 1654712443
transform 1 0 230200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2679
timestamp 1654712443
transform 1 0 233200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2779
timestamp 1654712443
transform 1 0 233200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2680
timestamp 1654712443
transform 1 0 236200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2780
timestamp 1654712443
transform 1 0 236200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2681
timestamp 1654712443
transform 1 0 239200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2781
timestamp 1654712443
transform 1 0 239200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2683
timestamp 1654712443
transform 1 0 245200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2682
timestamp 1654712443
transform 1 0 242200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2783
timestamp 1654712443
transform 1 0 245200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2782
timestamp 1654712443
transform 1 0 242200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2684
timestamp 1654712443
transform 1 0 248200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2784
timestamp 1654712443
transform 1 0 248200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2685
timestamp 1654712443
transform 1 0 251200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2785
timestamp 1654712443
transform 1 0 251200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2686
timestamp 1654712443
transform 1 0 254200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2786
timestamp 1654712443
transform 1 0 254200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2687
timestamp 1654712443
transform 1 0 257200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2787
timestamp 1654712443
transform 1 0 257200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2688
timestamp 1654712443
transform 1 0 260200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2788
timestamp 1654712443
transform 1 0 260200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2689
timestamp 1654712443
transform 1 0 263200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2789
timestamp 1654712443
transform 1 0 263200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2690
timestamp 1654712443
transform 1 0 266200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2790
timestamp 1654712443
transform 1 0 266200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2691
timestamp 1654712443
transform 1 0 269200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2791
timestamp 1654712443
transform 1 0 269200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2692
timestamp 1654712443
transform 1 0 272200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2792
timestamp 1654712443
transform 1 0 272200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2694
timestamp 1654712443
transform 1 0 278200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2693
timestamp 1654712443
transform 1 0 275200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2794
timestamp 1654712443
transform 1 0 278200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2793
timestamp 1654712443
transform 1 0 275200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2695
timestamp 1654712443
transform 1 0 281200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2795
timestamp 1654712443
transform 1 0 281200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2696
timestamp 1654712443
transform 1 0 284200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2796
timestamp 1654712443
transform 1 0 284200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2697
timestamp 1654712443
transform 1 0 287200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2797
timestamp 1654712443
transform 1 0 287200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2698
timestamp 1654712443
transform 1 0 290200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2798
timestamp 1654712443
transform 1 0 290200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2699
timestamp 1654712443
transform 1 0 293200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_2799
timestamp 1654712443
transform 1 0 293200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_2501
timestamp 1654712443
transform 1 0 -800 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2500
timestamp 1654712443
transform 1 0 -3800 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2502
timestamp 1654712443
transform 1 0 2200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2503
timestamp 1654712443
transform 1 0 5200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2504
timestamp 1654712443
transform 1 0 8200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2505
timestamp 1654712443
transform 1 0 11200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2506
timestamp 1654712443
transform 1 0 14200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2507
timestamp 1654712443
transform 1 0 17200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2508
timestamp 1654712443
transform 1 0 20200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2509
timestamp 1654712443
transform 1 0 23200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2511
timestamp 1654712443
transform 1 0 29200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2510
timestamp 1654712443
transform 1 0 26200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2512
timestamp 1654712443
transform 1 0 32200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2513
timestamp 1654712443
transform 1 0 35200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2514
timestamp 1654712443
transform 1 0 38200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2515
timestamp 1654712443
transform 1 0 41200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2516
timestamp 1654712443
transform 1 0 44200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2517
timestamp 1654712443
transform 1 0 47200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2518
timestamp 1654712443
transform 1 0 50200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2519
timestamp 1654712443
transform 1 0 53200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2521
timestamp 1654712443
transform 1 0 59200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2520
timestamp 1654712443
transform 1 0 56200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2522
timestamp 1654712443
transform 1 0 62200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2523
timestamp 1654712443
transform 1 0 65200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2524
timestamp 1654712443
transform 1 0 68200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2525
timestamp 1654712443
transform 1 0 71200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2526
timestamp 1654712443
transform 1 0 74200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2527
timestamp 1654712443
transform 1 0 77200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2528
timestamp 1654712443
transform 1 0 80200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2529
timestamp 1654712443
transform 1 0 83200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2530
timestamp 1654712443
transform 1 0 86200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2532
timestamp 1654712443
transform 1 0 92200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2531
timestamp 1654712443
transform 1 0 89200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2533
timestamp 1654712443
transform 1 0 95200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2534
timestamp 1654712443
transform 1 0 98200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2535
timestamp 1654712443
transform 1 0 101200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2536
timestamp 1654712443
transform 1 0 104200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2537
timestamp 1654712443
transform 1 0 107200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2538
timestamp 1654712443
transform 1 0 110200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2539
timestamp 1654712443
transform 1 0 113200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2540
timestamp 1654712443
transform 1 0 116200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2542
timestamp 1654712443
transform 1 0 122200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2541
timestamp 1654712443
transform 1 0 119200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2543
timestamp 1654712443
transform 1 0 125200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2544
timestamp 1654712443
transform 1 0 128200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2545
timestamp 1654712443
transform 1 0 131200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2546
timestamp 1654712443
transform 1 0 134200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2547
timestamp 1654712443
transform 1 0 137200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2548
timestamp 1654712443
transform 1 0 140200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2549
timestamp 1654712443
transform 1 0 143200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2550
timestamp 1654712443
transform 1 0 146200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2552
timestamp 1654712443
transform 1 0 152200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2551
timestamp 1654712443
transform 1 0 149200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2553
timestamp 1654712443
transform 1 0 155200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2554
timestamp 1654712443
transform 1 0 158200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2555
timestamp 1654712443
transform 1 0 161200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2556
timestamp 1654712443
transform 1 0 164200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2557
timestamp 1654712443
transform 1 0 167200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2558
timestamp 1654712443
transform 1 0 170200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2559
timestamp 1654712443
transform 1 0 173200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2560
timestamp 1654712443
transform 1 0 176200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2561
timestamp 1654712443
transform 1 0 179200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2563
timestamp 1654712443
transform 1 0 185200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2562
timestamp 1654712443
transform 1 0 182200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2564
timestamp 1654712443
transform 1 0 188200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2565
timestamp 1654712443
transform 1 0 191200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2566
timestamp 1654712443
transform 1 0 194200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2567
timestamp 1654712443
transform 1 0 197200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2568
timestamp 1654712443
transform 1 0 200200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2569
timestamp 1654712443
transform 1 0 203200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2570
timestamp 1654712443
transform 1 0 206200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2571
timestamp 1654712443
transform 1 0 209200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2573
timestamp 1654712443
transform 1 0 215200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2572
timestamp 1654712443
transform 1 0 212200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2574
timestamp 1654712443
transform 1 0 218200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2575
timestamp 1654712443
transform 1 0 221200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2576
timestamp 1654712443
transform 1 0 224200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2577
timestamp 1654712443
transform 1 0 227200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2578
timestamp 1654712443
transform 1 0 230200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2579
timestamp 1654712443
transform 1 0 233200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2580
timestamp 1654712443
transform 1 0 236200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2581
timestamp 1654712443
transform 1 0 239200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2583
timestamp 1654712443
transform 1 0 245200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2582
timestamp 1654712443
transform 1 0 242200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2584
timestamp 1654712443
transform 1 0 248200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2585
timestamp 1654712443
transform 1 0 251200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2586
timestamp 1654712443
transform 1 0 254200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2587
timestamp 1654712443
transform 1 0 257200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2588
timestamp 1654712443
transform 1 0 260200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2589
timestamp 1654712443
transform 1 0 263200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2590
timestamp 1654712443
transform 1 0 266200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2591
timestamp 1654712443
transform 1 0 269200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2592
timestamp 1654712443
transform 1 0 272200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2594
timestamp 1654712443
transform 1 0 278200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2593
timestamp 1654712443
transform 1 0 275200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2595
timestamp 1654712443
transform 1 0 281200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2596
timestamp 1654712443
transform 1 0 284200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2597
timestamp 1654712443
transform 1 0 287200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2598
timestamp 1654712443
transform 1 0 290200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2599
timestamp 1654712443
transform 1 0 293200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_2401
timestamp 1654712443
transform 1 0 -800 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2400
timestamp 1654712443
transform 1 0 -3800 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2402
timestamp 1654712443
transform 1 0 2200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2403
timestamp 1654712443
transform 1 0 5200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2404
timestamp 1654712443
transform 1 0 8200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2405
timestamp 1654712443
transform 1 0 11200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2406
timestamp 1654712443
transform 1 0 14200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2407
timestamp 1654712443
transform 1 0 17200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2408
timestamp 1654712443
transform 1 0 20200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2409
timestamp 1654712443
transform 1 0 23200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2411
timestamp 1654712443
transform 1 0 29200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2410
timestamp 1654712443
transform 1 0 26200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2412
timestamp 1654712443
transform 1 0 32200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2413
timestamp 1654712443
transform 1 0 35200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2414
timestamp 1654712443
transform 1 0 38200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2415
timestamp 1654712443
transform 1 0 41200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2416
timestamp 1654712443
transform 1 0 44200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2417
timestamp 1654712443
transform 1 0 47200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2418
timestamp 1654712443
transform 1 0 50200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2419
timestamp 1654712443
transform 1 0 53200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2421
timestamp 1654712443
transform 1 0 59200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2420
timestamp 1654712443
transform 1 0 56200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2422
timestamp 1654712443
transform 1 0 62200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2423
timestamp 1654712443
transform 1 0 65200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2424
timestamp 1654712443
transform 1 0 68200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2425
timestamp 1654712443
transform 1 0 71200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2426
timestamp 1654712443
transform 1 0 74200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2427
timestamp 1654712443
transform 1 0 77200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2428
timestamp 1654712443
transform 1 0 80200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2429
timestamp 1654712443
transform 1 0 83200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2430
timestamp 1654712443
transform 1 0 86200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2432
timestamp 1654712443
transform 1 0 92200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2431
timestamp 1654712443
transform 1 0 89200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2433
timestamp 1654712443
transform 1 0 95200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2434
timestamp 1654712443
transform 1 0 98200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2435
timestamp 1654712443
transform 1 0 101200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2436
timestamp 1654712443
transform 1 0 104200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2437
timestamp 1654712443
transform 1 0 107200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2438
timestamp 1654712443
transform 1 0 110200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2439
timestamp 1654712443
transform 1 0 113200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2440
timestamp 1654712443
transform 1 0 116200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2442
timestamp 1654712443
transform 1 0 122200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2441
timestamp 1654712443
transform 1 0 119200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2443
timestamp 1654712443
transform 1 0 125200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2444
timestamp 1654712443
transform 1 0 128200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2445
timestamp 1654712443
transform 1 0 131200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2446
timestamp 1654712443
transform 1 0 134200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2447
timestamp 1654712443
transform 1 0 137200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2448
timestamp 1654712443
transform 1 0 140200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2449
timestamp 1654712443
transform 1 0 143200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2450
timestamp 1654712443
transform 1 0 146200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2452
timestamp 1654712443
transform 1 0 152200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2451
timestamp 1654712443
transform 1 0 149200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2453
timestamp 1654712443
transform 1 0 155200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2454
timestamp 1654712443
transform 1 0 158200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2455
timestamp 1654712443
transform 1 0 161200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2456
timestamp 1654712443
transform 1 0 164200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2457
timestamp 1654712443
transform 1 0 167200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2458
timestamp 1654712443
transform 1 0 170200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2459
timestamp 1654712443
transform 1 0 173200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2460
timestamp 1654712443
transform 1 0 176200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2461
timestamp 1654712443
transform 1 0 179200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2463
timestamp 1654712443
transform 1 0 185200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2462
timestamp 1654712443
transform 1 0 182200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2464
timestamp 1654712443
transform 1 0 188200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2465
timestamp 1654712443
transform 1 0 191200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2466
timestamp 1654712443
transform 1 0 194200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2467
timestamp 1654712443
transform 1 0 197200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2468
timestamp 1654712443
transform 1 0 200200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2469
timestamp 1654712443
transform 1 0 203200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2470
timestamp 1654712443
transform 1 0 206200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2471
timestamp 1654712443
transform 1 0 209200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2473
timestamp 1654712443
transform 1 0 215200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2472
timestamp 1654712443
transform 1 0 212200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2474
timestamp 1654712443
transform 1 0 218200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2475
timestamp 1654712443
transform 1 0 221200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2476
timestamp 1654712443
transform 1 0 224200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2477
timestamp 1654712443
transform 1 0 227200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2478
timestamp 1654712443
transform 1 0 230200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2479
timestamp 1654712443
transform 1 0 233200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2480
timestamp 1654712443
transform 1 0 236200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2481
timestamp 1654712443
transform 1 0 239200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2483
timestamp 1654712443
transform 1 0 245200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2482
timestamp 1654712443
transform 1 0 242200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2484
timestamp 1654712443
transform 1 0 248200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2485
timestamp 1654712443
transform 1 0 251200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2486
timestamp 1654712443
transform 1 0 254200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2487
timestamp 1654712443
transform 1 0 257200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2488
timestamp 1654712443
transform 1 0 260200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2489
timestamp 1654712443
transform 1 0 263200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2490
timestamp 1654712443
transform 1 0 266200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2491
timestamp 1654712443
transform 1 0 269200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2492
timestamp 1654712443
transform 1 0 272200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2494
timestamp 1654712443
transform 1 0 278200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2493
timestamp 1654712443
transform 1 0 275200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2495
timestamp 1654712443
transform 1 0 281200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2496
timestamp 1654712443
transform 1 0 284200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2497
timestamp 1654712443
transform 1 0 287200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2498
timestamp 1654712443
transform 1 0 290200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2499
timestamp 1654712443
transform 1 0 293200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_2301
timestamp 1654712443
transform 1 0 -800 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2300
timestamp 1654712443
transform 1 0 -3800 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2302
timestamp 1654712443
transform 1 0 2200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2303
timestamp 1654712443
transform 1 0 5200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2304
timestamp 1654712443
transform 1 0 8200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2305
timestamp 1654712443
transform 1 0 11200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2306
timestamp 1654712443
transform 1 0 14200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2307
timestamp 1654712443
transform 1 0 17200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2308
timestamp 1654712443
transform 1 0 20200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2309
timestamp 1654712443
transform 1 0 23200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2311
timestamp 1654712443
transform 1 0 29200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2310
timestamp 1654712443
transform 1 0 26200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2312
timestamp 1654712443
transform 1 0 32200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2313
timestamp 1654712443
transform 1 0 35200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2314
timestamp 1654712443
transform 1 0 38200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2315
timestamp 1654712443
transform 1 0 41200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2316
timestamp 1654712443
transform 1 0 44200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2317
timestamp 1654712443
transform 1 0 47200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2318
timestamp 1654712443
transform 1 0 50200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2319
timestamp 1654712443
transform 1 0 53200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2321
timestamp 1654712443
transform 1 0 59200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2320
timestamp 1654712443
transform 1 0 56200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2322
timestamp 1654712443
transform 1 0 62200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2323
timestamp 1654712443
transform 1 0 65200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2324
timestamp 1654712443
transform 1 0 68200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2325
timestamp 1654712443
transform 1 0 71200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2326
timestamp 1654712443
transform 1 0 74200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2327
timestamp 1654712443
transform 1 0 77200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2328
timestamp 1654712443
transform 1 0 80200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2329
timestamp 1654712443
transform 1 0 83200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2330
timestamp 1654712443
transform 1 0 86200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2332
timestamp 1654712443
transform 1 0 92200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2331
timestamp 1654712443
transform 1 0 89200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2333
timestamp 1654712443
transform 1 0 95200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2334
timestamp 1654712443
transform 1 0 98200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2335
timestamp 1654712443
transform 1 0 101200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2336
timestamp 1654712443
transform 1 0 104200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2337
timestamp 1654712443
transform 1 0 107200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2338
timestamp 1654712443
transform 1 0 110200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2339
timestamp 1654712443
transform 1 0 113200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2340
timestamp 1654712443
transform 1 0 116200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2342
timestamp 1654712443
transform 1 0 122200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2341
timestamp 1654712443
transform 1 0 119200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2343
timestamp 1654712443
transform 1 0 125200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2344
timestamp 1654712443
transform 1 0 128200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2345
timestamp 1654712443
transform 1 0 131200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2346
timestamp 1654712443
transform 1 0 134200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2347
timestamp 1654712443
transform 1 0 137200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2348
timestamp 1654712443
transform 1 0 140200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2349
timestamp 1654712443
transform 1 0 143200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2350
timestamp 1654712443
transform 1 0 146200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2352
timestamp 1654712443
transform 1 0 152200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2351
timestamp 1654712443
transform 1 0 149200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2353
timestamp 1654712443
transform 1 0 155200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2354
timestamp 1654712443
transform 1 0 158200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2355
timestamp 1654712443
transform 1 0 161200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2356
timestamp 1654712443
transform 1 0 164200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2357
timestamp 1654712443
transform 1 0 167200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2358
timestamp 1654712443
transform 1 0 170200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2359
timestamp 1654712443
transform 1 0 173200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2360
timestamp 1654712443
transform 1 0 176200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2361
timestamp 1654712443
transform 1 0 179200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2363
timestamp 1654712443
transform 1 0 185200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2362
timestamp 1654712443
transform 1 0 182200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2364
timestamp 1654712443
transform 1 0 188200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2365
timestamp 1654712443
transform 1 0 191200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2366
timestamp 1654712443
transform 1 0 194200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2367
timestamp 1654712443
transform 1 0 197200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2368
timestamp 1654712443
transform 1 0 200200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2369
timestamp 1654712443
transform 1 0 203200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2370
timestamp 1654712443
transform 1 0 206200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2371
timestamp 1654712443
transform 1 0 209200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2373
timestamp 1654712443
transform 1 0 215200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2372
timestamp 1654712443
transform 1 0 212200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2374
timestamp 1654712443
transform 1 0 218200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2375
timestamp 1654712443
transform 1 0 221200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2376
timestamp 1654712443
transform 1 0 224200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2377
timestamp 1654712443
transform 1 0 227200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2378
timestamp 1654712443
transform 1 0 230200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2379
timestamp 1654712443
transform 1 0 233200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2380
timestamp 1654712443
transform 1 0 236200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2381
timestamp 1654712443
transform 1 0 239200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2383
timestamp 1654712443
transform 1 0 245200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2382
timestamp 1654712443
transform 1 0 242200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2384
timestamp 1654712443
transform 1 0 248200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2385
timestamp 1654712443
transform 1 0 251200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2386
timestamp 1654712443
transform 1 0 254200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2387
timestamp 1654712443
transform 1 0 257200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2388
timestamp 1654712443
transform 1 0 260200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2389
timestamp 1654712443
transform 1 0 263200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2390
timestamp 1654712443
transform 1 0 266200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2391
timestamp 1654712443
transform 1 0 269200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2392
timestamp 1654712443
transform 1 0 272200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2394
timestamp 1654712443
transform 1 0 278200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2393
timestamp 1654712443
transform 1 0 275200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2395
timestamp 1654712443
transform 1 0 281200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2396
timestamp 1654712443
transform 1 0 284200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2397
timestamp 1654712443
transform 1 0 287200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2398
timestamp 1654712443
transform 1 0 290200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2399
timestamp 1654712443
transform 1 0 293200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_2201
timestamp 1654712443
transform 1 0 -800 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2200
timestamp 1654712443
transform 1 0 -3800 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2202
timestamp 1654712443
transform 1 0 2200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2203
timestamp 1654712443
transform 1 0 5200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2204
timestamp 1654712443
transform 1 0 8200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2205
timestamp 1654712443
transform 1 0 11200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2206
timestamp 1654712443
transform 1 0 14200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2207
timestamp 1654712443
transform 1 0 17200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2208
timestamp 1654712443
transform 1 0 20200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2209
timestamp 1654712443
transform 1 0 23200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2211
timestamp 1654712443
transform 1 0 29200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2210
timestamp 1654712443
transform 1 0 26200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2212
timestamp 1654712443
transform 1 0 32200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2213
timestamp 1654712443
transform 1 0 35200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2214
timestamp 1654712443
transform 1 0 38200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2215
timestamp 1654712443
transform 1 0 41200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2216
timestamp 1654712443
transform 1 0 44200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2217
timestamp 1654712443
transform 1 0 47200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2218
timestamp 1654712443
transform 1 0 50200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2219
timestamp 1654712443
transform 1 0 53200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2221
timestamp 1654712443
transform 1 0 59200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2220
timestamp 1654712443
transform 1 0 56200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2222
timestamp 1654712443
transform 1 0 62200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2223
timestamp 1654712443
transform 1 0 65200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2224
timestamp 1654712443
transform 1 0 68200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2225
timestamp 1654712443
transform 1 0 71200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2226
timestamp 1654712443
transform 1 0 74200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2227
timestamp 1654712443
transform 1 0 77200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2228
timestamp 1654712443
transform 1 0 80200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2229
timestamp 1654712443
transform 1 0 83200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2230
timestamp 1654712443
transform 1 0 86200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2232
timestamp 1654712443
transform 1 0 92200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2231
timestamp 1654712443
transform 1 0 89200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2233
timestamp 1654712443
transform 1 0 95200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2234
timestamp 1654712443
transform 1 0 98200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2235
timestamp 1654712443
transform 1 0 101200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2236
timestamp 1654712443
transform 1 0 104200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2237
timestamp 1654712443
transform 1 0 107200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2238
timestamp 1654712443
transform 1 0 110200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2239
timestamp 1654712443
transform 1 0 113200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2240
timestamp 1654712443
transform 1 0 116200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2242
timestamp 1654712443
transform 1 0 122200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2241
timestamp 1654712443
transform 1 0 119200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2243
timestamp 1654712443
transform 1 0 125200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2244
timestamp 1654712443
transform 1 0 128200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2245
timestamp 1654712443
transform 1 0 131200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2246
timestamp 1654712443
transform 1 0 134200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2247
timestamp 1654712443
transform 1 0 137200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2248
timestamp 1654712443
transform 1 0 140200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2249
timestamp 1654712443
transform 1 0 143200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2250
timestamp 1654712443
transform 1 0 146200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2252
timestamp 1654712443
transform 1 0 152200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2251
timestamp 1654712443
transform 1 0 149200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2253
timestamp 1654712443
transform 1 0 155200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2254
timestamp 1654712443
transform 1 0 158200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2255
timestamp 1654712443
transform 1 0 161200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2256
timestamp 1654712443
transform 1 0 164200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2257
timestamp 1654712443
transform 1 0 167200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2258
timestamp 1654712443
transform 1 0 170200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2259
timestamp 1654712443
transform 1 0 173200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2260
timestamp 1654712443
transform 1 0 176200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2261
timestamp 1654712443
transform 1 0 179200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2263
timestamp 1654712443
transform 1 0 185200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2262
timestamp 1654712443
transform 1 0 182200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2264
timestamp 1654712443
transform 1 0 188200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2265
timestamp 1654712443
transform 1 0 191200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2266
timestamp 1654712443
transform 1 0 194200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2267
timestamp 1654712443
transform 1 0 197200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2268
timestamp 1654712443
transform 1 0 200200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2269
timestamp 1654712443
transform 1 0 203200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2270
timestamp 1654712443
transform 1 0 206200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2271
timestamp 1654712443
transform 1 0 209200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2273
timestamp 1654712443
transform 1 0 215200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2272
timestamp 1654712443
transform 1 0 212200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2274
timestamp 1654712443
transform 1 0 218200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2275
timestamp 1654712443
transform 1 0 221200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2276
timestamp 1654712443
transform 1 0 224200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2277
timestamp 1654712443
transform 1 0 227200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2278
timestamp 1654712443
transform 1 0 230200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2279
timestamp 1654712443
transform 1 0 233200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2280
timestamp 1654712443
transform 1 0 236200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2281
timestamp 1654712443
transform 1 0 239200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2283
timestamp 1654712443
transform 1 0 245200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2282
timestamp 1654712443
transform 1 0 242200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2284
timestamp 1654712443
transform 1 0 248200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2285
timestamp 1654712443
transform 1 0 251200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2286
timestamp 1654712443
transform 1 0 254200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2287
timestamp 1654712443
transform 1 0 257200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2288
timestamp 1654712443
transform 1 0 260200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2289
timestamp 1654712443
transform 1 0 263200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2290
timestamp 1654712443
transform 1 0 266200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2291
timestamp 1654712443
transform 1 0 269200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2292
timestamp 1654712443
transform 1 0 272200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2294
timestamp 1654712443
transform 1 0 278200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2293
timestamp 1654712443
transform 1 0 275200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2295
timestamp 1654712443
transform 1 0 281200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2296
timestamp 1654712443
transform 1 0 284200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2297
timestamp 1654712443
transform 1 0 287200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2298
timestamp 1654712443
transform 1 0 290200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2299
timestamp 1654712443
transform 1 0 293200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_2101
timestamp 1654712443
transform 1 0 -800 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2100
timestamp 1654712443
transform 1 0 -3800 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2102
timestamp 1654712443
transform 1 0 2200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2103
timestamp 1654712443
transform 1 0 5200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2104
timestamp 1654712443
transform 1 0 8200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2105
timestamp 1654712443
transform 1 0 11200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2106
timestamp 1654712443
transform 1 0 14200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2107
timestamp 1654712443
transform 1 0 17200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2108
timestamp 1654712443
transform 1 0 20200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2109
timestamp 1654712443
transform 1 0 23200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2111
timestamp 1654712443
transform 1 0 29200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2110
timestamp 1654712443
transform 1 0 26200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2112
timestamp 1654712443
transform 1 0 32200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2113
timestamp 1654712443
transform 1 0 35200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2114
timestamp 1654712443
transform 1 0 38200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2115
timestamp 1654712443
transform 1 0 41200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2116
timestamp 1654712443
transform 1 0 44200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2117
timestamp 1654712443
transform 1 0 47200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2118
timestamp 1654712443
transform 1 0 50200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2119
timestamp 1654712443
transform 1 0 53200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2121
timestamp 1654712443
transform 1 0 59200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2120
timestamp 1654712443
transform 1 0 56200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2122
timestamp 1654712443
transform 1 0 62200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2123
timestamp 1654712443
transform 1 0 65200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2124
timestamp 1654712443
transform 1 0 68200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2125
timestamp 1654712443
transform 1 0 71200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2126
timestamp 1654712443
transform 1 0 74200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2127
timestamp 1654712443
transform 1 0 77200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2128
timestamp 1654712443
transform 1 0 80200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2129
timestamp 1654712443
transform 1 0 83200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2130
timestamp 1654712443
transform 1 0 86200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2132
timestamp 1654712443
transform 1 0 92200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2131
timestamp 1654712443
transform 1 0 89200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2133
timestamp 1654712443
transform 1 0 95200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2134
timestamp 1654712443
transform 1 0 98200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2135
timestamp 1654712443
transform 1 0 101200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2136
timestamp 1654712443
transform 1 0 104200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2137
timestamp 1654712443
transform 1 0 107200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2138
timestamp 1654712443
transform 1 0 110200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2139
timestamp 1654712443
transform 1 0 113200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2140
timestamp 1654712443
transform 1 0 116200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2142
timestamp 1654712443
transform 1 0 122200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2141
timestamp 1654712443
transform 1 0 119200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2143
timestamp 1654712443
transform 1 0 125200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2144
timestamp 1654712443
transform 1 0 128200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2145
timestamp 1654712443
transform 1 0 131200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2146
timestamp 1654712443
transform 1 0 134200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2147
timestamp 1654712443
transform 1 0 137200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2148
timestamp 1654712443
transform 1 0 140200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2149
timestamp 1654712443
transform 1 0 143200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2150
timestamp 1654712443
transform 1 0 146200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2152
timestamp 1654712443
transform 1 0 152200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2151
timestamp 1654712443
transform 1 0 149200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2153
timestamp 1654712443
transform 1 0 155200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2154
timestamp 1654712443
transform 1 0 158200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2155
timestamp 1654712443
transform 1 0 161200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2156
timestamp 1654712443
transform 1 0 164200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2157
timestamp 1654712443
transform 1 0 167200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2158
timestamp 1654712443
transform 1 0 170200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2159
timestamp 1654712443
transform 1 0 173200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2160
timestamp 1654712443
transform 1 0 176200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2161
timestamp 1654712443
transform 1 0 179200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2163
timestamp 1654712443
transform 1 0 185200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2162
timestamp 1654712443
transform 1 0 182200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2164
timestamp 1654712443
transform 1 0 188200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2165
timestamp 1654712443
transform 1 0 191200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2166
timestamp 1654712443
transform 1 0 194200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2167
timestamp 1654712443
transform 1 0 197200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2168
timestamp 1654712443
transform 1 0 200200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2169
timestamp 1654712443
transform 1 0 203200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2170
timestamp 1654712443
transform 1 0 206200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2171
timestamp 1654712443
transform 1 0 209200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2173
timestamp 1654712443
transform 1 0 215200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2172
timestamp 1654712443
transform 1 0 212200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2174
timestamp 1654712443
transform 1 0 218200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2175
timestamp 1654712443
transform 1 0 221200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2176
timestamp 1654712443
transform 1 0 224200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2177
timestamp 1654712443
transform 1 0 227200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2178
timestamp 1654712443
transform 1 0 230200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2179
timestamp 1654712443
transform 1 0 233200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2180
timestamp 1654712443
transform 1 0 236200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2181
timestamp 1654712443
transform 1 0 239200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2183
timestamp 1654712443
transform 1 0 245200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2182
timestamp 1654712443
transform 1 0 242200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2184
timestamp 1654712443
transform 1 0 248200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2185
timestamp 1654712443
transform 1 0 251200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2186
timestamp 1654712443
transform 1 0 254200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2187
timestamp 1654712443
transform 1 0 257200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2188
timestamp 1654712443
transform 1 0 260200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2189
timestamp 1654712443
transform 1 0 263200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2190
timestamp 1654712443
transform 1 0 266200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2191
timestamp 1654712443
transform 1 0 269200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2192
timestamp 1654712443
transform 1 0 272200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2194
timestamp 1654712443
transform 1 0 278200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2193
timestamp 1654712443
transform 1 0 275200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2195
timestamp 1654712443
transform 1 0 281200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2196
timestamp 1654712443
transform 1 0 284200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2197
timestamp 1654712443
transform 1 0 287200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2198
timestamp 1654712443
transform 1 0 290200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2199
timestamp 1654712443
transform 1 0 293200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_2001
timestamp 1654712443
transform 1 0 -800 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2000
timestamp 1654712443
transform 1 0 -3800 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2002
timestamp 1654712443
transform 1 0 2200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2003
timestamp 1654712443
transform 1 0 5200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2004
timestamp 1654712443
transform 1 0 8200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2005
timestamp 1654712443
transform 1 0 11200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2006
timestamp 1654712443
transform 1 0 14200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2007
timestamp 1654712443
transform 1 0 17200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2008
timestamp 1654712443
transform 1 0 20200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2009
timestamp 1654712443
transform 1 0 23200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2011
timestamp 1654712443
transform 1 0 29200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2010
timestamp 1654712443
transform 1 0 26200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2012
timestamp 1654712443
transform 1 0 32200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2013
timestamp 1654712443
transform 1 0 35200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2014
timestamp 1654712443
transform 1 0 38200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2015
timestamp 1654712443
transform 1 0 41200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2016
timestamp 1654712443
transform 1 0 44200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2017
timestamp 1654712443
transform 1 0 47200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2018
timestamp 1654712443
transform 1 0 50200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2019
timestamp 1654712443
transform 1 0 53200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2021
timestamp 1654712443
transform 1 0 59200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2020
timestamp 1654712443
transform 1 0 56200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2022
timestamp 1654712443
transform 1 0 62200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2023
timestamp 1654712443
transform 1 0 65200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2024
timestamp 1654712443
transform 1 0 68200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2025
timestamp 1654712443
transform 1 0 71200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2026
timestamp 1654712443
transform 1 0 74200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2027
timestamp 1654712443
transform 1 0 77200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2028
timestamp 1654712443
transform 1 0 80200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2029
timestamp 1654712443
transform 1 0 83200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2030
timestamp 1654712443
transform 1 0 86200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2032
timestamp 1654712443
transform 1 0 92200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2031
timestamp 1654712443
transform 1 0 89200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2033
timestamp 1654712443
transform 1 0 95200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2034
timestamp 1654712443
transform 1 0 98200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2035
timestamp 1654712443
transform 1 0 101200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2036
timestamp 1654712443
transform 1 0 104200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2037
timestamp 1654712443
transform 1 0 107200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2038
timestamp 1654712443
transform 1 0 110200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2039
timestamp 1654712443
transform 1 0 113200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2040
timestamp 1654712443
transform 1 0 116200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2042
timestamp 1654712443
transform 1 0 122200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2041
timestamp 1654712443
transform 1 0 119200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2043
timestamp 1654712443
transform 1 0 125200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2044
timestamp 1654712443
transform 1 0 128200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2045
timestamp 1654712443
transform 1 0 131200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2046
timestamp 1654712443
transform 1 0 134200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2047
timestamp 1654712443
transform 1 0 137200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2048
timestamp 1654712443
transform 1 0 140200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2049
timestamp 1654712443
transform 1 0 143200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2050
timestamp 1654712443
transform 1 0 146200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2052
timestamp 1654712443
transform 1 0 152200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2051
timestamp 1654712443
transform 1 0 149200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2053
timestamp 1654712443
transform 1 0 155200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2054
timestamp 1654712443
transform 1 0 158200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2055
timestamp 1654712443
transform 1 0 161200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2056
timestamp 1654712443
transform 1 0 164200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2057
timestamp 1654712443
transform 1 0 167200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2058
timestamp 1654712443
transform 1 0 170200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2059
timestamp 1654712443
transform 1 0 173200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2060
timestamp 1654712443
transform 1 0 176200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2061
timestamp 1654712443
transform 1 0 179200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2063
timestamp 1654712443
transform 1 0 185200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2062
timestamp 1654712443
transform 1 0 182200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2064
timestamp 1654712443
transform 1 0 188200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2065
timestamp 1654712443
transform 1 0 191200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2066
timestamp 1654712443
transform 1 0 194200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2067
timestamp 1654712443
transform 1 0 197200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2068
timestamp 1654712443
transform 1 0 200200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2069
timestamp 1654712443
transform 1 0 203200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2070
timestamp 1654712443
transform 1 0 206200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2071
timestamp 1654712443
transform 1 0 209200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2073
timestamp 1654712443
transform 1 0 215200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2072
timestamp 1654712443
transform 1 0 212200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2074
timestamp 1654712443
transform 1 0 218200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2075
timestamp 1654712443
transform 1 0 221200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2076
timestamp 1654712443
transform 1 0 224200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2077
timestamp 1654712443
transform 1 0 227200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2078
timestamp 1654712443
transform 1 0 230200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2079
timestamp 1654712443
transform 1 0 233200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2080
timestamp 1654712443
transform 1 0 236200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2081
timestamp 1654712443
transform 1 0 239200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2083
timestamp 1654712443
transform 1 0 245200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2082
timestamp 1654712443
transform 1 0 242200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2084
timestamp 1654712443
transform 1 0 248200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2085
timestamp 1654712443
transform 1 0 251200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2086
timestamp 1654712443
transform 1 0 254200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2087
timestamp 1654712443
transform 1 0 257200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2088
timestamp 1654712443
transform 1 0 260200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2089
timestamp 1654712443
transform 1 0 263200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2090
timestamp 1654712443
transform 1 0 266200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2091
timestamp 1654712443
transform 1 0 269200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2092
timestamp 1654712443
transform 1 0 272200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2094
timestamp 1654712443
transform 1 0 278200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2093
timestamp 1654712443
transform 1 0 275200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2095
timestamp 1654712443
transform 1 0 281200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2096
timestamp 1654712443
transform 1 0 284200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2097
timestamp 1654712443
transform 1 0 287200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2098
timestamp 1654712443
transform 1 0 290200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_2099
timestamp 1654712443
transform 1 0 293200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_1901
timestamp 1654712443
transform 1 0 -800 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1900
timestamp 1654712443
transform 1 0 -3800 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1902
timestamp 1654712443
transform 1 0 2200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1903
timestamp 1654712443
transform 1 0 5200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1904
timestamp 1654712443
transform 1 0 8200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1905
timestamp 1654712443
transform 1 0 11200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1906
timestamp 1654712443
transform 1 0 14200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1907
timestamp 1654712443
transform 1 0 17200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1908
timestamp 1654712443
transform 1 0 20200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1909
timestamp 1654712443
transform 1 0 23200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1911
timestamp 1654712443
transform 1 0 29200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1910
timestamp 1654712443
transform 1 0 26200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1912
timestamp 1654712443
transform 1 0 32200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1913
timestamp 1654712443
transform 1 0 35200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1914
timestamp 1654712443
transform 1 0 38200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1915
timestamp 1654712443
transform 1 0 41200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1916
timestamp 1654712443
transform 1 0 44200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1917
timestamp 1654712443
transform 1 0 47200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1918
timestamp 1654712443
transform 1 0 50200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1919
timestamp 1654712443
transform 1 0 53200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1921
timestamp 1654712443
transform 1 0 59200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1920
timestamp 1654712443
transform 1 0 56200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1922
timestamp 1654712443
transform 1 0 62200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1923
timestamp 1654712443
transform 1 0 65200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1924
timestamp 1654712443
transform 1 0 68200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1925
timestamp 1654712443
transform 1 0 71200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1926
timestamp 1654712443
transform 1 0 74200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1927
timestamp 1654712443
transform 1 0 77200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1928
timestamp 1654712443
transform 1 0 80200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1929
timestamp 1654712443
transform 1 0 83200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1930
timestamp 1654712443
transform 1 0 86200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1932
timestamp 1654712443
transform 1 0 92200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1931
timestamp 1654712443
transform 1 0 89200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1933
timestamp 1654712443
transform 1 0 95200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1934
timestamp 1654712443
transform 1 0 98200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1935
timestamp 1654712443
transform 1 0 101200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1936
timestamp 1654712443
transform 1 0 104200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1937
timestamp 1654712443
transform 1 0 107200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1938
timestamp 1654712443
transform 1 0 110200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1939
timestamp 1654712443
transform 1 0 113200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1940
timestamp 1654712443
transform 1 0 116200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1942
timestamp 1654712443
transform 1 0 122200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1941
timestamp 1654712443
transform 1 0 119200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1943
timestamp 1654712443
transform 1 0 125200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1944
timestamp 1654712443
transform 1 0 128200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1945
timestamp 1654712443
transform 1 0 131200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1946
timestamp 1654712443
transform 1 0 134200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1947
timestamp 1654712443
transform 1 0 137200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1948
timestamp 1654712443
transform 1 0 140200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1949
timestamp 1654712443
transform 1 0 143200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1950
timestamp 1654712443
transform 1 0 146200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1952
timestamp 1654712443
transform 1 0 152200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1951
timestamp 1654712443
transform 1 0 149200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1953
timestamp 1654712443
transform 1 0 155200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1954
timestamp 1654712443
transform 1 0 158200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1955
timestamp 1654712443
transform 1 0 161200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1956
timestamp 1654712443
transform 1 0 164200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1957
timestamp 1654712443
transform 1 0 167200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1958
timestamp 1654712443
transform 1 0 170200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1959
timestamp 1654712443
transform 1 0 173200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1960
timestamp 1654712443
transform 1 0 176200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1961
timestamp 1654712443
transform 1 0 179200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1963
timestamp 1654712443
transform 1 0 185200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1962
timestamp 1654712443
transform 1 0 182200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1964
timestamp 1654712443
transform 1 0 188200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1965
timestamp 1654712443
transform 1 0 191200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1966
timestamp 1654712443
transform 1 0 194200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1967
timestamp 1654712443
transform 1 0 197200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1968
timestamp 1654712443
transform 1 0 200200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1969
timestamp 1654712443
transform 1 0 203200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1970
timestamp 1654712443
transform 1 0 206200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1971
timestamp 1654712443
transform 1 0 209200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1973
timestamp 1654712443
transform 1 0 215200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1972
timestamp 1654712443
transform 1 0 212200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1974
timestamp 1654712443
transform 1 0 218200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1975
timestamp 1654712443
transform 1 0 221200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1976
timestamp 1654712443
transform 1 0 224200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1977
timestamp 1654712443
transform 1 0 227200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1978
timestamp 1654712443
transform 1 0 230200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1979
timestamp 1654712443
transform 1 0 233200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1980
timestamp 1654712443
transform 1 0 236200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1981
timestamp 1654712443
transform 1 0 239200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1983
timestamp 1654712443
transform 1 0 245200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1982
timestamp 1654712443
transform 1 0 242200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1984
timestamp 1654712443
transform 1 0 248200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1985
timestamp 1654712443
transform 1 0 251200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1986
timestamp 1654712443
transform 1 0 254200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1987
timestamp 1654712443
transform 1 0 257200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1988
timestamp 1654712443
transform 1 0 260200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1989
timestamp 1654712443
transform 1 0 263200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1990
timestamp 1654712443
transform 1 0 266200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1991
timestamp 1654712443
transform 1 0 269200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1992
timestamp 1654712443
transform 1 0 272200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1994
timestamp 1654712443
transform 1 0 278200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1993
timestamp 1654712443
transform 1 0 275200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1995
timestamp 1654712443
transform 1 0 281200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1996
timestamp 1654712443
transform 1 0 284200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1997
timestamp 1654712443
transform 1 0 287200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1998
timestamp 1654712443
transform 1 0 290200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1999
timestamp 1654712443
transform 1 0 293200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1801
timestamp 1654712443
transform 1 0 -800 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1800
timestamp 1654712443
transform 1 0 -3800 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1802
timestamp 1654712443
transform 1 0 2200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1803
timestamp 1654712443
transform 1 0 5200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1804
timestamp 1654712443
transform 1 0 8200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1805
timestamp 1654712443
transform 1 0 11200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1806
timestamp 1654712443
transform 1 0 14200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1807
timestamp 1654712443
transform 1 0 17200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1808
timestamp 1654712443
transform 1 0 20200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1809
timestamp 1654712443
transform 1 0 23200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1811
timestamp 1654712443
transform 1 0 29200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1810
timestamp 1654712443
transform 1 0 26200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1812
timestamp 1654712443
transform 1 0 32200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1813
timestamp 1654712443
transform 1 0 35200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1814
timestamp 1654712443
transform 1 0 38200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1815
timestamp 1654712443
transform 1 0 41200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1816
timestamp 1654712443
transform 1 0 44200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1817
timestamp 1654712443
transform 1 0 47200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1818
timestamp 1654712443
transform 1 0 50200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1819
timestamp 1654712443
transform 1 0 53200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1821
timestamp 1654712443
transform 1 0 59200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1820
timestamp 1654712443
transform 1 0 56200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1822
timestamp 1654712443
transform 1 0 62200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1823
timestamp 1654712443
transform 1 0 65200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1824
timestamp 1654712443
transform 1 0 68200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1825
timestamp 1654712443
transform 1 0 71200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1826
timestamp 1654712443
transform 1 0 74200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1827
timestamp 1654712443
transform 1 0 77200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1828
timestamp 1654712443
transform 1 0 80200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1829
timestamp 1654712443
transform 1 0 83200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1830
timestamp 1654712443
transform 1 0 86200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1832
timestamp 1654712443
transform 1 0 92200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1831
timestamp 1654712443
transform 1 0 89200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1833
timestamp 1654712443
transform 1 0 95200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1834
timestamp 1654712443
transform 1 0 98200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1835
timestamp 1654712443
transform 1 0 101200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1836
timestamp 1654712443
transform 1 0 104200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1837
timestamp 1654712443
transform 1 0 107200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1838
timestamp 1654712443
transform 1 0 110200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1839
timestamp 1654712443
transform 1 0 113200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1840
timestamp 1654712443
transform 1 0 116200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1842
timestamp 1654712443
transform 1 0 122200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1841
timestamp 1654712443
transform 1 0 119200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1843
timestamp 1654712443
transform 1 0 125200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1844
timestamp 1654712443
transform 1 0 128200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1845
timestamp 1654712443
transform 1 0 131200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1846
timestamp 1654712443
transform 1 0 134200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1847
timestamp 1654712443
transform 1 0 137200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1848
timestamp 1654712443
transform 1 0 140200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1849
timestamp 1654712443
transform 1 0 143200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1850
timestamp 1654712443
transform 1 0 146200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1852
timestamp 1654712443
transform 1 0 152200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1851
timestamp 1654712443
transform 1 0 149200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1853
timestamp 1654712443
transform 1 0 155200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1854
timestamp 1654712443
transform 1 0 158200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1855
timestamp 1654712443
transform 1 0 161200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1856
timestamp 1654712443
transform 1 0 164200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1857
timestamp 1654712443
transform 1 0 167200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1858
timestamp 1654712443
transform 1 0 170200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1859
timestamp 1654712443
transform 1 0 173200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1860
timestamp 1654712443
transform 1 0 176200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1861
timestamp 1654712443
transform 1 0 179200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1863
timestamp 1654712443
transform 1 0 185200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1862
timestamp 1654712443
transform 1 0 182200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1864
timestamp 1654712443
transform 1 0 188200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1865
timestamp 1654712443
transform 1 0 191200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1866
timestamp 1654712443
transform 1 0 194200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1867
timestamp 1654712443
transform 1 0 197200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1868
timestamp 1654712443
transform 1 0 200200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1869
timestamp 1654712443
transform 1 0 203200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1870
timestamp 1654712443
transform 1 0 206200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1871
timestamp 1654712443
transform 1 0 209200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1873
timestamp 1654712443
transform 1 0 215200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1872
timestamp 1654712443
transform 1 0 212200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1874
timestamp 1654712443
transform 1 0 218200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1875
timestamp 1654712443
transform 1 0 221200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1876
timestamp 1654712443
transform 1 0 224200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1877
timestamp 1654712443
transform 1 0 227200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1878
timestamp 1654712443
transform 1 0 230200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1879
timestamp 1654712443
transform 1 0 233200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1880
timestamp 1654712443
transform 1 0 236200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1881
timestamp 1654712443
transform 1 0 239200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1883
timestamp 1654712443
transform 1 0 245200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1882
timestamp 1654712443
transform 1 0 242200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1884
timestamp 1654712443
transform 1 0 248200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1885
timestamp 1654712443
transform 1 0 251200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1886
timestamp 1654712443
transform 1 0 254200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1887
timestamp 1654712443
transform 1 0 257200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1888
timestamp 1654712443
transform 1 0 260200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1889
timestamp 1654712443
transform 1 0 263200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1890
timestamp 1654712443
transform 1 0 266200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1891
timestamp 1654712443
transform 1 0 269200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1892
timestamp 1654712443
transform 1 0 272200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1894
timestamp 1654712443
transform 1 0 278200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1893
timestamp 1654712443
transform 1 0 275200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1895
timestamp 1654712443
transform 1 0 281200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1896
timestamp 1654712443
transform 1 0 284200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1897
timestamp 1654712443
transform 1 0 287200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1898
timestamp 1654712443
transform 1 0 290200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1899
timestamp 1654712443
transform 1 0 293200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_1601
timestamp 1654712443
transform 1 0 -800 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1600
timestamp 1654712443
transform 1 0 -3800 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1701
timestamp 1654712443
transform 1 0 -800 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1700
timestamp 1654712443
transform 1 0 -3800 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1602
timestamp 1654712443
transform 1 0 2200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1702
timestamp 1654712443
transform 1 0 2200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1603
timestamp 1654712443
transform 1 0 5200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1703
timestamp 1654712443
transform 1 0 5200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1604
timestamp 1654712443
transform 1 0 8200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1704
timestamp 1654712443
transform 1 0 8200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1605
timestamp 1654712443
transform 1 0 11200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1705
timestamp 1654712443
transform 1 0 11200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1606
timestamp 1654712443
transform 1 0 14200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1706
timestamp 1654712443
transform 1 0 14200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1607
timestamp 1654712443
transform 1 0 17200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1707
timestamp 1654712443
transform 1 0 17200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1608
timestamp 1654712443
transform 1 0 20200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1708
timestamp 1654712443
transform 1 0 20200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1609
timestamp 1654712443
transform 1 0 23200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1709
timestamp 1654712443
transform 1 0 23200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1611
timestamp 1654712443
transform 1 0 29200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1610
timestamp 1654712443
transform 1 0 26200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1711
timestamp 1654712443
transform 1 0 29200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1710
timestamp 1654712443
transform 1 0 26200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1612
timestamp 1654712443
transform 1 0 32200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1712
timestamp 1654712443
transform 1 0 32200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1613
timestamp 1654712443
transform 1 0 35200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1713
timestamp 1654712443
transform 1 0 35200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1614
timestamp 1654712443
transform 1 0 38200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1714
timestamp 1654712443
transform 1 0 38200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1615
timestamp 1654712443
transform 1 0 41200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1715
timestamp 1654712443
transform 1 0 41200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1616
timestamp 1654712443
transform 1 0 44200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1716
timestamp 1654712443
transform 1 0 44200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1617
timestamp 1654712443
transform 1 0 47200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1717
timestamp 1654712443
transform 1 0 47200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1618
timestamp 1654712443
transform 1 0 50200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1718
timestamp 1654712443
transform 1 0 50200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1619
timestamp 1654712443
transform 1 0 53200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1719
timestamp 1654712443
transform 1 0 53200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1621
timestamp 1654712443
transform 1 0 59200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1620
timestamp 1654712443
transform 1 0 56200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1721
timestamp 1654712443
transform 1 0 59200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1720
timestamp 1654712443
transform 1 0 56200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1622
timestamp 1654712443
transform 1 0 62200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1722
timestamp 1654712443
transform 1 0 62200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1623
timestamp 1654712443
transform 1 0 65200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1723
timestamp 1654712443
transform 1 0 65200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1624
timestamp 1654712443
transform 1 0 68200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1724
timestamp 1654712443
transform 1 0 68200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1625
timestamp 1654712443
transform 1 0 71200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1725
timestamp 1654712443
transform 1 0 71200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1626
timestamp 1654712443
transform 1 0 74200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1726
timestamp 1654712443
transform 1 0 74200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1627
timestamp 1654712443
transform 1 0 77200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1727
timestamp 1654712443
transform 1 0 77200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1628
timestamp 1654712443
transform 1 0 80200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1728
timestamp 1654712443
transform 1 0 80200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1629
timestamp 1654712443
transform 1 0 83200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1729
timestamp 1654712443
transform 1 0 83200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1630
timestamp 1654712443
transform 1 0 86200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1730
timestamp 1654712443
transform 1 0 86200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1632
timestamp 1654712443
transform 1 0 92200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1631
timestamp 1654712443
transform 1 0 89200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1732
timestamp 1654712443
transform 1 0 92200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1731
timestamp 1654712443
transform 1 0 89200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1633
timestamp 1654712443
transform 1 0 95200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1733
timestamp 1654712443
transform 1 0 95200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1634
timestamp 1654712443
transform 1 0 98200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1734
timestamp 1654712443
transform 1 0 98200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1635
timestamp 1654712443
transform 1 0 101200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1735
timestamp 1654712443
transform 1 0 101200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1636
timestamp 1654712443
transform 1 0 104200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1736
timestamp 1654712443
transform 1 0 104200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1637
timestamp 1654712443
transform 1 0 107200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1737
timestamp 1654712443
transform 1 0 107200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1638
timestamp 1654712443
transform 1 0 110200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1738
timestamp 1654712443
transform 1 0 110200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1639
timestamp 1654712443
transform 1 0 113200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1739
timestamp 1654712443
transform 1 0 113200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1640
timestamp 1654712443
transform 1 0 116200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1740
timestamp 1654712443
transform 1 0 116200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1642
timestamp 1654712443
transform 1 0 122200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1641
timestamp 1654712443
transform 1 0 119200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1742
timestamp 1654712443
transform 1 0 122200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1741
timestamp 1654712443
transform 1 0 119200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1643
timestamp 1654712443
transform 1 0 125200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1743
timestamp 1654712443
transform 1 0 125200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1644
timestamp 1654712443
transform 1 0 128200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1744
timestamp 1654712443
transform 1 0 128200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1645
timestamp 1654712443
transform 1 0 131200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1745
timestamp 1654712443
transform 1 0 131200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1646
timestamp 1654712443
transform 1 0 134200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1746
timestamp 1654712443
transform 1 0 134200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1647
timestamp 1654712443
transform 1 0 137200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1747
timestamp 1654712443
transform 1 0 137200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1648
timestamp 1654712443
transform 1 0 140200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1748
timestamp 1654712443
transform 1 0 140200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1649
timestamp 1654712443
transform 1 0 143200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1749
timestamp 1654712443
transform 1 0 143200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1650
timestamp 1654712443
transform 1 0 146200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1750
timestamp 1654712443
transform 1 0 146200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1652
timestamp 1654712443
transform 1 0 152200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1651
timestamp 1654712443
transform 1 0 149200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1752
timestamp 1654712443
transform 1 0 152200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1751
timestamp 1654712443
transform 1 0 149200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1653
timestamp 1654712443
transform 1 0 155200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1753
timestamp 1654712443
transform 1 0 155200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1654
timestamp 1654712443
transform 1 0 158200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1754
timestamp 1654712443
transform 1 0 158200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1655
timestamp 1654712443
transform 1 0 161200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1755
timestamp 1654712443
transform 1 0 161200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1656
timestamp 1654712443
transform 1 0 164200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1756
timestamp 1654712443
transform 1 0 164200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1657
timestamp 1654712443
transform 1 0 167200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1757
timestamp 1654712443
transform 1 0 167200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1658
timestamp 1654712443
transform 1 0 170200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1758
timestamp 1654712443
transform 1 0 170200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1659
timestamp 1654712443
transform 1 0 173200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1759
timestamp 1654712443
transform 1 0 173200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1660
timestamp 1654712443
transform 1 0 176200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1760
timestamp 1654712443
transform 1 0 176200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1661
timestamp 1654712443
transform 1 0 179200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1761
timestamp 1654712443
transform 1 0 179200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1663
timestamp 1654712443
transform 1 0 185200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1662
timestamp 1654712443
transform 1 0 182200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1763
timestamp 1654712443
transform 1 0 185200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1762
timestamp 1654712443
transform 1 0 182200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1664
timestamp 1654712443
transform 1 0 188200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1764
timestamp 1654712443
transform 1 0 188200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1665
timestamp 1654712443
transform 1 0 191200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1765
timestamp 1654712443
transform 1 0 191200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1666
timestamp 1654712443
transform 1 0 194200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1766
timestamp 1654712443
transform 1 0 194200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1667
timestamp 1654712443
transform 1 0 197200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1767
timestamp 1654712443
transform 1 0 197200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1668
timestamp 1654712443
transform 1 0 200200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1768
timestamp 1654712443
transform 1 0 200200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1669
timestamp 1654712443
transform 1 0 203200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1769
timestamp 1654712443
transform 1 0 203200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1670
timestamp 1654712443
transform 1 0 206200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1770
timestamp 1654712443
transform 1 0 206200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1671
timestamp 1654712443
transform 1 0 209200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1771
timestamp 1654712443
transform 1 0 209200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1673
timestamp 1654712443
transform 1 0 215200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1672
timestamp 1654712443
transform 1 0 212200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1773
timestamp 1654712443
transform 1 0 215200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1772
timestamp 1654712443
transform 1 0 212200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1674
timestamp 1654712443
transform 1 0 218200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1774
timestamp 1654712443
transform 1 0 218200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1675
timestamp 1654712443
transform 1 0 221200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1775
timestamp 1654712443
transform 1 0 221200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1676
timestamp 1654712443
transform 1 0 224200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1776
timestamp 1654712443
transform 1 0 224200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1677
timestamp 1654712443
transform 1 0 227200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1777
timestamp 1654712443
transform 1 0 227200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1678
timestamp 1654712443
transform 1 0 230200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1778
timestamp 1654712443
transform 1 0 230200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1679
timestamp 1654712443
transform 1 0 233200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1779
timestamp 1654712443
transform 1 0 233200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1680
timestamp 1654712443
transform 1 0 236200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1780
timestamp 1654712443
transform 1 0 236200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1681
timestamp 1654712443
transform 1 0 239200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1781
timestamp 1654712443
transform 1 0 239200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1683
timestamp 1654712443
transform 1 0 245200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1682
timestamp 1654712443
transform 1 0 242200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1783
timestamp 1654712443
transform 1 0 245200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1782
timestamp 1654712443
transform 1 0 242200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1684
timestamp 1654712443
transform 1 0 248200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1784
timestamp 1654712443
transform 1 0 248200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1685
timestamp 1654712443
transform 1 0 251200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1785
timestamp 1654712443
transform 1 0 251200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1686
timestamp 1654712443
transform 1 0 254200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1786
timestamp 1654712443
transform 1 0 254200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1687
timestamp 1654712443
transform 1 0 257200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1787
timestamp 1654712443
transform 1 0 257200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1688
timestamp 1654712443
transform 1 0 260200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1788
timestamp 1654712443
transform 1 0 260200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1689
timestamp 1654712443
transform 1 0 263200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1789
timestamp 1654712443
transform 1 0 263200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1690
timestamp 1654712443
transform 1 0 266200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1790
timestamp 1654712443
transform 1 0 266200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1691
timestamp 1654712443
transform 1 0 269200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1791
timestamp 1654712443
transform 1 0 269200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1692
timestamp 1654712443
transform 1 0 272200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1792
timestamp 1654712443
transform 1 0 272200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1694
timestamp 1654712443
transform 1 0 278200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1693
timestamp 1654712443
transform 1 0 275200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1794
timestamp 1654712443
transform 1 0 278200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1793
timestamp 1654712443
transform 1 0 275200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1695
timestamp 1654712443
transform 1 0 281200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1795
timestamp 1654712443
transform 1 0 281200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1696
timestamp 1654712443
transform 1 0 284200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1796
timestamp 1654712443
transform 1 0 284200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1697
timestamp 1654712443
transform 1 0 287200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1797
timestamp 1654712443
transform 1 0 287200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1698
timestamp 1654712443
transform 1 0 290200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1798
timestamp 1654712443
transform 1 0 290200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1699
timestamp 1654712443
transform 1 0 293200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_1799
timestamp 1654712443
transform 1 0 293200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_1501
timestamp 1654712443
transform 1 0 -800 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1500
timestamp 1654712443
transform 1 0 -3800 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1502
timestamp 1654712443
transform 1 0 2200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1503
timestamp 1654712443
transform 1 0 5200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1504
timestamp 1654712443
transform 1 0 8200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1505
timestamp 1654712443
transform 1 0 11200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1506
timestamp 1654712443
transform 1 0 14200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1507
timestamp 1654712443
transform 1 0 17200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1508
timestamp 1654712443
transform 1 0 20200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1509
timestamp 1654712443
transform 1 0 23200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1511
timestamp 1654712443
transform 1 0 29200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1510
timestamp 1654712443
transform 1 0 26200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1512
timestamp 1654712443
transform 1 0 32200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1513
timestamp 1654712443
transform 1 0 35200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1514
timestamp 1654712443
transform 1 0 38200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1515
timestamp 1654712443
transform 1 0 41200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1516
timestamp 1654712443
transform 1 0 44200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1517
timestamp 1654712443
transform 1 0 47200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1518
timestamp 1654712443
transform 1 0 50200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1519
timestamp 1654712443
transform 1 0 53200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1521
timestamp 1654712443
transform 1 0 59200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1520
timestamp 1654712443
transform 1 0 56200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1522
timestamp 1654712443
transform 1 0 62200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1523
timestamp 1654712443
transform 1 0 65200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1524
timestamp 1654712443
transform 1 0 68200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1525
timestamp 1654712443
transform 1 0 71200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1526
timestamp 1654712443
transform 1 0 74200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1527
timestamp 1654712443
transform 1 0 77200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1528
timestamp 1654712443
transform 1 0 80200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1529
timestamp 1654712443
transform 1 0 83200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1530
timestamp 1654712443
transform 1 0 86200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1532
timestamp 1654712443
transform 1 0 92200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1531
timestamp 1654712443
transform 1 0 89200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1533
timestamp 1654712443
transform 1 0 95200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1534
timestamp 1654712443
transform 1 0 98200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1535
timestamp 1654712443
transform 1 0 101200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1536
timestamp 1654712443
transform 1 0 104200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1537
timestamp 1654712443
transform 1 0 107200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1538
timestamp 1654712443
transform 1 0 110200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1539
timestamp 1654712443
transform 1 0 113200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1540
timestamp 1654712443
transform 1 0 116200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1542
timestamp 1654712443
transform 1 0 122200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1541
timestamp 1654712443
transform 1 0 119200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1543
timestamp 1654712443
transform 1 0 125200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1544
timestamp 1654712443
transform 1 0 128200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1545
timestamp 1654712443
transform 1 0 131200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1546
timestamp 1654712443
transform 1 0 134200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1547
timestamp 1654712443
transform 1 0 137200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1548
timestamp 1654712443
transform 1 0 140200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1549
timestamp 1654712443
transform 1 0 143200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1550
timestamp 1654712443
transform 1 0 146200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1552
timestamp 1654712443
transform 1 0 152200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1551
timestamp 1654712443
transform 1 0 149200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1553
timestamp 1654712443
transform 1 0 155200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1554
timestamp 1654712443
transform 1 0 158200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1555
timestamp 1654712443
transform 1 0 161200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1556
timestamp 1654712443
transform 1 0 164200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1557
timestamp 1654712443
transform 1 0 167200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1558
timestamp 1654712443
transform 1 0 170200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1559
timestamp 1654712443
transform 1 0 173200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1560
timestamp 1654712443
transform 1 0 176200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1561
timestamp 1654712443
transform 1 0 179200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1563
timestamp 1654712443
transform 1 0 185200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1562
timestamp 1654712443
transform 1 0 182200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1564
timestamp 1654712443
transform 1 0 188200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1565
timestamp 1654712443
transform 1 0 191200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1566
timestamp 1654712443
transform 1 0 194200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1567
timestamp 1654712443
transform 1 0 197200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1568
timestamp 1654712443
transform 1 0 200200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1569
timestamp 1654712443
transform 1 0 203200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1570
timestamp 1654712443
transform 1 0 206200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1571
timestamp 1654712443
transform 1 0 209200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1573
timestamp 1654712443
transform 1 0 215200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1572
timestamp 1654712443
transform 1 0 212200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1574
timestamp 1654712443
transform 1 0 218200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1575
timestamp 1654712443
transform 1 0 221200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1576
timestamp 1654712443
transform 1 0 224200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1577
timestamp 1654712443
transform 1 0 227200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1578
timestamp 1654712443
transform 1 0 230200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1579
timestamp 1654712443
transform 1 0 233200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1580
timestamp 1654712443
transform 1 0 236200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1581
timestamp 1654712443
transform 1 0 239200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1583
timestamp 1654712443
transform 1 0 245200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1582
timestamp 1654712443
transform 1 0 242200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1584
timestamp 1654712443
transform 1 0 248200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1585
timestamp 1654712443
transform 1 0 251200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1586
timestamp 1654712443
transform 1 0 254200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1587
timestamp 1654712443
transform 1 0 257200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1588
timestamp 1654712443
transform 1 0 260200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1589
timestamp 1654712443
transform 1 0 263200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1590
timestamp 1654712443
transform 1 0 266200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1591
timestamp 1654712443
transform 1 0 269200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1592
timestamp 1654712443
transform 1 0 272200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1594
timestamp 1654712443
transform 1 0 278200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1593
timestamp 1654712443
transform 1 0 275200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1595
timestamp 1654712443
transform 1 0 281200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1596
timestamp 1654712443
transform 1 0 284200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1597
timestamp 1654712443
transform 1 0 287200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1598
timestamp 1654712443
transform 1 0 290200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1599
timestamp 1654712443
transform 1 0 293200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_1401
timestamp 1654712443
transform 1 0 -800 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1400
timestamp 1654712443
transform 1 0 -3800 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1402
timestamp 1654712443
transform 1 0 2200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1403
timestamp 1654712443
transform 1 0 5200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1404
timestamp 1654712443
transform 1 0 8200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1405
timestamp 1654712443
transform 1 0 11200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1406
timestamp 1654712443
transform 1 0 14200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1407
timestamp 1654712443
transform 1 0 17200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1408
timestamp 1654712443
transform 1 0 20200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1409
timestamp 1654712443
transform 1 0 23200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1411
timestamp 1654712443
transform 1 0 29200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1410
timestamp 1654712443
transform 1 0 26200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1412
timestamp 1654712443
transform 1 0 32200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1413
timestamp 1654712443
transform 1 0 35200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1414
timestamp 1654712443
transform 1 0 38200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1415
timestamp 1654712443
transform 1 0 41200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1416
timestamp 1654712443
transform 1 0 44200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1417
timestamp 1654712443
transform 1 0 47200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1418
timestamp 1654712443
transform 1 0 50200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1419
timestamp 1654712443
transform 1 0 53200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1421
timestamp 1654712443
transform 1 0 59200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1420
timestamp 1654712443
transform 1 0 56200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1422
timestamp 1654712443
transform 1 0 62200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1423
timestamp 1654712443
transform 1 0 65200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1424
timestamp 1654712443
transform 1 0 68200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1425
timestamp 1654712443
transform 1 0 71200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1426
timestamp 1654712443
transform 1 0 74200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1427
timestamp 1654712443
transform 1 0 77200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1428
timestamp 1654712443
transform 1 0 80200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1429
timestamp 1654712443
transform 1 0 83200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1430
timestamp 1654712443
transform 1 0 86200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1432
timestamp 1654712443
transform 1 0 92200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1431
timestamp 1654712443
transform 1 0 89200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1433
timestamp 1654712443
transform 1 0 95200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1434
timestamp 1654712443
transform 1 0 98200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1435
timestamp 1654712443
transform 1 0 101200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1436
timestamp 1654712443
transform 1 0 104200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1437
timestamp 1654712443
transform 1 0 107200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1438
timestamp 1654712443
transform 1 0 110200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1439
timestamp 1654712443
transform 1 0 113200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1440
timestamp 1654712443
transform 1 0 116200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1442
timestamp 1654712443
transform 1 0 122200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1441
timestamp 1654712443
transform 1 0 119200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1443
timestamp 1654712443
transform 1 0 125200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1444
timestamp 1654712443
transform 1 0 128200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1445
timestamp 1654712443
transform 1 0 131200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1446
timestamp 1654712443
transform 1 0 134200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1447
timestamp 1654712443
transform 1 0 137200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1448
timestamp 1654712443
transform 1 0 140200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1449
timestamp 1654712443
transform 1 0 143200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1450
timestamp 1654712443
transform 1 0 146200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1452
timestamp 1654712443
transform 1 0 152200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1451
timestamp 1654712443
transform 1 0 149200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1453
timestamp 1654712443
transform 1 0 155200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1454
timestamp 1654712443
transform 1 0 158200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1455
timestamp 1654712443
transform 1 0 161200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1456
timestamp 1654712443
transform 1 0 164200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1457
timestamp 1654712443
transform 1 0 167200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1458
timestamp 1654712443
transform 1 0 170200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1459
timestamp 1654712443
transform 1 0 173200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1460
timestamp 1654712443
transform 1 0 176200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1461
timestamp 1654712443
transform 1 0 179200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1463
timestamp 1654712443
transform 1 0 185200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1462
timestamp 1654712443
transform 1 0 182200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1464
timestamp 1654712443
transform 1 0 188200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1465
timestamp 1654712443
transform 1 0 191200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1466
timestamp 1654712443
transform 1 0 194200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1467
timestamp 1654712443
transform 1 0 197200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1468
timestamp 1654712443
transform 1 0 200200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1469
timestamp 1654712443
transform 1 0 203200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1470
timestamp 1654712443
transform 1 0 206200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1471
timestamp 1654712443
transform 1 0 209200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1473
timestamp 1654712443
transform 1 0 215200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1472
timestamp 1654712443
transform 1 0 212200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1474
timestamp 1654712443
transform 1 0 218200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1475
timestamp 1654712443
transform 1 0 221200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1476
timestamp 1654712443
transform 1 0 224200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1477
timestamp 1654712443
transform 1 0 227200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1478
timestamp 1654712443
transform 1 0 230200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1479
timestamp 1654712443
transform 1 0 233200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1480
timestamp 1654712443
transform 1 0 236200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1481
timestamp 1654712443
transform 1 0 239200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1483
timestamp 1654712443
transform 1 0 245200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1482
timestamp 1654712443
transform 1 0 242200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1484
timestamp 1654712443
transform 1 0 248200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1485
timestamp 1654712443
transform 1 0 251200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1486
timestamp 1654712443
transform 1 0 254200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1487
timestamp 1654712443
transform 1 0 257200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1488
timestamp 1654712443
transform 1 0 260200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1489
timestamp 1654712443
transform 1 0 263200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1490
timestamp 1654712443
transform 1 0 266200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1491
timestamp 1654712443
transform 1 0 269200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1492
timestamp 1654712443
transform 1 0 272200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1494
timestamp 1654712443
transform 1 0 278200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1493
timestamp 1654712443
transform 1 0 275200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1495
timestamp 1654712443
transform 1 0 281200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1496
timestamp 1654712443
transform 1 0 284200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1497
timestamp 1654712443
transform 1 0 287200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1498
timestamp 1654712443
transform 1 0 290200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1499
timestamp 1654712443
transform 1 0 293200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_1301
timestamp 1654712443
transform 1 0 -800 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1300
timestamp 1654712443
transform 1 0 -3800 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1302
timestamp 1654712443
transform 1 0 2200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1303
timestamp 1654712443
transform 1 0 5200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1304
timestamp 1654712443
transform 1 0 8200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1305
timestamp 1654712443
transform 1 0 11200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1306
timestamp 1654712443
transform 1 0 14200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1307
timestamp 1654712443
transform 1 0 17200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1308
timestamp 1654712443
transform 1 0 20200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1309
timestamp 1654712443
transform 1 0 23200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1311
timestamp 1654712443
transform 1 0 29200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1310
timestamp 1654712443
transform 1 0 26200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1312
timestamp 1654712443
transform 1 0 32200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1313
timestamp 1654712443
transform 1 0 35200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1314
timestamp 1654712443
transform 1 0 38200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1315
timestamp 1654712443
transform 1 0 41200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1316
timestamp 1654712443
transform 1 0 44200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1317
timestamp 1654712443
transform 1 0 47200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1318
timestamp 1654712443
transform 1 0 50200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1319
timestamp 1654712443
transform 1 0 53200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1321
timestamp 1654712443
transform 1 0 59200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1320
timestamp 1654712443
transform 1 0 56200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1322
timestamp 1654712443
transform 1 0 62200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1323
timestamp 1654712443
transform 1 0 65200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1324
timestamp 1654712443
transform 1 0 68200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1325
timestamp 1654712443
transform 1 0 71200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1326
timestamp 1654712443
transform 1 0 74200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1327
timestamp 1654712443
transform 1 0 77200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1328
timestamp 1654712443
transform 1 0 80200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1329
timestamp 1654712443
transform 1 0 83200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1330
timestamp 1654712443
transform 1 0 86200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1332
timestamp 1654712443
transform 1 0 92200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1331
timestamp 1654712443
transform 1 0 89200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1333
timestamp 1654712443
transform 1 0 95200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1334
timestamp 1654712443
transform 1 0 98200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1335
timestamp 1654712443
transform 1 0 101200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1336
timestamp 1654712443
transform 1 0 104200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1337
timestamp 1654712443
transform 1 0 107200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1338
timestamp 1654712443
transform 1 0 110200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1339
timestamp 1654712443
transform 1 0 113200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1340
timestamp 1654712443
transform 1 0 116200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1342
timestamp 1654712443
transform 1 0 122200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1341
timestamp 1654712443
transform 1 0 119200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1343
timestamp 1654712443
transform 1 0 125200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1344
timestamp 1654712443
transform 1 0 128200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1345
timestamp 1654712443
transform 1 0 131200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1346
timestamp 1654712443
transform 1 0 134200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1347
timestamp 1654712443
transform 1 0 137200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1348
timestamp 1654712443
transform 1 0 140200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1349
timestamp 1654712443
transform 1 0 143200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1350
timestamp 1654712443
transform 1 0 146200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1352
timestamp 1654712443
transform 1 0 152200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1351
timestamp 1654712443
transform 1 0 149200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1353
timestamp 1654712443
transform 1 0 155200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1354
timestamp 1654712443
transform 1 0 158200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1355
timestamp 1654712443
transform 1 0 161200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1356
timestamp 1654712443
transform 1 0 164200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1357
timestamp 1654712443
transform 1 0 167200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1358
timestamp 1654712443
transform 1 0 170200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1359
timestamp 1654712443
transform 1 0 173200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1360
timestamp 1654712443
transform 1 0 176200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1361
timestamp 1654712443
transform 1 0 179200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1363
timestamp 1654712443
transform 1 0 185200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1362
timestamp 1654712443
transform 1 0 182200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1364
timestamp 1654712443
transform 1 0 188200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1365
timestamp 1654712443
transform 1 0 191200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1366
timestamp 1654712443
transform 1 0 194200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1367
timestamp 1654712443
transform 1 0 197200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1368
timestamp 1654712443
transform 1 0 200200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1369
timestamp 1654712443
transform 1 0 203200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1370
timestamp 1654712443
transform 1 0 206200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1371
timestamp 1654712443
transform 1 0 209200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1373
timestamp 1654712443
transform 1 0 215200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1372
timestamp 1654712443
transform 1 0 212200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1374
timestamp 1654712443
transform 1 0 218200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1375
timestamp 1654712443
transform 1 0 221200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1376
timestamp 1654712443
transform 1 0 224200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1377
timestamp 1654712443
transform 1 0 227200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1378
timestamp 1654712443
transform 1 0 230200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1379
timestamp 1654712443
transform 1 0 233200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1380
timestamp 1654712443
transform 1 0 236200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1381
timestamp 1654712443
transform 1 0 239200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1383
timestamp 1654712443
transform 1 0 245200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1382
timestamp 1654712443
transform 1 0 242200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1384
timestamp 1654712443
transform 1 0 248200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1385
timestamp 1654712443
transform 1 0 251200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1386
timestamp 1654712443
transform 1 0 254200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1387
timestamp 1654712443
transform 1 0 257200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1388
timestamp 1654712443
transform 1 0 260200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1389
timestamp 1654712443
transform 1 0 263200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1390
timestamp 1654712443
transform 1 0 266200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1391
timestamp 1654712443
transform 1 0 269200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1392
timestamp 1654712443
transform 1 0 272200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1394
timestamp 1654712443
transform 1 0 278200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1393
timestamp 1654712443
transform 1 0 275200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1395
timestamp 1654712443
transform 1 0 281200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1396
timestamp 1654712443
transform 1 0 284200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1397
timestamp 1654712443
transform 1 0 287200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1398
timestamp 1654712443
transform 1 0 290200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1399
timestamp 1654712443
transform 1 0 293200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_1201
timestamp 1654712443
transform 1 0 -800 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1200
timestamp 1654712443
transform 1 0 -3800 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1202
timestamp 1654712443
transform 1 0 2200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1203
timestamp 1654712443
transform 1 0 5200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1204
timestamp 1654712443
transform 1 0 8200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1205
timestamp 1654712443
transform 1 0 11200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1206
timestamp 1654712443
transform 1 0 14200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1207
timestamp 1654712443
transform 1 0 17200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1208
timestamp 1654712443
transform 1 0 20200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1209
timestamp 1654712443
transform 1 0 23200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1211
timestamp 1654712443
transform 1 0 29200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1210
timestamp 1654712443
transform 1 0 26200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1212
timestamp 1654712443
transform 1 0 32200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1213
timestamp 1654712443
transform 1 0 35200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1214
timestamp 1654712443
transform 1 0 38200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1215
timestamp 1654712443
transform 1 0 41200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1216
timestamp 1654712443
transform 1 0 44200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1217
timestamp 1654712443
transform 1 0 47200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1218
timestamp 1654712443
transform 1 0 50200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1219
timestamp 1654712443
transform 1 0 53200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1221
timestamp 1654712443
transform 1 0 59200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1220
timestamp 1654712443
transform 1 0 56200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1222
timestamp 1654712443
transform 1 0 62200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1223
timestamp 1654712443
transform 1 0 65200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1224
timestamp 1654712443
transform 1 0 68200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1225
timestamp 1654712443
transform 1 0 71200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1226
timestamp 1654712443
transform 1 0 74200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1227
timestamp 1654712443
transform 1 0 77200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1228
timestamp 1654712443
transform 1 0 80200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1229
timestamp 1654712443
transform 1 0 83200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1230
timestamp 1654712443
transform 1 0 86200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1232
timestamp 1654712443
transform 1 0 92200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1231
timestamp 1654712443
transform 1 0 89200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1233
timestamp 1654712443
transform 1 0 95200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1234
timestamp 1654712443
transform 1 0 98200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1235
timestamp 1654712443
transform 1 0 101200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1236
timestamp 1654712443
transform 1 0 104200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1237
timestamp 1654712443
transform 1 0 107200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1238
timestamp 1654712443
transform 1 0 110200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1239
timestamp 1654712443
transform 1 0 113200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1240
timestamp 1654712443
transform 1 0 116200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1242
timestamp 1654712443
transform 1 0 122200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1241
timestamp 1654712443
transform 1 0 119200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1243
timestamp 1654712443
transform 1 0 125200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1244
timestamp 1654712443
transform 1 0 128200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1245
timestamp 1654712443
transform 1 0 131200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1246
timestamp 1654712443
transform 1 0 134200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1247
timestamp 1654712443
transform 1 0 137200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1248
timestamp 1654712443
transform 1 0 140200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1249
timestamp 1654712443
transform 1 0 143200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1250
timestamp 1654712443
transform 1 0 146200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1252
timestamp 1654712443
transform 1 0 152200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1251
timestamp 1654712443
transform 1 0 149200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1253
timestamp 1654712443
transform 1 0 155200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1254
timestamp 1654712443
transform 1 0 158200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1255
timestamp 1654712443
transform 1 0 161200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1256
timestamp 1654712443
transform 1 0 164200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1257
timestamp 1654712443
transform 1 0 167200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1258
timestamp 1654712443
transform 1 0 170200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1259
timestamp 1654712443
transform 1 0 173200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1260
timestamp 1654712443
transform 1 0 176200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1261
timestamp 1654712443
transform 1 0 179200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1263
timestamp 1654712443
transform 1 0 185200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1262
timestamp 1654712443
transform 1 0 182200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1264
timestamp 1654712443
transform 1 0 188200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1265
timestamp 1654712443
transform 1 0 191200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1266
timestamp 1654712443
transform 1 0 194200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1267
timestamp 1654712443
transform 1 0 197200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1268
timestamp 1654712443
transform 1 0 200200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1269
timestamp 1654712443
transform 1 0 203200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1270
timestamp 1654712443
transform 1 0 206200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1271
timestamp 1654712443
transform 1 0 209200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1273
timestamp 1654712443
transform 1 0 215200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1272
timestamp 1654712443
transform 1 0 212200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1274
timestamp 1654712443
transform 1 0 218200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1275
timestamp 1654712443
transform 1 0 221200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1276
timestamp 1654712443
transform 1 0 224200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1277
timestamp 1654712443
transform 1 0 227200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1278
timestamp 1654712443
transform 1 0 230200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1279
timestamp 1654712443
transform 1 0 233200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1280
timestamp 1654712443
transform 1 0 236200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1281
timestamp 1654712443
transform 1 0 239200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1283
timestamp 1654712443
transform 1 0 245200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1282
timestamp 1654712443
transform 1 0 242200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1284
timestamp 1654712443
transform 1 0 248200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1285
timestamp 1654712443
transform 1 0 251200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1286
timestamp 1654712443
transform 1 0 254200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1287
timestamp 1654712443
transform 1 0 257200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1288
timestamp 1654712443
transform 1 0 260200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1289
timestamp 1654712443
transform 1 0 263200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1290
timestamp 1654712443
transform 1 0 266200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1291
timestamp 1654712443
transform 1 0 269200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1292
timestamp 1654712443
transform 1 0 272200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1294
timestamp 1654712443
transform 1 0 278200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1293
timestamp 1654712443
transform 1 0 275200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1295
timestamp 1654712443
transform 1 0 281200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1296
timestamp 1654712443
transform 1 0 284200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1297
timestamp 1654712443
transform 1 0 287200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1298
timestamp 1654712443
transform 1 0 290200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1299
timestamp 1654712443
transform 1 0 293200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_1101
timestamp 1654712443
transform 1 0 -800 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1100
timestamp 1654712443
transform 1 0 -3800 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1102
timestamp 1654712443
transform 1 0 2200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1103
timestamp 1654712443
transform 1 0 5200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1104
timestamp 1654712443
transform 1 0 8200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1105
timestamp 1654712443
transform 1 0 11200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1106
timestamp 1654712443
transform 1 0 14200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1107
timestamp 1654712443
transform 1 0 17200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1108
timestamp 1654712443
transform 1 0 20200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1109
timestamp 1654712443
transform 1 0 23200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1111
timestamp 1654712443
transform 1 0 29200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1110
timestamp 1654712443
transform 1 0 26200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1112
timestamp 1654712443
transform 1 0 32200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1113
timestamp 1654712443
transform 1 0 35200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1114
timestamp 1654712443
transform 1 0 38200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1115
timestamp 1654712443
transform 1 0 41200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1116
timestamp 1654712443
transform 1 0 44200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1117
timestamp 1654712443
transform 1 0 47200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1118
timestamp 1654712443
transform 1 0 50200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1119
timestamp 1654712443
transform 1 0 53200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1121
timestamp 1654712443
transform 1 0 59200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1120
timestamp 1654712443
transform 1 0 56200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1122
timestamp 1654712443
transform 1 0 62200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1123
timestamp 1654712443
transform 1 0 65200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1124
timestamp 1654712443
transform 1 0 68200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1125
timestamp 1654712443
transform 1 0 71200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1126
timestamp 1654712443
transform 1 0 74200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1127
timestamp 1654712443
transform 1 0 77200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1128
timestamp 1654712443
transform 1 0 80200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1129
timestamp 1654712443
transform 1 0 83200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1130
timestamp 1654712443
transform 1 0 86200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1132
timestamp 1654712443
transform 1 0 92200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1131
timestamp 1654712443
transform 1 0 89200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1133
timestamp 1654712443
transform 1 0 95200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1134
timestamp 1654712443
transform 1 0 98200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1135
timestamp 1654712443
transform 1 0 101200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1136
timestamp 1654712443
transform 1 0 104200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1137
timestamp 1654712443
transform 1 0 107200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1138
timestamp 1654712443
transform 1 0 110200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1139
timestamp 1654712443
transform 1 0 113200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1140
timestamp 1654712443
transform 1 0 116200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1142
timestamp 1654712443
transform 1 0 122200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1141
timestamp 1654712443
transform 1 0 119200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1143
timestamp 1654712443
transform 1 0 125200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1144
timestamp 1654712443
transform 1 0 128200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1145
timestamp 1654712443
transform 1 0 131200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1146
timestamp 1654712443
transform 1 0 134200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1147
timestamp 1654712443
transform 1 0 137200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1148
timestamp 1654712443
transform 1 0 140200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1149
timestamp 1654712443
transform 1 0 143200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1150
timestamp 1654712443
transform 1 0 146200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1152
timestamp 1654712443
transform 1 0 152200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1151
timestamp 1654712443
transform 1 0 149200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1153
timestamp 1654712443
transform 1 0 155200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1154
timestamp 1654712443
transform 1 0 158200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1155
timestamp 1654712443
transform 1 0 161200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1156
timestamp 1654712443
transform 1 0 164200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1157
timestamp 1654712443
transform 1 0 167200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1158
timestamp 1654712443
transform 1 0 170200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1159
timestamp 1654712443
transform 1 0 173200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1160
timestamp 1654712443
transform 1 0 176200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1161
timestamp 1654712443
transform 1 0 179200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1163
timestamp 1654712443
transform 1 0 185200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1162
timestamp 1654712443
transform 1 0 182200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1164
timestamp 1654712443
transform 1 0 188200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1165
timestamp 1654712443
transform 1 0 191200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1166
timestamp 1654712443
transform 1 0 194200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1167
timestamp 1654712443
transform 1 0 197200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1168
timestamp 1654712443
transform 1 0 200200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1169
timestamp 1654712443
transform 1 0 203200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1170
timestamp 1654712443
transform 1 0 206200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1171
timestamp 1654712443
transform 1 0 209200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1173
timestamp 1654712443
transform 1 0 215200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1172
timestamp 1654712443
transform 1 0 212200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1174
timestamp 1654712443
transform 1 0 218200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1175
timestamp 1654712443
transform 1 0 221200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1176
timestamp 1654712443
transform 1 0 224200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1177
timestamp 1654712443
transform 1 0 227200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1178
timestamp 1654712443
transform 1 0 230200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1179
timestamp 1654712443
transform 1 0 233200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1180
timestamp 1654712443
transform 1 0 236200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1181
timestamp 1654712443
transform 1 0 239200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1183
timestamp 1654712443
transform 1 0 245200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1182
timestamp 1654712443
transform 1 0 242200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1184
timestamp 1654712443
transform 1 0 248200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1185
timestamp 1654712443
transform 1 0 251200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1186
timestamp 1654712443
transform 1 0 254200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1187
timestamp 1654712443
transform 1 0 257200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1188
timestamp 1654712443
transform 1 0 260200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1189
timestamp 1654712443
transform 1 0 263200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1190
timestamp 1654712443
transform 1 0 266200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1191
timestamp 1654712443
transform 1 0 269200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1192
timestamp 1654712443
transform 1 0 272200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1194
timestamp 1654712443
transform 1 0 278200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1193
timestamp 1654712443
transform 1 0 275200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1195
timestamp 1654712443
transform 1 0 281200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1196
timestamp 1654712443
transform 1 0 284200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1197
timestamp 1654712443
transform 1 0 287200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1198
timestamp 1654712443
transform 1 0 290200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1199
timestamp 1654712443
transform 1 0 293200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_1001
timestamp 1654712443
transform 1 0 -800 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1000
timestamp 1654712443
transform 1 0 -3800 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1002
timestamp 1654712443
transform 1 0 2200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1003
timestamp 1654712443
transform 1 0 5200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1004
timestamp 1654712443
transform 1 0 8200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1005
timestamp 1654712443
transform 1 0 11200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1006
timestamp 1654712443
transform 1 0 14200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1007
timestamp 1654712443
transform 1 0 17200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1008
timestamp 1654712443
transform 1 0 20200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1009
timestamp 1654712443
transform 1 0 23200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1011
timestamp 1654712443
transform 1 0 29200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1010
timestamp 1654712443
transform 1 0 26200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1012
timestamp 1654712443
transform 1 0 32200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1013
timestamp 1654712443
transform 1 0 35200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1014
timestamp 1654712443
transform 1 0 38200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1015
timestamp 1654712443
transform 1 0 41200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1016
timestamp 1654712443
transform 1 0 44200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1017
timestamp 1654712443
transform 1 0 47200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1018
timestamp 1654712443
transform 1 0 50200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1019
timestamp 1654712443
transform 1 0 53200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1021
timestamp 1654712443
transform 1 0 59200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1020
timestamp 1654712443
transform 1 0 56200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1022
timestamp 1654712443
transform 1 0 62200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1023
timestamp 1654712443
transform 1 0 65200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1024
timestamp 1654712443
transform 1 0 68200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1025
timestamp 1654712443
transform 1 0 71200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1026
timestamp 1654712443
transform 1 0 74200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1027
timestamp 1654712443
transform 1 0 77200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1028
timestamp 1654712443
transform 1 0 80200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1029
timestamp 1654712443
transform 1 0 83200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1030
timestamp 1654712443
transform 1 0 86200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1032
timestamp 1654712443
transform 1 0 92200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1031
timestamp 1654712443
transform 1 0 89200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1033
timestamp 1654712443
transform 1 0 95200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1034
timestamp 1654712443
transform 1 0 98200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1035
timestamp 1654712443
transform 1 0 101200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1036
timestamp 1654712443
transform 1 0 104200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1037
timestamp 1654712443
transform 1 0 107200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1038
timestamp 1654712443
transform 1 0 110200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1039
timestamp 1654712443
transform 1 0 113200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1040
timestamp 1654712443
transform 1 0 116200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1042
timestamp 1654712443
transform 1 0 122200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1041
timestamp 1654712443
transform 1 0 119200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1043
timestamp 1654712443
transform 1 0 125200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1044
timestamp 1654712443
transform 1 0 128200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1045
timestamp 1654712443
transform 1 0 131200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1046
timestamp 1654712443
transform 1 0 134200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1047
timestamp 1654712443
transform 1 0 137200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1048
timestamp 1654712443
transform 1 0 140200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1049
timestamp 1654712443
transform 1 0 143200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1050
timestamp 1654712443
transform 1 0 146200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1052
timestamp 1654712443
transform 1 0 152200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1051
timestamp 1654712443
transform 1 0 149200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1053
timestamp 1654712443
transform 1 0 155200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1054
timestamp 1654712443
transform 1 0 158200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1055
timestamp 1654712443
transform 1 0 161200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1056
timestamp 1654712443
transform 1 0 164200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1057
timestamp 1654712443
transform 1 0 167200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1058
timestamp 1654712443
transform 1 0 170200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1059
timestamp 1654712443
transform 1 0 173200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1060
timestamp 1654712443
transform 1 0 176200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1061
timestamp 1654712443
transform 1 0 179200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1063
timestamp 1654712443
transform 1 0 185200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1062
timestamp 1654712443
transform 1 0 182200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1064
timestamp 1654712443
transform 1 0 188200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1065
timestamp 1654712443
transform 1 0 191200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1066
timestamp 1654712443
transform 1 0 194200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1067
timestamp 1654712443
transform 1 0 197200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1068
timestamp 1654712443
transform 1 0 200200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1069
timestamp 1654712443
transform 1 0 203200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1070
timestamp 1654712443
transform 1 0 206200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1071
timestamp 1654712443
transform 1 0 209200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1073
timestamp 1654712443
transform 1 0 215200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1072
timestamp 1654712443
transform 1 0 212200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1074
timestamp 1654712443
transform 1 0 218200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1075
timestamp 1654712443
transform 1 0 221200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1076
timestamp 1654712443
transform 1 0 224200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1077
timestamp 1654712443
transform 1 0 227200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1078
timestamp 1654712443
transform 1 0 230200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1079
timestamp 1654712443
transform 1 0 233200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1080
timestamp 1654712443
transform 1 0 236200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1081
timestamp 1654712443
transform 1 0 239200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1083
timestamp 1654712443
transform 1 0 245200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1082
timestamp 1654712443
transform 1 0 242200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1084
timestamp 1654712443
transform 1 0 248200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1085
timestamp 1654712443
transform 1 0 251200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1086
timestamp 1654712443
transform 1 0 254200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1087
timestamp 1654712443
transform 1 0 257200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1088
timestamp 1654712443
transform 1 0 260200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1089
timestamp 1654712443
transform 1 0 263200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1090
timestamp 1654712443
transform 1 0 266200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1091
timestamp 1654712443
transform 1 0 269200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1092
timestamp 1654712443
transform 1 0 272200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1094
timestamp 1654712443
transform 1 0 278200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1093
timestamp 1654712443
transform 1 0 275200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1095
timestamp 1654712443
transform 1 0 281200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1096
timestamp 1654712443
transform 1 0 284200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1097
timestamp 1654712443
transform 1 0 287200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1098
timestamp 1654712443
transform 1 0 290200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_1099
timestamp 1654712443
transform 1 0 293200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_901
timestamp 1654712443
transform 1 0 -800 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_900
timestamp 1654712443
transform 1 0 -3800 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_902
timestamp 1654712443
transform 1 0 2200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_903
timestamp 1654712443
transform 1 0 5200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_904
timestamp 1654712443
transform 1 0 8200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_905
timestamp 1654712443
transform 1 0 11200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_906
timestamp 1654712443
transform 1 0 14200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_907
timestamp 1654712443
transform 1 0 17200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_908
timestamp 1654712443
transform 1 0 20200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_909
timestamp 1654712443
transform 1 0 23200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_911
timestamp 1654712443
transform 1 0 29200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_910
timestamp 1654712443
transform 1 0 26200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_912
timestamp 1654712443
transform 1 0 32200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_913
timestamp 1654712443
transform 1 0 35200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_914
timestamp 1654712443
transform 1 0 38200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_915
timestamp 1654712443
transform 1 0 41200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_916
timestamp 1654712443
transform 1 0 44200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_917
timestamp 1654712443
transform 1 0 47200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_918
timestamp 1654712443
transform 1 0 50200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_919
timestamp 1654712443
transform 1 0 53200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_921
timestamp 1654712443
transform 1 0 59200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_920
timestamp 1654712443
transform 1 0 56200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_922
timestamp 1654712443
transform 1 0 62200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_923
timestamp 1654712443
transform 1 0 65200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_924
timestamp 1654712443
transform 1 0 68200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_925
timestamp 1654712443
transform 1 0 71200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_926
timestamp 1654712443
transform 1 0 74200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_927
timestamp 1654712443
transform 1 0 77200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_928
timestamp 1654712443
transform 1 0 80200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_929
timestamp 1654712443
transform 1 0 83200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_930
timestamp 1654712443
transform 1 0 86200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_932
timestamp 1654712443
transform 1 0 92200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_931
timestamp 1654712443
transform 1 0 89200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_933
timestamp 1654712443
transform 1 0 95200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_934
timestamp 1654712443
transform 1 0 98200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_935
timestamp 1654712443
transform 1 0 101200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_936
timestamp 1654712443
transform 1 0 104200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_937
timestamp 1654712443
transform 1 0 107200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_938
timestamp 1654712443
transform 1 0 110200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_939
timestamp 1654712443
transform 1 0 113200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_940
timestamp 1654712443
transform 1 0 116200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_942
timestamp 1654712443
transform 1 0 122200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_941
timestamp 1654712443
transform 1 0 119200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_943
timestamp 1654712443
transform 1 0 125200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_944
timestamp 1654712443
transform 1 0 128200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_945
timestamp 1654712443
transform 1 0 131200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_946
timestamp 1654712443
transform 1 0 134200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_947
timestamp 1654712443
transform 1 0 137200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_948
timestamp 1654712443
transform 1 0 140200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_949
timestamp 1654712443
transform 1 0 143200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_950
timestamp 1654712443
transform 1 0 146200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_952
timestamp 1654712443
transform 1 0 152200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_951
timestamp 1654712443
transform 1 0 149200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_953
timestamp 1654712443
transform 1 0 155200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_954
timestamp 1654712443
transform 1 0 158200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_955
timestamp 1654712443
transform 1 0 161200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_956
timestamp 1654712443
transform 1 0 164200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_957
timestamp 1654712443
transform 1 0 167200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_958
timestamp 1654712443
transform 1 0 170200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_959
timestamp 1654712443
transform 1 0 173200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_960
timestamp 1654712443
transform 1 0 176200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_961
timestamp 1654712443
transform 1 0 179200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_963
timestamp 1654712443
transform 1 0 185200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_962
timestamp 1654712443
transform 1 0 182200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_964
timestamp 1654712443
transform 1 0 188200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_965
timestamp 1654712443
transform 1 0 191200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_966
timestamp 1654712443
transform 1 0 194200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_967
timestamp 1654712443
transform 1 0 197200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_968
timestamp 1654712443
transform 1 0 200200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_969
timestamp 1654712443
transform 1 0 203200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_970
timestamp 1654712443
transform 1 0 206200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_971
timestamp 1654712443
transform 1 0 209200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_973
timestamp 1654712443
transform 1 0 215200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_972
timestamp 1654712443
transform 1 0 212200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_974
timestamp 1654712443
transform 1 0 218200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_975
timestamp 1654712443
transform 1 0 221200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_976
timestamp 1654712443
transform 1 0 224200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_977
timestamp 1654712443
transform 1 0 227200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_978
timestamp 1654712443
transform 1 0 230200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_979
timestamp 1654712443
transform 1 0 233200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_980
timestamp 1654712443
transform 1 0 236200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_981
timestamp 1654712443
transform 1 0 239200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_983
timestamp 1654712443
transform 1 0 245200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_982
timestamp 1654712443
transform 1 0 242200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_984
timestamp 1654712443
transform 1 0 248200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_985
timestamp 1654712443
transform 1 0 251200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_986
timestamp 1654712443
transform 1 0 254200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_987
timestamp 1654712443
transform 1 0 257200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_988
timestamp 1654712443
transform 1 0 260200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_989
timestamp 1654712443
transform 1 0 263200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_990
timestamp 1654712443
transform 1 0 266200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_991
timestamp 1654712443
transform 1 0 269200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_992
timestamp 1654712443
transform 1 0 272200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_994
timestamp 1654712443
transform 1 0 278200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_993
timestamp 1654712443
transform 1 0 275200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_995
timestamp 1654712443
transform 1 0 281200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_996
timestamp 1654712443
transform 1 0 284200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_997
timestamp 1654712443
transform 1 0 287200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_998
timestamp 1654712443
transform 1 0 290200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_999
timestamp 1654712443
transform 1 0 293200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_801
timestamp 1654712443
transform 1 0 -800 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_800
timestamp 1654712443
transform 1 0 -3800 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_802
timestamp 1654712443
transform 1 0 2200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_803
timestamp 1654712443
transform 1 0 5200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_804
timestamp 1654712443
transform 1 0 8200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_805
timestamp 1654712443
transform 1 0 11200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_806
timestamp 1654712443
transform 1 0 14200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_807
timestamp 1654712443
transform 1 0 17200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_808
timestamp 1654712443
transform 1 0 20200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_809
timestamp 1654712443
transform 1 0 23200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_811
timestamp 1654712443
transform 1 0 29200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_810
timestamp 1654712443
transform 1 0 26200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_812
timestamp 1654712443
transform 1 0 32200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_813
timestamp 1654712443
transform 1 0 35200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_814
timestamp 1654712443
transform 1 0 38200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_815
timestamp 1654712443
transform 1 0 41200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_816
timestamp 1654712443
transform 1 0 44200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_817
timestamp 1654712443
transform 1 0 47200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_818
timestamp 1654712443
transform 1 0 50200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_819
timestamp 1654712443
transform 1 0 53200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_821
timestamp 1654712443
transform 1 0 59200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_820
timestamp 1654712443
transform 1 0 56200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_822
timestamp 1654712443
transform 1 0 62200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_823
timestamp 1654712443
transform 1 0 65200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_824
timestamp 1654712443
transform 1 0 68200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_825
timestamp 1654712443
transform 1 0 71200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_826
timestamp 1654712443
transform 1 0 74200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_827
timestamp 1654712443
transform 1 0 77200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_828
timestamp 1654712443
transform 1 0 80200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_829
timestamp 1654712443
transform 1 0 83200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_830
timestamp 1654712443
transform 1 0 86200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_832
timestamp 1654712443
transform 1 0 92200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_831
timestamp 1654712443
transform 1 0 89200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_833
timestamp 1654712443
transform 1 0 95200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_834
timestamp 1654712443
transform 1 0 98200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_835
timestamp 1654712443
transform 1 0 101200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_836
timestamp 1654712443
transform 1 0 104200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_837
timestamp 1654712443
transform 1 0 107200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_838
timestamp 1654712443
transform 1 0 110200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_839
timestamp 1654712443
transform 1 0 113200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_840
timestamp 1654712443
transform 1 0 116200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_842
timestamp 1654712443
transform 1 0 122200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_841
timestamp 1654712443
transform 1 0 119200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_843
timestamp 1654712443
transform 1 0 125200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_844
timestamp 1654712443
transform 1 0 128200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_845
timestamp 1654712443
transform 1 0 131200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_846
timestamp 1654712443
transform 1 0 134200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_847
timestamp 1654712443
transform 1 0 137200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_848
timestamp 1654712443
transform 1 0 140200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_849
timestamp 1654712443
transform 1 0 143200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_850
timestamp 1654712443
transform 1 0 146200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_852
timestamp 1654712443
transform 1 0 152200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_851
timestamp 1654712443
transform 1 0 149200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_853
timestamp 1654712443
transform 1 0 155200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_854
timestamp 1654712443
transform 1 0 158200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_855
timestamp 1654712443
transform 1 0 161200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_856
timestamp 1654712443
transform 1 0 164200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_857
timestamp 1654712443
transform 1 0 167200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_858
timestamp 1654712443
transform 1 0 170200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_859
timestamp 1654712443
transform 1 0 173200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_860
timestamp 1654712443
transform 1 0 176200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_861
timestamp 1654712443
transform 1 0 179200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_863
timestamp 1654712443
transform 1 0 185200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_862
timestamp 1654712443
transform 1 0 182200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_864
timestamp 1654712443
transform 1 0 188200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_865
timestamp 1654712443
transform 1 0 191200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_866
timestamp 1654712443
transform 1 0 194200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_867
timestamp 1654712443
transform 1 0 197200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_868
timestamp 1654712443
transform 1 0 200200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_869
timestamp 1654712443
transform 1 0 203200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_870
timestamp 1654712443
transform 1 0 206200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_871
timestamp 1654712443
transform 1 0 209200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_873
timestamp 1654712443
transform 1 0 215200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_872
timestamp 1654712443
transform 1 0 212200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_874
timestamp 1654712443
transform 1 0 218200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_875
timestamp 1654712443
transform 1 0 221200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_876
timestamp 1654712443
transform 1 0 224200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_877
timestamp 1654712443
transform 1 0 227200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_878
timestamp 1654712443
transform 1 0 230200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_879
timestamp 1654712443
transform 1 0 233200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_880
timestamp 1654712443
transform 1 0 236200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_881
timestamp 1654712443
transform 1 0 239200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_883
timestamp 1654712443
transform 1 0 245200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_882
timestamp 1654712443
transform 1 0 242200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_884
timestamp 1654712443
transform 1 0 248200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_885
timestamp 1654712443
transform 1 0 251200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_886
timestamp 1654712443
transform 1 0 254200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_887
timestamp 1654712443
transform 1 0 257200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_888
timestamp 1654712443
transform 1 0 260200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_889
timestamp 1654712443
transform 1 0 263200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_890
timestamp 1654712443
transform 1 0 266200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_891
timestamp 1654712443
transform 1 0 269200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_892
timestamp 1654712443
transform 1 0 272200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_894
timestamp 1654712443
transform 1 0 278200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_893
timestamp 1654712443
transform 1 0 275200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_895
timestamp 1654712443
transform 1 0 281200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_896
timestamp 1654712443
transform 1 0 284200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_897
timestamp 1654712443
transform 1 0 287200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_898
timestamp 1654712443
transform 1 0 290200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_899
timestamp 1654712443
transform 1 0 293200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_701
timestamp 1654712443
transform 1 0 -800 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_700
timestamp 1654712443
transform 1 0 -3800 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_702
timestamp 1654712443
transform 1 0 2200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_703
timestamp 1654712443
transform 1 0 5200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_704
timestamp 1654712443
transform 1 0 8200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_705
timestamp 1654712443
transform 1 0 11200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_706
timestamp 1654712443
transform 1 0 14200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_707
timestamp 1654712443
transform 1 0 17200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_708
timestamp 1654712443
transform 1 0 20200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_709
timestamp 1654712443
transform 1 0 23200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_711
timestamp 1654712443
transform 1 0 29200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_710
timestamp 1654712443
transform 1 0 26200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_712
timestamp 1654712443
transform 1 0 32200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_713
timestamp 1654712443
transform 1 0 35200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_714
timestamp 1654712443
transform 1 0 38200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_715
timestamp 1654712443
transform 1 0 41200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_716
timestamp 1654712443
transform 1 0 44200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_717
timestamp 1654712443
transform 1 0 47200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_718
timestamp 1654712443
transform 1 0 50200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_719
timestamp 1654712443
transform 1 0 53200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_721
timestamp 1654712443
transform 1 0 59200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_720
timestamp 1654712443
transform 1 0 56200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_722
timestamp 1654712443
transform 1 0 62200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_723
timestamp 1654712443
transform 1 0 65200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_724
timestamp 1654712443
transform 1 0 68200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_725
timestamp 1654712443
transform 1 0 71200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_726
timestamp 1654712443
transform 1 0 74200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_727
timestamp 1654712443
transform 1 0 77200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_728
timestamp 1654712443
transform 1 0 80200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_729
timestamp 1654712443
transform 1 0 83200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_730
timestamp 1654712443
transform 1 0 86200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_732
timestamp 1654712443
transform 1 0 92200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_731
timestamp 1654712443
transform 1 0 89200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_733
timestamp 1654712443
transform 1 0 95200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_734
timestamp 1654712443
transform 1 0 98200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_735
timestamp 1654712443
transform 1 0 101200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_736
timestamp 1654712443
transform 1 0 104200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_737
timestamp 1654712443
transform 1 0 107200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_738
timestamp 1654712443
transform 1 0 110200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_739
timestamp 1654712443
transform 1 0 113200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_740
timestamp 1654712443
transform 1 0 116200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_742
timestamp 1654712443
transform 1 0 122200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_741
timestamp 1654712443
transform 1 0 119200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_743
timestamp 1654712443
transform 1 0 125200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_744
timestamp 1654712443
transform 1 0 128200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_745
timestamp 1654712443
transform 1 0 131200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_746
timestamp 1654712443
transform 1 0 134200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_747
timestamp 1654712443
transform 1 0 137200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_748
timestamp 1654712443
transform 1 0 140200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_749
timestamp 1654712443
transform 1 0 143200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_750
timestamp 1654712443
transform 1 0 146200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_752
timestamp 1654712443
transform 1 0 152200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_751
timestamp 1654712443
transform 1 0 149200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_753
timestamp 1654712443
transform 1 0 155200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_754
timestamp 1654712443
transform 1 0 158200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_755
timestamp 1654712443
transform 1 0 161200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_756
timestamp 1654712443
transform 1 0 164200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_757
timestamp 1654712443
transform 1 0 167200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_758
timestamp 1654712443
transform 1 0 170200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_759
timestamp 1654712443
transform 1 0 173200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_760
timestamp 1654712443
transform 1 0 176200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_761
timestamp 1654712443
transform 1 0 179200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_763
timestamp 1654712443
transform 1 0 185200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_762
timestamp 1654712443
transform 1 0 182200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_764
timestamp 1654712443
transform 1 0 188200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_765
timestamp 1654712443
transform 1 0 191200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_766
timestamp 1654712443
transform 1 0 194200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_767
timestamp 1654712443
transform 1 0 197200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_768
timestamp 1654712443
transform 1 0 200200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_769
timestamp 1654712443
transform 1 0 203200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_770
timestamp 1654712443
transform 1 0 206200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_771
timestamp 1654712443
transform 1 0 209200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_773
timestamp 1654712443
transform 1 0 215200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_772
timestamp 1654712443
transform 1 0 212200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_774
timestamp 1654712443
transform 1 0 218200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_775
timestamp 1654712443
transform 1 0 221200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_776
timestamp 1654712443
transform 1 0 224200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_777
timestamp 1654712443
transform 1 0 227200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_778
timestamp 1654712443
transform 1 0 230200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_779
timestamp 1654712443
transform 1 0 233200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_780
timestamp 1654712443
transform 1 0 236200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_781
timestamp 1654712443
transform 1 0 239200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_783
timestamp 1654712443
transform 1 0 245200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_782
timestamp 1654712443
transform 1 0 242200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_784
timestamp 1654712443
transform 1 0 248200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_785
timestamp 1654712443
transform 1 0 251200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_786
timestamp 1654712443
transform 1 0 254200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_787
timestamp 1654712443
transform 1 0 257200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_788
timestamp 1654712443
transform 1 0 260200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_789
timestamp 1654712443
transform 1 0 263200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_790
timestamp 1654712443
transform 1 0 266200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_791
timestamp 1654712443
transform 1 0 269200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_792
timestamp 1654712443
transform 1 0 272200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_794
timestamp 1654712443
transform 1 0 278200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_793
timestamp 1654712443
transform 1 0 275200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_795
timestamp 1654712443
transform 1 0 281200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_796
timestamp 1654712443
transform 1 0 284200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_797
timestamp 1654712443
transform 1 0 287200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_798
timestamp 1654712443
transform 1 0 290200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_799
timestamp 1654712443
transform 1 0 293200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_501
timestamp 1654712443
transform 1 0 -800 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_601
timestamp 1654712443
transform 1 0 -800 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_500
timestamp 1654712443
transform 1 0 -3800 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_600
timestamp 1654712443
transform 1 0 -3800 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_502
timestamp 1654712443
transform 1 0 2200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_602
timestamp 1654712443
transform 1 0 2200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_503
timestamp 1654712443
transform 1 0 5200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_603
timestamp 1654712443
transform 1 0 5200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_504
timestamp 1654712443
transform 1 0 8200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_604
timestamp 1654712443
transform 1 0 8200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_505
timestamp 1654712443
transform 1 0 11200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_605
timestamp 1654712443
transform 1 0 11200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_506
timestamp 1654712443
transform 1 0 14200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_606
timestamp 1654712443
transform 1 0 14200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_507
timestamp 1654712443
transform 1 0 17200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_607
timestamp 1654712443
transform 1 0 17200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_508
timestamp 1654712443
transform 1 0 20200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_608
timestamp 1654712443
transform 1 0 20200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_509
timestamp 1654712443
transform 1 0 23200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_609
timestamp 1654712443
transform 1 0 23200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_511
timestamp 1654712443
transform 1 0 29200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_611
timestamp 1654712443
transform 1 0 29200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_510
timestamp 1654712443
transform 1 0 26200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_610
timestamp 1654712443
transform 1 0 26200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_512
timestamp 1654712443
transform 1 0 32200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_612
timestamp 1654712443
transform 1 0 32200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_513
timestamp 1654712443
transform 1 0 35200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_613
timestamp 1654712443
transform 1 0 35200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_514
timestamp 1654712443
transform 1 0 38200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_614
timestamp 1654712443
transform 1 0 38200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_515
timestamp 1654712443
transform 1 0 41200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_615
timestamp 1654712443
transform 1 0 41200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_516
timestamp 1654712443
transform 1 0 44200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_616
timestamp 1654712443
transform 1 0 44200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_517
timestamp 1654712443
transform 1 0 47200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_617
timestamp 1654712443
transform 1 0 47200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_518
timestamp 1654712443
transform 1 0 50200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_618
timestamp 1654712443
transform 1 0 50200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_519
timestamp 1654712443
transform 1 0 53200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_619
timestamp 1654712443
transform 1 0 53200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_521
timestamp 1654712443
transform 1 0 59200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_621
timestamp 1654712443
transform 1 0 59200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_520
timestamp 1654712443
transform 1 0 56200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_620
timestamp 1654712443
transform 1 0 56200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_522
timestamp 1654712443
transform 1 0 62200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_622
timestamp 1654712443
transform 1 0 62200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_523
timestamp 1654712443
transform 1 0 65200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_623
timestamp 1654712443
transform 1 0 65200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_524
timestamp 1654712443
transform 1 0 68200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_624
timestamp 1654712443
transform 1 0 68200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_525
timestamp 1654712443
transform 1 0 71200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_625
timestamp 1654712443
transform 1 0 71200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_526
timestamp 1654712443
transform 1 0 74200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_626
timestamp 1654712443
transform 1 0 74200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_527
timestamp 1654712443
transform 1 0 77200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_627
timestamp 1654712443
transform 1 0 77200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_528
timestamp 1654712443
transform 1 0 80200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_628
timestamp 1654712443
transform 1 0 80200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_529
timestamp 1654712443
transform 1 0 83200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_629
timestamp 1654712443
transform 1 0 83200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_530
timestamp 1654712443
transform 1 0 86200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_630
timestamp 1654712443
transform 1 0 86200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_532
timestamp 1654712443
transform 1 0 92200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_531
timestamp 1654712443
transform 1 0 89200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_632
timestamp 1654712443
transform 1 0 92200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_631
timestamp 1654712443
transform 1 0 89200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_533
timestamp 1654712443
transform 1 0 95200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_633
timestamp 1654712443
transform 1 0 95200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_534
timestamp 1654712443
transform 1 0 98200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_634
timestamp 1654712443
transform 1 0 98200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_535
timestamp 1654712443
transform 1 0 101200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_635
timestamp 1654712443
transform 1 0 101200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_536
timestamp 1654712443
transform 1 0 104200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_636
timestamp 1654712443
transform 1 0 104200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_537
timestamp 1654712443
transform 1 0 107200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_637
timestamp 1654712443
transform 1 0 107200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_538
timestamp 1654712443
transform 1 0 110200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_638
timestamp 1654712443
transform 1 0 110200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_539
timestamp 1654712443
transform 1 0 113200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_639
timestamp 1654712443
transform 1 0 113200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_540
timestamp 1654712443
transform 1 0 116200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_640
timestamp 1654712443
transform 1 0 116200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_542
timestamp 1654712443
transform 1 0 122200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_541
timestamp 1654712443
transform 1 0 119200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_642
timestamp 1654712443
transform 1 0 122200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_641
timestamp 1654712443
transform 1 0 119200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_543
timestamp 1654712443
transform 1 0 125200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_643
timestamp 1654712443
transform 1 0 125200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_544
timestamp 1654712443
transform 1 0 128200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_644
timestamp 1654712443
transform 1 0 128200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_545
timestamp 1654712443
transform 1 0 131200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_645
timestamp 1654712443
transform 1 0 131200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_546
timestamp 1654712443
transform 1 0 134200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_646
timestamp 1654712443
transform 1 0 134200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_547
timestamp 1654712443
transform 1 0 137200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_647
timestamp 1654712443
transform 1 0 137200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_548
timestamp 1654712443
transform 1 0 140200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_648
timestamp 1654712443
transform 1 0 140200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_549
timestamp 1654712443
transform 1 0 143200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_649
timestamp 1654712443
transform 1 0 143200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_550
timestamp 1654712443
transform 1 0 146200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_650
timestamp 1654712443
transform 1 0 146200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_552
timestamp 1654712443
transform 1 0 152200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_551
timestamp 1654712443
transform 1 0 149200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_652
timestamp 1654712443
transform 1 0 152200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_651
timestamp 1654712443
transform 1 0 149200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_553
timestamp 1654712443
transform 1 0 155200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_653
timestamp 1654712443
transform 1 0 155200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_554
timestamp 1654712443
transform 1 0 158200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_654
timestamp 1654712443
transform 1 0 158200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_555
timestamp 1654712443
transform 1 0 161200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_655
timestamp 1654712443
transform 1 0 161200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_556
timestamp 1654712443
transform 1 0 164200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_656
timestamp 1654712443
transform 1 0 164200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_557
timestamp 1654712443
transform 1 0 167200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_657
timestamp 1654712443
transform 1 0 167200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_558
timestamp 1654712443
transform 1 0 170200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_658
timestamp 1654712443
transform 1 0 170200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_559
timestamp 1654712443
transform 1 0 173200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_659
timestamp 1654712443
transform 1 0 173200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_560
timestamp 1654712443
transform 1 0 176200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_660
timestamp 1654712443
transform 1 0 176200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_561
timestamp 1654712443
transform 1 0 179200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_661
timestamp 1654712443
transform 1 0 179200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_563
timestamp 1654712443
transform 1 0 185200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_663
timestamp 1654712443
transform 1 0 185200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_562
timestamp 1654712443
transform 1 0 182200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_662
timestamp 1654712443
transform 1 0 182200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_564
timestamp 1654712443
transform 1 0 188200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_664
timestamp 1654712443
transform 1 0 188200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_565
timestamp 1654712443
transform 1 0 191200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_665
timestamp 1654712443
transform 1 0 191200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_566
timestamp 1654712443
transform 1 0 194200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_666
timestamp 1654712443
transform 1 0 194200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_567
timestamp 1654712443
transform 1 0 197200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_667
timestamp 1654712443
transform 1 0 197200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_568
timestamp 1654712443
transform 1 0 200200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_668
timestamp 1654712443
transform 1 0 200200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_569
timestamp 1654712443
transform 1 0 203200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_669
timestamp 1654712443
transform 1 0 203200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_570
timestamp 1654712443
transform 1 0 206200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_670
timestamp 1654712443
transform 1 0 206200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_571
timestamp 1654712443
transform 1 0 209200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_671
timestamp 1654712443
transform 1 0 209200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_573
timestamp 1654712443
transform 1 0 215200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_673
timestamp 1654712443
transform 1 0 215200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_572
timestamp 1654712443
transform 1 0 212200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_672
timestamp 1654712443
transform 1 0 212200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_574
timestamp 1654712443
transform 1 0 218200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_674
timestamp 1654712443
transform 1 0 218200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_575
timestamp 1654712443
transform 1 0 221200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_675
timestamp 1654712443
transform 1 0 221200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_576
timestamp 1654712443
transform 1 0 224200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_676
timestamp 1654712443
transform 1 0 224200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_577
timestamp 1654712443
transform 1 0 227200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_677
timestamp 1654712443
transform 1 0 227200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_578
timestamp 1654712443
transform 1 0 230200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_678
timestamp 1654712443
transform 1 0 230200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_579
timestamp 1654712443
transform 1 0 233200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_679
timestamp 1654712443
transform 1 0 233200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_580
timestamp 1654712443
transform 1 0 236200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_680
timestamp 1654712443
transform 1 0 236200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_581
timestamp 1654712443
transform 1 0 239200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_681
timestamp 1654712443
transform 1 0 239200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_583
timestamp 1654712443
transform 1 0 245200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_683
timestamp 1654712443
transform 1 0 245200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_582
timestamp 1654712443
transform 1 0 242200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_682
timestamp 1654712443
transform 1 0 242200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_584
timestamp 1654712443
transform 1 0 248200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_684
timestamp 1654712443
transform 1 0 248200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_585
timestamp 1654712443
transform 1 0 251200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_685
timestamp 1654712443
transform 1 0 251200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_586
timestamp 1654712443
transform 1 0 254200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_686
timestamp 1654712443
transform 1 0 254200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_587
timestamp 1654712443
transform 1 0 257200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_687
timestamp 1654712443
transform 1 0 257200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_588
timestamp 1654712443
transform 1 0 260200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_688
timestamp 1654712443
transform 1 0 260200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_589
timestamp 1654712443
transform 1 0 263200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_689
timestamp 1654712443
transform 1 0 263200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_590
timestamp 1654712443
transform 1 0 266200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_690
timestamp 1654712443
transform 1 0 266200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_591
timestamp 1654712443
transform 1 0 269200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_691
timestamp 1654712443
transform 1 0 269200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_592
timestamp 1654712443
transform 1 0 272200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_692
timestamp 1654712443
transform 1 0 272200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_594
timestamp 1654712443
transform 1 0 278200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_593
timestamp 1654712443
transform 1 0 275200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_694
timestamp 1654712443
transform 1 0 278200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_693
timestamp 1654712443
transform 1 0 275200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_595
timestamp 1654712443
transform 1 0 281200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_695
timestamp 1654712443
transform 1 0 281200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_596
timestamp 1654712443
transform 1 0 284200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_696
timestamp 1654712443
transform 1 0 284200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_597
timestamp 1654712443
transform 1 0 287200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_697
timestamp 1654712443
transform 1 0 287200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_598
timestamp 1654712443
transform 1 0 290200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_698
timestamp 1654712443
transform 1 0 290200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_599
timestamp 1654712443
transform 1 0 293200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_699
timestamp 1654712443
transform 1 0 293200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_401
timestamp 1654712443
transform 1 0 -800 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_400
timestamp 1654712443
transform 1 0 -3800 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_402
timestamp 1654712443
transform 1 0 2200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_403
timestamp 1654712443
transform 1 0 5200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_404
timestamp 1654712443
transform 1 0 8200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_405
timestamp 1654712443
transform 1 0 11200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_406
timestamp 1654712443
transform 1 0 14200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_407
timestamp 1654712443
transform 1 0 17200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_408
timestamp 1654712443
transform 1 0 20200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_409
timestamp 1654712443
transform 1 0 23200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_411
timestamp 1654712443
transform 1 0 29200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_410
timestamp 1654712443
transform 1 0 26200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_412
timestamp 1654712443
transform 1 0 32200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_413
timestamp 1654712443
transform 1 0 35200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_414
timestamp 1654712443
transform 1 0 38200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_415
timestamp 1654712443
transform 1 0 41200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_416
timestamp 1654712443
transform 1 0 44200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_417
timestamp 1654712443
transform 1 0 47200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_418
timestamp 1654712443
transform 1 0 50200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_419
timestamp 1654712443
transform 1 0 53200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_421
timestamp 1654712443
transform 1 0 59200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_420
timestamp 1654712443
transform 1 0 56200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_422
timestamp 1654712443
transform 1 0 62200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_423
timestamp 1654712443
transform 1 0 65200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_424
timestamp 1654712443
transform 1 0 68200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_425
timestamp 1654712443
transform 1 0 71200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_426
timestamp 1654712443
transform 1 0 74200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_427
timestamp 1654712443
transform 1 0 77200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_428
timestamp 1654712443
transform 1 0 80200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_429
timestamp 1654712443
transform 1 0 83200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_430
timestamp 1654712443
transform 1 0 86200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_432
timestamp 1654712443
transform 1 0 92200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_431
timestamp 1654712443
transform 1 0 89200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_433
timestamp 1654712443
transform 1 0 95200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_434
timestamp 1654712443
transform 1 0 98200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_435
timestamp 1654712443
transform 1 0 101200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_436
timestamp 1654712443
transform 1 0 104200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_437
timestamp 1654712443
transform 1 0 107200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_438
timestamp 1654712443
transform 1 0 110200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_439
timestamp 1654712443
transform 1 0 113200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_440
timestamp 1654712443
transform 1 0 116200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_442
timestamp 1654712443
transform 1 0 122200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_441
timestamp 1654712443
transform 1 0 119200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_443
timestamp 1654712443
transform 1 0 125200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_444
timestamp 1654712443
transform 1 0 128200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_445
timestamp 1654712443
transform 1 0 131200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_446
timestamp 1654712443
transform 1 0 134200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_447
timestamp 1654712443
transform 1 0 137200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_448
timestamp 1654712443
transform 1 0 140200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_449
timestamp 1654712443
transform 1 0 143200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_450
timestamp 1654712443
transform 1 0 146200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_452
timestamp 1654712443
transform 1 0 152200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_451
timestamp 1654712443
transform 1 0 149200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_453
timestamp 1654712443
transform 1 0 155200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_454
timestamp 1654712443
transform 1 0 158200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_455
timestamp 1654712443
transform 1 0 161200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_456
timestamp 1654712443
transform 1 0 164200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_457
timestamp 1654712443
transform 1 0 167200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_458
timestamp 1654712443
transform 1 0 170200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_459
timestamp 1654712443
transform 1 0 173200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_460
timestamp 1654712443
transform 1 0 176200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_461
timestamp 1654712443
transform 1 0 179200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_463
timestamp 1654712443
transform 1 0 185200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_462
timestamp 1654712443
transform 1 0 182200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_464
timestamp 1654712443
transform 1 0 188200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_465
timestamp 1654712443
transform 1 0 191200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_466
timestamp 1654712443
transform 1 0 194200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_467
timestamp 1654712443
transform 1 0 197200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_468
timestamp 1654712443
transform 1 0 200200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_469
timestamp 1654712443
transform 1 0 203200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_470
timestamp 1654712443
transform 1 0 206200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_471
timestamp 1654712443
transform 1 0 209200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_473
timestamp 1654712443
transform 1 0 215200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_472
timestamp 1654712443
transform 1 0 212200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_474
timestamp 1654712443
transform 1 0 218200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_475
timestamp 1654712443
transform 1 0 221200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_476
timestamp 1654712443
transform 1 0 224200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_477
timestamp 1654712443
transform 1 0 227200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_478
timestamp 1654712443
transform 1 0 230200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_479
timestamp 1654712443
transform 1 0 233200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_480
timestamp 1654712443
transform 1 0 236200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_481
timestamp 1654712443
transform 1 0 239200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_483
timestamp 1654712443
transform 1 0 245200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_482
timestamp 1654712443
transform 1 0 242200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_484
timestamp 1654712443
transform 1 0 248200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_485
timestamp 1654712443
transform 1 0 251200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_486
timestamp 1654712443
transform 1 0 254200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_487
timestamp 1654712443
transform 1 0 257200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_488
timestamp 1654712443
transform 1 0 260200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_489
timestamp 1654712443
transform 1 0 263200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_490
timestamp 1654712443
transform 1 0 266200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_491
timestamp 1654712443
transform 1 0 269200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_492
timestamp 1654712443
transform 1 0 272200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_494
timestamp 1654712443
transform 1 0 278200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_493
timestamp 1654712443
transform 1 0 275200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_495
timestamp 1654712443
transform 1 0 281200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_496
timestamp 1654712443
transform 1 0 284200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_497
timestamp 1654712443
transform 1 0 287200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_498
timestamp 1654712443
transform 1 0 290200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_499
timestamp 1654712443
transform 1 0 293200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_301
timestamp 1654712443
transform 1 0 -800 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_300
timestamp 1654712443
transform 1 0 -3800 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_302
timestamp 1654712443
transform 1 0 2200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_303
timestamp 1654712443
transform 1 0 5200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_304
timestamp 1654712443
transform 1 0 8200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_305
timestamp 1654712443
transform 1 0 11200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_306
timestamp 1654712443
transform 1 0 14200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_307
timestamp 1654712443
transform 1 0 17200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_308
timestamp 1654712443
transform 1 0 20200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_309
timestamp 1654712443
transform 1 0 23200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_311
timestamp 1654712443
transform 1 0 29200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_310
timestamp 1654712443
transform 1 0 26200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_312
timestamp 1654712443
transform 1 0 32200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_313
timestamp 1654712443
transform 1 0 35200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_314
timestamp 1654712443
transform 1 0 38200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_315
timestamp 1654712443
transform 1 0 41200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_316
timestamp 1654712443
transform 1 0 44200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_317
timestamp 1654712443
transform 1 0 47200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_318
timestamp 1654712443
transform 1 0 50200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_319
timestamp 1654712443
transform 1 0 53200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_321
timestamp 1654712443
transform 1 0 59200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_320
timestamp 1654712443
transform 1 0 56200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_322
timestamp 1654712443
transform 1 0 62200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_323
timestamp 1654712443
transform 1 0 65200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_324
timestamp 1654712443
transform 1 0 68200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_325
timestamp 1654712443
transform 1 0 71200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_326
timestamp 1654712443
transform 1 0 74200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_327
timestamp 1654712443
transform 1 0 77200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_328
timestamp 1654712443
transform 1 0 80200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_329
timestamp 1654712443
transform 1 0 83200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_330
timestamp 1654712443
transform 1 0 86200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_332
timestamp 1654712443
transform 1 0 92200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_331
timestamp 1654712443
transform 1 0 89200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_333
timestamp 1654712443
transform 1 0 95200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_334
timestamp 1654712443
transform 1 0 98200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_335
timestamp 1654712443
transform 1 0 101200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_336
timestamp 1654712443
transform 1 0 104200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_337
timestamp 1654712443
transform 1 0 107200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_338
timestamp 1654712443
transform 1 0 110200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_339
timestamp 1654712443
transform 1 0 113200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_340
timestamp 1654712443
transform 1 0 116200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_342
timestamp 1654712443
transform 1 0 122200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_341
timestamp 1654712443
transform 1 0 119200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_343
timestamp 1654712443
transform 1 0 125200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_344
timestamp 1654712443
transform 1 0 128200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_345
timestamp 1654712443
transform 1 0 131200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_346
timestamp 1654712443
transform 1 0 134200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_347
timestamp 1654712443
transform 1 0 137200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_348
timestamp 1654712443
transform 1 0 140200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_349
timestamp 1654712443
transform 1 0 143200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_350
timestamp 1654712443
transform 1 0 146200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_352
timestamp 1654712443
transform 1 0 152200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_351
timestamp 1654712443
transform 1 0 149200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_353
timestamp 1654712443
transform 1 0 155200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_354
timestamp 1654712443
transform 1 0 158200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_355
timestamp 1654712443
transform 1 0 161200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_356
timestamp 1654712443
transform 1 0 164200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_357
timestamp 1654712443
transform 1 0 167200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_358
timestamp 1654712443
transform 1 0 170200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_359
timestamp 1654712443
transform 1 0 173200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_360
timestamp 1654712443
transform 1 0 176200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_361
timestamp 1654712443
transform 1 0 179200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_363
timestamp 1654712443
transform 1 0 185200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_362
timestamp 1654712443
transform 1 0 182200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_364
timestamp 1654712443
transform 1 0 188200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_365
timestamp 1654712443
transform 1 0 191200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_366
timestamp 1654712443
transform 1 0 194200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_367
timestamp 1654712443
transform 1 0 197200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_368
timestamp 1654712443
transform 1 0 200200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_369
timestamp 1654712443
transform 1 0 203200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_370
timestamp 1654712443
transform 1 0 206200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_371
timestamp 1654712443
transform 1 0 209200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_373
timestamp 1654712443
transform 1 0 215200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_372
timestamp 1654712443
transform 1 0 212200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_374
timestamp 1654712443
transform 1 0 218200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_375
timestamp 1654712443
transform 1 0 221200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_376
timestamp 1654712443
transform 1 0 224200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_377
timestamp 1654712443
transform 1 0 227200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_378
timestamp 1654712443
transform 1 0 230200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_379
timestamp 1654712443
transform 1 0 233200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_380
timestamp 1654712443
transform 1 0 236200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_381
timestamp 1654712443
transform 1 0 239200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_383
timestamp 1654712443
transform 1 0 245200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_382
timestamp 1654712443
transform 1 0 242200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_384
timestamp 1654712443
transform 1 0 248200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_385
timestamp 1654712443
transform 1 0 251200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_386
timestamp 1654712443
transform 1 0 254200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_387
timestamp 1654712443
transform 1 0 257200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_388
timestamp 1654712443
transform 1 0 260200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_389
timestamp 1654712443
transform 1 0 263200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_390
timestamp 1654712443
transform 1 0 266200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_391
timestamp 1654712443
transform 1 0 269200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_392
timestamp 1654712443
transform 1 0 272200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_394
timestamp 1654712443
transform 1 0 278200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_393
timestamp 1654712443
transform 1 0 275200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_395
timestamp 1654712443
transform 1 0 281200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_396
timestamp 1654712443
transform 1 0 284200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_397
timestamp 1654712443
transform 1 0 287200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_398
timestamp 1654712443
transform 1 0 290200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_399
timestamp 1654712443
transform 1 0 293200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_201
timestamp 1654712443
transform 1 0 -800 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_200
timestamp 1654712443
transform 1 0 -3800 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_202
timestamp 1654712443
transform 1 0 2200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_203
timestamp 1654712443
transform 1 0 5200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_204
timestamp 1654712443
transform 1 0 8200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_205
timestamp 1654712443
transform 1 0 11200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_206
timestamp 1654712443
transform 1 0 14200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_207
timestamp 1654712443
transform 1 0 17200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_208
timestamp 1654712443
transform 1 0 20200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_209
timestamp 1654712443
transform 1 0 23200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_211
timestamp 1654712443
transform 1 0 29200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_210
timestamp 1654712443
transform 1 0 26200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_212
timestamp 1654712443
transform 1 0 32200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_213
timestamp 1654712443
transform 1 0 35200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_214
timestamp 1654712443
transform 1 0 38200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_215
timestamp 1654712443
transform 1 0 41200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_216
timestamp 1654712443
transform 1 0 44200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_217
timestamp 1654712443
transform 1 0 47200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_218
timestamp 1654712443
transform 1 0 50200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_219
timestamp 1654712443
transform 1 0 53200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_221
timestamp 1654712443
transform 1 0 59200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_220
timestamp 1654712443
transform 1 0 56200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_222
timestamp 1654712443
transform 1 0 62200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_223
timestamp 1654712443
transform 1 0 65200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_224
timestamp 1654712443
transform 1 0 68200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_225
timestamp 1654712443
transform 1 0 71200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_226
timestamp 1654712443
transform 1 0 74200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_227
timestamp 1654712443
transform 1 0 77200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_228
timestamp 1654712443
transform 1 0 80200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_229
timestamp 1654712443
transform 1 0 83200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_230
timestamp 1654712443
transform 1 0 86200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_232
timestamp 1654712443
transform 1 0 92200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_231
timestamp 1654712443
transform 1 0 89200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_233
timestamp 1654712443
transform 1 0 95200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_234
timestamp 1654712443
transform 1 0 98200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_235
timestamp 1654712443
transform 1 0 101200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_236
timestamp 1654712443
transform 1 0 104200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_237
timestamp 1654712443
transform 1 0 107200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_238
timestamp 1654712443
transform 1 0 110200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_239
timestamp 1654712443
transform 1 0 113200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_240
timestamp 1654712443
transform 1 0 116200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_242
timestamp 1654712443
transform 1 0 122200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_241
timestamp 1654712443
transform 1 0 119200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_243
timestamp 1654712443
transform 1 0 125200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_244
timestamp 1654712443
transform 1 0 128200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_245
timestamp 1654712443
transform 1 0 131200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_246
timestamp 1654712443
transform 1 0 134200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_247
timestamp 1654712443
transform 1 0 137200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_248
timestamp 1654712443
transform 1 0 140200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_249
timestamp 1654712443
transform 1 0 143200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_250
timestamp 1654712443
transform 1 0 146200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_252
timestamp 1654712443
transform 1 0 152200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_251
timestamp 1654712443
transform 1 0 149200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_253
timestamp 1654712443
transform 1 0 155200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_254
timestamp 1654712443
transform 1 0 158200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_255
timestamp 1654712443
transform 1 0 161200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_256
timestamp 1654712443
transform 1 0 164200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_257
timestamp 1654712443
transform 1 0 167200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_258
timestamp 1654712443
transform 1 0 170200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_259
timestamp 1654712443
transform 1 0 173200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_260
timestamp 1654712443
transform 1 0 176200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_261
timestamp 1654712443
transform 1 0 179200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_263
timestamp 1654712443
transform 1 0 185200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_262
timestamp 1654712443
transform 1 0 182200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_264
timestamp 1654712443
transform 1 0 188200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_265
timestamp 1654712443
transform 1 0 191200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_266
timestamp 1654712443
transform 1 0 194200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_267
timestamp 1654712443
transform 1 0 197200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_268
timestamp 1654712443
transform 1 0 200200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_269
timestamp 1654712443
transform 1 0 203200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_270
timestamp 1654712443
transform 1 0 206200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_271
timestamp 1654712443
transform 1 0 209200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_273
timestamp 1654712443
transform 1 0 215200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_272
timestamp 1654712443
transform 1 0 212200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_274
timestamp 1654712443
transform 1 0 218200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_275
timestamp 1654712443
transform 1 0 221200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_276
timestamp 1654712443
transform 1 0 224200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_277
timestamp 1654712443
transform 1 0 227200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_278
timestamp 1654712443
transform 1 0 230200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_279
timestamp 1654712443
transform 1 0 233200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_280
timestamp 1654712443
transform 1 0 236200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_281
timestamp 1654712443
transform 1 0 239200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_283
timestamp 1654712443
transform 1 0 245200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_282
timestamp 1654712443
transform 1 0 242200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_284
timestamp 1654712443
transform 1 0 248200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_285
timestamp 1654712443
transform 1 0 251200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_286
timestamp 1654712443
transform 1 0 254200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_287
timestamp 1654712443
transform 1 0 257200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_288
timestamp 1654712443
transform 1 0 260200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_289
timestamp 1654712443
transform 1 0 263200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_290
timestamp 1654712443
transform 1 0 266200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_291
timestamp 1654712443
transform 1 0 269200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_292
timestamp 1654712443
transform 1 0 272200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_294
timestamp 1654712443
transform 1 0 278200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_293
timestamp 1654712443
transform 1 0 275200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_295
timestamp 1654712443
transform 1 0 281200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_296
timestamp 1654712443
transform 1 0 284200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_297
timestamp 1654712443
transform 1 0 287200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_298
timestamp 1654712443
transform 1 0 290200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_299
timestamp 1654712443
transform 1 0 293200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_101
timestamp 1654712443
transform 1 0 -800 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_100
timestamp 1654712443
transform 1 0 -3800 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_102
timestamp 1654712443
transform 1 0 2200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_103
timestamp 1654712443
transform 1 0 5200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_104
timestamp 1654712443
transform 1 0 8200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_105
timestamp 1654712443
transform 1 0 11200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_106
timestamp 1654712443
transform 1 0 14200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_107
timestamp 1654712443
transform 1 0 17200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_108
timestamp 1654712443
transform 1 0 20200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_109
timestamp 1654712443
transform 1 0 23200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_111
timestamp 1654712443
transform 1 0 29200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_110
timestamp 1654712443
transform 1 0 26200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_112
timestamp 1654712443
transform 1 0 32200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_113
timestamp 1654712443
transform 1 0 35200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_114
timestamp 1654712443
transform 1 0 38200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_115
timestamp 1654712443
transform 1 0 41200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_116
timestamp 1654712443
transform 1 0 44200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_117
timestamp 1654712443
transform 1 0 47200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_118
timestamp 1654712443
transform 1 0 50200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_119
timestamp 1654712443
transform 1 0 53200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_121
timestamp 1654712443
transform 1 0 59200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_120
timestamp 1654712443
transform 1 0 56200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_122
timestamp 1654712443
transform 1 0 62200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_123
timestamp 1654712443
transform 1 0 65200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_124
timestamp 1654712443
transform 1 0 68200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_125
timestamp 1654712443
transform 1 0 71200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_126
timestamp 1654712443
transform 1 0 74200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_127
timestamp 1654712443
transform 1 0 77200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_128
timestamp 1654712443
transform 1 0 80200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_129
timestamp 1654712443
transform 1 0 83200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_130
timestamp 1654712443
transform 1 0 86200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_132
timestamp 1654712443
transform 1 0 92200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_131
timestamp 1654712443
transform 1 0 89200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_133
timestamp 1654712443
transform 1 0 95200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_134
timestamp 1654712443
transform 1 0 98200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_135
timestamp 1654712443
transform 1 0 101200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_136
timestamp 1654712443
transform 1 0 104200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_137
timestamp 1654712443
transform 1 0 107200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_138
timestamp 1654712443
transform 1 0 110200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_139
timestamp 1654712443
transform 1 0 113200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_140
timestamp 1654712443
transform 1 0 116200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_142
timestamp 1654712443
transform 1 0 122200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_141
timestamp 1654712443
transform 1 0 119200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_143
timestamp 1654712443
transform 1 0 125200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_144
timestamp 1654712443
transform 1 0 128200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_145
timestamp 1654712443
transform 1 0 131200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_146
timestamp 1654712443
transform 1 0 134200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_147
timestamp 1654712443
transform 1 0 137200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_148
timestamp 1654712443
transform 1 0 140200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_149
timestamp 1654712443
transform 1 0 143200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_150
timestamp 1654712443
transform 1 0 146200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_152
timestamp 1654712443
transform 1 0 152200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_151
timestamp 1654712443
transform 1 0 149200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_153
timestamp 1654712443
transform 1 0 155200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_154
timestamp 1654712443
transform 1 0 158200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_155
timestamp 1654712443
transform 1 0 161200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_156
timestamp 1654712443
transform 1 0 164200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_157
timestamp 1654712443
transform 1 0 167200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_158
timestamp 1654712443
transform 1 0 170200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_159
timestamp 1654712443
transform 1 0 173200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_160
timestamp 1654712443
transform 1 0 176200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_161
timestamp 1654712443
transform 1 0 179200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_163
timestamp 1654712443
transform 1 0 185200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_162
timestamp 1654712443
transform 1 0 182200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_164
timestamp 1654712443
transform 1 0 188200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_165
timestamp 1654712443
transform 1 0 191200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_166
timestamp 1654712443
transform 1 0 194200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_167
timestamp 1654712443
transform 1 0 197200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_168
timestamp 1654712443
transform 1 0 200200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_169
timestamp 1654712443
transform 1 0 203200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_170
timestamp 1654712443
transform 1 0 206200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_171
timestamp 1654712443
transform 1 0 209200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_173
timestamp 1654712443
transform 1 0 215200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_172
timestamp 1654712443
transform 1 0 212200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_174
timestamp 1654712443
transform 1 0 218200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_175
timestamp 1654712443
transform 1 0 221200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_176
timestamp 1654712443
transform 1 0 224200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_177
timestamp 1654712443
transform 1 0 227200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_178
timestamp 1654712443
transform 1 0 230200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_179
timestamp 1654712443
transform 1 0 233200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_180
timestamp 1654712443
transform 1 0 236200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_181
timestamp 1654712443
transform 1 0 239200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_183
timestamp 1654712443
transform 1 0 245200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_182
timestamp 1654712443
transform 1 0 242200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_184
timestamp 1654712443
transform 1 0 248200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_185
timestamp 1654712443
transform 1 0 251200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_186
timestamp 1654712443
transform 1 0 254200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_187
timestamp 1654712443
transform 1 0 257200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_188
timestamp 1654712443
transform 1 0 260200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_189
timestamp 1654712443
transform 1 0 263200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_190
timestamp 1654712443
transform 1 0 266200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_191
timestamp 1654712443
transform 1 0 269200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_192
timestamp 1654712443
transform 1 0 272200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_194
timestamp 1654712443
transform 1 0 278200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_193
timestamp 1654712443
transform 1 0 275200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_195
timestamp 1654712443
transform 1 0 281200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_196
timestamp 1654712443
transform 1 0 284200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_197
timestamp 1654712443
transform 1 0 287200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_198
timestamp 1654712443
transform 1 0 290200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_199
timestamp 1654712443
transform 1 0 293200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_1
timestamp 1654712443
transform 1 0 -800 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_0
timestamp 1654712443
transform 1 0 -3800 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_2
timestamp 1654712443
transform 1 0 2200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_3
timestamp 1654712443
transform 1 0 5200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_4
timestamp 1654712443
transform 1 0 8200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_5
timestamp 1654712443
transform 1 0 11200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_6
timestamp 1654712443
transform 1 0 14200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_7
timestamp 1654712443
transform 1 0 17200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_8
timestamp 1654712443
transform 1 0 20200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_9
timestamp 1654712443
transform 1 0 23200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_11
timestamp 1654712443
transform 1 0 29200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_10
timestamp 1654712443
transform 1 0 26200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_12
timestamp 1654712443
transform 1 0 32200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_13
timestamp 1654712443
transform 1 0 35200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_14
timestamp 1654712443
transform 1 0 38200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_15
timestamp 1654712443
transform 1 0 41200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_16
timestamp 1654712443
transform 1 0 44200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_17
timestamp 1654712443
transform 1 0 47200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_18
timestamp 1654712443
transform 1 0 50200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_19
timestamp 1654712443
transform 1 0 53200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_21
timestamp 1654712443
transform 1 0 59200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_20
timestamp 1654712443
transform 1 0 56200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_22
timestamp 1654712443
transform 1 0 62200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_23
timestamp 1654712443
transform 1 0 65200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_24
timestamp 1654712443
transform 1 0 68200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_25
timestamp 1654712443
transform 1 0 71200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_26
timestamp 1654712443
transform 1 0 74200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_27
timestamp 1654712443
transform 1 0 77200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_28
timestamp 1654712443
transform 1 0 80200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_29
timestamp 1654712443
transform 1 0 83200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_30
timestamp 1654712443
transform 1 0 86200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_32
timestamp 1654712443
transform 1 0 92200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_31
timestamp 1654712443
transform 1 0 89200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_33
timestamp 1654712443
transform 1 0 95200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_34
timestamp 1654712443
transform 1 0 98200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_35
timestamp 1654712443
transform 1 0 101200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_36
timestamp 1654712443
transform 1 0 104200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_37
timestamp 1654712443
transform 1 0 107200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_38
timestamp 1654712443
transform 1 0 110200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_39
timestamp 1654712443
transform 1 0 113200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_40
timestamp 1654712443
transform 1 0 116200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_42
timestamp 1654712443
transform 1 0 122200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_41
timestamp 1654712443
transform 1 0 119200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_43
timestamp 1654712443
transform 1 0 125200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_44
timestamp 1654712443
transform 1 0 128200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_45
timestamp 1654712443
transform 1 0 131200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_46
timestamp 1654712443
transform 1 0 134200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_47
timestamp 1654712443
transform 1 0 137200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_48
timestamp 1654712443
transform 1 0 140200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_49
timestamp 1654712443
transform 1 0 143200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_50
timestamp 1654712443
transform 1 0 146200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_52
timestamp 1654712443
transform 1 0 152200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_51
timestamp 1654712443
transform 1 0 149200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_53
timestamp 1654712443
transform 1 0 155200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_54
timestamp 1654712443
transform 1 0 158200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_55
timestamp 1654712443
transform 1 0 161200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_56
timestamp 1654712443
transform 1 0 164200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_57
timestamp 1654712443
transform 1 0 167200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_58
timestamp 1654712443
transform 1 0 170200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_59
timestamp 1654712443
transform 1 0 173200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_60
timestamp 1654712443
transform 1 0 176200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_61
timestamp 1654712443
transform 1 0 179200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_63
timestamp 1654712443
transform 1 0 185200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_62
timestamp 1654712443
transform 1 0 182200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_64
timestamp 1654712443
transform 1 0 188200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_65
timestamp 1654712443
transform 1 0 191200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_66
timestamp 1654712443
transform 1 0 194200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_67
timestamp 1654712443
transform 1 0 197200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_68
timestamp 1654712443
transform 1 0 200200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_69
timestamp 1654712443
transform 1 0 203200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_70
timestamp 1654712443
transform 1 0 206200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_71
timestamp 1654712443
transform 1 0 209200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_73
timestamp 1654712443
transform 1 0 215200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_72
timestamp 1654712443
transform 1 0 212200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_74
timestamp 1654712443
transform 1 0 218200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_75
timestamp 1654712443
transform 1 0 221200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_76
timestamp 1654712443
transform 1 0 224200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_77
timestamp 1654712443
transform 1 0 227200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_78
timestamp 1654712443
transform 1 0 230200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_79
timestamp 1654712443
transform 1 0 233200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_80
timestamp 1654712443
transform 1 0 236200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_81
timestamp 1654712443
transform 1 0 239200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_83
timestamp 1654712443
transform 1 0 245200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_82
timestamp 1654712443
transform 1 0 242200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_84
timestamp 1654712443
transform 1 0 248200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_85
timestamp 1654712443
transform 1 0 251200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_86
timestamp 1654712443
transform 1 0 254200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_87
timestamp 1654712443
transform 1 0 257200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_88
timestamp 1654712443
transform 1 0 260200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_89
timestamp 1654712443
transform 1 0 263200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_90
timestamp 1654712443
transform 1 0 266200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_91
timestamp 1654712443
transform 1 0 269200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_92
timestamp 1654712443
transform 1 0 272200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_94
timestamp 1654712443
transform 1 0 278200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_93
timestamp 1654712443
transform 1 0 275200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_95
timestamp 1654712443
transform 1 0 281200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_96
timestamp 1654712443
transform 1 0 284200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_97
timestamp 1654712443
transform 1 0 287200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_98
timestamp 1654712443
transform 1 0 290200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_99
timestamp 1654712443
transform 1 0 293200 0 1 2700
box 3640 -2860 6960 460
<< labels >>
rlabel metal4 -3000 3550 -3000 3660 1 VBIAS
port 2 n
rlabel metal2 -3000 3350 -3000 3450 3 VREF
port 3 e
rlabel metal2 0 4040 0 4040 1 NB2
port 4 n
rlabel metal1 -2000 0 -2000 0 1 VDD
port 5 n
rlabel space -1160 5750 -1160 5750 5 SF_IB
port 6 s
rlabel metal2 -740 3560 -740 3560 1 NB1
port 7 n
rlabel metal2 -3000 1480 -3000 1570 3 ROW_SEL[0]
port 8 e
rlabel metal5 -2000 2840 -2000 2840 1 GRING
port 9 n
rlabel metal1 300400 30 300400 30 1 GND
port 109 n
rlabel metal2 -3000 -1520 -3000 -1430 3 ROW_SEL[1]
port 111 e
rlabel metal2 -3000 -4520 -3000 -4430 3 ROW_SEL[2]
port 212 e
rlabel metal2 -3000 -7520 -3000 -7430 3 ROW_SEL[3]
port 313 e
rlabel metal2 -3000 -10520 -3000 -10430 3 ROW_SEL[4]
port 414 e
rlabel metal2 -3000 -13520 -3000 -13430 3 ROW_SEL[5]
port 515 e
rlabel metal2 -3000 -16520 -3000 -16430 3 ROW_SEL[6]
port 616 e
rlabel metal2 -3000 -19520 -3000 -19430 3 ROW_SEL[7]
port 717 e
rlabel metal2 -3000 -22520 -3000 -22430 3 ROW_SEL[8]
port 818 e
rlabel metal2 -3000 -25520 -3000 -25430 3 ROW_SEL[9]
port 919 e
rlabel metal2 -3000 -28520 -3000 -28430 3 ROW_SEL[10]
port 1020 e
rlabel metal2 -3000 -31520 -3000 -31430 3 ROW_SEL[11]
port 1121 e
rlabel metal2 -3000 -34520 -3000 -34430 3 ROW_SEL[12]
port 1222 e
rlabel metal2 -3000 -37520 -3000 -37430 3 ROW_SEL[13]
port 1323 e
rlabel metal2 -3000 -40520 -3000 -40430 3 ROW_SEL[14]
port 1424 e
rlabel metal2 -3000 -43520 -3000 -43430 3 ROW_SEL[15]
port 1525 e
rlabel metal2 -3000 -46520 -3000 -46430 3 ROW_SEL[16]
port 1626 e
rlabel metal2 -3000 -49520 -3000 -49430 3 ROW_SEL[17]
port 1727 e
rlabel metal2 -3000 -52520 -3000 -52430 3 ROW_SEL[18]
port 1828 e
rlabel metal2 -3000 -55520 -3000 -55430 3 ROW_SEL[19]
port 1929 e
rlabel metal2 -3000 -58520 -3000 -58430 3 ROW_SEL[20]
port 2030 e
rlabel metal2 -3000 -61520 -3000 -61430 3 ROW_SEL[21]
port 2131 e
rlabel metal2 -3000 -64520 -3000 -64430 3 ROW_SEL[22]
port 2232 e
rlabel metal2 -3000 -67520 -3000 -67430 3 ROW_SEL[23]
port 2333 e
rlabel metal2 -3000 -70520 -3000 -70430 3 ROW_SEL[24]
port 2434 e
rlabel metal2 -3000 -73520 -3000 -73430 3 ROW_SEL[25]
port 2535 e
rlabel metal2 -3000 -76520 -3000 -76430 3 ROW_SEL[26]
port 2636 e
rlabel metal2 -3000 -79520 -3000 -79430 3 ROW_SEL[27]
port 2737 e
rlabel metal2 -3000 -82520 -3000 -82430 3 ROW_SEL[28]
port 2838 e
rlabel metal2 -3000 -85520 -3000 -85430 3 ROW_SEL[29]
port 2939 e
rlabel metal2 -3000 -88520 -3000 -88430 3 ROW_SEL[30]
port 3040 e
rlabel metal2 -3000 -91520 -3000 -91430 3 ROW_SEL[31]
port 3141 e
rlabel metal2 -3000 -94520 -3000 -94430 3 ROW_SEL[32]
port 3242 e
rlabel metal2 -3000 -97520 -3000 -97430 3 ROW_SEL[33]
port 3343 e
rlabel metal2 -3000 -100520 -3000 -100430 3 ROW_SEL[34]
port 3444 e
rlabel metal2 -3000 -103520 -3000 -103430 3 ROW_SEL[35]
port 3545 e
rlabel metal2 -3000 -106520 -3000 -106430 3 ROW_SEL[36]
port 3646 e
rlabel metal2 -3000 -109520 -3000 -109430 3 ROW_SEL[37]
port 3747 e
rlabel metal2 -3000 -112520 -3000 -112430 3 ROW_SEL[38]
port 3848 e
rlabel metal2 -3000 -115520 -3000 -115430 3 ROW_SEL[39]
port 3949 e
rlabel metal2 -3000 -118520 -3000 -118430 3 ROW_SEL[40]
port 4050 e
rlabel metal2 -3000 -121520 -3000 -121430 3 ROW_SEL[41]
port 4151 e
rlabel metal2 -3000 -124520 -3000 -124430 3 ROW_SEL[42]
port 4252 e
rlabel metal2 -3000 -127520 -3000 -127430 3 ROW_SEL[43]
port 4353 e
rlabel metal2 -3000 -130520 -3000 -130430 3 ROW_SEL[44]
port 4454 e
rlabel metal2 -3000 -133520 -3000 -133430 3 ROW_SEL[45]
port 4555 e
rlabel metal2 -3000 -136520 -3000 -136430 3 ROW_SEL[46]
port 4656 e
rlabel metal2 -3000 -139520 -3000 -139430 3 ROW_SEL[47]
port 4757 e
rlabel metal2 -3000 -142520 -3000 -142430 3 ROW_SEL[48]
port 4858 e
rlabel metal2 -3000 -145520 -3000 -145430 3 ROW_SEL[49]
port 4959 e
rlabel metal2 -3000 -148520 -3000 -148430 3 ROW_SEL[50]
port 5060 e
rlabel metal2 -3000 -151520 -3000 -151430 3 ROW_SEL[51]
port 5161 e
rlabel metal2 -3000 -154520 -3000 -154430 3 ROW_SEL[52]
port 5262 e
rlabel metal2 -3000 -157520 -3000 -157430 3 ROW_SEL[53]
port 5363 e
rlabel metal2 -3000 -160520 -3000 -160430 3 ROW_SEL[54]
port 5464 e
rlabel metal2 -3000 -163520 -3000 -163430 3 ROW_SEL[55]
port 5565 e
rlabel metal2 -3000 -166520 -3000 -166430 3 ROW_SEL[56]
port 5666 e
rlabel metal2 -3000 -169520 -3000 -169430 3 ROW_SEL[57]
port 5767 e
rlabel metal2 -3000 -172520 -3000 -172430 3 ROW_SEL[58]
port 5868 e
rlabel metal2 -3000 -175520 -3000 -175430 3 ROW_SEL[59]
port 5969 e
rlabel metal2 -3000 -178520 -3000 -178430 3 ROW_SEL[60]
port 6070 e
rlabel metal2 -3000 -181520 -3000 -181430 3 ROW_SEL[61]
port 6171 e
rlabel metal2 -3000 -184520 -3000 -184430 3 ROW_SEL[62]
port 6272 e
rlabel metal2 -3000 -187520 -3000 -187430 3 ROW_SEL[63]
port 6373 e
rlabel metal2 -3000 -190520 -3000 -190430 3 ROW_SEL[64]
port 6474 e
rlabel metal2 -3000 -193520 -3000 -193430 3 ROW_SEL[65]
port 6575 e
rlabel metal2 -3000 -196520 -3000 -196430 3 ROW_SEL[66]
port 6676 e
rlabel metal2 -3000 -199520 -3000 -199430 3 ROW_SEL[67]
port 6777 e
rlabel metal2 -3000 -202520 -3000 -202430 3 ROW_SEL[68]
port 6878 e
rlabel metal2 -3000 -205520 -3000 -205430 3 ROW_SEL[69]
port 6979 e
rlabel metal2 -3000 -208520 -3000 -208430 3 ROW_SEL[70]
port 7080 e
rlabel metal2 -3000 -211520 -3000 -211430 3 ROW_SEL[71]
port 7181 e
rlabel metal2 -3000 -214520 -3000 -214430 3 ROW_SEL[72]
port 7282 e
rlabel metal2 -3000 -217520 -3000 -217430 3 ROW_SEL[73]
port 7383 e
rlabel metal2 -3000 -220520 -3000 -220430 3 ROW_SEL[74]
port 7484 e
rlabel metal2 -3000 -223520 -3000 -223430 3 ROW_SEL[75]
port 7585 e
rlabel metal2 -3000 -226520 -3000 -226430 3 ROW_SEL[76]
port 7686 e
rlabel metal2 -3000 -229520 -3000 -229430 3 ROW_SEL[77]
port 7787 e
rlabel metal2 -3000 -232520 -3000 -232430 3 ROW_SEL[78]
port 7888 e
rlabel metal2 -3000 -235520 -3000 -235430 3 ROW_SEL[79]
port 7989 e
rlabel metal2 -3000 -238520 -3000 -238430 3 ROW_SEL[80]
port 8090 e
rlabel metal2 -3000 -241520 -3000 -241430 3 ROW_SEL[81]
port 8191 e
rlabel metal2 -3000 -244520 -3000 -244430 3 ROW_SEL[82]
port 8292 e
rlabel metal2 -3000 -247520 -3000 -247430 3 ROW_SEL[83]
port 8393 e
rlabel metal2 -3000 -250520 -3000 -250430 3 ROW_SEL[84]
port 8494 e
rlabel metal2 -3000 -253520 -3000 -253430 3 ROW_SEL[85]
port 8595 e
rlabel metal2 -3000 -256520 -3000 -256430 3 ROW_SEL[86]
port 8696 e
rlabel metal2 -3000 -259520 -3000 -259430 3 ROW_SEL[87]
port 8797 e
rlabel metal2 -3000 -262520 -3000 -262430 3 ROW_SEL[88]
port 8898 e
rlabel metal2 -3000 -265520 -3000 -265430 3 ROW_SEL[89]
port 8999 e
rlabel metal2 -3000 -268520 -3000 -268430 3 ROW_SEL[90]
port 9100 e
rlabel metal2 -3000 -271520 -3000 -271430 3 ROW_SEL[91]
port 9201 e
rlabel metal2 -3000 -274520 -3000 -274430 3 ROW_SEL[92]
port 9302 e
rlabel metal2 -3000 -277520 -3000 -277430 3 ROW_SEL[93]
port 9403 e
rlabel metal2 -3000 -280520 -3000 -280430 3 ROW_SEL[94]
port 9504 e
rlabel metal2 -3000 -283520 -3000 -283430 3 ROW_SEL[95]
port 9605 e
rlabel metal2 -3000 -286520 -3000 -286430 3 ROW_SEL[96]
port 9706 e
rlabel metal2 -3000 -289520 -3000 -289430 3 ROW_SEL[97]
port 9807 e
rlabel metal2 -3000 -292520 -3000 -292430 3 ROW_SEL[98]
port 9908 e
rlabel metal4 2630 -297200 2780 -297000 1 PIX_OUT0
port 10009 n
rlabel metal4 220 -298100 440 -298100 1 COL_SEL[0]
port 10010 n
rlabel metal4 -480 -298600 -480 -298600 1 CSA_VREF
port 10011 n
rlabel metal2 -3000 -295520 -3000 -295430 3 ROW_SEL[99]
port 10012 e
rlabel metal4 5630 -297200 5780 -297000 1 PIX_OUT1
port 10014 n
rlabel metal4 3220 -298100 3440 -298100 1 COL_SEL[1]
port 10015 n
rlabel metal4 8630 -297200 8780 -297000 1 PIX_OUT2
port 10017 n
rlabel metal4 6220 -298100 6440 -298100 1 COL_SEL[2]
port 10018 n
rlabel metal4 11630 -297200 11780 -297000 1 PIX_OUT3
port 10020 n
rlabel metal4 9220 -298100 9440 -298100 1 COL_SEL[3]
port 10021 n
rlabel metal4 14630 -297200 14780 -297000 1 PIX_OUT4
port 10023 n
rlabel metal4 12220 -298100 12440 -298100 1 COL_SEL[4]
port 10024 n
rlabel metal4 17630 -297200 17780 -297000 1 PIX_OUT5
port 10026 n
rlabel metal4 15220 -298100 15440 -298100 1 COL_SEL[5]
port 10027 n
rlabel metal4 20630 -297200 20780 -297000 1 PIX_OUT6
port 10029 n
rlabel metal4 18220 -298100 18440 -298100 1 COL_SEL[6]
port 10030 n
rlabel metal4 23630 -297200 23780 -297000 1 PIX_OUT7
port 10032 n
rlabel metal4 21220 -298100 21440 -298100 1 COL_SEL[7]
port 10033 n
rlabel metal4 26630 -297200 26780 -297000 1 PIX_OUT8
port 10035 n
rlabel metal4 24220 -298100 24440 -298100 1 COL_SEL[8]
port 10036 n
rlabel metal4 29630 -297200 29780 -297000 1 PIX_OUT9
port 10038 n
rlabel metal4 27220 -298100 27440 -298100 1 COL_SEL[9]
port 10039 n
rlabel metal4 32630 -297200 32780 -297000 1 PIX_OUT10
port 10041 n
rlabel metal4 30220 -298100 30440 -298100 1 COL_SEL[10]
port 10042 n
rlabel metal4 35630 -297200 35780 -297000 1 PIX_OUT11
port 10044 n
rlabel metal4 33220 -298100 33440 -298100 1 COL_SEL[11]
port 10045 n
rlabel metal4 38630 -297200 38780 -297000 1 PIX_OUT12
port 10047 n
rlabel metal4 36220 -298100 36440 -298100 1 COL_SEL[12]
port 10048 n
rlabel metal4 41630 -297200 41780 -297000 1 PIX_OUT13
port 10050 n
rlabel metal4 39220 -298100 39440 -298100 1 COL_SEL[13]
port 10051 n
rlabel metal4 44630 -297200 44780 -297000 1 PIX_OUT14
port 10053 n
rlabel metal4 42220 -298100 42440 -298100 1 COL_SEL[14]
port 10054 n
rlabel metal4 47630 -297200 47780 -297000 1 PIX_OUT15
port 10056 n
rlabel metal4 45220 -298100 45440 -298100 1 COL_SEL[15]
port 10057 n
rlabel metal4 50630 -297200 50780 -297000 1 PIX_OUT16
port 10059 n
rlabel metal4 48220 -298100 48440 -298100 1 COL_SEL[16]
port 10060 n
rlabel metal4 53630 -297200 53780 -297000 1 PIX_OUT17
port 10062 n
rlabel metal4 51220 -298100 51440 -298100 1 COL_SEL[17]
port 10063 n
rlabel metal4 56630 -297200 56780 -297000 1 PIX_OUT18
port 10065 n
rlabel metal4 54220 -298100 54440 -298100 1 COL_SEL[18]
port 10066 n
rlabel metal4 59630 -297200 59780 -297000 1 PIX_OUT19
port 10068 n
rlabel metal4 57220 -298100 57440 -298100 1 COL_SEL[19]
port 10069 n
rlabel metal4 62630 -297200 62780 -297000 1 PIX_OUT20
port 10071 n
rlabel metal4 60220 -298100 60440 -298100 1 COL_SEL[20]
port 10072 n
rlabel metal4 65630 -297200 65780 -297000 1 PIX_OUT21
port 10074 n
rlabel metal4 63220 -298100 63440 -298100 1 COL_SEL[21]
port 10075 n
rlabel metal4 68630 -297200 68780 -297000 1 PIX_OUT22
port 10077 n
rlabel metal4 66220 -298100 66440 -298100 1 COL_SEL[22]
port 10078 n
rlabel metal4 71630 -297200 71780 -297000 1 PIX_OUT23
port 10080 n
rlabel metal4 69220 -298100 69440 -298100 1 COL_SEL[23]
port 10081 n
rlabel metal4 74630 -297200 74780 -297000 1 PIX_OUT24
port 10083 n
rlabel metal4 72220 -298100 72440 -298100 1 COL_SEL[24]
port 10084 n
rlabel metal4 77630 -297200 77780 -297000 1 PIX_OUT25
port 10086 n
rlabel metal4 75220 -298100 75440 -298100 1 COL_SEL[25]
port 10087 n
rlabel metal4 80630 -297200 80780 -297000 1 PIX_OUT26
port 10089 n
rlabel metal4 78220 -298100 78440 -298100 1 COL_SEL[26]
port 10090 n
rlabel metal4 83630 -297200 83780 -297000 1 PIX_OUT27
port 10092 n
rlabel metal4 81220 -298100 81440 -298100 1 COL_SEL[27]
port 10093 n
rlabel metal4 86630 -297200 86780 -297000 1 PIX_OUT28
port 10095 n
rlabel metal4 84220 -298100 84440 -298100 1 COL_SEL[28]
port 10096 n
rlabel metal4 89630 -297200 89780 -297000 1 PIX_OUT29
port 10098 n
rlabel metal4 87220 -298100 87440 -298100 1 COL_SEL[29]
port 10099 n
rlabel metal4 92630 -297200 92780 -297000 1 PIX_OUT30
port 10101 n
rlabel metal4 90220 -298100 90440 -298100 1 COL_SEL[30]
port 10102 n
rlabel metal4 95630 -297200 95780 -297000 1 PIX_OUT31
port 10104 n
rlabel metal4 93220 -298100 93440 -298100 1 COL_SEL[31]
port 10105 n
rlabel metal4 98630 -297200 98780 -297000 1 PIX_OUT32
port 10107 n
rlabel metal4 96220 -298100 96440 -298100 1 COL_SEL[32]
port 10108 n
rlabel metal4 101630 -297200 101780 -297000 1 PIX_OUT33
port 10110 n
rlabel metal4 99220 -298100 99440 -298100 1 COL_SEL[33]
port 10111 n
rlabel metal4 104630 -297200 104780 -297000 1 PIX_OUT34
port 10113 n
rlabel metal4 102220 -298100 102440 -298100 1 COL_SEL[34]
port 10114 n
rlabel metal4 107630 -297200 107780 -297000 1 PIX_OUT35
port 10116 n
rlabel metal4 105220 -298100 105440 -298100 1 COL_SEL[35]
port 10117 n
rlabel metal4 110630 -297200 110780 -297000 1 PIX_OUT36
port 10119 n
rlabel metal4 108220 -298100 108440 -298100 1 COL_SEL[36]
port 10120 n
rlabel metal4 113630 -297200 113780 -297000 1 PIX_OUT37
port 10122 n
rlabel metal4 111220 -298100 111440 -298100 1 COL_SEL[37]
port 10123 n
rlabel metal4 116630 -297200 116780 -297000 1 PIX_OUT38
port 10125 n
rlabel metal4 114220 -298100 114440 -298100 1 COL_SEL[38]
port 10126 n
rlabel metal4 119630 -297200 119780 -297000 1 PIX_OUT39
port 10128 n
rlabel metal4 117220 -298100 117440 -298100 1 COL_SEL[39]
port 10129 n
rlabel metal4 122630 -297200 122780 -297000 1 PIX_OUT40
port 10131 n
rlabel metal4 120220 -298100 120440 -298100 1 COL_SEL[40]
port 10132 n
rlabel metal4 125630 -297200 125780 -297000 1 PIX_OUT41
port 10134 n
rlabel metal4 123220 -298100 123440 -298100 1 COL_SEL[41]
port 10135 n
rlabel metal4 128630 -297200 128780 -297000 1 PIX_OUT42
port 10137 n
rlabel metal4 126220 -298100 126440 -298100 1 COL_SEL[42]
port 10138 n
rlabel metal4 131630 -297200 131780 -297000 1 PIX_OUT43
port 10140 n
rlabel metal4 129220 -298100 129440 -298100 1 COL_SEL[43]
port 10141 n
rlabel metal4 134630 -297200 134780 -297000 1 PIX_OUT44
port 10143 n
rlabel metal4 132220 -298100 132440 -298100 1 COL_SEL[44]
port 10144 n
rlabel metal4 137630 -297200 137780 -297000 1 PIX_OUT45
port 10146 n
rlabel metal4 135220 -298100 135440 -298100 1 COL_SEL[45]
port 10147 n
rlabel metal4 140630 -297200 140780 -297000 1 PIX_OUT46
port 10149 n
rlabel metal4 138220 -298100 138440 -298100 1 COL_SEL[46]
port 10150 n
rlabel metal4 143630 -297200 143780 -297000 1 PIX_OUT47
port 10152 n
rlabel metal4 141220 -298100 141440 -298100 1 COL_SEL[47]
port 10153 n
rlabel metal4 146630 -297200 146780 -297000 1 PIX_OUT48
port 10155 n
rlabel metal4 144220 -298100 144440 -298100 1 COL_SEL[48]
port 10156 n
rlabel metal4 149630 -297200 149780 -297000 1 PIX_OUT49
port 10158 n
rlabel metal4 147220 -298100 147440 -298100 1 COL_SEL[49]
port 10159 n
rlabel metal4 152630 -297200 152780 -297000 1 PIX_OUT50
port 10161 n
rlabel metal4 150220 -298100 150440 -298100 1 COL_SEL[50]
port 10162 n
rlabel metal4 155630 -297200 155780 -297000 1 PIX_OUT51
port 10164 n
rlabel metal4 153220 -298100 153440 -298100 1 COL_SEL[51]
port 10165 n
rlabel metal4 158630 -297200 158780 -297000 1 PIX_OUT52
port 10167 n
rlabel metal4 156220 -298100 156440 -298100 1 COL_SEL[52]
port 10168 n
rlabel metal4 161630 -297200 161780 -297000 1 PIX_OUT53
port 10170 n
rlabel metal4 159220 -298100 159440 -298100 1 COL_SEL[53]
port 10171 n
rlabel metal4 164630 -297200 164780 -297000 1 PIX_OUT54
port 10173 n
rlabel metal4 162220 -298100 162440 -298100 1 COL_SEL[54]
port 10174 n
rlabel metal4 167630 -297200 167780 -297000 1 PIX_OUT55
port 10176 n
rlabel metal4 165220 -298100 165440 -298100 1 COL_SEL[55]
port 10177 n
rlabel metal4 170630 -297200 170780 -297000 1 PIX_OUT56
port 10179 n
rlabel metal4 168220 -298100 168440 -298100 1 COL_SEL[56]
port 10180 n
rlabel metal4 173630 -297200 173780 -297000 1 PIX_OUT57
port 10182 n
rlabel metal4 171220 -298100 171440 -298100 1 COL_SEL[57]
port 10183 n
rlabel metal4 176630 -297200 176780 -297000 1 PIX_OUT58
port 10185 n
rlabel metal4 174220 -298100 174440 -298100 1 COL_SEL[58]
port 10186 n
rlabel metal4 179630 -297200 179780 -297000 1 PIX_OUT59
port 10188 n
rlabel metal4 177220 -298100 177440 -298100 1 COL_SEL[59]
port 10189 n
rlabel metal4 182630 -297200 182780 -297000 1 PIX_OUT60
port 10191 n
rlabel metal4 180220 -298100 180440 -298100 1 COL_SEL[60]
port 10192 n
rlabel metal4 185630 -297200 185780 -297000 1 PIX_OUT61
port 10194 n
rlabel metal4 183220 -298100 183440 -298100 1 COL_SEL[61]
port 10195 n
rlabel metal4 188630 -297200 188780 -297000 1 PIX_OUT62
port 10197 n
rlabel metal4 186220 -298100 186440 -298100 1 COL_SEL[62]
port 10198 n
rlabel metal4 191630 -297200 191780 -297000 1 PIX_OUT63
port 10200 n
rlabel metal4 189220 -298100 189440 -298100 1 COL_SEL[63]
port 10201 n
rlabel metal4 194630 -297200 194780 -297000 1 PIX_OUT64
port 10203 n
rlabel metal4 192220 -298100 192440 -298100 1 COL_SEL[64]
port 10204 n
rlabel metal4 197630 -297200 197780 -297000 1 PIX_OUT65
port 10206 n
rlabel metal4 195220 -298100 195440 -298100 1 COL_SEL[65]
port 10207 n
rlabel metal4 200630 -297200 200780 -297000 1 PIX_OUT66
port 10209 n
rlabel metal4 198220 -298100 198440 -298100 1 COL_SEL[66]
port 10210 n
rlabel metal4 203630 -297200 203780 -297000 1 PIX_OUT67
port 10212 n
rlabel metal4 201220 -298100 201440 -298100 1 COL_SEL[67]
port 10213 n
rlabel metal4 206630 -297200 206780 -297000 1 PIX_OUT68
port 10215 n
rlabel metal4 204220 -298100 204440 -298100 1 COL_SEL[68]
port 10216 n
rlabel metal4 209630 -297200 209780 -297000 1 PIX_OUT69
port 10218 n
rlabel metal4 207220 -298100 207440 -298100 1 COL_SEL[69]
port 10219 n
rlabel metal4 212630 -297200 212780 -297000 1 PIX_OUT70
port 10221 n
rlabel metal4 210220 -298100 210440 -298100 1 COL_SEL[70]
port 10222 n
rlabel metal4 215630 -297200 215780 -297000 1 PIX_OUT71
port 10224 n
rlabel metal4 213220 -298100 213440 -298100 1 COL_SEL[71]
port 10225 n
rlabel metal4 218630 -297200 218780 -297000 1 PIX_OUT72
port 10227 n
rlabel metal4 216220 -298100 216440 -298100 1 COL_SEL[72]
port 10228 n
rlabel metal4 221630 -297200 221780 -297000 1 PIX_OUT73
port 10230 n
rlabel metal4 219220 -298100 219440 -298100 1 COL_SEL[73]
port 10231 n
rlabel metal4 224630 -297200 224780 -297000 1 PIX_OUT74
port 10233 n
rlabel metal4 222220 -298100 222440 -298100 1 COL_SEL[74]
port 10234 n
rlabel metal4 227630 -297200 227780 -297000 1 PIX_OUT75
port 10236 n
rlabel metal4 225220 -298100 225440 -298100 1 COL_SEL[75]
port 10237 n
rlabel metal4 230630 -297200 230780 -297000 1 PIX_OUT76
port 10239 n
rlabel metal4 228220 -298100 228440 -298100 1 COL_SEL[76]
port 10240 n
rlabel metal4 233630 -297200 233780 -297000 1 PIX_OUT77
port 10242 n
rlabel metal4 231220 -298100 231440 -298100 1 COL_SEL[77]
port 10243 n
rlabel metal4 236630 -297200 236780 -297000 1 PIX_OUT78
port 10245 n
rlabel metal4 234220 -298100 234440 -298100 1 COL_SEL[78]
port 10246 n
rlabel metal4 239630 -297200 239780 -297000 1 PIX_OUT79
port 10248 n
rlabel metal4 237220 -298100 237440 -298100 1 COL_SEL[79]
port 10249 n
rlabel metal4 242630 -297200 242780 -297000 1 PIX_OUT80
port 10251 n
rlabel metal4 240220 -298100 240440 -298100 1 COL_SEL[80]
port 10252 n
rlabel metal4 245630 -297200 245780 -297000 1 PIX_OUT81
port 10254 n
rlabel metal4 243220 -298100 243440 -298100 1 COL_SEL[81]
port 10255 n
rlabel metal4 248630 -297200 248780 -297000 1 PIX_OUT82
port 10257 n
rlabel metal4 246220 -298100 246440 -298100 1 COL_SEL[82]
port 10258 n
rlabel metal4 251630 -297200 251780 -297000 1 PIX_OUT83
port 10260 n
rlabel metal4 249220 -298100 249440 -298100 1 COL_SEL[83]
port 10261 n
rlabel metal4 254630 -297200 254780 -297000 1 PIX_OUT84
port 10263 n
rlabel metal4 252220 -298100 252440 -298100 1 COL_SEL[84]
port 10264 n
rlabel metal4 257630 -297200 257780 -297000 1 PIX_OUT85
port 10266 n
rlabel metal4 255220 -298100 255440 -298100 1 COL_SEL[85]
port 10267 n
rlabel metal4 260630 -297200 260780 -297000 1 PIX_OUT86
port 10269 n
rlabel metal4 258220 -298100 258440 -298100 1 COL_SEL[86]
port 10270 n
rlabel metal4 263630 -297200 263780 -297000 1 PIX_OUT87
port 10272 n
rlabel metal4 261220 -298100 261440 -298100 1 COL_SEL[87]
port 10273 n
rlabel metal4 266630 -297200 266780 -297000 1 PIX_OUT88
port 10275 n
rlabel metal4 264220 -298100 264440 -298100 1 COL_SEL[88]
port 10276 n
rlabel metal4 269630 -297200 269780 -297000 1 PIX_OUT89
port 10278 n
rlabel metal4 267220 -298100 267440 -298100 1 COL_SEL[89]
port 10279 n
rlabel metal4 272630 -297200 272780 -297000 1 PIX_OUT90
port 10281 n
rlabel metal4 270220 -298100 270440 -298100 1 COL_SEL[90]
port 10282 n
rlabel metal4 275630 -297200 275780 -297000 1 PIX_OUT91
port 10284 n
rlabel metal4 273220 -298100 273440 -298100 1 COL_SEL[91]
port 10285 n
rlabel metal4 278630 -297200 278780 -297000 1 PIX_OUT92
port 10287 n
rlabel metal4 276220 -298100 276440 -298100 1 COL_SEL[92]
port 10288 n
rlabel metal4 281630 -297200 281780 -297000 1 PIX_OUT93
port 10290 n
rlabel metal4 279220 -298100 279440 -298100 1 COL_SEL[93]
port 10291 n
rlabel metal4 284630 -297200 284780 -297000 1 PIX_OUT94
port 10293 n
rlabel metal4 282220 -298100 282440 -298100 1 COL_SEL[94]
port 10294 n
rlabel metal4 287630 -297200 287780 -297000 1 PIX_OUT95
port 10296 n
rlabel metal4 285220 -298100 285440 -298100 1 COL_SEL[95]
port 10297 n
rlabel metal4 290630 -297200 290780 -297000 1 PIX_OUT96
port 10299 n
rlabel metal4 288220 -298100 288440 -298100 1 COL_SEL[96]
port 10300 n
rlabel metal4 293630 -297200 293780 -297000 1 PIX_OUT97
port 10302 n
rlabel metal4 291220 -298100 291440 -298100 1 COL_SEL[97]
port 10303 n
rlabel metal4 296630 -297200 296780 -297000 1 PIX_OUT98
port 10305 n
rlabel metal4 294220 -298100 294440 -298100 1 COL_SEL[98]
port 10306 n
rlabel metal4 299630 -297200 299780 -297000 1 PIX_OUT99
port 10308 n
rlabel metal2 299940 -298100 299940 -298100 1 ARRAY_OUT
port 10309 n
rlabel metal4 297220 -298100 297440 -298100 1 COL_SEL[99]
port 10310 n
<< end >>
