magic
tech sky130A
magscale 1 2
timestamp 1608345554
<< nwell >>
rect 3563 672 3809 1469
rect 3572 -1405 3818 -608
<< pwell >>
rect 3626 75 3793 614
rect 3626 67 3650 75
rect 3588 -550 3755 55
rect 5692 -3274 6579 -2442
<< metal1 >>
rect -186 1368 675 1370
rect -278 1185 675 1368
rect 2942 1190 4485 1375
rect -278 -1126 -97 1185
rect 6464 233 7624 257
rect 64 -203 7624 233
rect 7437 -224 7624 -203
rect -278 -1160 2469 -1126
rect 2915 -1160 4402 -1126
rect 4748 -1160 6543 -1121
rect -278 -1654 6543 -1160
rect -278 -1676 2469 -1654
rect -218 -1679 2469 -1676
rect 4748 -1679 6543 -1654
rect -222 -2258 -212 -2144
rect -56 -2157 -46 -2144
rect -56 -2173 1869 -2157
rect -56 -2236 2008 -2173
rect -56 -2251 1869 -2236
rect -56 -2258 -46 -2251
rect 5539 -2480 5549 -2266
rect 5751 -2480 5761 -2266
rect 1848 -3022 5350 -2683
rect 7437 -3022 7626 -224
rect 1834 -3211 7626 -3022
<< via1 >>
rect -212 -2258 -56 -2144
rect 5549 -2480 5751 -2266
<< metal2 >>
rect 6 722 96 732
rect 6 588 96 598
rect 7359 539 7473 549
rect 7332 401 7359 493
rect 7332 391 7473 401
rect -208 -338 -88 -328
rect -208 -498 -88 -488
rect -204 -692 -96 -498
rect -203 -2134 -96 -692
rect 7332 -717 7465 391
rect -212 -2144 -56 -2134
rect -212 -2268 -56 -2258
rect 5549 -2266 5751 -2256
rect -203 -2272 -96 -2268
rect 5549 -2490 5751 -2480
rect 6358 -2496 7323 -2266
<< via2 >>
rect 6 598 96 722
rect 7359 401 7473 539
rect -208 -488 -88 -338
rect 5574 -2470 5724 -2286
<< metal3 >>
rect -10 732 116 926
rect -296 722 116 732
rect -296 610 6 722
rect -10 598 6 610
rect 96 598 116 722
rect -10 442 116 598
rect 7349 539 7483 544
rect 7349 401 7359 539
rect 7473 401 7483 539
rect 7349 396 7483 401
rect -218 -338 -78 -333
rect -218 -488 -208 -338
rect -88 -488 -78 -338
rect -218 -493 -78 -488
rect 5550 -2286 5750 -2266
rect 5550 -2337 5574 -2286
rect 5415 -2447 5574 -2337
rect 5550 -2470 5574 -2447
rect 5724 -2470 5750 -2286
rect 5550 -2480 5750 -2470
use inverter_out  inverter_out_0
timestamp 1608344763
transform 1 0 5270 0 1 -3032
box 408 -247 1342 1692
use freq_div  freq_div_2
timestamp 1608334096
transform -1 0 2955 0 -1 49
box -710 -10 3151 1455
use freq_div  freq_div_3
timestamp 1608334096
transform -1 0 6671 0 -1 54
box -710 -10 3151 1455
use freq_div  freq_div_1
timestamp 1608334096
transform 1 0 4426 0 1 15
box -710 -10 3151 1455
use freq_div  freq_div_0
timestamp 1608334096
transform 1 0 710 0 1 10
box -710 -10 3151 1455
use freq_div  freq_div_4
timestamp 1608334096
transform 1 0 2484 0 1 -2854
box -710 -10 3151 1455
<< labels >>
rlabel metal3 -296 610 116 732 1 in
rlabel space 1904 -2801 7626 -2612 1 vss
rlabel space 2942 1190 7273 1375 1 vdd
rlabel metal2 7093 -2496 7323 -2266 1 out
<< end >>
