magic
tech sky130A
magscale 1 2
timestamp 1654708041
<< error_p >>
rect 159959 -136004 159993 -135428
rect 165297 -136005 165331 -135429
rect 165415 -136005 165449 -135429
rect 165533 -136005 165567 -135429
rect 165651 -136005 165685 -135429
rect 165769 -136005 165803 -135429
rect 165887 -136005 165921 -135429
rect 166005 -136005 166039 -135429
rect 166123 -136005 166157 -135429
rect 166241 -136005 166275 -135429
rect 166359 -136005 166393 -135429
rect 166477 -136005 166511 -135429
rect 166595 -136005 166629 -135429
rect 166713 -136005 166747 -135429
rect 166831 -136005 166865 -135429
rect 166949 -136005 166983 -135429
rect 167067 -136005 167101 -135429
rect 167185 -136005 167219 -135429
rect 167303 -136005 167337 -135429
rect 167421 -136005 167455 -135429
rect 167539 -136005 167573 -135429
rect 167657 -136005 167691 -135429
rect 167775 -136005 167809 -135429
rect 167893 -136005 167927 -135429
rect 168011 -136005 168045 -135429
rect 169420 -136005 169454 -135429
rect 169538 -136005 169572 -135429
rect 169656 -136005 169690 -135429
rect 169774 -136005 169808 -135429
rect 169892 -136005 169926 -135429
rect 170010 -136005 170044 -135429
rect 170128 -136005 170162 -135429
rect 170246 -136005 170280 -135429
rect 170364 -136005 170398 -135429
rect 170482 -136005 170516 -135429
rect 170600 -136005 170634 -135429
rect 170718 -136005 170752 -135429
rect 170836 -136005 170870 -135429
rect 170954 -136005 170988 -135429
rect 171072 -136005 171106 -135429
rect 171190 -136005 171224 -135429
rect 171308 -136005 171342 -135429
rect 171426 -136005 171460 -135429
rect 171544 -136005 171578 -135429
rect 171662 -136005 171696 -135429
rect 171780 -136005 171814 -135429
rect 171898 -136005 171932 -135429
rect 172016 -136005 172050 -135429
rect 172134 -136005 172168 -135429
rect 173543 -136005 173577 -135429
rect 173661 -136005 173695 -135429
rect 173779 -136005 173813 -135429
rect 173897 -136005 173931 -135429
rect 174015 -136005 174049 -135429
rect 174133 -136005 174167 -135429
rect 174251 -136005 174285 -135429
rect 174369 -136005 174403 -135429
rect 174487 -136005 174521 -135429
rect 174605 -136005 174639 -135429
rect 174723 -136005 174757 -135429
rect 174841 -136005 174875 -135429
rect 174959 -136005 174993 -135429
rect 175077 -136005 175111 -135429
rect 175195 -136005 175229 -135429
rect 175313 -136005 175347 -135429
rect 175431 -136005 175465 -135429
rect 175549 -136005 175583 -135429
rect 175667 -136005 175701 -135429
rect 175785 -136005 175819 -135429
rect 175903 -136005 175937 -135429
rect 176021 -136005 176055 -135429
rect 176139 -136005 176173 -135429
rect 176257 -136005 176291 -135429
rect 157353 -136764 163323 -136730
rect 157257 -138436 157291 -136826
rect 157371 -137501 157405 -136925
rect 157489 -137501 157523 -136925
rect 157607 -137501 157641 -136925
rect 157725 -137501 157759 -136925
rect 157843 -137501 157877 -136925
rect 157961 -137501 157995 -136925
rect 158079 -137501 158113 -136925
rect 158197 -137501 158231 -136925
rect 158315 -137501 158349 -136925
rect 158433 -137501 158467 -136925
rect 158551 -137501 158585 -136925
rect 158669 -137501 158703 -136925
rect 158787 -137501 158821 -136925
rect 158905 -137501 158939 -136925
rect 159023 -137501 159057 -136925
rect 159141 -137501 159175 -136925
rect 159259 -137501 159293 -136925
rect 159377 -137501 159411 -136925
rect 159495 -137501 159529 -136925
rect 159613 -137501 159647 -136925
rect 159731 -137501 159765 -136925
rect 159849 -137501 159883 -136925
rect 159967 -137501 160001 -136925
rect 160085 -137501 160119 -136925
rect 160203 -137501 160237 -136925
rect 160321 -137501 160355 -136925
rect 160439 -137501 160473 -136925
rect 160557 -137501 160591 -136925
rect 160675 -137501 160709 -136925
rect 160793 -137501 160827 -136925
rect 160911 -137501 160945 -136925
rect 161029 -137501 161063 -136925
rect 161147 -137501 161181 -136925
rect 161265 -137501 161299 -136925
rect 161383 -137501 161417 -136925
rect 161501 -137501 161535 -136925
rect 161619 -137501 161653 -136925
rect 161737 -137501 161771 -136925
rect 161855 -137501 161889 -136925
rect 161973 -137501 162007 -136925
rect 162091 -137501 162125 -136925
rect 162209 -137501 162243 -136925
rect 162327 -137501 162361 -136925
rect 162445 -137501 162479 -136925
rect 162563 -137501 162597 -136925
rect 162681 -137501 162715 -136925
rect 162799 -137501 162833 -136925
rect 162917 -137501 162951 -136925
rect 163035 -137501 163069 -136925
rect 163153 -137501 163187 -136925
rect 163271 -137501 163305 -136925
rect 157371 -138337 157405 -137761
rect 157489 -138337 157523 -137761
rect 157607 -138337 157641 -137761
rect 157725 -138337 157759 -137761
rect 157843 -138337 157877 -137761
rect 157961 -138337 157995 -137761
rect 158079 -138337 158113 -137761
rect 158197 -138337 158231 -137761
rect 158315 -138337 158349 -137761
rect 158433 -138337 158467 -137761
rect 158551 -138337 158585 -137761
rect 158669 -138337 158703 -137761
rect 158787 -138337 158821 -137761
rect 158905 -138337 158939 -137761
rect 159023 -138337 159057 -137761
rect 159141 -138337 159175 -137761
rect 159259 -138337 159293 -137761
rect 159377 -138337 159411 -137761
rect 159495 -138337 159529 -137761
rect 159613 -138337 159647 -137761
rect 159731 -138337 159765 -137761
rect 159849 -138337 159883 -137761
rect 159967 -138337 160001 -137761
rect 160085 -138337 160119 -137761
rect 160203 -138337 160237 -137761
rect 160321 -138337 160355 -137761
rect 160439 -138337 160473 -137761
rect 160557 -138337 160591 -137761
rect 160675 -138337 160709 -137761
rect 160793 -138337 160827 -137761
rect 160911 -138337 160945 -137761
rect 161029 -138337 161063 -137761
rect 161147 -138337 161181 -137761
rect 161265 -138337 161299 -137761
rect 161383 -138337 161417 -137761
rect 161501 -138337 161535 -137761
rect 161619 -138337 161653 -137761
rect 161737 -138337 161771 -137761
rect 161855 -138337 161889 -137761
rect 161973 -138337 162007 -137761
rect 162091 -138337 162125 -137761
rect 162209 -138337 162243 -137761
rect 162327 -138337 162361 -137761
rect 162445 -138337 162479 -137761
rect 162563 -138337 162597 -137761
rect 162681 -138337 162715 -137761
rect 162799 -138337 162833 -137761
rect 162917 -138337 162951 -137761
rect 163035 -138337 163069 -137761
rect 163153 -138337 163187 -137761
rect 163271 -138337 163305 -137761
rect 163385 -138436 163419 -136826
rect 165061 -136841 165095 -136265
rect 165179 -136841 165213 -136265
rect 165297 -136841 165331 -136265
rect 165415 -136841 165449 -136265
rect 165533 -136841 165567 -136265
rect 165651 -136841 165685 -136265
rect 165769 -136841 165803 -136265
rect 165887 -136841 165921 -136265
rect 166005 -136841 166039 -136265
rect 166123 -136841 166157 -136265
rect 166241 -136841 166275 -136265
rect 166359 -136841 166393 -136265
rect 166477 -136841 166511 -136265
rect 166595 -136841 166629 -136265
rect 166713 -136841 166747 -136265
rect 166831 -136841 166865 -136265
rect 166949 -136841 166983 -136265
rect 167067 -136841 167101 -136265
rect 167185 -136841 167219 -136265
rect 167303 -136841 167337 -136265
rect 167421 -136841 167455 -136265
rect 167539 -136841 167573 -136265
rect 167657 -136841 167691 -136265
rect 167775 -136841 167809 -136265
rect 167893 -136841 167927 -136265
rect 168011 -136841 168045 -136265
rect 169184 -136841 169218 -136265
rect 169302 -136841 169336 -136265
rect 169420 -136841 169454 -136265
rect 169538 -136841 169572 -136265
rect 169656 -136841 169690 -136265
rect 169774 -136841 169808 -136265
rect 169892 -136841 169926 -136265
rect 170010 -136841 170044 -136265
rect 170128 -136841 170162 -136265
rect 170246 -136841 170280 -136265
rect 170364 -136841 170398 -136265
rect 170482 -136841 170516 -136265
rect 170600 -136841 170634 -136265
rect 170718 -136841 170752 -136265
rect 170836 -136841 170870 -136265
rect 170954 -136841 170988 -136265
rect 171072 -136841 171106 -136265
rect 171190 -136841 171224 -136265
rect 171308 -136841 171342 -136265
rect 171426 -136841 171460 -136265
rect 171544 -136841 171578 -136265
rect 171662 -136841 171696 -136265
rect 171780 -136841 171814 -136265
rect 171898 -136841 171932 -136265
rect 172016 -136841 172050 -136265
rect 172134 -136841 172168 -136265
rect 173307 -136841 173341 -136265
rect 173425 -136841 173459 -136265
rect 173543 -136841 173577 -136265
rect 173661 -136841 173695 -136265
rect 173779 -136841 173813 -136265
rect 173897 -136841 173931 -136265
rect 174015 -136841 174049 -136265
rect 174133 -136841 174167 -136265
rect 174251 -136841 174285 -136265
rect 174369 -136841 174403 -136265
rect 174487 -136841 174521 -136265
rect 174605 -136841 174639 -136265
rect 174723 -136841 174757 -136265
rect 174841 -136841 174875 -136265
rect 174959 -136841 174993 -136265
rect 175077 -136841 175111 -136265
rect 175195 -136841 175229 -136265
rect 175313 -136841 175347 -136265
rect 175431 -136841 175465 -136265
rect 175549 -136841 175583 -136265
rect 175667 -136841 175701 -136265
rect 175785 -136841 175819 -136265
rect 175903 -136841 175937 -136265
rect 176021 -136841 176055 -136265
rect 176139 -136841 176173 -136265
rect 176257 -136841 176291 -136265
rect 157353 -138532 163323 -138498
rect 157353 -138814 163323 -138780
rect 157257 -140486 157291 -138876
rect 157371 -139551 157405 -138975
rect 157489 -139551 157523 -138975
rect 157607 -139551 157641 -138975
rect 157725 -139551 157759 -138975
rect 157843 -139551 157877 -138975
rect 157961 -139551 157995 -138975
rect 158079 -139551 158113 -138975
rect 158197 -139551 158231 -138975
rect 158315 -139551 158349 -138975
rect 158433 -139551 158467 -138975
rect 158551 -139551 158585 -138975
rect 158669 -139551 158703 -138975
rect 158787 -139551 158821 -138975
rect 158905 -139551 158939 -138975
rect 159023 -139551 159057 -138975
rect 159141 -139551 159175 -138975
rect 159259 -139551 159293 -138975
rect 159377 -139551 159411 -138975
rect 159495 -139551 159529 -138975
rect 159613 -139551 159647 -138975
rect 159731 -139551 159765 -138975
rect 159849 -139551 159883 -138975
rect 159967 -139551 160001 -138975
rect 160085 -139551 160119 -138975
rect 160203 -139551 160237 -138975
rect 160321 -139551 160355 -138975
rect 160439 -139551 160473 -138975
rect 160557 -139551 160591 -138975
rect 160675 -139551 160709 -138975
rect 160793 -139551 160827 -138975
rect 160911 -139551 160945 -138975
rect 161029 -139551 161063 -138975
rect 161147 -139551 161181 -138975
rect 161265 -139551 161299 -138975
rect 161383 -139551 161417 -138975
rect 161501 -139551 161535 -138975
rect 161619 -139551 161653 -138975
rect 161737 -139551 161771 -138975
rect 161855 -139551 161889 -138975
rect 161973 -139551 162007 -138975
rect 162091 -139551 162125 -138975
rect 162209 -139551 162243 -138975
rect 162327 -139551 162361 -138975
rect 162445 -139551 162479 -138975
rect 162563 -139551 162597 -138975
rect 162681 -139551 162715 -138975
rect 162799 -139551 162833 -138975
rect 162917 -139551 162951 -138975
rect 163035 -139551 163069 -138975
rect 163153 -139551 163187 -138975
rect 163271 -139551 163305 -138975
rect 157371 -140387 157405 -139811
rect 157489 -140387 157523 -139811
rect 157607 -140387 157641 -139811
rect 157725 -140387 157759 -139811
rect 157843 -140387 157877 -139811
rect 157961 -140387 157995 -139811
rect 158079 -140387 158113 -139811
rect 158197 -140387 158231 -139811
rect 158315 -140387 158349 -139811
rect 158433 -140387 158467 -139811
rect 158551 -140387 158585 -139811
rect 158669 -140387 158703 -139811
rect 158787 -140387 158821 -139811
rect 158905 -140387 158939 -139811
rect 159023 -140387 159057 -139811
rect 159141 -140387 159175 -139811
rect 159259 -140387 159293 -139811
rect 159377 -140387 159411 -139811
rect 159495 -140387 159529 -139811
rect 159613 -140387 159647 -139811
rect 159731 -140387 159765 -139811
rect 159849 -140387 159883 -139811
rect 159967 -140387 160001 -139811
rect 160085 -140387 160119 -139811
rect 160203 -140387 160237 -139811
rect 160321 -140387 160355 -139811
rect 160439 -140387 160473 -139811
rect 160557 -140387 160591 -139811
rect 160675 -140387 160709 -139811
rect 160793 -140387 160827 -139811
rect 160911 -140387 160945 -139811
rect 161029 -140387 161063 -139811
rect 161147 -140387 161181 -139811
rect 161265 -140387 161299 -139811
rect 161383 -140387 161417 -139811
rect 161501 -140387 161535 -139811
rect 161619 -140387 161653 -139811
rect 161737 -140387 161771 -139811
rect 161855 -140387 161889 -139811
rect 161973 -140387 162007 -139811
rect 162091 -140387 162125 -139811
rect 162209 -140387 162243 -139811
rect 162327 -140387 162361 -139811
rect 162445 -140387 162479 -139811
rect 162563 -140387 162597 -139811
rect 162681 -140387 162715 -139811
rect 162799 -140387 162833 -139811
rect 162917 -140387 162951 -139811
rect 163035 -140387 163069 -139811
rect 163153 -140387 163187 -139811
rect 163271 -140387 163305 -139811
rect 163385 -140486 163419 -138876
rect 157353 -140582 163323 -140548
rect 157353 -140864 163323 -140830
rect 157257 -142536 157291 -140926
rect 157371 -141601 157405 -141025
rect 157489 -141601 157523 -141025
rect 157607 -141601 157641 -141025
rect 157725 -141601 157759 -141025
rect 157843 -141601 157877 -141025
rect 157961 -141601 157995 -141025
rect 158079 -141601 158113 -141025
rect 158197 -141601 158231 -141025
rect 158315 -141601 158349 -141025
rect 158433 -141601 158467 -141025
rect 158551 -141601 158585 -141025
rect 158669 -141601 158703 -141025
rect 158787 -141601 158821 -141025
rect 158905 -141601 158939 -141025
rect 159023 -141601 159057 -141025
rect 159141 -141601 159175 -141025
rect 159259 -141601 159293 -141025
rect 159377 -141601 159411 -141025
rect 159495 -141601 159529 -141025
rect 159613 -141601 159647 -141025
rect 159731 -141601 159765 -141025
rect 159849 -141601 159883 -141025
rect 159967 -141601 160001 -141025
rect 160085 -141601 160119 -141025
rect 160203 -141601 160237 -141025
rect 160321 -141601 160355 -141025
rect 160439 -141601 160473 -141025
rect 160557 -141601 160591 -141025
rect 160675 -141601 160709 -141025
rect 160793 -141601 160827 -141025
rect 160911 -141601 160945 -141025
rect 161029 -141601 161063 -141025
rect 161147 -141601 161181 -141025
rect 161265 -141601 161299 -141025
rect 161383 -141601 161417 -141025
rect 161501 -141601 161535 -141025
rect 161619 -141601 161653 -141025
rect 161737 -141601 161771 -141025
rect 161855 -141601 161889 -141025
rect 161973 -141601 162007 -141025
rect 162091 -141601 162125 -141025
rect 162209 -141601 162243 -141025
rect 162327 -141601 162361 -141025
rect 162445 -141601 162479 -141025
rect 162563 -141601 162597 -141025
rect 162681 -141601 162715 -141025
rect 162799 -141601 162833 -141025
rect 162917 -141601 162951 -141025
rect 163035 -141601 163069 -141025
rect 163153 -141601 163187 -141025
rect 163271 -141601 163305 -141025
rect 157371 -142437 157405 -141861
rect 157489 -142437 157523 -141861
rect 157607 -142437 157641 -141861
rect 157725 -142437 157759 -141861
rect 157843 -142437 157877 -141861
rect 157961 -142437 157995 -141861
rect 158079 -142437 158113 -141861
rect 158197 -142437 158231 -141861
rect 158315 -142437 158349 -141861
rect 158433 -142437 158467 -141861
rect 158551 -142437 158585 -141861
rect 158669 -142437 158703 -141861
rect 158787 -142437 158821 -141861
rect 158905 -142437 158939 -141861
rect 159023 -142437 159057 -141861
rect 159141 -142437 159175 -141861
rect 159259 -142437 159293 -141861
rect 159377 -142437 159411 -141861
rect 159495 -142437 159529 -141861
rect 159613 -142437 159647 -141861
rect 159731 -142437 159765 -141861
rect 159849 -142437 159883 -141861
rect 159967 -142437 160001 -141861
rect 160085 -142437 160119 -141861
rect 160203 -142437 160237 -141861
rect 160321 -142437 160355 -141861
rect 160439 -142437 160473 -141861
rect 160557 -142437 160591 -141861
rect 160675 -142437 160709 -141861
rect 160793 -142437 160827 -141861
rect 160911 -142437 160945 -141861
rect 161029 -142437 161063 -141861
rect 161147 -142437 161181 -141861
rect 161265 -142437 161299 -141861
rect 161383 -142437 161417 -141861
rect 161501 -142437 161535 -141861
rect 161619 -142437 161653 -141861
rect 161737 -142437 161771 -141861
rect 161855 -142437 161889 -141861
rect 161973 -142437 162007 -141861
rect 162091 -142437 162125 -141861
rect 162209 -142437 162243 -141861
rect 162327 -142437 162361 -141861
rect 162445 -142437 162479 -141861
rect 162563 -142437 162597 -141861
rect 162681 -142437 162715 -141861
rect 162799 -142437 162833 -141861
rect 162917 -142437 162951 -141861
rect 163035 -142437 163069 -141861
rect 163153 -142437 163187 -141861
rect 163271 -142437 163305 -141861
rect 163385 -142536 163419 -140926
rect 157353 -142632 163323 -142598
rect 157607 -143651 157641 -143075
rect 157725 -143651 157759 -143075
rect 157843 -143651 157877 -143075
rect 157961 -143651 157995 -143075
rect 158079 -143651 158113 -143075
rect 158197 -143651 158231 -143075
rect 158315 -143651 158349 -143075
rect 158433 -143651 158467 -143075
rect 158551 -143651 158585 -143075
rect 158669 -143651 158703 -143075
rect 158787 -143651 158821 -143075
rect 158905 -143651 158939 -143075
rect 159023 -143651 159057 -143075
rect 159141 -143651 159175 -143075
rect 159259 -143651 159293 -143075
rect 159377 -143651 159411 -143075
rect 159495 -143651 159529 -143075
rect 159613 -143651 159647 -143075
rect 159731 -143651 159765 -143075
rect 159849 -143651 159883 -143075
rect 159967 -143651 160001 -143075
rect 160085 -143651 160119 -143075
rect 160203 -143651 160237 -143075
rect 160321 -143651 160355 -143075
rect 160439 -143651 160473 -143075
rect 160557 -143651 160591 -143075
rect 160675 -143651 160709 -143075
rect 160793 -143651 160827 -143075
rect 160911 -143651 160945 -143075
rect 161029 -143651 161063 -143075
rect 161147 -143651 161181 -143075
rect 161265 -143651 161299 -143075
rect 161383 -143651 161417 -143075
rect 161501 -143651 161535 -143075
rect 161619 -143651 161653 -143075
rect 161737 -143651 161771 -143075
rect 161855 -143651 161889 -143075
rect 161973 -143651 162007 -143075
rect 162091 -143651 162125 -143075
rect 162209 -143651 162243 -143075
rect 162327 -143651 162361 -143075
rect 162445 -143651 162479 -143075
rect 162563 -143651 162597 -143075
rect 162681 -143651 162715 -143075
rect 162799 -143651 162833 -143075
rect 162917 -143651 162951 -143075
rect 163035 -143651 163069 -143075
rect 163153 -143651 163187 -143075
rect 163271 -143651 163305 -143075
rect 157371 -144487 157405 -143911
rect 157489 -144487 157523 -143911
rect 157607 -144487 157641 -143911
rect 157725 -144487 157759 -143911
rect 157843 -144487 157877 -143911
rect 157961 -144487 157995 -143911
rect 158079 -144487 158113 -143911
rect 158197 -144487 158231 -143911
rect 158315 -144487 158349 -143911
rect 158433 -144487 158467 -143911
rect 158551 -144487 158585 -143911
rect 158669 -144487 158703 -143911
rect 158787 -144487 158821 -143911
rect 158905 -144487 158939 -143911
rect 159023 -144487 159057 -143911
rect 159141 -144487 159175 -143911
rect 159259 -144487 159293 -143911
rect 159377 -144487 159411 -143911
rect 159495 -144487 159529 -143911
rect 159613 -144487 159647 -143911
rect 159731 -144487 159765 -143911
rect 159849 -144487 159883 -143911
rect 159967 -144487 160001 -143911
rect 160085 -144487 160119 -143911
rect 160203 -144487 160237 -143911
rect 160321 -144487 160355 -143911
rect 160439 -144487 160473 -143911
rect 160557 -144487 160591 -143911
rect 160675 -144487 160709 -143911
rect 160793 -144487 160827 -143911
rect 160911 -144487 160945 -143911
rect 161029 -144487 161063 -143911
rect 161147 -144487 161181 -143911
rect 161265 -144487 161299 -143911
rect 161383 -144487 161417 -143911
rect 161501 -144487 161535 -143911
rect 161619 -144487 161653 -143911
rect 161737 -144487 161771 -143911
rect 161855 -144487 161889 -143911
rect 161973 -144487 162007 -143911
rect 162091 -144487 162125 -143911
rect 162209 -144487 162243 -143911
rect 162327 -144487 162361 -143911
rect 162445 -144487 162479 -143911
rect 162563 -144487 162597 -143911
rect 162681 -144487 162715 -143911
rect 162799 -144487 162833 -143911
rect 162917 -144487 162951 -143911
rect 163035 -144487 163069 -143911
rect 163153 -144487 163187 -143911
rect 163271 -144487 163305 -143911
rect 158673 -145894 158707 -145318
rect 158791 -145894 158825 -145318
rect 158909 -145894 158943 -145318
rect 159027 -145894 159061 -145318
rect 159145 -145894 159179 -145318
rect 159263 -145894 159297 -145318
rect 159381 -145894 159415 -145318
rect 159499 -145894 159533 -145318
rect 159617 -145894 159651 -145318
rect 159735 -145894 159769 -145318
rect 159853 -145894 159887 -145318
rect 159971 -145894 160005 -145318
rect 160089 -145894 160123 -145318
rect 160207 -145894 160241 -145318
rect 160435 -145894 160469 -145318
rect 160553 -145894 160587 -145318
rect 160671 -145894 160705 -145318
rect 160789 -145894 160823 -145318
rect 160907 -145894 160941 -145318
rect 161025 -145894 161059 -145318
rect 161143 -145894 161177 -145318
rect 161261 -145894 161295 -145318
rect 161379 -145894 161413 -145318
rect 161497 -145894 161531 -145318
rect 161615 -145894 161649 -145318
rect 161733 -145894 161767 -145318
rect 161851 -145894 161885 -145318
rect 161969 -145894 162003 -145318
rect 162087 -145894 162121 -145318
rect 162205 -145894 162239 -145318
rect 163298 -145696 163332 -145390
rect 163412 -145606 163446 -145480
rect 163500 -145606 163534 -145480
rect 163614 -145696 163648 -145390
rect 163728 -145606 163762 -145480
rect 163816 -145606 163850 -145480
rect 163930 -145696 163964 -145390
rect 164044 -145606 164078 -145480
rect 164132 -145606 164166 -145480
rect 164246 -145696 164280 -145390
rect 164360 -145606 164394 -145480
rect 164448 -145606 164482 -145480
rect 164562 -145696 164596 -145390
rect 164676 -145606 164710 -145480
rect 164764 -145606 164798 -145480
rect 164878 -145696 164912 -145390
rect 158437 -146712 158471 -146136
rect 158555 -146712 158589 -146136
rect 158673 -146712 158707 -146136
rect 158791 -146712 158825 -146136
rect 158909 -146712 158943 -146136
rect 159027 -146712 159061 -146136
rect 159145 -146712 159179 -146136
rect 159263 -146712 159297 -146136
rect 159381 -146712 159415 -146136
rect 159499 -146712 159533 -146136
rect 159617 -146712 159651 -146136
rect 159735 -146712 159769 -146136
rect 159853 -146712 159887 -146136
rect 159971 -146712 160005 -146136
rect 160089 -146712 160123 -146136
rect 160207 -146712 160241 -146136
rect 160435 -146712 160469 -146136
rect 160553 -146712 160587 -146136
rect 160671 -146712 160705 -146136
rect 160789 -146712 160823 -146136
rect 160907 -146712 160941 -146136
rect 161025 -146712 161059 -146136
rect 161143 -146712 161177 -146136
rect 161261 -146712 161295 -146136
rect 161379 -146712 161413 -146136
rect 161497 -146712 161531 -146136
rect 161615 -146712 161649 -146136
rect 161733 -146712 161767 -146136
rect 161851 -146712 161885 -146136
rect 161969 -146712 162003 -146136
rect 162087 -146712 162121 -146136
rect 162205 -146712 162239 -146136
rect 165095 -146194 165129 -145318
rect 165243 -146194 165277 -145318
rect 165391 -146194 165425 -145318
rect 165539 -146194 165573 -145318
rect 165687 -146194 165721 -145318
rect 165835 -146194 165869 -145318
rect 165983 -146194 166017 -145318
rect 166131 -146194 166165 -145318
rect 166279 -146194 166313 -145318
rect 166427 -146194 166461 -145318
rect 166575 -146194 166609 -145318
rect 166723 -146194 166757 -145318
rect 166871 -146194 166905 -145318
rect 167019 -146194 167053 -145318
rect 167167 -146194 167201 -145318
rect 167315 -146194 167349 -145318
rect 167463 -146194 167497 -145318
rect 167611 -146194 167645 -145318
rect 167759 -146194 167793 -145318
rect 167907 -146194 167941 -145318
rect 168055 -146194 168089 -145318
rect 168203 -146194 168237 -145318
rect 168351 -146194 168385 -145318
rect 168499 -146194 168533 -145318
rect 168647 -146194 168681 -145318
rect 168795 -146194 168829 -145318
rect 168943 -146194 168977 -145318
rect 169091 -146194 169125 -145318
rect 169239 -146194 169273 -145318
rect 169387 -146194 169421 -145318
rect 169535 -146194 169569 -145318
rect 169683 -146194 169717 -145318
rect 169831 -146194 169865 -145318
rect 169979 -146194 170013 -145318
rect 170127 -146194 170161 -145318
rect 170275 -146194 170309 -145318
rect 170423 -146194 170457 -145318
rect 170571 -146194 170605 -145318
rect 170719 -146194 170753 -145318
rect 170867 -146194 170901 -145318
rect 171015 -146194 171049 -145318
rect 171163 -146194 171197 -145318
rect 171311 -146194 171345 -145318
rect 171459 -146194 171493 -145318
rect 171607 -146194 171641 -145318
rect 171755 -146194 171789 -145318
rect 171903 -146194 171937 -145318
rect 172051 -146194 172085 -145318
rect 172199 -146194 172233 -145318
rect 172347 -146194 172381 -145318
rect 172495 -146194 172529 -145318
rect 172643 -146194 172677 -145318
rect 172791 -146194 172825 -145318
rect 172939 -146194 172973 -145318
rect 173087 -146194 173121 -145318
rect 173235 -146194 173269 -145318
rect 173383 -146194 173417 -145318
rect 173531 -146194 173565 -145318
rect 173679 -146194 173713 -145318
rect 173827 -146194 173861 -145318
rect 173975 -146194 174009 -145318
rect 174123 -146194 174157 -145318
rect 174271 -146194 174305 -145318
rect 174419 -146194 174453 -145318
rect 174567 -146194 174601 -145318
rect 174715 -146194 174749 -145318
rect 174863 -146194 174897 -145318
rect 175011 -146194 175045 -145318
rect 175159 -146194 175193 -145318
rect 175307 -146194 175341 -145318
rect 175455 -146194 175489 -145318
rect 175603 -146194 175637 -145318
rect 175751 -146194 175785 -145318
rect 175899 -146194 175933 -145318
rect 176195 -146194 176229 -145318
rect 165305 -146278 165363 -146244
rect 165453 -146278 165511 -146244
rect 165601 -146278 165659 -146244
rect 165749 -146278 165807 -146244
rect 165897 -146278 165955 -146244
rect 166045 -146278 166103 -146244
rect 166193 -146278 166251 -146244
rect 166341 -146278 166399 -146244
rect 166489 -146278 166547 -146244
rect 166637 -146278 166695 -146244
rect 166785 -146278 166843 -146244
rect 166933 -146278 166991 -146244
rect 167081 -146278 167139 -146244
rect 167229 -146278 167287 -146244
rect 167377 -146278 167435 -146244
rect 167525 -146278 167583 -146244
rect 167673 -146278 167731 -146244
rect 167821 -146278 167879 -146244
rect 167969 -146278 168027 -146244
rect 168117 -146278 168175 -146244
rect 168265 -146278 168323 -146244
rect 168413 -146278 168471 -146244
rect 168561 -146278 168619 -146244
rect 168709 -146278 168767 -146244
rect 168857 -146278 168915 -146244
rect 169005 -146278 169063 -146244
rect 169153 -146278 169211 -146244
rect 169301 -146278 169359 -146244
rect 169449 -146278 169507 -146244
rect 169597 -146278 169655 -146244
rect 169745 -146278 169803 -146244
rect 169893 -146278 169951 -146244
rect 170041 -146278 170099 -146244
rect 170189 -146278 170247 -146244
rect 170337 -146278 170395 -146244
rect 170485 -146278 170543 -146244
rect 170633 -146278 170691 -146244
rect 170781 -146278 170839 -146244
rect 170929 -146278 170987 -146244
rect 171077 -146278 171135 -146244
rect 171225 -146278 171283 -146244
rect 171373 -146278 171431 -146244
rect 171521 -146278 171579 -146244
rect 171669 -146278 171727 -146244
rect 171817 -146278 171875 -146244
rect 171965 -146278 172023 -146244
rect 172113 -146278 172171 -146244
rect 172261 -146278 172319 -146244
rect 172409 -146278 172467 -146244
rect 172557 -146278 172615 -146244
rect 172705 -146278 172763 -146244
rect 172853 -146278 172911 -146244
rect 173001 -146278 173059 -146244
rect 173149 -146278 173207 -146244
rect 173297 -146278 173355 -146244
rect 173445 -146278 173503 -146244
rect 173593 -146278 173651 -146244
rect 173741 -146278 173799 -146244
rect 173889 -146278 173947 -146244
rect 174037 -146278 174095 -146244
rect 174185 -146278 174243 -146244
rect 174333 -146278 174391 -146244
rect 174481 -146278 174539 -146244
rect 174629 -146278 174687 -146244
rect 174777 -146278 174835 -146244
rect 174925 -146278 174983 -146244
rect 175073 -146278 175131 -146244
rect 175221 -146278 175279 -146244
rect 175369 -146278 175427 -146244
rect 175517 -146278 175575 -146244
rect 175665 -146278 175723 -146244
rect 175813 -146278 175871 -146244
rect 175961 -146278 176019 -146244
rect 176109 -146278 176167 -146244
rect 165305 -146386 165363 -146352
rect 165453 -146386 165511 -146352
rect 165601 -146386 165659 -146352
rect 165749 -146386 165807 -146352
rect 165897 -146386 165955 -146352
rect 166045 -146386 166103 -146352
rect 166193 -146386 166251 -146352
rect 166341 -146386 166399 -146352
rect 166489 -146386 166547 -146352
rect 166637 -146386 166695 -146352
rect 166785 -146386 166843 -146352
rect 166933 -146386 166991 -146352
rect 167081 -146386 167139 -146352
rect 167229 -146386 167287 -146352
rect 167377 -146386 167435 -146352
rect 167525 -146386 167583 -146352
rect 167673 -146386 167731 -146352
rect 167821 -146386 167879 -146352
rect 167969 -146386 168027 -146352
rect 168117 -146386 168175 -146352
rect 168265 -146386 168323 -146352
rect 168413 -146386 168471 -146352
rect 168561 -146386 168619 -146352
rect 168709 -146386 168767 -146352
rect 168857 -146386 168915 -146352
rect 169005 -146386 169063 -146352
rect 169153 -146386 169211 -146352
rect 169301 -146386 169359 -146352
rect 169449 -146386 169507 -146352
rect 169597 -146386 169655 -146352
rect 169745 -146386 169803 -146352
rect 169893 -146386 169951 -146352
rect 170041 -146386 170099 -146352
rect 170189 -146386 170247 -146352
rect 170337 -146386 170395 -146352
rect 170485 -146386 170543 -146352
rect 170633 -146386 170691 -146352
rect 170781 -146386 170839 -146352
rect 170929 -146386 170987 -146352
rect 171077 -146386 171135 -146352
rect 171225 -146386 171283 -146352
rect 171373 -146386 171431 -146352
rect 171521 -146386 171579 -146352
rect 171669 -146386 171727 -146352
rect 171817 -146386 171875 -146352
rect 171965 -146386 172023 -146352
rect 172113 -146386 172171 -146352
rect 172261 -146386 172319 -146352
rect 172409 -146386 172467 -146352
rect 172557 -146386 172615 -146352
rect 172705 -146386 172763 -146352
rect 172853 -146386 172911 -146352
rect 173001 -146386 173059 -146352
rect 173149 -146386 173207 -146352
rect 173297 -146386 173355 -146352
rect 173445 -146386 173503 -146352
rect 173593 -146386 173651 -146352
rect 173741 -146386 173799 -146352
rect 173889 -146386 173947 -146352
rect 174037 -146386 174095 -146352
rect 174185 -146386 174243 -146352
rect 174333 -146386 174391 -146352
rect 174481 -146386 174539 -146352
rect 174629 -146386 174687 -146352
rect 174777 -146386 174835 -146352
rect 174925 -146386 174983 -146352
rect 175073 -146386 175131 -146352
rect 175221 -146386 175279 -146352
rect 175369 -146386 175427 -146352
rect 175517 -146386 175575 -146352
rect 175665 -146386 175723 -146352
rect 175813 -146386 175871 -146352
rect 175961 -146386 176019 -146352
rect 176109 -146386 176167 -146352
rect 165095 -147312 165129 -146436
rect 165243 -147312 165277 -146436
rect 165391 -147312 165425 -146436
rect 165539 -147312 165573 -146436
rect 165687 -147312 165721 -146436
rect 165835 -147312 165869 -146436
rect 165983 -147312 166017 -146436
rect 166131 -147312 166165 -146436
rect 166279 -147312 166313 -146436
rect 166427 -147312 166461 -146436
rect 166575 -147312 166609 -146436
rect 166723 -147312 166757 -146436
rect 166871 -147312 166905 -146436
rect 167019 -147312 167053 -146436
rect 167167 -147312 167201 -146436
rect 167315 -147312 167349 -146436
rect 167463 -147312 167497 -146436
rect 167611 -147312 167645 -146436
rect 167759 -147312 167793 -146436
rect 167907 -147312 167941 -146436
rect 168055 -147312 168089 -146436
rect 168203 -147312 168237 -146436
rect 168351 -147312 168385 -146436
rect 168499 -147312 168533 -146436
rect 168647 -147312 168681 -146436
rect 168795 -147312 168829 -146436
rect 168943 -147312 168977 -146436
rect 169091 -147312 169125 -146436
rect 169239 -147312 169273 -146436
rect 169387 -147312 169421 -146436
rect 169535 -147312 169569 -146436
rect 169683 -147312 169717 -146436
rect 169831 -147312 169865 -146436
rect 169979 -147312 170013 -146436
rect 170127 -147312 170161 -146436
rect 170275 -147312 170309 -146436
rect 170423 -147312 170457 -146436
rect 170571 -147312 170605 -146436
rect 170719 -147312 170753 -146436
rect 170867 -147312 170901 -146436
rect 171015 -147312 171049 -146436
rect 171163 -147312 171197 -146436
rect 171311 -147312 171345 -146436
rect 171459 -147312 171493 -146436
rect 171607 -147312 171641 -146436
rect 171755 -147312 171789 -146436
rect 171903 -147312 171937 -146436
rect 172051 -147312 172085 -146436
rect 172199 -147312 172233 -146436
rect 172347 -147312 172381 -146436
rect 172495 -147312 172529 -146436
rect 172643 -147312 172677 -146436
rect 172791 -147312 172825 -146436
rect 172939 -147312 172973 -146436
rect 173087 -147312 173121 -146436
rect 173235 -147312 173269 -146436
rect 173383 -147312 173417 -146436
rect 173531 -147312 173565 -146436
rect 173679 -147312 173713 -146436
rect 173827 -147312 173861 -146436
rect 173975 -147312 174009 -146436
rect 174123 -147312 174157 -146436
rect 174271 -147312 174305 -146436
rect 174419 -147312 174453 -146436
rect 174567 -147312 174601 -146436
rect 174715 -147312 174749 -146436
rect 174863 -147312 174897 -146436
rect 175011 -147312 175045 -146436
rect 175159 -147312 175193 -146436
rect 175307 -147312 175341 -146436
rect 175455 -147312 175489 -146436
rect 175603 -147312 175637 -146436
rect 175751 -147312 175785 -146436
rect 175899 -147312 175933 -146436
<< nmoslvt >>
rect 540 -147800 2140 -147400
rect 3540 -147800 5140 -147400
rect 6540 -147800 8140 -147400
rect 9540 -147800 11140 -147400
rect 12540 -147800 14140 -147400
rect 15540 -147800 17140 -147400
rect 18540 -147800 20140 -147400
rect 21540 -147800 23140 -147400
rect 24540 -147800 26140 -147400
rect 27540 -147800 29140 -147400
rect 30540 -147800 32140 -147400
rect 33540 -147800 35140 -147400
rect 36540 -147800 38140 -147400
rect 39540 -147800 41140 -147400
rect 42540 -147800 44140 -147400
rect 45540 -147800 47140 -147400
rect 48540 -147800 50140 -147400
rect 51540 -147800 53140 -147400
rect 54540 -147800 56140 -147400
rect 57540 -147800 59140 -147400
rect 60540 -147800 62140 -147400
rect 63540 -147800 65140 -147400
rect 66540 -147800 68140 -147400
rect 69540 -147800 71140 -147400
rect 72540 -147800 74140 -147400
rect 75540 -147800 77140 -147400
rect 78540 -147800 80140 -147400
rect 81540 -147800 83140 -147400
rect 84540 -147800 86140 -147400
rect 87540 -147800 89140 -147400
rect 90540 -147800 92140 -147400
rect 93540 -147800 95140 -147400
rect 96540 -147800 98140 -147400
rect 99540 -147800 101140 -147400
rect 102540 -147800 104140 -147400
rect 105540 -147800 107140 -147400
rect 108540 -147800 110140 -147400
rect 111540 -147800 113140 -147400
rect 114540 -147800 116140 -147400
rect 117540 -147800 119140 -147400
rect 120540 -147800 122140 -147400
rect 123540 -147800 125140 -147400
rect 126540 -147800 128140 -147400
rect 129540 -147800 131140 -147400
rect 132540 -147800 134140 -147400
rect 135540 -147800 137140 -147400
rect 138540 -147800 140140 -147400
rect 141540 -147800 143140 -147400
rect 144540 -147800 146140 -147400
rect 147540 -147800 149140 -147400
<< ndiff >>
rect 540 -147320 2140 -147300
rect 540 -147380 560 -147320
rect 2120 -147380 2140 -147320
rect 540 -147400 2140 -147380
rect 3540 -147320 5140 -147300
rect 3540 -147380 3560 -147320
rect 5120 -147380 5140 -147320
rect 3540 -147400 5140 -147380
rect 6540 -147320 8140 -147300
rect 6540 -147380 6560 -147320
rect 8120 -147380 8140 -147320
rect 6540 -147400 8140 -147380
rect 9540 -147320 11140 -147300
rect 9540 -147380 9560 -147320
rect 11120 -147380 11140 -147320
rect 9540 -147400 11140 -147380
rect 12540 -147320 14140 -147300
rect 12540 -147380 12560 -147320
rect 14120 -147380 14140 -147320
rect 12540 -147400 14140 -147380
rect 15540 -147320 17140 -147300
rect 15540 -147380 15560 -147320
rect 17120 -147380 17140 -147320
rect 15540 -147400 17140 -147380
rect 18540 -147320 20140 -147300
rect 18540 -147380 18560 -147320
rect 20120 -147380 20140 -147320
rect 18540 -147400 20140 -147380
rect 21540 -147320 23140 -147300
rect 21540 -147380 21560 -147320
rect 23120 -147380 23140 -147320
rect 21540 -147400 23140 -147380
rect 24540 -147320 26140 -147300
rect 24540 -147380 24560 -147320
rect 26120 -147380 26140 -147320
rect 24540 -147400 26140 -147380
rect 27540 -147320 29140 -147300
rect 27540 -147380 27560 -147320
rect 29120 -147380 29140 -147320
rect 27540 -147400 29140 -147380
rect 30540 -147320 32140 -147300
rect 30540 -147380 30560 -147320
rect 32120 -147380 32140 -147320
rect 30540 -147400 32140 -147380
rect 33540 -147320 35140 -147300
rect 33540 -147380 33560 -147320
rect 35120 -147380 35140 -147320
rect 33540 -147400 35140 -147380
rect 36540 -147320 38140 -147300
rect 36540 -147380 36560 -147320
rect 38120 -147380 38140 -147320
rect 36540 -147400 38140 -147380
rect 39540 -147320 41140 -147300
rect 39540 -147380 39560 -147320
rect 41120 -147380 41140 -147320
rect 39540 -147400 41140 -147380
rect 42540 -147320 44140 -147300
rect 42540 -147380 42560 -147320
rect 44120 -147380 44140 -147320
rect 42540 -147400 44140 -147380
rect 45540 -147320 47140 -147300
rect 45540 -147380 45560 -147320
rect 47120 -147380 47140 -147320
rect 45540 -147400 47140 -147380
rect 48540 -147320 50140 -147300
rect 48540 -147380 48560 -147320
rect 50120 -147380 50140 -147320
rect 48540 -147400 50140 -147380
rect 51540 -147320 53140 -147300
rect 51540 -147380 51560 -147320
rect 53120 -147380 53140 -147320
rect 51540 -147400 53140 -147380
rect 54540 -147320 56140 -147300
rect 54540 -147380 54560 -147320
rect 56120 -147380 56140 -147320
rect 54540 -147400 56140 -147380
rect 57540 -147320 59140 -147300
rect 57540 -147380 57560 -147320
rect 59120 -147380 59140 -147320
rect 57540 -147400 59140 -147380
rect 60540 -147320 62140 -147300
rect 60540 -147380 60560 -147320
rect 62120 -147380 62140 -147320
rect 60540 -147400 62140 -147380
rect 63540 -147320 65140 -147300
rect 63540 -147380 63560 -147320
rect 65120 -147380 65140 -147320
rect 63540 -147400 65140 -147380
rect 66540 -147320 68140 -147300
rect 66540 -147380 66560 -147320
rect 68120 -147380 68140 -147320
rect 66540 -147400 68140 -147380
rect 69540 -147320 71140 -147300
rect 69540 -147380 69560 -147320
rect 71120 -147380 71140 -147320
rect 69540 -147400 71140 -147380
rect 72540 -147320 74140 -147300
rect 72540 -147380 72560 -147320
rect 74120 -147380 74140 -147320
rect 72540 -147400 74140 -147380
rect 75540 -147320 77140 -147300
rect 75540 -147380 75560 -147320
rect 77120 -147380 77140 -147320
rect 75540 -147400 77140 -147380
rect 78540 -147320 80140 -147300
rect 78540 -147380 78560 -147320
rect 80120 -147380 80140 -147320
rect 78540 -147400 80140 -147380
rect 81540 -147320 83140 -147300
rect 81540 -147380 81560 -147320
rect 83120 -147380 83140 -147320
rect 81540 -147400 83140 -147380
rect 84540 -147320 86140 -147300
rect 84540 -147380 84560 -147320
rect 86120 -147380 86140 -147320
rect 84540 -147400 86140 -147380
rect 87540 -147320 89140 -147300
rect 87540 -147380 87560 -147320
rect 89120 -147380 89140 -147320
rect 87540 -147400 89140 -147380
rect 90540 -147320 92140 -147300
rect 90540 -147380 90560 -147320
rect 92120 -147380 92140 -147320
rect 90540 -147400 92140 -147380
rect 93540 -147320 95140 -147300
rect 93540 -147380 93560 -147320
rect 95120 -147380 95140 -147320
rect 93540 -147400 95140 -147380
rect 96540 -147320 98140 -147300
rect 96540 -147380 96560 -147320
rect 98120 -147380 98140 -147320
rect 96540 -147400 98140 -147380
rect 99540 -147320 101140 -147300
rect 99540 -147380 99560 -147320
rect 101120 -147380 101140 -147320
rect 99540 -147400 101140 -147380
rect 102540 -147320 104140 -147300
rect 102540 -147380 102560 -147320
rect 104120 -147380 104140 -147320
rect 102540 -147400 104140 -147380
rect 105540 -147320 107140 -147300
rect 105540 -147380 105560 -147320
rect 107120 -147380 107140 -147320
rect 105540 -147400 107140 -147380
rect 108540 -147320 110140 -147300
rect 108540 -147380 108560 -147320
rect 110120 -147380 110140 -147320
rect 108540 -147400 110140 -147380
rect 111540 -147320 113140 -147300
rect 111540 -147380 111560 -147320
rect 113120 -147380 113140 -147320
rect 111540 -147400 113140 -147380
rect 114540 -147320 116140 -147300
rect 114540 -147380 114560 -147320
rect 116120 -147380 116140 -147320
rect 114540 -147400 116140 -147380
rect 117540 -147320 119140 -147300
rect 117540 -147380 117560 -147320
rect 119120 -147380 119140 -147320
rect 117540 -147400 119140 -147380
rect 120540 -147320 122140 -147300
rect 120540 -147380 120560 -147320
rect 122120 -147380 122140 -147320
rect 120540 -147400 122140 -147380
rect 123540 -147320 125140 -147300
rect 123540 -147380 123560 -147320
rect 125120 -147380 125140 -147320
rect 123540 -147400 125140 -147380
rect 126540 -147320 128140 -147300
rect 126540 -147380 126560 -147320
rect 128120 -147380 128140 -147320
rect 126540 -147400 128140 -147380
rect 129540 -147320 131140 -147300
rect 129540 -147380 129560 -147320
rect 131120 -147380 131140 -147320
rect 129540 -147400 131140 -147380
rect 132540 -147320 134140 -147300
rect 132540 -147380 132560 -147320
rect 134120 -147380 134140 -147320
rect 132540 -147400 134140 -147380
rect 135540 -147320 137140 -147300
rect 135540 -147380 135560 -147320
rect 137120 -147380 137140 -147320
rect 135540 -147400 137140 -147380
rect 138540 -147320 140140 -147300
rect 138540 -147380 138560 -147320
rect 140120 -147380 140140 -147320
rect 138540 -147400 140140 -147380
rect 141540 -147320 143140 -147300
rect 141540 -147380 141560 -147320
rect 143120 -147380 143140 -147320
rect 141540 -147400 143140 -147380
rect 144540 -147320 146140 -147300
rect 144540 -147380 144560 -147320
rect 146120 -147380 146140 -147320
rect 144540 -147400 146140 -147380
rect 147540 -147320 149140 -147300
rect 147540 -147380 147560 -147320
rect 149120 -147380 149140 -147320
rect 147540 -147400 149140 -147380
rect 540 -147830 2140 -147800
rect 540 -147870 560 -147830
rect 2120 -147870 2140 -147830
rect 540 -147880 2140 -147870
rect 3540 -147830 5140 -147800
rect 3540 -147870 3560 -147830
rect 5120 -147870 5140 -147830
rect 3540 -147880 5140 -147870
rect 6540 -147830 8140 -147800
rect 6540 -147870 6560 -147830
rect 8120 -147870 8140 -147830
rect 6540 -147880 8140 -147870
rect 9540 -147830 11140 -147800
rect 9540 -147870 9560 -147830
rect 11120 -147870 11140 -147830
rect 9540 -147880 11140 -147870
rect 12540 -147830 14140 -147800
rect 12540 -147870 12560 -147830
rect 14120 -147870 14140 -147830
rect 12540 -147880 14140 -147870
rect 15540 -147830 17140 -147800
rect 15540 -147870 15560 -147830
rect 17120 -147870 17140 -147830
rect 15540 -147880 17140 -147870
rect 18540 -147830 20140 -147800
rect 18540 -147870 18560 -147830
rect 20120 -147870 20140 -147830
rect 18540 -147880 20140 -147870
rect 21540 -147830 23140 -147800
rect 21540 -147870 21560 -147830
rect 23120 -147870 23140 -147830
rect 21540 -147880 23140 -147870
rect 24540 -147830 26140 -147800
rect 24540 -147870 24560 -147830
rect 26120 -147870 26140 -147830
rect 24540 -147880 26140 -147870
rect 27540 -147830 29140 -147800
rect 27540 -147870 27560 -147830
rect 29120 -147870 29140 -147830
rect 27540 -147880 29140 -147870
rect 30540 -147830 32140 -147800
rect 30540 -147870 30560 -147830
rect 32120 -147870 32140 -147830
rect 30540 -147880 32140 -147870
rect 33540 -147830 35140 -147800
rect 33540 -147870 33560 -147830
rect 35120 -147870 35140 -147830
rect 33540 -147880 35140 -147870
rect 36540 -147830 38140 -147800
rect 36540 -147870 36560 -147830
rect 38120 -147870 38140 -147830
rect 36540 -147880 38140 -147870
rect 39540 -147830 41140 -147800
rect 39540 -147870 39560 -147830
rect 41120 -147870 41140 -147830
rect 39540 -147880 41140 -147870
rect 42540 -147830 44140 -147800
rect 42540 -147870 42560 -147830
rect 44120 -147870 44140 -147830
rect 42540 -147880 44140 -147870
rect 45540 -147830 47140 -147800
rect 45540 -147870 45560 -147830
rect 47120 -147870 47140 -147830
rect 45540 -147880 47140 -147870
rect 48540 -147830 50140 -147800
rect 48540 -147870 48560 -147830
rect 50120 -147870 50140 -147830
rect 48540 -147880 50140 -147870
rect 51540 -147830 53140 -147800
rect 51540 -147870 51560 -147830
rect 53120 -147870 53140 -147830
rect 51540 -147880 53140 -147870
rect 54540 -147830 56140 -147800
rect 54540 -147870 54560 -147830
rect 56120 -147870 56140 -147830
rect 54540 -147880 56140 -147870
rect 57540 -147830 59140 -147800
rect 57540 -147870 57560 -147830
rect 59120 -147870 59140 -147830
rect 57540 -147880 59140 -147870
rect 60540 -147830 62140 -147800
rect 60540 -147870 60560 -147830
rect 62120 -147870 62140 -147830
rect 60540 -147880 62140 -147870
rect 63540 -147830 65140 -147800
rect 63540 -147870 63560 -147830
rect 65120 -147870 65140 -147830
rect 63540 -147880 65140 -147870
rect 66540 -147830 68140 -147800
rect 66540 -147870 66560 -147830
rect 68120 -147870 68140 -147830
rect 66540 -147880 68140 -147870
rect 69540 -147830 71140 -147800
rect 69540 -147870 69560 -147830
rect 71120 -147870 71140 -147830
rect 69540 -147880 71140 -147870
rect 72540 -147830 74140 -147800
rect 72540 -147870 72560 -147830
rect 74120 -147870 74140 -147830
rect 72540 -147880 74140 -147870
rect 75540 -147830 77140 -147800
rect 75540 -147870 75560 -147830
rect 77120 -147870 77140 -147830
rect 75540 -147880 77140 -147870
rect 78540 -147830 80140 -147800
rect 78540 -147870 78560 -147830
rect 80120 -147870 80140 -147830
rect 78540 -147880 80140 -147870
rect 81540 -147830 83140 -147800
rect 81540 -147870 81560 -147830
rect 83120 -147870 83140 -147830
rect 81540 -147880 83140 -147870
rect 84540 -147830 86140 -147800
rect 84540 -147870 84560 -147830
rect 86120 -147870 86140 -147830
rect 84540 -147880 86140 -147870
rect 87540 -147830 89140 -147800
rect 87540 -147870 87560 -147830
rect 89120 -147870 89140 -147830
rect 87540 -147880 89140 -147870
rect 90540 -147830 92140 -147800
rect 90540 -147870 90560 -147830
rect 92120 -147870 92140 -147830
rect 90540 -147880 92140 -147870
rect 93540 -147830 95140 -147800
rect 93540 -147870 93560 -147830
rect 95120 -147870 95140 -147830
rect 93540 -147880 95140 -147870
rect 96540 -147830 98140 -147800
rect 96540 -147870 96560 -147830
rect 98120 -147870 98140 -147830
rect 96540 -147880 98140 -147870
rect 99540 -147830 101140 -147800
rect 99540 -147870 99560 -147830
rect 101120 -147870 101140 -147830
rect 99540 -147880 101140 -147870
rect 102540 -147830 104140 -147800
rect 102540 -147870 102560 -147830
rect 104120 -147870 104140 -147830
rect 102540 -147880 104140 -147870
rect 105540 -147830 107140 -147800
rect 105540 -147870 105560 -147830
rect 107120 -147870 107140 -147830
rect 105540 -147880 107140 -147870
rect 108540 -147830 110140 -147800
rect 108540 -147870 108560 -147830
rect 110120 -147870 110140 -147830
rect 108540 -147880 110140 -147870
rect 111540 -147830 113140 -147800
rect 111540 -147870 111560 -147830
rect 113120 -147870 113140 -147830
rect 111540 -147880 113140 -147870
rect 114540 -147830 116140 -147800
rect 114540 -147870 114560 -147830
rect 116120 -147870 116140 -147830
rect 114540 -147880 116140 -147870
rect 117540 -147830 119140 -147800
rect 117540 -147870 117560 -147830
rect 119120 -147870 119140 -147830
rect 117540 -147880 119140 -147870
rect 120540 -147830 122140 -147800
rect 120540 -147870 120560 -147830
rect 122120 -147870 122140 -147830
rect 120540 -147880 122140 -147870
rect 123540 -147830 125140 -147800
rect 123540 -147870 123560 -147830
rect 125120 -147870 125140 -147830
rect 123540 -147880 125140 -147870
rect 126540 -147830 128140 -147800
rect 126540 -147870 126560 -147830
rect 128120 -147870 128140 -147830
rect 126540 -147880 128140 -147870
rect 129540 -147830 131140 -147800
rect 129540 -147870 129560 -147830
rect 131120 -147870 131140 -147830
rect 129540 -147880 131140 -147870
rect 132540 -147830 134140 -147800
rect 132540 -147870 132560 -147830
rect 134120 -147870 134140 -147830
rect 132540 -147880 134140 -147870
rect 135540 -147830 137140 -147800
rect 135540 -147870 135560 -147830
rect 137120 -147870 137140 -147830
rect 135540 -147880 137140 -147870
rect 138540 -147830 140140 -147800
rect 138540 -147870 138560 -147830
rect 140120 -147870 140140 -147830
rect 138540 -147880 140140 -147870
rect 141540 -147830 143140 -147800
rect 141540 -147870 141560 -147830
rect 143120 -147870 143140 -147830
rect 141540 -147880 143140 -147870
rect 144540 -147830 146140 -147800
rect 144540 -147870 144560 -147830
rect 146120 -147870 146140 -147830
rect 144540 -147880 146140 -147870
rect 147540 -147830 149140 -147800
rect 147540 -147870 147560 -147830
rect 149120 -147870 149140 -147830
rect 147540 -147880 149140 -147870
<< ndiffc >>
rect 560 -147380 2120 -147320
rect 3560 -147380 5120 -147320
rect 6560 -147380 8120 -147320
rect 9560 -147380 11120 -147320
rect 12560 -147380 14120 -147320
rect 15560 -147380 17120 -147320
rect 18560 -147380 20120 -147320
rect 21560 -147380 23120 -147320
rect 24560 -147380 26120 -147320
rect 27560 -147380 29120 -147320
rect 30560 -147380 32120 -147320
rect 33560 -147380 35120 -147320
rect 36560 -147380 38120 -147320
rect 39560 -147380 41120 -147320
rect 42560 -147380 44120 -147320
rect 45560 -147380 47120 -147320
rect 48560 -147380 50120 -147320
rect 51560 -147380 53120 -147320
rect 54560 -147380 56120 -147320
rect 57560 -147380 59120 -147320
rect 60560 -147380 62120 -147320
rect 63560 -147380 65120 -147320
rect 66560 -147380 68120 -147320
rect 69560 -147380 71120 -147320
rect 72560 -147380 74120 -147320
rect 75560 -147380 77120 -147320
rect 78560 -147380 80120 -147320
rect 81560 -147380 83120 -147320
rect 84560 -147380 86120 -147320
rect 87560 -147380 89120 -147320
rect 90560 -147380 92120 -147320
rect 93560 -147380 95120 -147320
rect 96560 -147380 98120 -147320
rect 99560 -147380 101120 -147320
rect 102560 -147380 104120 -147320
rect 105560 -147380 107120 -147320
rect 108560 -147380 110120 -147320
rect 111560 -147380 113120 -147320
rect 114560 -147380 116120 -147320
rect 117560 -147380 119120 -147320
rect 120560 -147380 122120 -147320
rect 123560 -147380 125120 -147320
rect 126560 -147380 128120 -147320
rect 129560 -147380 131120 -147320
rect 132560 -147380 134120 -147320
rect 135560 -147380 137120 -147320
rect 138560 -147380 140120 -147320
rect 141560 -147380 143120 -147320
rect 144560 -147380 146120 -147320
rect 147560 -147380 149120 -147320
rect 560 -147870 2120 -147830
rect 3560 -147870 5120 -147830
rect 6560 -147870 8120 -147830
rect 9560 -147870 11120 -147830
rect 12560 -147870 14120 -147830
rect 15560 -147870 17120 -147830
rect 18560 -147870 20120 -147830
rect 21560 -147870 23120 -147830
rect 24560 -147870 26120 -147830
rect 27560 -147870 29120 -147830
rect 30560 -147870 32120 -147830
rect 33560 -147870 35120 -147830
rect 36560 -147870 38120 -147830
rect 39560 -147870 41120 -147830
rect 42560 -147870 44120 -147830
rect 45560 -147870 47120 -147830
rect 48560 -147870 50120 -147830
rect 51560 -147870 53120 -147830
rect 54560 -147870 56120 -147830
rect 57560 -147870 59120 -147830
rect 60560 -147870 62120 -147830
rect 63560 -147870 65120 -147830
rect 66560 -147870 68120 -147830
rect 69560 -147870 71120 -147830
rect 72560 -147870 74120 -147830
rect 75560 -147870 77120 -147830
rect 78560 -147870 80120 -147830
rect 81560 -147870 83120 -147830
rect 84560 -147870 86120 -147830
rect 87560 -147870 89120 -147830
rect 90560 -147870 92120 -147830
rect 93560 -147870 95120 -147830
rect 96560 -147870 98120 -147830
rect 99560 -147870 101120 -147830
rect 102560 -147870 104120 -147830
rect 105560 -147870 107120 -147830
rect 108560 -147870 110120 -147830
rect 111560 -147870 113120 -147830
rect 114560 -147870 116120 -147830
rect 117560 -147870 119120 -147830
rect 120560 -147870 122120 -147830
rect 123560 -147870 125120 -147830
rect 126560 -147870 128120 -147830
rect 129560 -147870 131120 -147830
rect 132560 -147870 134120 -147830
rect 135560 -147870 137120 -147830
rect 138560 -147870 140120 -147830
rect 141560 -147870 143120 -147830
rect 144560 -147870 146120 -147830
rect 147560 -147870 149120 -147830
<< poly >>
rect 510 -147490 540 -147400
rect 220 -147500 540 -147490
rect 220 -147700 240 -147500
rect 420 -147700 540 -147500
rect 220 -147710 540 -147700
rect 510 -147800 540 -147710
rect 2140 -147800 2170 -147400
rect 3510 -147490 3540 -147400
rect 3220 -147500 3540 -147490
rect 3220 -147700 3240 -147500
rect 3420 -147700 3540 -147500
rect 3220 -147710 3540 -147700
rect 3510 -147800 3540 -147710
rect 5140 -147800 5170 -147400
rect 6510 -147490 6540 -147400
rect 6220 -147500 6540 -147490
rect 6220 -147700 6240 -147500
rect 6420 -147700 6540 -147500
rect 6220 -147710 6540 -147700
rect 6510 -147800 6540 -147710
rect 8140 -147800 8170 -147400
rect 9510 -147490 9540 -147400
rect 9220 -147500 9540 -147490
rect 9220 -147700 9240 -147500
rect 9420 -147700 9540 -147500
rect 9220 -147710 9540 -147700
rect 9510 -147800 9540 -147710
rect 11140 -147800 11170 -147400
rect 12510 -147490 12540 -147400
rect 12220 -147500 12540 -147490
rect 12220 -147700 12240 -147500
rect 12420 -147700 12540 -147500
rect 12220 -147710 12540 -147700
rect 12510 -147800 12540 -147710
rect 14140 -147800 14170 -147400
rect 15510 -147490 15540 -147400
rect 15220 -147500 15540 -147490
rect 15220 -147700 15240 -147500
rect 15420 -147700 15540 -147500
rect 15220 -147710 15540 -147700
rect 15510 -147800 15540 -147710
rect 17140 -147800 17170 -147400
rect 18510 -147490 18540 -147400
rect 18220 -147500 18540 -147490
rect 18220 -147700 18240 -147500
rect 18420 -147700 18540 -147500
rect 18220 -147710 18540 -147700
rect 18510 -147800 18540 -147710
rect 20140 -147800 20170 -147400
rect 21510 -147490 21540 -147400
rect 21220 -147500 21540 -147490
rect 21220 -147700 21240 -147500
rect 21420 -147700 21540 -147500
rect 21220 -147710 21540 -147700
rect 21510 -147800 21540 -147710
rect 23140 -147800 23170 -147400
rect 24510 -147490 24540 -147400
rect 24220 -147500 24540 -147490
rect 24220 -147700 24240 -147500
rect 24420 -147700 24540 -147500
rect 24220 -147710 24540 -147700
rect 24510 -147800 24540 -147710
rect 26140 -147800 26170 -147400
rect 27510 -147490 27540 -147400
rect 27220 -147500 27540 -147490
rect 27220 -147700 27240 -147500
rect 27420 -147700 27540 -147500
rect 27220 -147710 27540 -147700
rect 27510 -147800 27540 -147710
rect 29140 -147800 29170 -147400
rect 30510 -147490 30540 -147400
rect 30220 -147500 30540 -147490
rect 30220 -147700 30240 -147500
rect 30420 -147700 30540 -147500
rect 30220 -147710 30540 -147700
rect 30510 -147800 30540 -147710
rect 32140 -147800 32170 -147400
rect 33510 -147490 33540 -147400
rect 33220 -147500 33540 -147490
rect 33220 -147700 33240 -147500
rect 33420 -147700 33540 -147500
rect 33220 -147710 33540 -147700
rect 33510 -147800 33540 -147710
rect 35140 -147800 35170 -147400
rect 36510 -147490 36540 -147400
rect 36220 -147500 36540 -147490
rect 36220 -147700 36240 -147500
rect 36420 -147700 36540 -147500
rect 36220 -147710 36540 -147700
rect 36510 -147800 36540 -147710
rect 38140 -147800 38170 -147400
rect 39510 -147490 39540 -147400
rect 39220 -147500 39540 -147490
rect 39220 -147700 39240 -147500
rect 39420 -147700 39540 -147500
rect 39220 -147710 39540 -147700
rect 39510 -147800 39540 -147710
rect 41140 -147800 41170 -147400
rect 42510 -147490 42540 -147400
rect 42220 -147500 42540 -147490
rect 42220 -147700 42240 -147500
rect 42420 -147700 42540 -147500
rect 42220 -147710 42540 -147700
rect 42510 -147800 42540 -147710
rect 44140 -147800 44170 -147400
rect 45510 -147490 45540 -147400
rect 45220 -147500 45540 -147490
rect 45220 -147700 45240 -147500
rect 45420 -147700 45540 -147500
rect 45220 -147710 45540 -147700
rect 45510 -147800 45540 -147710
rect 47140 -147800 47170 -147400
rect 48510 -147490 48540 -147400
rect 48220 -147500 48540 -147490
rect 48220 -147700 48240 -147500
rect 48420 -147700 48540 -147500
rect 48220 -147710 48540 -147700
rect 48510 -147800 48540 -147710
rect 50140 -147800 50170 -147400
rect 51510 -147490 51540 -147400
rect 51220 -147500 51540 -147490
rect 51220 -147700 51240 -147500
rect 51420 -147700 51540 -147500
rect 51220 -147710 51540 -147700
rect 51510 -147800 51540 -147710
rect 53140 -147800 53170 -147400
rect 54510 -147490 54540 -147400
rect 54220 -147500 54540 -147490
rect 54220 -147700 54240 -147500
rect 54420 -147700 54540 -147500
rect 54220 -147710 54540 -147700
rect 54510 -147800 54540 -147710
rect 56140 -147800 56170 -147400
rect 57510 -147490 57540 -147400
rect 57220 -147500 57540 -147490
rect 57220 -147700 57240 -147500
rect 57420 -147700 57540 -147500
rect 57220 -147710 57540 -147700
rect 57510 -147800 57540 -147710
rect 59140 -147800 59170 -147400
rect 60510 -147490 60540 -147400
rect 60220 -147500 60540 -147490
rect 60220 -147700 60240 -147500
rect 60420 -147700 60540 -147500
rect 60220 -147710 60540 -147700
rect 60510 -147800 60540 -147710
rect 62140 -147800 62170 -147400
rect 63510 -147490 63540 -147400
rect 63220 -147500 63540 -147490
rect 63220 -147700 63240 -147500
rect 63420 -147700 63540 -147500
rect 63220 -147710 63540 -147700
rect 63510 -147800 63540 -147710
rect 65140 -147800 65170 -147400
rect 66510 -147490 66540 -147400
rect 66220 -147500 66540 -147490
rect 66220 -147700 66240 -147500
rect 66420 -147700 66540 -147500
rect 66220 -147710 66540 -147700
rect 66510 -147800 66540 -147710
rect 68140 -147800 68170 -147400
rect 69510 -147490 69540 -147400
rect 69220 -147500 69540 -147490
rect 69220 -147700 69240 -147500
rect 69420 -147700 69540 -147500
rect 69220 -147710 69540 -147700
rect 69510 -147800 69540 -147710
rect 71140 -147800 71170 -147400
rect 72510 -147490 72540 -147400
rect 72220 -147500 72540 -147490
rect 72220 -147700 72240 -147500
rect 72420 -147700 72540 -147500
rect 72220 -147710 72540 -147700
rect 72510 -147800 72540 -147710
rect 74140 -147800 74170 -147400
rect 75510 -147490 75540 -147400
rect 75220 -147500 75540 -147490
rect 75220 -147700 75240 -147500
rect 75420 -147700 75540 -147500
rect 75220 -147710 75540 -147700
rect 75510 -147800 75540 -147710
rect 77140 -147800 77170 -147400
rect 78510 -147490 78540 -147400
rect 78220 -147500 78540 -147490
rect 78220 -147700 78240 -147500
rect 78420 -147700 78540 -147500
rect 78220 -147710 78540 -147700
rect 78510 -147800 78540 -147710
rect 80140 -147800 80170 -147400
rect 81510 -147490 81540 -147400
rect 81220 -147500 81540 -147490
rect 81220 -147700 81240 -147500
rect 81420 -147700 81540 -147500
rect 81220 -147710 81540 -147700
rect 81510 -147800 81540 -147710
rect 83140 -147800 83170 -147400
rect 84510 -147490 84540 -147400
rect 84220 -147500 84540 -147490
rect 84220 -147700 84240 -147500
rect 84420 -147700 84540 -147500
rect 84220 -147710 84540 -147700
rect 84510 -147800 84540 -147710
rect 86140 -147800 86170 -147400
rect 87510 -147490 87540 -147400
rect 87220 -147500 87540 -147490
rect 87220 -147700 87240 -147500
rect 87420 -147700 87540 -147500
rect 87220 -147710 87540 -147700
rect 87510 -147800 87540 -147710
rect 89140 -147800 89170 -147400
rect 90510 -147490 90540 -147400
rect 90220 -147500 90540 -147490
rect 90220 -147700 90240 -147500
rect 90420 -147700 90540 -147500
rect 90220 -147710 90540 -147700
rect 90510 -147800 90540 -147710
rect 92140 -147800 92170 -147400
rect 93510 -147490 93540 -147400
rect 93220 -147500 93540 -147490
rect 93220 -147700 93240 -147500
rect 93420 -147700 93540 -147500
rect 93220 -147710 93540 -147700
rect 93510 -147800 93540 -147710
rect 95140 -147800 95170 -147400
rect 96510 -147490 96540 -147400
rect 96220 -147500 96540 -147490
rect 96220 -147700 96240 -147500
rect 96420 -147700 96540 -147500
rect 96220 -147710 96540 -147700
rect 96510 -147800 96540 -147710
rect 98140 -147800 98170 -147400
rect 99510 -147490 99540 -147400
rect 99220 -147500 99540 -147490
rect 99220 -147700 99240 -147500
rect 99420 -147700 99540 -147500
rect 99220 -147710 99540 -147700
rect 99510 -147800 99540 -147710
rect 101140 -147800 101170 -147400
rect 102510 -147490 102540 -147400
rect 102220 -147500 102540 -147490
rect 102220 -147700 102240 -147500
rect 102420 -147700 102540 -147500
rect 102220 -147710 102540 -147700
rect 102510 -147800 102540 -147710
rect 104140 -147800 104170 -147400
rect 105510 -147490 105540 -147400
rect 105220 -147500 105540 -147490
rect 105220 -147700 105240 -147500
rect 105420 -147700 105540 -147500
rect 105220 -147710 105540 -147700
rect 105510 -147800 105540 -147710
rect 107140 -147800 107170 -147400
rect 108510 -147490 108540 -147400
rect 108220 -147500 108540 -147490
rect 108220 -147700 108240 -147500
rect 108420 -147700 108540 -147500
rect 108220 -147710 108540 -147700
rect 108510 -147800 108540 -147710
rect 110140 -147800 110170 -147400
rect 111510 -147490 111540 -147400
rect 111220 -147500 111540 -147490
rect 111220 -147700 111240 -147500
rect 111420 -147700 111540 -147500
rect 111220 -147710 111540 -147700
rect 111510 -147800 111540 -147710
rect 113140 -147800 113170 -147400
rect 114510 -147490 114540 -147400
rect 114220 -147500 114540 -147490
rect 114220 -147700 114240 -147500
rect 114420 -147700 114540 -147500
rect 114220 -147710 114540 -147700
rect 114510 -147800 114540 -147710
rect 116140 -147800 116170 -147400
rect 117510 -147490 117540 -147400
rect 117220 -147500 117540 -147490
rect 117220 -147700 117240 -147500
rect 117420 -147700 117540 -147500
rect 117220 -147710 117540 -147700
rect 117510 -147800 117540 -147710
rect 119140 -147800 119170 -147400
rect 120510 -147490 120540 -147400
rect 120220 -147500 120540 -147490
rect 120220 -147700 120240 -147500
rect 120420 -147700 120540 -147500
rect 120220 -147710 120540 -147700
rect 120510 -147800 120540 -147710
rect 122140 -147800 122170 -147400
rect 123510 -147490 123540 -147400
rect 123220 -147500 123540 -147490
rect 123220 -147700 123240 -147500
rect 123420 -147700 123540 -147500
rect 123220 -147710 123540 -147700
rect 123510 -147800 123540 -147710
rect 125140 -147800 125170 -147400
rect 126510 -147490 126540 -147400
rect 126220 -147500 126540 -147490
rect 126220 -147700 126240 -147500
rect 126420 -147700 126540 -147500
rect 126220 -147710 126540 -147700
rect 126510 -147800 126540 -147710
rect 128140 -147800 128170 -147400
rect 129510 -147490 129540 -147400
rect 129220 -147500 129540 -147490
rect 129220 -147700 129240 -147500
rect 129420 -147700 129540 -147500
rect 129220 -147710 129540 -147700
rect 129510 -147800 129540 -147710
rect 131140 -147800 131170 -147400
rect 132510 -147490 132540 -147400
rect 132220 -147500 132540 -147490
rect 132220 -147700 132240 -147500
rect 132420 -147700 132540 -147500
rect 132220 -147710 132540 -147700
rect 132510 -147800 132540 -147710
rect 134140 -147800 134170 -147400
rect 135510 -147490 135540 -147400
rect 135220 -147500 135540 -147490
rect 135220 -147700 135240 -147500
rect 135420 -147700 135540 -147500
rect 135220 -147710 135540 -147700
rect 135510 -147800 135540 -147710
rect 137140 -147800 137170 -147400
rect 138510 -147490 138540 -147400
rect 138220 -147500 138540 -147490
rect 138220 -147700 138240 -147500
rect 138420 -147700 138540 -147500
rect 138220 -147710 138540 -147700
rect 138510 -147800 138540 -147710
rect 140140 -147800 140170 -147400
rect 141510 -147490 141540 -147400
rect 141220 -147500 141540 -147490
rect 141220 -147700 141240 -147500
rect 141420 -147700 141540 -147500
rect 141220 -147710 141540 -147700
rect 141510 -147800 141540 -147710
rect 143140 -147800 143170 -147400
rect 144510 -147490 144540 -147400
rect 144220 -147500 144540 -147490
rect 144220 -147700 144240 -147500
rect 144420 -147700 144540 -147500
rect 144220 -147710 144540 -147700
rect 144510 -147800 144540 -147710
rect 146140 -147800 146170 -147400
rect 147510 -147490 147540 -147400
rect 147220 -147500 147540 -147490
rect 147220 -147700 147240 -147500
rect 147420 -147700 147540 -147500
rect 147220 -147710 147540 -147700
rect 147510 -147800 147540 -147710
rect 149140 -147800 149170 -147400
<< polycont >>
rect 240 -147700 420 -147500
rect 3240 -147700 3420 -147500
rect 6240 -147700 6420 -147500
rect 9240 -147700 9420 -147500
rect 12240 -147700 12420 -147500
rect 15240 -147700 15420 -147500
rect 18240 -147700 18420 -147500
rect 21240 -147700 21420 -147500
rect 24240 -147700 24420 -147500
rect 27240 -147700 27420 -147500
rect 30240 -147700 30420 -147500
rect 33240 -147700 33420 -147500
rect 36240 -147700 36420 -147500
rect 39240 -147700 39420 -147500
rect 42240 -147700 42420 -147500
rect 45240 -147700 45420 -147500
rect 48240 -147700 48420 -147500
rect 51240 -147700 51420 -147500
rect 54240 -147700 54420 -147500
rect 57240 -147700 57420 -147500
rect 60240 -147700 60420 -147500
rect 63240 -147700 63420 -147500
rect 66240 -147700 66420 -147500
rect 69240 -147700 69420 -147500
rect 72240 -147700 72420 -147500
rect 75240 -147700 75420 -147500
rect 78240 -147700 78420 -147500
rect 81240 -147700 81420 -147500
rect 84240 -147700 84420 -147500
rect 87240 -147700 87420 -147500
rect 90240 -147700 90420 -147500
rect 93240 -147700 93420 -147500
rect 96240 -147700 96420 -147500
rect 99240 -147700 99420 -147500
rect 102240 -147700 102420 -147500
rect 105240 -147700 105420 -147500
rect 108240 -147700 108420 -147500
rect 111240 -147700 111420 -147500
rect 114240 -147700 114420 -147500
rect 117240 -147700 117420 -147500
rect 120240 -147700 120420 -147500
rect 123240 -147700 123420 -147500
rect 126240 -147700 126420 -147500
rect 129240 -147700 129420 -147500
rect 132240 -147700 132420 -147500
rect 135240 -147700 135420 -147500
rect 138240 -147700 138420 -147500
rect 141240 -147700 141420 -147500
rect 144240 -147700 144420 -147500
rect 147240 -147700 147420 -147500
<< locali >>
rect 540 -147290 560 -147230
rect 2120 -147290 2140 -147230
rect 540 -147320 2140 -147290
rect 540 -147380 560 -147320
rect 2120 -147380 2140 -147320
rect 3540 -147290 3560 -147230
rect 5120 -147290 5140 -147230
rect 3540 -147320 5140 -147290
rect 3540 -147380 3560 -147320
rect 5120 -147380 5140 -147320
rect 6540 -147290 6560 -147230
rect 8120 -147290 8140 -147230
rect 6540 -147320 8140 -147290
rect 6540 -147380 6560 -147320
rect 8120 -147380 8140 -147320
rect 9540 -147290 9560 -147230
rect 11120 -147290 11140 -147230
rect 9540 -147320 11140 -147290
rect 9540 -147380 9560 -147320
rect 11120 -147380 11140 -147320
rect 12540 -147290 12560 -147230
rect 14120 -147290 14140 -147230
rect 12540 -147320 14140 -147290
rect 12540 -147380 12560 -147320
rect 14120 -147380 14140 -147320
rect 15540 -147290 15560 -147230
rect 17120 -147290 17140 -147230
rect 15540 -147320 17140 -147290
rect 15540 -147380 15560 -147320
rect 17120 -147380 17140 -147320
rect 18540 -147290 18560 -147230
rect 20120 -147290 20140 -147230
rect 18540 -147320 20140 -147290
rect 18540 -147380 18560 -147320
rect 20120 -147380 20140 -147320
rect 21540 -147290 21560 -147230
rect 23120 -147290 23140 -147230
rect 21540 -147320 23140 -147290
rect 21540 -147380 21560 -147320
rect 23120 -147380 23140 -147320
rect 24540 -147290 24560 -147230
rect 26120 -147290 26140 -147230
rect 24540 -147320 26140 -147290
rect 24540 -147380 24560 -147320
rect 26120 -147380 26140 -147320
rect 27540 -147290 27560 -147230
rect 29120 -147290 29140 -147230
rect 27540 -147320 29140 -147290
rect 27540 -147380 27560 -147320
rect 29120 -147380 29140 -147320
rect 30540 -147290 30560 -147230
rect 32120 -147290 32140 -147230
rect 30540 -147320 32140 -147290
rect 30540 -147380 30560 -147320
rect 32120 -147380 32140 -147320
rect 33540 -147290 33560 -147230
rect 35120 -147290 35140 -147230
rect 33540 -147320 35140 -147290
rect 33540 -147380 33560 -147320
rect 35120 -147380 35140 -147320
rect 36540 -147290 36560 -147230
rect 38120 -147290 38140 -147230
rect 36540 -147320 38140 -147290
rect 36540 -147380 36560 -147320
rect 38120 -147380 38140 -147320
rect 39540 -147290 39560 -147230
rect 41120 -147290 41140 -147230
rect 39540 -147320 41140 -147290
rect 39540 -147380 39560 -147320
rect 41120 -147380 41140 -147320
rect 42540 -147290 42560 -147230
rect 44120 -147290 44140 -147230
rect 42540 -147320 44140 -147290
rect 42540 -147380 42560 -147320
rect 44120 -147380 44140 -147320
rect 45540 -147290 45560 -147230
rect 47120 -147290 47140 -147230
rect 45540 -147320 47140 -147290
rect 45540 -147380 45560 -147320
rect 47120 -147380 47140 -147320
rect 48540 -147290 48560 -147230
rect 50120 -147290 50140 -147230
rect 48540 -147320 50140 -147290
rect 48540 -147380 48560 -147320
rect 50120 -147380 50140 -147320
rect 51540 -147290 51560 -147230
rect 53120 -147290 53140 -147230
rect 51540 -147320 53140 -147290
rect 51540 -147380 51560 -147320
rect 53120 -147380 53140 -147320
rect 54540 -147290 54560 -147230
rect 56120 -147290 56140 -147230
rect 54540 -147320 56140 -147290
rect 54540 -147380 54560 -147320
rect 56120 -147380 56140 -147320
rect 57540 -147290 57560 -147230
rect 59120 -147290 59140 -147230
rect 57540 -147320 59140 -147290
rect 57540 -147380 57560 -147320
rect 59120 -147380 59140 -147320
rect 60540 -147290 60560 -147230
rect 62120 -147290 62140 -147230
rect 60540 -147320 62140 -147290
rect 60540 -147380 60560 -147320
rect 62120 -147380 62140 -147320
rect 63540 -147290 63560 -147230
rect 65120 -147290 65140 -147230
rect 63540 -147320 65140 -147290
rect 63540 -147380 63560 -147320
rect 65120 -147380 65140 -147320
rect 66540 -147290 66560 -147230
rect 68120 -147290 68140 -147230
rect 66540 -147320 68140 -147290
rect 66540 -147380 66560 -147320
rect 68120 -147380 68140 -147320
rect 69540 -147290 69560 -147230
rect 71120 -147290 71140 -147230
rect 69540 -147320 71140 -147290
rect 69540 -147380 69560 -147320
rect 71120 -147380 71140 -147320
rect 72540 -147290 72560 -147230
rect 74120 -147290 74140 -147230
rect 72540 -147320 74140 -147290
rect 72540 -147380 72560 -147320
rect 74120 -147380 74140 -147320
rect 75540 -147290 75560 -147230
rect 77120 -147290 77140 -147230
rect 75540 -147320 77140 -147290
rect 75540 -147380 75560 -147320
rect 77120 -147380 77140 -147320
rect 78540 -147290 78560 -147230
rect 80120 -147290 80140 -147230
rect 78540 -147320 80140 -147290
rect 78540 -147380 78560 -147320
rect 80120 -147380 80140 -147320
rect 81540 -147290 81560 -147230
rect 83120 -147290 83140 -147230
rect 81540 -147320 83140 -147290
rect 81540 -147380 81560 -147320
rect 83120 -147380 83140 -147320
rect 84540 -147290 84560 -147230
rect 86120 -147290 86140 -147230
rect 84540 -147320 86140 -147290
rect 84540 -147380 84560 -147320
rect 86120 -147380 86140 -147320
rect 87540 -147290 87560 -147230
rect 89120 -147290 89140 -147230
rect 87540 -147320 89140 -147290
rect 87540 -147380 87560 -147320
rect 89120 -147380 89140 -147320
rect 90540 -147290 90560 -147230
rect 92120 -147290 92140 -147230
rect 90540 -147320 92140 -147290
rect 90540 -147380 90560 -147320
rect 92120 -147380 92140 -147320
rect 93540 -147290 93560 -147230
rect 95120 -147290 95140 -147230
rect 93540 -147320 95140 -147290
rect 93540 -147380 93560 -147320
rect 95120 -147380 95140 -147320
rect 96540 -147290 96560 -147230
rect 98120 -147290 98140 -147230
rect 96540 -147320 98140 -147290
rect 96540 -147380 96560 -147320
rect 98120 -147380 98140 -147320
rect 99540 -147290 99560 -147230
rect 101120 -147290 101140 -147230
rect 99540 -147320 101140 -147290
rect 99540 -147380 99560 -147320
rect 101120 -147380 101140 -147320
rect 102540 -147290 102560 -147230
rect 104120 -147290 104140 -147230
rect 102540 -147320 104140 -147290
rect 102540 -147380 102560 -147320
rect 104120 -147380 104140 -147320
rect 105540 -147290 105560 -147230
rect 107120 -147290 107140 -147230
rect 105540 -147320 107140 -147290
rect 105540 -147380 105560 -147320
rect 107120 -147380 107140 -147320
rect 108540 -147290 108560 -147230
rect 110120 -147290 110140 -147230
rect 108540 -147320 110140 -147290
rect 108540 -147380 108560 -147320
rect 110120 -147380 110140 -147320
rect 111540 -147290 111560 -147230
rect 113120 -147290 113140 -147230
rect 111540 -147320 113140 -147290
rect 111540 -147380 111560 -147320
rect 113120 -147380 113140 -147320
rect 114540 -147290 114560 -147230
rect 116120 -147290 116140 -147230
rect 114540 -147320 116140 -147290
rect 114540 -147380 114560 -147320
rect 116120 -147380 116140 -147320
rect 117540 -147290 117560 -147230
rect 119120 -147290 119140 -147230
rect 117540 -147320 119140 -147290
rect 117540 -147380 117560 -147320
rect 119120 -147380 119140 -147320
rect 120540 -147290 120560 -147230
rect 122120 -147290 122140 -147230
rect 120540 -147320 122140 -147290
rect 120540 -147380 120560 -147320
rect 122120 -147380 122140 -147320
rect 123540 -147290 123560 -147230
rect 125120 -147290 125140 -147230
rect 123540 -147320 125140 -147290
rect 123540 -147380 123560 -147320
rect 125120 -147380 125140 -147320
rect 126540 -147290 126560 -147230
rect 128120 -147290 128140 -147230
rect 126540 -147320 128140 -147290
rect 126540 -147380 126560 -147320
rect 128120 -147380 128140 -147320
rect 129540 -147290 129560 -147230
rect 131120 -147290 131140 -147230
rect 129540 -147320 131140 -147290
rect 129540 -147380 129560 -147320
rect 131120 -147380 131140 -147320
rect 132540 -147290 132560 -147230
rect 134120 -147290 134140 -147230
rect 132540 -147320 134140 -147290
rect 132540 -147380 132560 -147320
rect 134120 -147380 134140 -147320
rect 135540 -147290 135560 -147230
rect 137120 -147290 137140 -147230
rect 135540 -147320 137140 -147290
rect 135540 -147380 135560 -147320
rect 137120 -147380 137140 -147320
rect 138540 -147290 138560 -147230
rect 140120 -147290 140140 -147230
rect 138540 -147320 140140 -147290
rect 138540 -147380 138560 -147320
rect 140120 -147380 140140 -147320
rect 141540 -147290 141560 -147230
rect 143120 -147290 143140 -147230
rect 141540 -147320 143140 -147290
rect 141540 -147380 141560 -147320
rect 143120 -147380 143140 -147320
rect 144540 -147290 144560 -147230
rect 146120 -147290 146140 -147230
rect 144540 -147320 146140 -147290
rect 144540 -147380 144560 -147320
rect 146120 -147380 146140 -147320
rect 147540 -147290 147560 -147230
rect 149120 -147290 149140 -147230
rect 147540 -147320 149140 -147290
rect 147540 -147380 147560 -147320
rect 149120 -147380 149140 -147320
rect 220 -147500 440 -147490
rect 220 -147700 240 -147500
rect 420 -147700 440 -147500
rect 220 -147710 440 -147700
rect 3220 -147500 3440 -147490
rect 3220 -147700 3240 -147500
rect 3420 -147700 3440 -147500
rect 3220 -147710 3440 -147700
rect 6220 -147500 6440 -147490
rect 6220 -147700 6240 -147500
rect 6420 -147700 6440 -147500
rect 6220 -147710 6440 -147700
rect 9220 -147500 9440 -147490
rect 9220 -147700 9240 -147500
rect 9420 -147700 9440 -147500
rect 9220 -147710 9440 -147700
rect 12220 -147500 12440 -147490
rect 12220 -147700 12240 -147500
rect 12420 -147700 12440 -147500
rect 12220 -147710 12440 -147700
rect 15220 -147500 15440 -147490
rect 15220 -147700 15240 -147500
rect 15420 -147700 15440 -147500
rect 15220 -147710 15440 -147700
rect 18220 -147500 18440 -147490
rect 18220 -147700 18240 -147500
rect 18420 -147700 18440 -147500
rect 18220 -147710 18440 -147700
rect 21220 -147500 21440 -147490
rect 21220 -147700 21240 -147500
rect 21420 -147700 21440 -147500
rect 21220 -147710 21440 -147700
rect 24220 -147500 24440 -147490
rect 24220 -147700 24240 -147500
rect 24420 -147700 24440 -147500
rect 24220 -147710 24440 -147700
rect 27220 -147500 27440 -147490
rect 27220 -147700 27240 -147500
rect 27420 -147700 27440 -147500
rect 27220 -147710 27440 -147700
rect 30220 -147500 30440 -147490
rect 30220 -147700 30240 -147500
rect 30420 -147700 30440 -147500
rect 30220 -147710 30440 -147700
rect 33220 -147500 33440 -147490
rect 33220 -147700 33240 -147500
rect 33420 -147700 33440 -147500
rect 33220 -147710 33440 -147700
rect 36220 -147500 36440 -147490
rect 36220 -147700 36240 -147500
rect 36420 -147700 36440 -147500
rect 36220 -147710 36440 -147700
rect 39220 -147500 39440 -147490
rect 39220 -147700 39240 -147500
rect 39420 -147700 39440 -147500
rect 39220 -147710 39440 -147700
rect 42220 -147500 42440 -147490
rect 42220 -147700 42240 -147500
rect 42420 -147700 42440 -147500
rect 42220 -147710 42440 -147700
rect 45220 -147500 45440 -147490
rect 45220 -147700 45240 -147500
rect 45420 -147700 45440 -147500
rect 45220 -147710 45440 -147700
rect 48220 -147500 48440 -147490
rect 48220 -147700 48240 -147500
rect 48420 -147700 48440 -147500
rect 48220 -147710 48440 -147700
rect 51220 -147500 51440 -147490
rect 51220 -147700 51240 -147500
rect 51420 -147700 51440 -147500
rect 51220 -147710 51440 -147700
rect 54220 -147500 54440 -147490
rect 54220 -147700 54240 -147500
rect 54420 -147700 54440 -147500
rect 54220 -147710 54440 -147700
rect 57220 -147500 57440 -147490
rect 57220 -147700 57240 -147500
rect 57420 -147700 57440 -147500
rect 57220 -147710 57440 -147700
rect 60220 -147500 60440 -147490
rect 60220 -147700 60240 -147500
rect 60420 -147700 60440 -147500
rect 60220 -147710 60440 -147700
rect 63220 -147500 63440 -147490
rect 63220 -147700 63240 -147500
rect 63420 -147700 63440 -147500
rect 63220 -147710 63440 -147700
rect 66220 -147500 66440 -147490
rect 66220 -147700 66240 -147500
rect 66420 -147700 66440 -147500
rect 66220 -147710 66440 -147700
rect 69220 -147500 69440 -147490
rect 69220 -147700 69240 -147500
rect 69420 -147700 69440 -147500
rect 69220 -147710 69440 -147700
rect 72220 -147500 72440 -147490
rect 72220 -147700 72240 -147500
rect 72420 -147700 72440 -147500
rect 72220 -147710 72440 -147700
rect 75220 -147500 75440 -147490
rect 75220 -147700 75240 -147500
rect 75420 -147700 75440 -147500
rect 75220 -147710 75440 -147700
rect 78220 -147500 78440 -147490
rect 78220 -147700 78240 -147500
rect 78420 -147700 78440 -147500
rect 78220 -147710 78440 -147700
rect 81220 -147500 81440 -147490
rect 81220 -147700 81240 -147500
rect 81420 -147700 81440 -147500
rect 81220 -147710 81440 -147700
rect 84220 -147500 84440 -147490
rect 84220 -147700 84240 -147500
rect 84420 -147700 84440 -147500
rect 84220 -147710 84440 -147700
rect 87220 -147500 87440 -147490
rect 87220 -147700 87240 -147500
rect 87420 -147700 87440 -147500
rect 87220 -147710 87440 -147700
rect 90220 -147500 90440 -147490
rect 90220 -147700 90240 -147500
rect 90420 -147700 90440 -147500
rect 90220 -147710 90440 -147700
rect 93220 -147500 93440 -147490
rect 93220 -147700 93240 -147500
rect 93420 -147700 93440 -147500
rect 93220 -147710 93440 -147700
rect 96220 -147500 96440 -147490
rect 96220 -147700 96240 -147500
rect 96420 -147700 96440 -147500
rect 96220 -147710 96440 -147700
rect 99220 -147500 99440 -147490
rect 99220 -147700 99240 -147500
rect 99420 -147700 99440 -147500
rect 99220 -147710 99440 -147700
rect 102220 -147500 102440 -147490
rect 102220 -147700 102240 -147500
rect 102420 -147700 102440 -147500
rect 102220 -147710 102440 -147700
rect 105220 -147500 105440 -147490
rect 105220 -147700 105240 -147500
rect 105420 -147700 105440 -147500
rect 105220 -147710 105440 -147700
rect 108220 -147500 108440 -147490
rect 108220 -147700 108240 -147500
rect 108420 -147700 108440 -147500
rect 108220 -147710 108440 -147700
rect 111220 -147500 111440 -147490
rect 111220 -147700 111240 -147500
rect 111420 -147700 111440 -147500
rect 111220 -147710 111440 -147700
rect 114220 -147500 114440 -147490
rect 114220 -147700 114240 -147500
rect 114420 -147700 114440 -147500
rect 114220 -147710 114440 -147700
rect 117220 -147500 117440 -147490
rect 117220 -147700 117240 -147500
rect 117420 -147700 117440 -147500
rect 117220 -147710 117440 -147700
rect 120220 -147500 120440 -147490
rect 120220 -147700 120240 -147500
rect 120420 -147700 120440 -147500
rect 120220 -147710 120440 -147700
rect 123220 -147500 123440 -147490
rect 123220 -147700 123240 -147500
rect 123420 -147700 123440 -147500
rect 123220 -147710 123440 -147700
rect 126220 -147500 126440 -147490
rect 126220 -147700 126240 -147500
rect 126420 -147700 126440 -147500
rect 126220 -147710 126440 -147700
rect 129220 -147500 129440 -147490
rect 129220 -147700 129240 -147500
rect 129420 -147700 129440 -147500
rect 129220 -147710 129440 -147700
rect 132220 -147500 132440 -147490
rect 132220 -147700 132240 -147500
rect 132420 -147700 132440 -147500
rect 132220 -147710 132440 -147700
rect 135220 -147500 135440 -147490
rect 135220 -147700 135240 -147500
rect 135420 -147700 135440 -147500
rect 135220 -147710 135440 -147700
rect 138220 -147500 138440 -147490
rect 138220 -147700 138240 -147500
rect 138420 -147700 138440 -147500
rect 138220 -147710 138440 -147700
rect 141220 -147500 141440 -147490
rect 141220 -147700 141240 -147500
rect 141420 -147700 141440 -147500
rect 141220 -147710 141440 -147700
rect 144220 -147500 144440 -147490
rect 144220 -147700 144240 -147500
rect 144420 -147700 144440 -147500
rect 144220 -147710 144440 -147700
rect 147220 -147500 147440 -147490
rect 147220 -147700 147240 -147500
rect 147420 -147700 147440 -147500
rect 147220 -147710 147440 -147700
rect 540 -147830 2140 -147800
rect 540 -147870 560 -147830
rect 2120 -147870 2140 -147830
rect 540 -147920 2140 -147870
rect 540 -147980 560 -147920
rect 2120 -147980 2140 -147920
rect 540 -148000 2140 -147980
rect 3540 -147830 5140 -147800
rect 3540 -147870 3560 -147830
rect 5120 -147870 5140 -147830
rect 3540 -147920 5140 -147870
rect 3540 -147980 3560 -147920
rect 5120 -147980 5140 -147920
rect 3540 -148000 5140 -147980
rect 6540 -147830 8140 -147800
rect 6540 -147870 6560 -147830
rect 8120 -147870 8140 -147830
rect 6540 -147920 8140 -147870
rect 6540 -147980 6560 -147920
rect 8120 -147980 8140 -147920
rect 6540 -148000 8140 -147980
rect 9540 -147830 11140 -147800
rect 9540 -147870 9560 -147830
rect 11120 -147870 11140 -147830
rect 9540 -147920 11140 -147870
rect 9540 -147980 9560 -147920
rect 11120 -147980 11140 -147920
rect 9540 -148000 11140 -147980
rect 12540 -147830 14140 -147800
rect 12540 -147870 12560 -147830
rect 14120 -147870 14140 -147830
rect 12540 -147920 14140 -147870
rect 12540 -147980 12560 -147920
rect 14120 -147980 14140 -147920
rect 12540 -148000 14140 -147980
rect 15540 -147830 17140 -147800
rect 15540 -147870 15560 -147830
rect 17120 -147870 17140 -147830
rect 15540 -147920 17140 -147870
rect 15540 -147980 15560 -147920
rect 17120 -147980 17140 -147920
rect 15540 -148000 17140 -147980
rect 18540 -147830 20140 -147800
rect 18540 -147870 18560 -147830
rect 20120 -147870 20140 -147830
rect 18540 -147920 20140 -147870
rect 18540 -147980 18560 -147920
rect 20120 -147980 20140 -147920
rect 18540 -148000 20140 -147980
rect 21540 -147830 23140 -147800
rect 21540 -147870 21560 -147830
rect 23120 -147870 23140 -147830
rect 21540 -147920 23140 -147870
rect 21540 -147980 21560 -147920
rect 23120 -147980 23140 -147920
rect 21540 -148000 23140 -147980
rect 24540 -147830 26140 -147800
rect 24540 -147870 24560 -147830
rect 26120 -147870 26140 -147830
rect 24540 -147920 26140 -147870
rect 24540 -147980 24560 -147920
rect 26120 -147980 26140 -147920
rect 24540 -148000 26140 -147980
rect 27540 -147830 29140 -147800
rect 27540 -147870 27560 -147830
rect 29120 -147870 29140 -147830
rect 27540 -147920 29140 -147870
rect 27540 -147980 27560 -147920
rect 29120 -147980 29140 -147920
rect 27540 -148000 29140 -147980
rect 30540 -147830 32140 -147800
rect 30540 -147870 30560 -147830
rect 32120 -147870 32140 -147830
rect 30540 -147920 32140 -147870
rect 30540 -147980 30560 -147920
rect 32120 -147980 32140 -147920
rect 30540 -148000 32140 -147980
rect 33540 -147830 35140 -147800
rect 33540 -147870 33560 -147830
rect 35120 -147870 35140 -147830
rect 33540 -147920 35140 -147870
rect 33540 -147980 33560 -147920
rect 35120 -147980 35140 -147920
rect 33540 -148000 35140 -147980
rect 36540 -147830 38140 -147800
rect 36540 -147870 36560 -147830
rect 38120 -147870 38140 -147830
rect 36540 -147920 38140 -147870
rect 36540 -147980 36560 -147920
rect 38120 -147980 38140 -147920
rect 36540 -148000 38140 -147980
rect 39540 -147830 41140 -147800
rect 39540 -147870 39560 -147830
rect 41120 -147870 41140 -147830
rect 39540 -147920 41140 -147870
rect 39540 -147980 39560 -147920
rect 41120 -147980 41140 -147920
rect 39540 -148000 41140 -147980
rect 42540 -147830 44140 -147800
rect 42540 -147870 42560 -147830
rect 44120 -147870 44140 -147830
rect 42540 -147920 44140 -147870
rect 42540 -147980 42560 -147920
rect 44120 -147980 44140 -147920
rect 42540 -148000 44140 -147980
rect 45540 -147830 47140 -147800
rect 45540 -147870 45560 -147830
rect 47120 -147870 47140 -147830
rect 45540 -147920 47140 -147870
rect 45540 -147980 45560 -147920
rect 47120 -147980 47140 -147920
rect 45540 -148000 47140 -147980
rect 48540 -147830 50140 -147800
rect 48540 -147870 48560 -147830
rect 50120 -147870 50140 -147830
rect 48540 -147920 50140 -147870
rect 48540 -147980 48560 -147920
rect 50120 -147980 50140 -147920
rect 48540 -148000 50140 -147980
rect 51540 -147830 53140 -147800
rect 51540 -147870 51560 -147830
rect 53120 -147870 53140 -147830
rect 51540 -147920 53140 -147870
rect 51540 -147980 51560 -147920
rect 53120 -147980 53140 -147920
rect 51540 -148000 53140 -147980
rect 54540 -147830 56140 -147800
rect 54540 -147870 54560 -147830
rect 56120 -147870 56140 -147830
rect 54540 -147920 56140 -147870
rect 54540 -147980 54560 -147920
rect 56120 -147980 56140 -147920
rect 54540 -148000 56140 -147980
rect 57540 -147830 59140 -147800
rect 57540 -147870 57560 -147830
rect 59120 -147870 59140 -147830
rect 57540 -147920 59140 -147870
rect 57540 -147980 57560 -147920
rect 59120 -147980 59140 -147920
rect 57540 -148000 59140 -147980
rect 60540 -147830 62140 -147800
rect 60540 -147870 60560 -147830
rect 62120 -147870 62140 -147830
rect 60540 -147920 62140 -147870
rect 60540 -147980 60560 -147920
rect 62120 -147980 62140 -147920
rect 60540 -148000 62140 -147980
rect 63540 -147830 65140 -147800
rect 63540 -147870 63560 -147830
rect 65120 -147870 65140 -147830
rect 63540 -147920 65140 -147870
rect 63540 -147980 63560 -147920
rect 65120 -147980 65140 -147920
rect 63540 -148000 65140 -147980
rect 66540 -147830 68140 -147800
rect 66540 -147870 66560 -147830
rect 68120 -147870 68140 -147830
rect 66540 -147920 68140 -147870
rect 66540 -147980 66560 -147920
rect 68120 -147980 68140 -147920
rect 66540 -148000 68140 -147980
rect 69540 -147830 71140 -147800
rect 69540 -147870 69560 -147830
rect 71120 -147870 71140 -147830
rect 69540 -147920 71140 -147870
rect 69540 -147980 69560 -147920
rect 71120 -147980 71140 -147920
rect 69540 -148000 71140 -147980
rect 72540 -147830 74140 -147800
rect 72540 -147870 72560 -147830
rect 74120 -147870 74140 -147830
rect 72540 -147920 74140 -147870
rect 72540 -147980 72560 -147920
rect 74120 -147980 74140 -147920
rect 72540 -148000 74140 -147980
rect 75540 -147830 77140 -147800
rect 75540 -147870 75560 -147830
rect 77120 -147870 77140 -147830
rect 75540 -147920 77140 -147870
rect 75540 -147980 75560 -147920
rect 77120 -147980 77140 -147920
rect 75540 -148000 77140 -147980
rect 78540 -147830 80140 -147800
rect 78540 -147870 78560 -147830
rect 80120 -147870 80140 -147830
rect 78540 -147920 80140 -147870
rect 78540 -147980 78560 -147920
rect 80120 -147980 80140 -147920
rect 78540 -148000 80140 -147980
rect 81540 -147830 83140 -147800
rect 81540 -147870 81560 -147830
rect 83120 -147870 83140 -147830
rect 81540 -147920 83140 -147870
rect 81540 -147980 81560 -147920
rect 83120 -147980 83140 -147920
rect 81540 -148000 83140 -147980
rect 84540 -147830 86140 -147800
rect 84540 -147870 84560 -147830
rect 86120 -147870 86140 -147830
rect 84540 -147920 86140 -147870
rect 84540 -147980 84560 -147920
rect 86120 -147980 86140 -147920
rect 84540 -148000 86140 -147980
rect 87540 -147830 89140 -147800
rect 87540 -147870 87560 -147830
rect 89120 -147870 89140 -147830
rect 87540 -147920 89140 -147870
rect 87540 -147980 87560 -147920
rect 89120 -147980 89140 -147920
rect 87540 -148000 89140 -147980
rect 90540 -147830 92140 -147800
rect 90540 -147870 90560 -147830
rect 92120 -147870 92140 -147830
rect 90540 -147920 92140 -147870
rect 90540 -147980 90560 -147920
rect 92120 -147980 92140 -147920
rect 90540 -148000 92140 -147980
rect 93540 -147830 95140 -147800
rect 93540 -147870 93560 -147830
rect 95120 -147870 95140 -147830
rect 93540 -147920 95140 -147870
rect 93540 -147980 93560 -147920
rect 95120 -147980 95140 -147920
rect 93540 -148000 95140 -147980
rect 96540 -147830 98140 -147800
rect 96540 -147870 96560 -147830
rect 98120 -147870 98140 -147830
rect 96540 -147920 98140 -147870
rect 96540 -147980 96560 -147920
rect 98120 -147980 98140 -147920
rect 96540 -148000 98140 -147980
rect 99540 -147830 101140 -147800
rect 99540 -147870 99560 -147830
rect 101120 -147870 101140 -147830
rect 99540 -147920 101140 -147870
rect 99540 -147980 99560 -147920
rect 101120 -147980 101140 -147920
rect 99540 -148000 101140 -147980
rect 102540 -147830 104140 -147800
rect 102540 -147870 102560 -147830
rect 104120 -147870 104140 -147830
rect 102540 -147920 104140 -147870
rect 102540 -147980 102560 -147920
rect 104120 -147980 104140 -147920
rect 102540 -148000 104140 -147980
rect 105540 -147830 107140 -147800
rect 105540 -147870 105560 -147830
rect 107120 -147870 107140 -147830
rect 105540 -147920 107140 -147870
rect 105540 -147980 105560 -147920
rect 107120 -147980 107140 -147920
rect 105540 -148000 107140 -147980
rect 108540 -147830 110140 -147800
rect 108540 -147870 108560 -147830
rect 110120 -147870 110140 -147830
rect 108540 -147920 110140 -147870
rect 108540 -147980 108560 -147920
rect 110120 -147980 110140 -147920
rect 108540 -148000 110140 -147980
rect 111540 -147830 113140 -147800
rect 111540 -147870 111560 -147830
rect 113120 -147870 113140 -147830
rect 111540 -147920 113140 -147870
rect 111540 -147980 111560 -147920
rect 113120 -147980 113140 -147920
rect 111540 -148000 113140 -147980
rect 114540 -147830 116140 -147800
rect 114540 -147870 114560 -147830
rect 116120 -147870 116140 -147830
rect 114540 -147920 116140 -147870
rect 114540 -147980 114560 -147920
rect 116120 -147980 116140 -147920
rect 114540 -148000 116140 -147980
rect 117540 -147830 119140 -147800
rect 117540 -147870 117560 -147830
rect 119120 -147870 119140 -147830
rect 117540 -147920 119140 -147870
rect 117540 -147980 117560 -147920
rect 119120 -147980 119140 -147920
rect 117540 -148000 119140 -147980
rect 120540 -147830 122140 -147800
rect 120540 -147870 120560 -147830
rect 122120 -147870 122140 -147830
rect 120540 -147920 122140 -147870
rect 120540 -147980 120560 -147920
rect 122120 -147980 122140 -147920
rect 120540 -148000 122140 -147980
rect 123540 -147830 125140 -147800
rect 123540 -147870 123560 -147830
rect 125120 -147870 125140 -147830
rect 123540 -147920 125140 -147870
rect 123540 -147980 123560 -147920
rect 125120 -147980 125140 -147920
rect 123540 -148000 125140 -147980
rect 126540 -147830 128140 -147800
rect 126540 -147870 126560 -147830
rect 128120 -147870 128140 -147830
rect 126540 -147920 128140 -147870
rect 126540 -147980 126560 -147920
rect 128120 -147980 128140 -147920
rect 126540 -148000 128140 -147980
rect 129540 -147830 131140 -147800
rect 129540 -147870 129560 -147830
rect 131120 -147870 131140 -147830
rect 129540 -147920 131140 -147870
rect 129540 -147980 129560 -147920
rect 131120 -147980 131140 -147920
rect 129540 -148000 131140 -147980
rect 132540 -147830 134140 -147800
rect 132540 -147870 132560 -147830
rect 134120 -147870 134140 -147830
rect 132540 -147920 134140 -147870
rect 132540 -147980 132560 -147920
rect 134120 -147980 134140 -147920
rect 132540 -148000 134140 -147980
rect 135540 -147830 137140 -147800
rect 135540 -147870 135560 -147830
rect 137120 -147870 137140 -147830
rect 135540 -147920 137140 -147870
rect 135540 -147980 135560 -147920
rect 137120 -147980 137140 -147920
rect 135540 -148000 137140 -147980
rect 138540 -147830 140140 -147800
rect 138540 -147870 138560 -147830
rect 140120 -147870 140140 -147830
rect 138540 -147920 140140 -147870
rect 138540 -147980 138560 -147920
rect 140120 -147980 140140 -147920
rect 138540 -148000 140140 -147980
rect 141540 -147830 143140 -147800
rect 141540 -147870 141560 -147830
rect 143120 -147870 143140 -147830
rect 141540 -147920 143140 -147870
rect 141540 -147980 141560 -147920
rect 143120 -147980 143140 -147920
rect 141540 -148000 143140 -147980
rect 144540 -147830 146140 -147800
rect 144540 -147870 144560 -147830
rect 146120 -147870 146140 -147830
rect 144540 -147920 146140 -147870
rect 144540 -147980 144560 -147920
rect 146120 -147980 146140 -147920
rect 144540 -148000 146140 -147980
rect 147540 -147830 149140 -147800
rect 147540 -147870 147560 -147830
rect 149120 -147870 149140 -147830
rect 147540 -147920 149140 -147870
rect 147540 -147980 147560 -147920
rect 149120 -147980 149140 -147920
rect 147540 -148000 149140 -147980
<< viali >>
rect 560 -147290 2120 -147230
rect 3560 -147290 5120 -147230
rect 6560 -147290 8120 -147230
rect 9560 -147290 11120 -147230
rect 12560 -147290 14120 -147230
rect 15560 -147290 17120 -147230
rect 18560 -147290 20120 -147230
rect 21560 -147290 23120 -147230
rect 24560 -147290 26120 -147230
rect 27560 -147290 29120 -147230
rect 30560 -147290 32120 -147230
rect 33560 -147290 35120 -147230
rect 36560 -147290 38120 -147230
rect 39560 -147290 41120 -147230
rect 42560 -147290 44120 -147230
rect 45560 -147290 47120 -147230
rect 48560 -147290 50120 -147230
rect 51560 -147290 53120 -147230
rect 54560 -147290 56120 -147230
rect 57560 -147290 59120 -147230
rect 60560 -147290 62120 -147230
rect 63560 -147290 65120 -147230
rect 66560 -147290 68120 -147230
rect 69560 -147290 71120 -147230
rect 72560 -147290 74120 -147230
rect 75560 -147290 77120 -147230
rect 78560 -147290 80120 -147230
rect 81560 -147290 83120 -147230
rect 84560 -147290 86120 -147230
rect 87560 -147290 89120 -147230
rect 90560 -147290 92120 -147230
rect 93560 -147290 95120 -147230
rect 96560 -147290 98120 -147230
rect 99560 -147290 101120 -147230
rect 102560 -147290 104120 -147230
rect 105560 -147290 107120 -147230
rect 108560 -147290 110120 -147230
rect 111560 -147290 113120 -147230
rect 114560 -147290 116120 -147230
rect 117560 -147290 119120 -147230
rect 120560 -147290 122120 -147230
rect 123560 -147290 125120 -147230
rect 126560 -147290 128120 -147230
rect 129560 -147290 131120 -147230
rect 132560 -147290 134120 -147230
rect 135560 -147290 137120 -147230
rect 138560 -147290 140120 -147230
rect 141560 -147290 143120 -147230
rect 144560 -147290 146120 -147230
rect 147560 -147290 149120 -147230
rect 240 -147700 420 -147500
rect 3240 -147700 3420 -147500
rect 6240 -147700 6420 -147500
rect 9240 -147700 9420 -147500
rect 12240 -147700 12420 -147500
rect 15240 -147700 15420 -147500
rect 18240 -147700 18420 -147500
rect 21240 -147700 21420 -147500
rect 24240 -147700 24420 -147500
rect 27240 -147700 27420 -147500
rect 30240 -147700 30420 -147500
rect 33240 -147700 33420 -147500
rect 36240 -147700 36420 -147500
rect 39240 -147700 39420 -147500
rect 42240 -147700 42420 -147500
rect 45240 -147700 45420 -147500
rect 48240 -147700 48420 -147500
rect 51240 -147700 51420 -147500
rect 54240 -147700 54420 -147500
rect 57240 -147700 57420 -147500
rect 60240 -147700 60420 -147500
rect 63240 -147700 63420 -147500
rect 66240 -147700 66420 -147500
rect 69240 -147700 69420 -147500
rect 72240 -147700 72420 -147500
rect 75240 -147700 75420 -147500
rect 78240 -147700 78420 -147500
rect 81240 -147700 81420 -147500
rect 84240 -147700 84420 -147500
rect 87240 -147700 87420 -147500
rect 90240 -147700 90420 -147500
rect 93240 -147700 93420 -147500
rect 96240 -147700 96420 -147500
rect 99240 -147700 99420 -147500
rect 102240 -147700 102420 -147500
rect 105240 -147700 105420 -147500
rect 108240 -147700 108420 -147500
rect 111240 -147700 111420 -147500
rect 114240 -147700 114420 -147500
rect 117240 -147700 117420 -147500
rect 120240 -147700 120420 -147500
rect 123240 -147700 123420 -147500
rect 126240 -147700 126420 -147500
rect 129240 -147700 129420 -147500
rect 132240 -147700 132420 -147500
rect 135240 -147700 135420 -147500
rect 138240 -147700 138420 -147500
rect 141240 -147700 141420 -147500
rect 144240 -147700 144420 -147500
rect 147240 -147700 147420 -147500
rect 560 -147980 2120 -147920
rect 3560 -147980 5120 -147920
rect 6560 -147980 8120 -147920
rect 9560 -147980 11120 -147920
rect 12560 -147980 14120 -147920
rect 15560 -147980 17120 -147920
rect 18560 -147980 20120 -147920
rect 21560 -147980 23120 -147920
rect 24560 -147980 26120 -147920
rect 27560 -147980 29120 -147920
rect 30560 -147980 32120 -147920
rect 33560 -147980 35120 -147920
rect 36560 -147980 38120 -147920
rect 39560 -147980 41120 -147920
rect 42560 -147980 44120 -147920
rect 45560 -147980 47120 -147920
rect 48560 -147980 50120 -147920
rect 51560 -147980 53120 -147920
rect 54560 -147980 56120 -147920
rect 57560 -147980 59120 -147920
rect 60560 -147980 62120 -147920
rect 63560 -147980 65120 -147920
rect 66560 -147980 68120 -147920
rect 69560 -147980 71120 -147920
rect 72560 -147980 74120 -147920
rect 75560 -147980 77120 -147920
rect 78560 -147980 80120 -147920
rect 81560 -147980 83120 -147920
rect 84560 -147980 86120 -147920
rect 87560 -147980 89120 -147920
rect 90560 -147980 92120 -147920
rect 93560 -147980 95120 -147920
rect 96560 -147980 98120 -147920
rect 99560 -147980 101120 -147920
rect 102560 -147980 104120 -147920
rect 105560 -147980 107120 -147920
rect 108560 -147980 110120 -147920
rect 111560 -147980 113120 -147920
rect 114560 -147980 116120 -147920
rect 117560 -147980 119120 -147920
rect 120560 -147980 122120 -147920
rect 123560 -147980 125120 -147920
rect 126560 -147980 128120 -147920
rect 129560 -147980 131120 -147920
rect 132560 -147980 134120 -147920
rect 135560 -147980 137120 -147920
rect 138560 -147980 140120 -147920
rect 141560 -147980 143120 -147920
rect 144560 -147980 146120 -147920
rect 147560 -147980 149120 -147920
<< metal1 >>
rect -1940 3450 149000 3460
rect -1940 3360 -1920 3450
rect -900 3360 50 3450
rect 140 3360 3050 3450
rect 3140 3360 6050 3450
rect 6140 3360 9050 3450
rect 9140 3360 12050 3450
rect 12140 3360 15050 3450
rect 15140 3360 18050 3450
rect 18140 3360 21050 3450
rect 21140 3360 24050 3450
rect 24140 3360 27050 3450
rect 27140 3360 30050 3450
rect 30140 3360 33050 3450
rect 33140 3360 36050 3450
rect 36140 3360 39050 3450
rect 39140 3360 42050 3450
rect 42140 3360 45050 3450
rect 45140 3360 48050 3450
rect 48140 3360 51050 3450
rect 51140 3360 54050 3450
rect 54140 3360 57050 3450
rect 57140 3360 60050 3450
rect 60140 3360 63050 3450
rect 63140 3360 66050 3450
rect 66140 3360 69050 3450
rect 69140 3360 72050 3450
rect 72140 3360 75050 3450
rect 75140 3360 78050 3450
rect 78140 3360 81050 3450
rect 81140 3360 84050 3450
rect 84140 3360 87050 3450
rect 87140 3360 90050 3450
rect 90140 3360 93050 3450
rect 93140 3360 96050 3450
rect 96140 3360 99050 3450
rect 99140 3360 102050 3450
rect 102140 3360 105050 3450
rect 105140 3360 108050 3450
rect 108140 3360 111050 3450
rect 111140 3360 114050 3450
rect 114140 3360 117050 3450
rect 117140 3360 120050 3450
rect 120140 3360 123050 3450
rect 123140 3360 126050 3450
rect 126140 3360 129050 3450
rect 129140 3360 132050 3450
rect 132140 3360 135050 3450
rect 135140 3360 138050 3450
rect 138140 3360 141050 3450
rect 141140 3360 144050 3450
rect 144140 3360 147050 3450
rect 147140 3360 149000 3450
rect -1940 3350 149000 3360
rect -2000 2970 -1800 3000
rect -2000 2820 0 2970
rect -2000 -30 -1800 2820
rect -1600 1560 0 1570
rect -1600 1490 -1580 1560
rect -1180 1490 -540 1560
rect -260 1490 0 1560
rect -1600 1480 0 1490
rect 150400 180 150600 3030
rect 150000 30 150600 180
rect -2000 -180 0 -30
rect -2000 -3030 -1800 -180
rect -1600 -1440 0 -1430
rect -1600 -1510 -1580 -1440
rect -1180 -1510 -540 -1440
rect -260 -1510 0 -1440
rect -1600 -1520 0 -1510
rect 150400 -2820 150600 30
rect 150000 -2970 150600 -2820
rect -2000 -3180 0 -3030
rect -2000 -6030 -1800 -3180
rect -1600 -4440 0 -4430
rect -1600 -4510 -1580 -4440
rect -1180 -4510 -540 -4440
rect -260 -4510 0 -4440
rect -1600 -4520 0 -4510
rect 150400 -5820 150600 -2970
rect 150000 -5970 150600 -5820
rect -2000 -6180 0 -6030
rect -2000 -9030 -1800 -6180
rect -1600 -7440 0 -7430
rect -1600 -7510 -1580 -7440
rect -1180 -7510 -540 -7440
rect -260 -7510 0 -7440
rect -1600 -7520 0 -7510
rect 150400 -8820 150600 -5970
rect 150000 -8970 150600 -8820
rect -2000 -9180 0 -9030
rect -2000 -12030 -1800 -9180
rect -1600 -10440 0 -10430
rect -1600 -10510 -1580 -10440
rect -1180 -10510 -540 -10440
rect -260 -10510 0 -10440
rect -1600 -10520 0 -10510
rect 150400 -11820 150600 -8970
rect 150000 -11970 150600 -11820
rect -2000 -12180 0 -12030
rect -2000 -15030 -1800 -12180
rect -1600 -13440 0 -13430
rect -1600 -13510 -1580 -13440
rect -1180 -13510 -540 -13440
rect -260 -13510 0 -13440
rect -1600 -13520 0 -13510
rect 150400 -14820 150600 -11970
rect 150000 -14970 150600 -14820
rect -2000 -15180 0 -15030
rect -2000 -18030 -1800 -15180
rect -1600 -16440 0 -16430
rect -1600 -16510 -1580 -16440
rect -1180 -16510 -540 -16440
rect -260 -16510 0 -16440
rect -1600 -16520 0 -16510
rect 150400 -17820 150600 -14970
rect 150000 -17970 150600 -17820
rect -2000 -18180 0 -18030
rect -2000 -21030 -1800 -18180
rect -1600 -19440 0 -19430
rect -1600 -19510 -1580 -19440
rect -1180 -19510 -540 -19440
rect -260 -19510 0 -19440
rect -1600 -19520 0 -19510
rect 150400 -20820 150600 -17970
rect 150000 -20970 150600 -20820
rect -2000 -21180 0 -21030
rect -2000 -24030 -1800 -21180
rect -1600 -22440 0 -22430
rect -1600 -22510 -1580 -22440
rect -1180 -22510 -540 -22440
rect -260 -22510 0 -22440
rect -1600 -22520 0 -22510
rect 150400 -23820 150600 -20970
rect 150000 -23970 150600 -23820
rect -2000 -24180 0 -24030
rect -2000 -27030 -1800 -24180
rect -1600 -25440 0 -25430
rect -1600 -25510 -1580 -25440
rect -1180 -25510 -540 -25440
rect -260 -25510 0 -25440
rect -1600 -25520 0 -25510
rect 150400 -26820 150600 -23970
rect 150000 -26970 150600 -26820
rect -2000 -27180 0 -27030
rect -2000 -30030 -1800 -27180
rect -1600 -28440 0 -28430
rect -1600 -28510 -1580 -28440
rect -1180 -28510 -540 -28440
rect -260 -28510 0 -28440
rect -1600 -28520 0 -28510
rect 150400 -29820 150600 -26970
rect 150000 -29970 150600 -29820
rect -2000 -30180 0 -30030
rect -2000 -33030 -1800 -30180
rect -1600 -31440 0 -31430
rect -1600 -31510 -1580 -31440
rect -1180 -31510 -540 -31440
rect -260 -31510 0 -31440
rect -1600 -31520 0 -31510
rect 150400 -32820 150600 -29970
rect 150000 -32970 150600 -32820
rect -2000 -33180 0 -33030
rect -2000 -36030 -1800 -33180
rect -1600 -34440 0 -34430
rect -1600 -34510 -1580 -34440
rect -1180 -34510 -540 -34440
rect -260 -34510 0 -34440
rect -1600 -34520 0 -34510
rect 150400 -35820 150600 -32970
rect 150000 -35970 150600 -35820
rect -2000 -36180 0 -36030
rect -2000 -39030 -1800 -36180
rect -1600 -37440 0 -37430
rect -1600 -37510 -1580 -37440
rect -1180 -37510 -540 -37440
rect -260 -37510 0 -37440
rect -1600 -37520 0 -37510
rect 150400 -38820 150600 -35970
rect 150000 -38970 150600 -38820
rect -2000 -39180 0 -39030
rect -2000 -42030 -1800 -39180
rect -1600 -40440 0 -40430
rect -1600 -40510 -1580 -40440
rect -1180 -40510 -540 -40440
rect -260 -40510 0 -40440
rect -1600 -40520 0 -40510
rect 150400 -41820 150600 -38970
rect 150000 -41970 150600 -41820
rect -2000 -42180 0 -42030
rect -2000 -45030 -1800 -42180
rect -1600 -43440 0 -43430
rect -1600 -43510 -1580 -43440
rect -1180 -43510 -540 -43440
rect -260 -43510 0 -43440
rect -1600 -43520 0 -43510
rect 150400 -44820 150600 -41970
rect 150000 -44970 150600 -44820
rect -2000 -45180 0 -45030
rect -2000 -48030 -1800 -45180
rect -1600 -46440 0 -46430
rect -1600 -46510 -1580 -46440
rect -1180 -46510 -540 -46440
rect -260 -46510 0 -46440
rect -1600 -46520 0 -46510
rect 150400 -47820 150600 -44970
rect 150000 -47970 150600 -47820
rect -2000 -48180 0 -48030
rect -2000 -51030 -1800 -48180
rect -1600 -49440 0 -49430
rect -1600 -49510 -1580 -49440
rect -1180 -49510 -540 -49440
rect -260 -49510 0 -49440
rect -1600 -49520 0 -49510
rect 150400 -50820 150600 -47970
rect 150000 -50970 150600 -50820
rect -2000 -51180 0 -51030
rect -2000 -54030 -1800 -51180
rect -1600 -52440 0 -52430
rect -1600 -52510 -1580 -52440
rect -1180 -52510 -540 -52440
rect -260 -52510 0 -52440
rect -1600 -52520 0 -52510
rect 150400 -53820 150600 -50970
rect 150000 -53970 150600 -53820
rect -2000 -54180 0 -54030
rect -2000 -57030 -1800 -54180
rect -1600 -55440 0 -55430
rect -1600 -55510 -1580 -55440
rect -1180 -55510 -540 -55440
rect -260 -55510 0 -55440
rect -1600 -55520 0 -55510
rect 150400 -56820 150600 -53970
rect 150000 -56970 150600 -56820
rect -2000 -57180 0 -57030
rect -2000 -60030 -1800 -57180
rect -1600 -58440 0 -58430
rect -1600 -58510 -1580 -58440
rect -1180 -58510 -540 -58440
rect -260 -58510 0 -58440
rect -1600 -58520 0 -58510
rect 150400 -59820 150600 -56970
rect 150000 -59970 150600 -59820
rect -2000 -60180 0 -60030
rect -2000 -63030 -1800 -60180
rect -1600 -61440 0 -61430
rect -1600 -61510 -1580 -61440
rect -1180 -61510 -540 -61440
rect -260 -61510 0 -61440
rect -1600 -61520 0 -61510
rect 150400 -62820 150600 -59970
rect 150000 -62970 150600 -62820
rect -2000 -63180 0 -63030
rect -2000 -66030 -1800 -63180
rect -1600 -64440 0 -64430
rect -1600 -64510 -1580 -64440
rect -1180 -64510 -540 -64440
rect -260 -64510 0 -64440
rect -1600 -64520 0 -64510
rect 150400 -65820 150600 -62970
rect 150000 -65970 150600 -65820
rect -2000 -66180 0 -66030
rect -2000 -69030 -1800 -66180
rect -1600 -67440 0 -67430
rect -1600 -67510 -1580 -67440
rect -1180 -67510 -540 -67440
rect -260 -67510 0 -67440
rect -1600 -67520 0 -67510
rect 150400 -68820 150600 -65970
rect 150000 -68970 150600 -68820
rect -2000 -69180 0 -69030
rect -2000 -72030 -1800 -69180
rect -1600 -70440 0 -70430
rect -1600 -70510 -1580 -70440
rect -1180 -70510 -540 -70440
rect -260 -70510 0 -70440
rect -1600 -70520 0 -70510
rect 150400 -71820 150600 -68970
rect 150000 -71970 150600 -71820
rect -2000 -72180 0 -72030
rect -2000 -75030 -1800 -72180
rect -1600 -73440 0 -73430
rect -1600 -73510 -1580 -73440
rect -1180 -73510 -540 -73440
rect -260 -73510 0 -73440
rect -1600 -73520 0 -73510
rect 150400 -74820 150600 -71970
rect 150000 -74970 150600 -74820
rect -2000 -75180 0 -75030
rect -2000 -78030 -1800 -75180
rect -1600 -76440 0 -76430
rect -1600 -76510 -1580 -76440
rect -1180 -76510 -540 -76440
rect -260 -76510 0 -76440
rect -1600 -76520 0 -76510
rect 150400 -77820 150600 -74970
rect 150000 -77970 150600 -77820
rect -2000 -78180 0 -78030
rect -2000 -81030 -1800 -78180
rect -1600 -79440 0 -79430
rect -1600 -79510 -1580 -79440
rect -1180 -79510 -540 -79440
rect -260 -79510 0 -79440
rect -1600 -79520 0 -79510
rect 150400 -80820 150600 -77970
rect 150000 -80970 150600 -80820
rect -2000 -81180 0 -81030
rect -2000 -84030 -1800 -81180
rect -1600 -82440 0 -82430
rect -1600 -82510 -1580 -82440
rect -1180 -82510 -540 -82440
rect -260 -82510 0 -82440
rect -1600 -82520 0 -82510
rect 150400 -83820 150600 -80970
rect 150000 -83970 150600 -83820
rect -2000 -84180 0 -84030
rect -2000 -87030 -1800 -84180
rect -1600 -85440 0 -85430
rect -1600 -85510 -1580 -85440
rect -1180 -85510 -540 -85440
rect -260 -85510 0 -85440
rect -1600 -85520 0 -85510
rect 150400 -86820 150600 -83970
rect 150000 -86970 150600 -86820
rect -2000 -87180 0 -87030
rect -2000 -90030 -1800 -87180
rect -1600 -88440 0 -88430
rect -1600 -88510 -1580 -88440
rect -1180 -88510 -540 -88440
rect -260 -88510 0 -88440
rect -1600 -88520 0 -88510
rect 150400 -89820 150600 -86970
rect 150000 -89970 150600 -89820
rect -2000 -90180 0 -90030
rect -2000 -93030 -1800 -90180
rect -1600 -91440 0 -91430
rect -1600 -91510 -1580 -91440
rect -1180 -91510 -540 -91440
rect -260 -91510 0 -91440
rect -1600 -91520 0 -91510
rect 150400 -92820 150600 -89970
rect 150000 -92970 150600 -92820
rect -2000 -93180 0 -93030
rect -2000 -96030 -1800 -93180
rect -1600 -94440 0 -94430
rect -1600 -94510 -1580 -94440
rect -1180 -94510 -540 -94440
rect -260 -94510 0 -94440
rect -1600 -94520 0 -94510
rect 150400 -95820 150600 -92970
rect 150000 -95970 150600 -95820
rect -2000 -96180 0 -96030
rect -2000 -99030 -1800 -96180
rect -1600 -97440 0 -97430
rect -1600 -97510 -1580 -97440
rect -1180 -97510 -540 -97440
rect -260 -97510 0 -97440
rect -1600 -97520 0 -97510
rect 150400 -98820 150600 -95970
rect 150000 -98970 150600 -98820
rect -2000 -99180 0 -99030
rect -2000 -102030 -1800 -99180
rect -1600 -100440 0 -100430
rect -1600 -100510 -1580 -100440
rect -1180 -100510 -540 -100440
rect -260 -100510 0 -100440
rect -1600 -100520 0 -100510
rect 150400 -101820 150600 -98970
rect 150000 -101970 150600 -101820
rect -2000 -102180 0 -102030
rect -2000 -105030 -1800 -102180
rect -1600 -103440 0 -103430
rect -1600 -103510 -1580 -103440
rect -1180 -103510 -540 -103440
rect -260 -103510 0 -103440
rect -1600 -103520 0 -103510
rect 150400 -104820 150600 -101970
rect 150000 -104970 150600 -104820
rect -2000 -105180 0 -105030
rect -2000 -108030 -1800 -105180
rect -1600 -106440 0 -106430
rect -1600 -106510 -1580 -106440
rect -1180 -106510 -540 -106440
rect -260 -106510 0 -106440
rect -1600 -106520 0 -106510
rect 150400 -107820 150600 -104970
rect 150000 -107970 150600 -107820
rect -2000 -108180 0 -108030
rect -2000 -111030 -1800 -108180
rect -1600 -109440 0 -109430
rect -1600 -109510 -1580 -109440
rect -1180 -109510 -540 -109440
rect -260 -109510 0 -109440
rect -1600 -109520 0 -109510
rect 150400 -110820 150600 -107970
rect 150000 -110970 150600 -110820
rect -2000 -111180 0 -111030
rect -2000 -114030 -1800 -111180
rect -1600 -112440 0 -112430
rect -1600 -112510 -1580 -112440
rect -1180 -112510 -540 -112440
rect -260 -112510 0 -112440
rect -1600 -112520 0 -112510
rect 150400 -113820 150600 -110970
rect 150000 -113970 150600 -113820
rect -2000 -114180 0 -114030
rect -2000 -117030 -1800 -114180
rect -1600 -115440 0 -115430
rect -1600 -115510 -1580 -115440
rect -1180 -115510 -540 -115440
rect -260 -115510 0 -115440
rect -1600 -115520 0 -115510
rect 150400 -116820 150600 -113970
rect 150000 -116970 150600 -116820
rect -2000 -117180 0 -117030
rect -2000 -120030 -1800 -117180
rect -1600 -118440 0 -118430
rect -1600 -118510 -1580 -118440
rect -1180 -118510 -540 -118440
rect -260 -118510 0 -118440
rect -1600 -118520 0 -118510
rect 150400 -119820 150600 -116970
rect 150000 -119970 150600 -119820
rect -2000 -120180 0 -120030
rect -2000 -123030 -1800 -120180
rect -1600 -121440 0 -121430
rect -1600 -121510 -1580 -121440
rect -1180 -121510 -540 -121440
rect -260 -121510 0 -121440
rect -1600 -121520 0 -121510
rect 150400 -122820 150600 -119970
rect 150000 -122970 150600 -122820
rect -2000 -123180 0 -123030
rect -2000 -126030 -1800 -123180
rect -1600 -124440 0 -124430
rect -1600 -124510 -1580 -124440
rect -1180 -124510 -540 -124440
rect -260 -124510 0 -124440
rect -1600 -124520 0 -124510
rect 150400 -125820 150600 -122970
rect 150000 -125970 150600 -125820
rect -2000 -126180 0 -126030
rect -2000 -129030 -1800 -126180
rect -1600 -127440 0 -127430
rect -1600 -127510 -1580 -127440
rect -1180 -127510 -540 -127440
rect -260 -127510 0 -127440
rect -1600 -127520 0 -127510
rect 150400 -128820 150600 -125970
rect 150000 -128970 150600 -128820
rect -2000 -129180 0 -129030
rect -2000 -132030 -1800 -129180
rect -1600 -130440 0 -130430
rect -1600 -130510 -1580 -130440
rect -1180 -130510 -540 -130440
rect -260 -130510 0 -130440
rect -1600 -130520 0 -130510
rect 150400 -131820 150600 -128970
rect 150000 -131970 150600 -131820
rect -2000 -132180 0 -132030
rect -2000 -135030 -1800 -132180
rect -1600 -133440 0 -133430
rect -1600 -133510 -1580 -133440
rect -1180 -133510 -540 -133440
rect -260 -133510 0 -133440
rect -1600 -133520 0 -133510
rect 150400 -134820 150600 -131970
rect 150000 -134970 150600 -134820
rect -2000 -135180 0 -135030
rect -2000 -138030 -1800 -135180
rect -1600 -136440 0 -136430
rect -1600 -136510 -1580 -136440
rect -1180 -136510 -540 -136440
rect -260 -136510 0 -136440
rect -1600 -136520 0 -136510
rect 150400 -137820 150600 -134970
rect 150000 -137970 150600 -137820
rect -2000 -138180 0 -138030
rect -2000 -141030 -1800 -138180
rect -1600 -139440 0 -139430
rect -1600 -139510 -1580 -139440
rect -1180 -139510 -540 -139440
rect -260 -139510 0 -139440
rect -1600 -139520 0 -139510
rect 150400 -140820 150600 -137970
rect 150000 -140970 150600 -140820
rect -2000 -141180 0 -141030
rect -2000 -144030 -1800 -141180
rect -1600 -142440 0 -142430
rect -1600 -142510 -1580 -142440
rect -1180 -142510 -540 -142440
rect -260 -142510 0 -142440
rect -1600 -142520 0 -142510
rect 150400 -143820 150600 -140970
rect 150000 -143970 150600 -143820
rect -2000 -144180 0 -144030
rect -2000 -147000 -1800 -144180
rect -1600 -145440 0 -145430
rect -1600 -145510 -1580 -145440
rect -1180 -145510 -540 -145440
rect -260 -145510 0 -145440
rect -1600 -145520 0 -145510
rect 150400 -146820 150600 -143970
rect 150000 -146970 150600 -146820
rect 540 -147200 560 -147130
rect 2120 -147200 2140 -147130
rect 540 -147230 2140 -147200
rect 540 -147290 560 -147230
rect 2120 -147290 2140 -147230
rect 540 -147300 2140 -147290
rect 3540 -147200 3560 -147130
rect 5120 -147200 5140 -147130
rect 3540 -147230 5140 -147200
rect 3540 -147290 3560 -147230
rect 5120 -147290 5140 -147230
rect 3540 -147300 5140 -147290
rect 6540 -147200 6560 -147130
rect 8120 -147200 8140 -147130
rect 6540 -147230 8140 -147200
rect 6540 -147290 6560 -147230
rect 8120 -147290 8140 -147230
rect 6540 -147300 8140 -147290
rect 9540 -147200 9560 -147130
rect 11120 -147200 11140 -147130
rect 9540 -147230 11140 -147200
rect 9540 -147290 9560 -147230
rect 11120 -147290 11140 -147230
rect 9540 -147300 11140 -147290
rect 12540 -147200 12560 -147130
rect 14120 -147200 14140 -147130
rect 12540 -147230 14140 -147200
rect 12540 -147290 12560 -147230
rect 14120 -147290 14140 -147230
rect 12540 -147300 14140 -147290
rect 15540 -147200 15560 -147130
rect 17120 -147200 17140 -147130
rect 15540 -147230 17140 -147200
rect 15540 -147290 15560 -147230
rect 17120 -147290 17140 -147230
rect 15540 -147300 17140 -147290
rect 18540 -147200 18560 -147130
rect 20120 -147200 20140 -147130
rect 18540 -147230 20140 -147200
rect 18540 -147290 18560 -147230
rect 20120 -147290 20140 -147230
rect 18540 -147300 20140 -147290
rect 21540 -147200 21560 -147130
rect 23120 -147200 23140 -147130
rect 21540 -147230 23140 -147200
rect 21540 -147290 21560 -147230
rect 23120 -147290 23140 -147230
rect 21540 -147300 23140 -147290
rect 24540 -147200 24560 -147130
rect 26120 -147200 26140 -147130
rect 24540 -147230 26140 -147200
rect 24540 -147290 24560 -147230
rect 26120 -147290 26140 -147230
rect 24540 -147300 26140 -147290
rect 27540 -147200 27560 -147130
rect 29120 -147200 29140 -147130
rect 27540 -147230 29140 -147200
rect 27540 -147290 27560 -147230
rect 29120 -147290 29140 -147230
rect 27540 -147300 29140 -147290
rect 30540 -147200 30560 -147130
rect 32120 -147200 32140 -147130
rect 30540 -147230 32140 -147200
rect 30540 -147290 30560 -147230
rect 32120 -147290 32140 -147230
rect 30540 -147300 32140 -147290
rect 33540 -147200 33560 -147130
rect 35120 -147200 35140 -147130
rect 33540 -147230 35140 -147200
rect 33540 -147290 33560 -147230
rect 35120 -147290 35140 -147230
rect 33540 -147300 35140 -147290
rect 36540 -147200 36560 -147130
rect 38120 -147200 38140 -147130
rect 36540 -147230 38140 -147200
rect 36540 -147290 36560 -147230
rect 38120 -147290 38140 -147230
rect 36540 -147300 38140 -147290
rect 39540 -147200 39560 -147130
rect 41120 -147200 41140 -147130
rect 39540 -147230 41140 -147200
rect 39540 -147290 39560 -147230
rect 41120 -147290 41140 -147230
rect 39540 -147300 41140 -147290
rect 42540 -147200 42560 -147130
rect 44120 -147200 44140 -147130
rect 42540 -147230 44140 -147200
rect 42540 -147290 42560 -147230
rect 44120 -147290 44140 -147230
rect 42540 -147300 44140 -147290
rect 45540 -147200 45560 -147130
rect 47120 -147200 47140 -147130
rect 45540 -147230 47140 -147200
rect 45540 -147290 45560 -147230
rect 47120 -147290 47140 -147230
rect 45540 -147300 47140 -147290
rect 48540 -147200 48560 -147130
rect 50120 -147200 50140 -147130
rect 48540 -147230 50140 -147200
rect 48540 -147290 48560 -147230
rect 50120 -147290 50140 -147230
rect 48540 -147300 50140 -147290
rect 51540 -147200 51560 -147130
rect 53120 -147200 53140 -147130
rect 51540 -147230 53140 -147200
rect 51540 -147290 51560 -147230
rect 53120 -147290 53140 -147230
rect 51540 -147300 53140 -147290
rect 54540 -147200 54560 -147130
rect 56120 -147200 56140 -147130
rect 54540 -147230 56140 -147200
rect 54540 -147290 54560 -147230
rect 56120 -147290 56140 -147230
rect 54540 -147300 56140 -147290
rect 57540 -147200 57560 -147130
rect 59120 -147200 59140 -147130
rect 57540 -147230 59140 -147200
rect 57540 -147290 57560 -147230
rect 59120 -147290 59140 -147230
rect 57540 -147300 59140 -147290
rect 60540 -147200 60560 -147130
rect 62120 -147200 62140 -147130
rect 60540 -147230 62140 -147200
rect 60540 -147290 60560 -147230
rect 62120 -147290 62140 -147230
rect 60540 -147300 62140 -147290
rect 63540 -147200 63560 -147130
rect 65120 -147200 65140 -147130
rect 63540 -147230 65140 -147200
rect 63540 -147290 63560 -147230
rect 65120 -147290 65140 -147230
rect 63540 -147300 65140 -147290
rect 66540 -147200 66560 -147130
rect 68120 -147200 68140 -147130
rect 66540 -147230 68140 -147200
rect 66540 -147290 66560 -147230
rect 68120 -147290 68140 -147230
rect 66540 -147300 68140 -147290
rect 69540 -147200 69560 -147130
rect 71120 -147200 71140 -147130
rect 69540 -147230 71140 -147200
rect 69540 -147290 69560 -147230
rect 71120 -147290 71140 -147230
rect 69540 -147300 71140 -147290
rect 72540 -147200 72560 -147130
rect 74120 -147200 74140 -147130
rect 72540 -147230 74140 -147200
rect 72540 -147290 72560 -147230
rect 74120 -147290 74140 -147230
rect 72540 -147300 74140 -147290
rect 75540 -147200 75560 -147130
rect 77120 -147200 77140 -147130
rect 75540 -147230 77140 -147200
rect 75540 -147290 75560 -147230
rect 77120 -147290 77140 -147230
rect 75540 -147300 77140 -147290
rect 78540 -147200 78560 -147130
rect 80120 -147200 80140 -147130
rect 78540 -147230 80140 -147200
rect 78540 -147290 78560 -147230
rect 80120 -147290 80140 -147230
rect 78540 -147300 80140 -147290
rect 81540 -147200 81560 -147130
rect 83120 -147200 83140 -147130
rect 81540 -147230 83140 -147200
rect 81540 -147290 81560 -147230
rect 83120 -147290 83140 -147230
rect 81540 -147300 83140 -147290
rect 84540 -147200 84560 -147130
rect 86120 -147200 86140 -147130
rect 84540 -147230 86140 -147200
rect 84540 -147290 84560 -147230
rect 86120 -147290 86140 -147230
rect 84540 -147300 86140 -147290
rect 87540 -147200 87560 -147130
rect 89120 -147200 89140 -147130
rect 87540 -147230 89140 -147200
rect 87540 -147290 87560 -147230
rect 89120 -147290 89140 -147230
rect 87540 -147300 89140 -147290
rect 90540 -147200 90560 -147130
rect 92120 -147200 92140 -147130
rect 90540 -147230 92140 -147200
rect 90540 -147290 90560 -147230
rect 92120 -147290 92140 -147230
rect 90540 -147300 92140 -147290
rect 93540 -147200 93560 -147130
rect 95120 -147200 95140 -147130
rect 93540 -147230 95140 -147200
rect 93540 -147290 93560 -147230
rect 95120 -147290 95140 -147230
rect 93540 -147300 95140 -147290
rect 96540 -147200 96560 -147130
rect 98120 -147200 98140 -147130
rect 96540 -147230 98140 -147200
rect 96540 -147290 96560 -147230
rect 98120 -147290 98140 -147230
rect 96540 -147300 98140 -147290
rect 99540 -147200 99560 -147130
rect 101120 -147200 101140 -147130
rect 99540 -147230 101140 -147200
rect 99540 -147290 99560 -147230
rect 101120 -147290 101140 -147230
rect 99540 -147300 101140 -147290
rect 102540 -147200 102560 -147130
rect 104120 -147200 104140 -147130
rect 102540 -147230 104140 -147200
rect 102540 -147290 102560 -147230
rect 104120 -147290 104140 -147230
rect 102540 -147300 104140 -147290
rect 105540 -147200 105560 -147130
rect 107120 -147200 107140 -147130
rect 105540 -147230 107140 -147200
rect 105540 -147290 105560 -147230
rect 107120 -147290 107140 -147230
rect 105540 -147300 107140 -147290
rect 108540 -147200 108560 -147130
rect 110120 -147200 110140 -147130
rect 108540 -147230 110140 -147200
rect 108540 -147290 108560 -147230
rect 110120 -147290 110140 -147230
rect 108540 -147300 110140 -147290
rect 111540 -147200 111560 -147130
rect 113120 -147200 113140 -147130
rect 111540 -147230 113140 -147200
rect 111540 -147290 111560 -147230
rect 113120 -147290 113140 -147230
rect 111540 -147300 113140 -147290
rect 114540 -147200 114560 -147130
rect 116120 -147200 116140 -147130
rect 114540 -147230 116140 -147200
rect 114540 -147290 114560 -147230
rect 116120 -147290 116140 -147230
rect 114540 -147300 116140 -147290
rect 117540 -147200 117560 -147130
rect 119120 -147200 119140 -147130
rect 117540 -147230 119140 -147200
rect 117540 -147290 117560 -147230
rect 119120 -147290 119140 -147230
rect 117540 -147300 119140 -147290
rect 120540 -147200 120560 -147130
rect 122120 -147200 122140 -147130
rect 120540 -147230 122140 -147200
rect 120540 -147290 120560 -147230
rect 122120 -147290 122140 -147230
rect 120540 -147300 122140 -147290
rect 123540 -147200 123560 -147130
rect 125120 -147200 125140 -147130
rect 123540 -147230 125140 -147200
rect 123540 -147290 123560 -147230
rect 125120 -147290 125140 -147230
rect 123540 -147300 125140 -147290
rect 126540 -147200 126560 -147130
rect 128120 -147200 128140 -147130
rect 126540 -147230 128140 -147200
rect 126540 -147290 126560 -147230
rect 128120 -147290 128140 -147230
rect 126540 -147300 128140 -147290
rect 129540 -147200 129560 -147130
rect 131120 -147200 131140 -147130
rect 129540 -147230 131140 -147200
rect 129540 -147290 129560 -147230
rect 131120 -147290 131140 -147230
rect 129540 -147300 131140 -147290
rect 132540 -147200 132560 -147130
rect 134120 -147200 134140 -147130
rect 132540 -147230 134140 -147200
rect 132540 -147290 132560 -147230
rect 134120 -147290 134140 -147230
rect 132540 -147300 134140 -147290
rect 135540 -147200 135560 -147130
rect 137120 -147200 137140 -147130
rect 135540 -147230 137140 -147200
rect 135540 -147290 135560 -147230
rect 137120 -147290 137140 -147230
rect 135540 -147300 137140 -147290
rect 138540 -147200 138560 -147130
rect 140120 -147200 140140 -147130
rect 138540 -147230 140140 -147200
rect 138540 -147290 138560 -147230
rect 140120 -147290 140140 -147230
rect 138540 -147300 140140 -147290
rect 141540 -147200 141560 -147130
rect 143120 -147200 143140 -147130
rect 141540 -147230 143140 -147200
rect 141540 -147290 141560 -147230
rect 143120 -147290 143140 -147230
rect 141540 -147300 143140 -147290
rect 144540 -147200 144560 -147130
rect 146120 -147200 146140 -147130
rect 144540 -147230 146140 -147200
rect 144540 -147290 144560 -147230
rect 146120 -147290 146140 -147230
rect 144540 -147300 146140 -147290
rect 147540 -147200 147560 -147130
rect 149120 -147200 149140 -147130
rect 147540 -147230 149140 -147200
rect 147540 -147290 147560 -147230
rect 149120 -147290 149140 -147230
rect 147540 -147300 149140 -147290
rect 220 -147500 440 -147490
rect 220 -147700 240 -147500
rect 420 -147700 440 -147500
rect 220 -147710 440 -147700
rect 3220 -147500 3440 -147490
rect 3220 -147700 3240 -147500
rect 3420 -147700 3440 -147500
rect 3220 -147710 3440 -147700
rect 6220 -147500 6440 -147490
rect 6220 -147700 6240 -147500
rect 6420 -147700 6440 -147500
rect 6220 -147710 6440 -147700
rect 9220 -147500 9440 -147490
rect 9220 -147700 9240 -147500
rect 9420 -147700 9440 -147500
rect 9220 -147710 9440 -147700
rect 12220 -147500 12440 -147490
rect 12220 -147700 12240 -147500
rect 12420 -147700 12440 -147500
rect 12220 -147710 12440 -147700
rect 15220 -147500 15440 -147490
rect 15220 -147700 15240 -147500
rect 15420 -147700 15440 -147500
rect 15220 -147710 15440 -147700
rect 18220 -147500 18440 -147490
rect 18220 -147700 18240 -147500
rect 18420 -147700 18440 -147500
rect 18220 -147710 18440 -147700
rect 21220 -147500 21440 -147490
rect 21220 -147700 21240 -147500
rect 21420 -147700 21440 -147500
rect 21220 -147710 21440 -147700
rect 24220 -147500 24440 -147490
rect 24220 -147700 24240 -147500
rect 24420 -147700 24440 -147500
rect 24220 -147710 24440 -147700
rect 27220 -147500 27440 -147490
rect 27220 -147700 27240 -147500
rect 27420 -147700 27440 -147500
rect 27220 -147710 27440 -147700
rect 30220 -147500 30440 -147490
rect 30220 -147700 30240 -147500
rect 30420 -147700 30440 -147500
rect 30220 -147710 30440 -147700
rect 33220 -147500 33440 -147490
rect 33220 -147700 33240 -147500
rect 33420 -147700 33440 -147500
rect 33220 -147710 33440 -147700
rect 36220 -147500 36440 -147490
rect 36220 -147700 36240 -147500
rect 36420 -147700 36440 -147500
rect 36220 -147710 36440 -147700
rect 39220 -147500 39440 -147490
rect 39220 -147700 39240 -147500
rect 39420 -147700 39440 -147500
rect 39220 -147710 39440 -147700
rect 42220 -147500 42440 -147490
rect 42220 -147700 42240 -147500
rect 42420 -147700 42440 -147500
rect 42220 -147710 42440 -147700
rect 45220 -147500 45440 -147490
rect 45220 -147700 45240 -147500
rect 45420 -147700 45440 -147500
rect 45220 -147710 45440 -147700
rect 48220 -147500 48440 -147490
rect 48220 -147700 48240 -147500
rect 48420 -147700 48440 -147500
rect 48220 -147710 48440 -147700
rect 51220 -147500 51440 -147490
rect 51220 -147700 51240 -147500
rect 51420 -147700 51440 -147500
rect 51220 -147710 51440 -147700
rect 54220 -147500 54440 -147490
rect 54220 -147700 54240 -147500
rect 54420 -147700 54440 -147500
rect 54220 -147710 54440 -147700
rect 57220 -147500 57440 -147490
rect 57220 -147700 57240 -147500
rect 57420 -147700 57440 -147500
rect 57220 -147710 57440 -147700
rect 60220 -147500 60440 -147490
rect 60220 -147700 60240 -147500
rect 60420 -147700 60440 -147500
rect 60220 -147710 60440 -147700
rect 63220 -147500 63440 -147490
rect 63220 -147700 63240 -147500
rect 63420 -147700 63440 -147500
rect 63220 -147710 63440 -147700
rect 66220 -147500 66440 -147490
rect 66220 -147700 66240 -147500
rect 66420 -147700 66440 -147500
rect 66220 -147710 66440 -147700
rect 69220 -147500 69440 -147490
rect 69220 -147700 69240 -147500
rect 69420 -147700 69440 -147500
rect 69220 -147710 69440 -147700
rect 72220 -147500 72440 -147490
rect 72220 -147700 72240 -147500
rect 72420 -147700 72440 -147500
rect 72220 -147710 72440 -147700
rect 75220 -147500 75440 -147490
rect 75220 -147700 75240 -147500
rect 75420 -147700 75440 -147500
rect 75220 -147710 75440 -147700
rect 78220 -147500 78440 -147490
rect 78220 -147700 78240 -147500
rect 78420 -147700 78440 -147500
rect 78220 -147710 78440 -147700
rect 81220 -147500 81440 -147490
rect 81220 -147700 81240 -147500
rect 81420 -147700 81440 -147500
rect 81220 -147710 81440 -147700
rect 84220 -147500 84440 -147490
rect 84220 -147700 84240 -147500
rect 84420 -147700 84440 -147500
rect 84220 -147710 84440 -147700
rect 87220 -147500 87440 -147490
rect 87220 -147700 87240 -147500
rect 87420 -147700 87440 -147500
rect 87220 -147710 87440 -147700
rect 90220 -147500 90440 -147490
rect 90220 -147700 90240 -147500
rect 90420 -147700 90440 -147500
rect 90220 -147710 90440 -147700
rect 93220 -147500 93440 -147490
rect 93220 -147700 93240 -147500
rect 93420 -147700 93440 -147500
rect 93220 -147710 93440 -147700
rect 96220 -147500 96440 -147490
rect 96220 -147700 96240 -147500
rect 96420 -147700 96440 -147500
rect 96220 -147710 96440 -147700
rect 99220 -147500 99440 -147490
rect 99220 -147700 99240 -147500
rect 99420 -147700 99440 -147500
rect 99220 -147710 99440 -147700
rect 102220 -147500 102440 -147490
rect 102220 -147700 102240 -147500
rect 102420 -147700 102440 -147500
rect 102220 -147710 102440 -147700
rect 105220 -147500 105440 -147490
rect 105220 -147700 105240 -147500
rect 105420 -147700 105440 -147500
rect 105220 -147710 105440 -147700
rect 108220 -147500 108440 -147490
rect 108220 -147700 108240 -147500
rect 108420 -147700 108440 -147500
rect 108220 -147710 108440 -147700
rect 111220 -147500 111440 -147490
rect 111220 -147700 111240 -147500
rect 111420 -147700 111440 -147500
rect 111220 -147710 111440 -147700
rect 114220 -147500 114440 -147490
rect 114220 -147700 114240 -147500
rect 114420 -147700 114440 -147500
rect 114220 -147710 114440 -147700
rect 117220 -147500 117440 -147490
rect 117220 -147700 117240 -147500
rect 117420 -147700 117440 -147500
rect 117220 -147710 117440 -147700
rect 120220 -147500 120440 -147490
rect 120220 -147700 120240 -147500
rect 120420 -147700 120440 -147500
rect 120220 -147710 120440 -147700
rect 123220 -147500 123440 -147490
rect 123220 -147700 123240 -147500
rect 123420 -147700 123440 -147500
rect 123220 -147710 123440 -147700
rect 126220 -147500 126440 -147490
rect 126220 -147700 126240 -147500
rect 126420 -147700 126440 -147500
rect 126220 -147710 126440 -147700
rect 129220 -147500 129440 -147490
rect 129220 -147700 129240 -147500
rect 129420 -147700 129440 -147500
rect 129220 -147710 129440 -147700
rect 132220 -147500 132440 -147490
rect 132220 -147700 132240 -147500
rect 132420 -147700 132440 -147500
rect 132220 -147710 132440 -147700
rect 135220 -147500 135440 -147490
rect 135220 -147700 135240 -147500
rect 135420 -147700 135440 -147500
rect 135220 -147710 135440 -147700
rect 138220 -147500 138440 -147490
rect 138220 -147700 138240 -147500
rect 138420 -147700 138440 -147500
rect 138220 -147710 138440 -147700
rect 141220 -147500 141440 -147490
rect 141220 -147700 141240 -147500
rect 141420 -147700 141440 -147500
rect 141220 -147710 141440 -147700
rect 144220 -147500 144440 -147490
rect 144220 -147700 144240 -147500
rect 144420 -147700 144440 -147500
rect 144220 -147710 144440 -147700
rect 147220 -147500 147440 -147490
rect 147220 -147700 147240 -147500
rect 147420 -147700 147440 -147500
rect 147220 -147710 147440 -147700
rect 540 -147920 150740 -147900
rect 540 -148080 560 -147920
rect 540 -148100 150740 -148080
<< via1 >>
rect -1920 3360 -900 3450
rect 50 3360 140 3450
rect 3050 3360 3140 3450
rect 6050 3360 6140 3450
rect 9050 3360 9140 3450
rect 12050 3360 12140 3450
rect 15050 3360 15140 3450
rect 18050 3360 18140 3450
rect 21050 3360 21140 3450
rect 24050 3360 24140 3450
rect 27050 3360 27140 3450
rect 30050 3360 30140 3450
rect 33050 3360 33140 3450
rect 36050 3360 36140 3450
rect 39050 3360 39140 3450
rect 42050 3360 42140 3450
rect 45050 3360 45140 3450
rect 48050 3360 48140 3450
rect 51050 3360 51140 3450
rect 54050 3360 54140 3450
rect 57050 3360 57140 3450
rect 60050 3360 60140 3450
rect 63050 3360 63140 3450
rect 66050 3360 66140 3450
rect 69050 3360 69140 3450
rect 72050 3360 72140 3450
rect 75050 3360 75140 3450
rect 78050 3360 78140 3450
rect 81050 3360 81140 3450
rect 84050 3360 84140 3450
rect 87050 3360 87140 3450
rect 90050 3360 90140 3450
rect 93050 3360 93140 3450
rect 96050 3360 96140 3450
rect 99050 3360 99140 3450
rect 102050 3360 102140 3450
rect 105050 3360 105140 3450
rect 108050 3360 108140 3450
rect 111050 3360 111140 3450
rect 114050 3360 114140 3450
rect 117050 3360 117140 3450
rect 120050 3360 120140 3450
rect 123050 3360 123140 3450
rect 126050 3360 126140 3450
rect 129050 3360 129140 3450
rect 132050 3360 132140 3450
rect 135050 3360 135140 3450
rect 138050 3360 138140 3450
rect 141050 3360 141140 3450
rect 144050 3360 144140 3450
rect 147050 3360 147140 3450
rect -1580 1490 -1180 1560
rect -540 1490 -260 1560
rect -1580 -1510 -1180 -1440
rect -540 -1510 -260 -1440
rect -1580 -4510 -1180 -4440
rect -540 -4510 -260 -4440
rect -1580 -7510 -1180 -7440
rect -540 -7510 -260 -7440
rect -1580 -10510 -1180 -10440
rect -540 -10510 -260 -10440
rect -1580 -13510 -1180 -13440
rect -540 -13510 -260 -13440
rect -1580 -16510 -1180 -16440
rect -540 -16510 -260 -16440
rect -1580 -19510 -1180 -19440
rect -540 -19510 -260 -19440
rect -1580 -22510 -1180 -22440
rect -540 -22510 -260 -22440
rect -1580 -25510 -1180 -25440
rect -540 -25510 -260 -25440
rect -1580 -28510 -1180 -28440
rect -540 -28510 -260 -28440
rect -1580 -31510 -1180 -31440
rect -540 -31510 -260 -31440
rect -1580 -34510 -1180 -34440
rect -540 -34510 -260 -34440
rect -1580 -37510 -1180 -37440
rect -540 -37510 -260 -37440
rect -1580 -40510 -1180 -40440
rect -540 -40510 -260 -40440
rect -1580 -43510 -1180 -43440
rect -540 -43510 -260 -43440
rect -1580 -46510 -1180 -46440
rect -540 -46510 -260 -46440
rect -1580 -49510 -1180 -49440
rect -540 -49510 -260 -49440
rect -1580 -52510 -1180 -52440
rect -540 -52510 -260 -52440
rect -1580 -55510 -1180 -55440
rect -540 -55510 -260 -55440
rect -1580 -58510 -1180 -58440
rect -540 -58510 -260 -58440
rect -1580 -61510 -1180 -61440
rect -540 -61510 -260 -61440
rect -1580 -64510 -1180 -64440
rect -540 -64510 -260 -64440
rect -1580 -67510 -1180 -67440
rect -540 -67510 -260 -67440
rect -1580 -70510 -1180 -70440
rect -540 -70510 -260 -70440
rect -1580 -73510 -1180 -73440
rect -540 -73510 -260 -73440
rect -1580 -76510 -1180 -76440
rect -540 -76510 -260 -76440
rect -1580 -79510 -1180 -79440
rect -540 -79510 -260 -79440
rect -1580 -82510 -1180 -82440
rect -540 -82510 -260 -82440
rect -1580 -85510 -1180 -85440
rect -540 -85510 -260 -85440
rect -1580 -88510 -1180 -88440
rect -540 -88510 -260 -88440
rect -1580 -91510 -1180 -91440
rect -540 -91510 -260 -91440
rect -1580 -94510 -1180 -94440
rect -540 -94510 -260 -94440
rect -1580 -97510 -1180 -97440
rect -540 -97510 -260 -97440
rect -1580 -100510 -1180 -100440
rect -540 -100510 -260 -100440
rect -1580 -103510 -1180 -103440
rect -540 -103510 -260 -103440
rect -1580 -106510 -1180 -106440
rect -540 -106510 -260 -106440
rect -1580 -109510 -1180 -109440
rect -540 -109510 -260 -109440
rect -1580 -112510 -1180 -112440
rect -540 -112510 -260 -112440
rect -1580 -115510 -1180 -115440
rect -540 -115510 -260 -115440
rect -1580 -118510 -1180 -118440
rect -540 -118510 -260 -118440
rect -1580 -121510 -1180 -121440
rect -540 -121510 -260 -121440
rect -1580 -124510 -1180 -124440
rect -540 -124510 -260 -124440
rect -1580 -127510 -1180 -127440
rect -540 -127510 -260 -127440
rect -1580 -130510 -1180 -130440
rect -540 -130510 -260 -130440
rect -1580 -133510 -1180 -133440
rect -540 -133510 -260 -133440
rect -1580 -136510 -1180 -136440
rect -540 -136510 -260 -136440
rect -1580 -139510 -1180 -139440
rect -540 -139510 -260 -139440
rect -1580 -142510 -1180 -142440
rect -540 -142510 -260 -142440
rect -1580 -145510 -1180 -145440
rect -540 -145510 -260 -145440
rect 560 -147200 2120 -147130
rect 3560 -147200 5120 -147130
rect 6560 -147200 8120 -147130
rect 9560 -147200 11120 -147130
rect 12560 -147200 14120 -147130
rect 15560 -147200 17120 -147130
rect 18560 -147200 20120 -147130
rect 21560 -147200 23120 -147130
rect 24560 -147200 26120 -147130
rect 27560 -147200 29120 -147130
rect 30560 -147200 32120 -147130
rect 33560 -147200 35120 -147130
rect 36560 -147200 38120 -147130
rect 39560 -147200 41120 -147130
rect 42560 -147200 44120 -147130
rect 45560 -147200 47120 -147130
rect 48560 -147200 50120 -147130
rect 51560 -147200 53120 -147130
rect 54560 -147200 56120 -147130
rect 57560 -147200 59120 -147130
rect 60560 -147200 62120 -147130
rect 63560 -147200 65120 -147130
rect 66560 -147200 68120 -147130
rect 69560 -147200 71120 -147130
rect 72560 -147200 74120 -147130
rect 75560 -147200 77120 -147130
rect 78560 -147200 80120 -147130
rect 81560 -147200 83120 -147130
rect 84560 -147200 86120 -147130
rect 87560 -147200 89120 -147130
rect 90560 -147200 92120 -147130
rect 93560 -147200 95120 -147130
rect 96560 -147200 98120 -147130
rect 99560 -147200 101120 -147130
rect 102560 -147200 104120 -147130
rect 105560 -147200 107120 -147130
rect 108560 -147200 110120 -147130
rect 111560 -147200 113120 -147130
rect 114560 -147200 116120 -147130
rect 117560 -147200 119120 -147130
rect 120560 -147200 122120 -147130
rect 123560 -147200 125120 -147130
rect 126560 -147200 128120 -147130
rect 129560 -147200 131120 -147130
rect 132560 -147200 134120 -147130
rect 135560 -147200 137120 -147130
rect 138560 -147200 140120 -147130
rect 141560 -147200 143120 -147130
rect 144560 -147200 146120 -147130
rect 147560 -147200 149120 -147130
rect 240 -147700 420 -147500
rect 3240 -147700 3420 -147500
rect 6240 -147700 6420 -147500
rect 9240 -147700 9420 -147500
rect 12240 -147700 12420 -147500
rect 15240 -147700 15420 -147500
rect 18240 -147700 18420 -147500
rect 21240 -147700 21420 -147500
rect 24240 -147700 24420 -147500
rect 27240 -147700 27420 -147500
rect 30240 -147700 30420 -147500
rect 33240 -147700 33420 -147500
rect 36240 -147700 36420 -147500
rect 39240 -147700 39420 -147500
rect 42240 -147700 42420 -147500
rect 45240 -147700 45420 -147500
rect 48240 -147700 48420 -147500
rect 51240 -147700 51420 -147500
rect 54240 -147700 54420 -147500
rect 57240 -147700 57420 -147500
rect 60240 -147700 60420 -147500
rect 63240 -147700 63420 -147500
rect 66240 -147700 66420 -147500
rect 69240 -147700 69420 -147500
rect 72240 -147700 72420 -147500
rect 75240 -147700 75420 -147500
rect 78240 -147700 78420 -147500
rect 81240 -147700 81420 -147500
rect 84240 -147700 84420 -147500
rect 87240 -147700 87420 -147500
rect 90240 -147700 90420 -147500
rect 93240 -147700 93420 -147500
rect 96240 -147700 96420 -147500
rect 99240 -147700 99420 -147500
rect 102240 -147700 102420 -147500
rect 105240 -147700 105420 -147500
rect 108240 -147700 108420 -147500
rect 111240 -147700 111420 -147500
rect 114240 -147700 114420 -147500
rect 117240 -147700 117420 -147500
rect 120240 -147700 120420 -147500
rect 123240 -147700 123420 -147500
rect 126240 -147700 126420 -147500
rect 129240 -147700 129420 -147500
rect 132240 -147700 132420 -147500
rect 135240 -147700 135420 -147500
rect 138240 -147700 138420 -147500
rect 141240 -147700 141420 -147500
rect 144240 -147700 144420 -147500
rect 147240 -147700 147420 -147500
rect 560 -147980 2120 -147920
rect 2120 -147980 3560 -147920
rect 3560 -147980 5120 -147920
rect 5120 -147980 6560 -147920
rect 6560 -147980 8120 -147920
rect 8120 -147980 9560 -147920
rect 9560 -147980 11120 -147920
rect 11120 -147980 12560 -147920
rect 12560 -147980 14120 -147920
rect 14120 -147980 15560 -147920
rect 15560 -147980 17120 -147920
rect 17120 -147980 18560 -147920
rect 18560 -147980 20120 -147920
rect 20120 -147980 21560 -147920
rect 21560 -147980 23120 -147920
rect 23120 -147980 24560 -147920
rect 24560 -147980 26120 -147920
rect 26120 -147980 27560 -147920
rect 27560 -147980 29120 -147920
rect 29120 -147980 30560 -147920
rect 30560 -147980 32120 -147920
rect 32120 -147980 33560 -147920
rect 33560 -147980 35120 -147920
rect 35120 -147980 36560 -147920
rect 36560 -147980 38120 -147920
rect 38120 -147980 39560 -147920
rect 39560 -147980 41120 -147920
rect 41120 -147980 42560 -147920
rect 42560 -147980 44120 -147920
rect 44120 -147980 45560 -147920
rect 45560 -147980 47120 -147920
rect 47120 -147980 48560 -147920
rect 48560 -147980 50120 -147920
rect 50120 -147980 51560 -147920
rect 51560 -147980 53120 -147920
rect 53120 -147980 54560 -147920
rect 54560 -147980 56120 -147920
rect 56120 -147980 57560 -147920
rect 57560 -147980 59120 -147920
rect 59120 -147980 60560 -147920
rect 60560 -147980 62120 -147920
rect 62120 -147980 63560 -147920
rect 63560 -147980 65120 -147920
rect 65120 -147980 66560 -147920
rect 66560 -147980 68120 -147920
rect 68120 -147980 69560 -147920
rect 69560 -147980 71120 -147920
rect 71120 -147980 72560 -147920
rect 72560 -147980 74120 -147920
rect 74120 -147980 75560 -147920
rect 75560 -147980 77120 -147920
rect 77120 -147980 78560 -147920
rect 78560 -147980 80120 -147920
rect 80120 -147980 81560 -147920
rect 81560 -147980 83120 -147920
rect 83120 -147980 84560 -147920
rect 84560 -147980 86120 -147920
rect 86120 -147980 87560 -147920
rect 87560 -147980 89120 -147920
rect 89120 -147980 90560 -147920
rect 90560 -147980 92120 -147920
rect 92120 -147980 93560 -147920
rect 93560 -147980 95120 -147920
rect 95120 -147980 96560 -147920
rect 96560 -147980 98120 -147920
rect 98120 -147980 99560 -147920
rect 99560 -147980 101120 -147920
rect 101120 -147980 102560 -147920
rect 102560 -147980 104120 -147920
rect 104120 -147980 105560 -147920
rect 105560 -147980 107120 -147920
rect 107120 -147980 108560 -147920
rect 108560 -147980 110120 -147920
rect 110120 -147980 111560 -147920
rect 111560 -147980 113120 -147920
rect 113120 -147980 114560 -147920
rect 114560 -147980 116120 -147920
rect 116120 -147980 117560 -147920
rect 117560 -147980 119120 -147920
rect 119120 -147980 120560 -147920
rect 120560 -147980 122120 -147920
rect 122120 -147980 123560 -147920
rect 123560 -147980 125120 -147920
rect 125120 -147980 126560 -147920
rect 126560 -147980 128120 -147920
rect 128120 -147980 129560 -147920
rect 129560 -147980 131120 -147920
rect 131120 -147980 132560 -147920
rect 132560 -147980 134120 -147920
rect 134120 -147980 135560 -147920
rect 135560 -147980 137120 -147920
rect 137120 -147980 138560 -147920
rect 138560 -147980 140120 -147920
rect 140120 -147980 141560 -147920
rect 141560 -147980 143120 -147920
rect 143120 -147980 144560 -147920
rect 144560 -147980 146120 -147920
rect 146120 -147980 147560 -147920
rect 147560 -147980 149120 -147920
rect 149120 -147980 150740 -147920
rect 560 -148080 150740 -147980
<< metal2 >>
rect 0 4040 150000 4150
rect -3000 3450 -890 3460
rect -3000 3360 -1920 3450
rect -900 3360 -890 3450
rect -3000 3350 -890 3360
rect -3000 1560 -1000 1570
rect -3000 1490 -1580 1560
rect -1180 1490 -1000 1560
rect -3000 1480 -1000 1490
rect -750 230 -640 4000
rect 480 3650 590 3660
rect 480 3560 490 3650
rect 580 3560 590 3650
rect 480 3550 590 3560
rect 40 3450 150 3460
rect 40 3360 50 3450
rect 140 3360 150 3450
rect 40 3350 150 3360
rect 60 3000 130 3350
rect 500 3000 570 3550
rect 1020 3000 1090 4040
rect 3480 3650 3590 3660
rect 3480 3560 3490 3650
rect 3580 3560 3590 3650
rect 3480 3550 3590 3560
rect 3040 3450 3150 3460
rect 3040 3360 3050 3450
rect 3140 3360 3150 3450
rect 3040 3350 3150 3360
rect 3060 3000 3130 3350
rect 3500 3000 3570 3550
rect 4020 3000 4090 4040
rect 6480 3650 6590 3660
rect 6480 3560 6490 3650
rect 6580 3560 6590 3650
rect 6480 3550 6590 3560
rect 6040 3450 6150 3460
rect 6040 3360 6050 3450
rect 6140 3360 6150 3450
rect 6040 3350 6150 3360
rect 6060 3000 6130 3350
rect 6500 3000 6570 3550
rect 7020 3000 7090 4040
rect 9480 3650 9590 3660
rect 9480 3560 9490 3650
rect 9580 3560 9590 3650
rect 9480 3550 9590 3560
rect 9040 3450 9150 3460
rect 9040 3360 9050 3450
rect 9140 3360 9150 3450
rect 9040 3350 9150 3360
rect 9060 3000 9130 3350
rect 9500 3000 9570 3550
rect 10020 3000 10090 4040
rect 12480 3650 12590 3660
rect 12480 3560 12490 3650
rect 12580 3560 12590 3650
rect 12480 3550 12590 3560
rect 12040 3450 12150 3460
rect 12040 3360 12050 3450
rect 12140 3360 12150 3450
rect 12040 3350 12150 3360
rect 12060 3000 12130 3350
rect 12500 3000 12570 3550
rect 13020 3000 13090 4040
rect 15480 3650 15590 3660
rect 15480 3560 15490 3650
rect 15580 3560 15590 3650
rect 15480 3550 15590 3560
rect 15040 3450 15150 3460
rect 15040 3360 15050 3450
rect 15140 3360 15150 3450
rect 15040 3350 15150 3360
rect 15060 3000 15130 3350
rect 15500 3000 15570 3550
rect 16020 3000 16090 4040
rect 18480 3650 18590 3660
rect 18480 3560 18490 3650
rect 18580 3560 18590 3650
rect 18480 3550 18590 3560
rect 18040 3450 18150 3460
rect 18040 3360 18050 3450
rect 18140 3360 18150 3450
rect 18040 3350 18150 3360
rect 18060 3000 18130 3350
rect 18500 3000 18570 3550
rect 19020 3000 19090 4040
rect 21480 3650 21590 3660
rect 21480 3560 21490 3650
rect 21580 3560 21590 3650
rect 21480 3550 21590 3560
rect 21040 3450 21150 3460
rect 21040 3360 21050 3450
rect 21140 3360 21150 3450
rect 21040 3350 21150 3360
rect 21060 3000 21130 3350
rect 21500 3000 21570 3550
rect 22020 3000 22090 4040
rect 24480 3650 24590 3660
rect 24480 3560 24490 3650
rect 24580 3560 24590 3650
rect 24480 3550 24590 3560
rect 24040 3450 24150 3460
rect 24040 3360 24050 3450
rect 24140 3360 24150 3450
rect 24040 3350 24150 3360
rect 24060 3000 24130 3350
rect 24500 3000 24570 3550
rect 25020 3000 25090 4040
rect 27480 3650 27590 3660
rect 27480 3560 27490 3650
rect 27580 3560 27590 3650
rect 27480 3550 27590 3560
rect 27040 3450 27150 3460
rect 27040 3360 27050 3450
rect 27140 3360 27150 3450
rect 27040 3350 27150 3360
rect 27060 3000 27130 3350
rect 27500 3000 27570 3550
rect 28020 3000 28090 4040
rect 30480 3650 30590 3660
rect 30480 3560 30490 3650
rect 30580 3560 30590 3650
rect 30480 3550 30590 3560
rect 30040 3450 30150 3460
rect 30040 3360 30050 3450
rect 30140 3360 30150 3450
rect 30040 3350 30150 3360
rect 30060 3000 30130 3350
rect 30500 3000 30570 3550
rect 31020 3000 31090 4040
rect 33480 3650 33590 3660
rect 33480 3560 33490 3650
rect 33580 3560 33590 3650
rect 33480 3550 33590 3560
rect 33040 3450 33150 3460
rect 33040 3360 33050 3450
rect 33140 3360 33150 3450
rect 33040 3350 33150 3360
rect 33060 3000 33130 3350
rect 33500 3000 33570 3550
rect 34020 3000 34090 4040
rect 36480 3650 36590 3660
rect 36480 3560 36490 3650
rect 36580 3560 36590 3650
rect 36480 3550 36590 3560
rect 36040 3450 36150 3460
rect 36040 3360 36050 3450
rect 36140 3360 36150 3450
rect 36040 3350 36150 3360
rect 36060 3000 36130 3350
rect 36500 3000 36570 3550
rect 37020 3000 37090 4040
rect 39480 3650 39590 3660
rect 39480 3560 39490 3650
rect 39580 3560 39590 3650
rect 39480 3550 39590 3560
rect 39040 3450 39150 3460
rect 39040 3360 39050 3450
rect 39140 3360 39150 3450
rect 39040 3350 39150 3360
rect 39060 3000 39130 3350
rect 39500 3000 39570 3550
rect 40020 3000 40090 4040
rect 42480 3650 42590 3660
rect 42480 3560 42490 3650
rect 42580 3560 42590 3650
rect 42480 3550 42590 3560
rect 42040 3450 42150 3460
rect 42040 3360 42050 3450
rect 42140 3360 42150 3450
rect 42040 3350 42150 3360
rect 42060 3000 42130 3350
rect 42500 3000 42570 3550
rect 43020 3000 43090 4040
rect 45480 3650 45590 3660
rect 45480 3560 45490 3650
rect 45580 3560 45590 3650
rect 45480 3550 45590 3560
rect 45040 3450 45150 3460
rect 45040 3360 45050 3450
rect 45140 3360 45150 3450
rect 45040 3350 45150 3360
rect 45060 3000 45130 3350
rect 45500 3000 45570 3550
rect 46020 3000 46090 4040
rect 48480 3650 48590 3660
rect 48480 3560 48490 3650
rect 48580 3560 48590 3650
rect 48480 3550 48590 3560
rect 48040 3450 48150 3460
rect 48040 3360 48050 3450
rect 48140 3360 48150 3450
rect 48040 3350 48150 3360
rect 48060 3000 48130 3350
rect 48500 3000 48570 3550
rect 49020 3000 49090 4040
rect 51480 3650 51590 3660
rect 51480 3560 51490 3650
rect 51580 3560 51590 3650
rect 51480 3550 51590 3560
rect 51040 3450 51150 3460
rect 51040 3360 51050 3450
rect 51140 3360 51150 3450
rect 51040 3350 51150 3360
rect 51060 3000 51130 3350
rect 51500 3000 51570 3550
rect 52020 3000 52090 4040
rect 54480 3650 54590 3660
rect 54480 3560 54490 3650
rect 54580 3560 54590 3650
rect 54480 3550 54590 3560
rect 54040 3450 54150 3460
rect 54040 3360 54050 3450
rect 54140 3360 54150 3450
rect 54040 3350 54150 3360
rect 54060 3000 54130 3350
rect 54500 3000 54570 3550
rect 55020 3000 55090 4040
rect 57480 3650 57590 3660
rect 57480 3560 57490 3650
rect 57580 3560 57590 3650
rect 57480 3550 57590 3560
rect 57040 3450 57150 3460
rect 57040 3360 57050 3450
rect 57140 3360 57150 3450
rect 57040 3350 57150 3360
rect 57060 3000 57130 3350
rect 57500 3000 57570 3550
rect 58020 3000 58090 4040
rect 60480 3650 60590 3660
rect 60480 3560 60490 3650
rect 60580 3560 60590 3650
rect 60480 3550 60590 3560
rect 60040 3450 60150 3460
rect 60040 3360 60050 3450
rect 60140 3360 60150 3450
rect 60040 3350 60150 3360
rect 60060 3000 60130 3350
rect 60500 3000 60570 3550
rect 61020 3000 61090 4040
rect 63480 3650 63590 3660
rect 63480 3560 63490 3650
rect 63580 3560 63590 3650
rect 63480 3550 63590 3560
rect 63040 3450 63150 3460
rect 63040 3360 63050 3450
rect 63140 3360 63150 3450
rect 63040 3350 63150 3360
rect 63060 3000 63130 3350
rect 63500 3000 63570 3550
rect 64020 3000 64090 4040
rect 66480 3650 66590 3660
rect 66480 3560 66490 3650
rect 66580 3560 66590 3650
rect 66480 3550 66590 3560
rect 66040 3450 66150 3460
rect 66040 3360 66050 3450
rect 66140 3360 66150 3450
rect 66040 3350 66150 3360
rect 66060 3000 66130 3350
rect 66500 3000 66570 3550
rect 67020 3000 67090 4040
rect 69480 3650 69590 3660
rect 69480 3560 69490 3650
rect 69580 3560 69590 3650
rect 69480 3550 69590 3560
rect 69040 3450 69150 3460
rect 69040 3360 69050 3450
rect 69140 3360 69150 3450
rect 69040 3350 69150 3360
rect 69060 3000 69130 3350
rect 69500 3000 69570 3550
rect 70020 3000 70090 4040
rect 72480 3650 72590 3660
rect 72480 3560 72490 3650
rect 72580 3560 72590 3650
rect 72480 3550 72590 3560
rect 72040 3450 72150 3460
rect 72040 3360 72050 3450
rect 72140 3360 72150 3450
rect 72040 3350 72150 3360
rect 72060 3000 72130 3350
rect 72500 3000 72570 3550
rect 73020 3000 73090 4040
rect 75480 3650 75590 3660
rect 75480 3560 75490 3650
rect 75580 3560 75590 3650
rect 75480 3550 75590 3560
rect 75040 3450 75150 3460
rect 75040 3360 75050 3450
rect 75140 3360 75150 3450
rect 75040 3350 75150 3360
rect 75060 3000 75130 3350
rect 75500 3000 75570 3550
rect 76020 3000 76090 4040
rect 78480 3650 78590 3660
rect 78480 3560 78490 3650
rect 78580 3560 78590 3650
rect 78480 3550 78590 3560
rect 78040 3450 78150 3460
rect 78040 3360 78050 3450
rect 78140 3360 78150 3450
rect 78040 3350 78150 3360
rect 78060 3000 78130 3350
rect 78500 3000 78570 3550
rect 79020 3000 79090 4040
rect 81480 3650 81590 3660
rect 81480 3560 81490 3650
rect 81580 3560 81590 3650
rect 81480 3550 81590 3560
rect 81040 3450 81150 3460
rect 81040 3360 81050 3450
rect 81140 3360 81150 3450
rect 81040 3350 81150 3360
rect 81060 3000 81130 3350
rect 81500 3000 81570 3550
rect 82020 3000 82090 4040
rect 84480 3650 84590 3660
rect 84480 3560 84490 3650
rect 84580 3560 84590 3650
rect 84480 3550 84590 3560
rect 84040 3450 84150 3460
rect 84040 3360 84050 3450
rect 84140 3360 84150 3450
rect 84040 3350 84150 3360
rect 84060 3000 84130 3350
rect 84500 3000 84570 3550
rect 85020 3000 85090 4040
rect 87480 3650 87590 3660
rect 87480 3560 87490 3650
rect 87580 3560 87590 3650
rect 87480 3550 87590 3560
rect 87040 3450 87150 3460
rect 87040 3360 87050 3450
rect 87140 3360 87150 3450
rect 87040 3350 87150 3360
rect 87060 3000 87130 3350
rect 87500 3000 87570 3550
rect 88020 3000 88090 4040
rect 90480 3650 90590 3660
rect 90480 3560 90490 3650
rect 90580 3560 90590 3650
rect 90480 3550 90590 3560
rect 90040 3450 90150 3460
rect 90040 3360 90050 3450
rect 90140 3360 90150 3450
rect 90040 3350 90150 3360
rect 90060 3000 90130 3350
rect 90500 3000 90570 3550
rect 91020 3000 91090 4040
rect 93480 3650 93590 3660
rect 93480 3560 93490 3650
rect 93580 3560 93590 3650
rect 93480 3550 93590 3560
rect 93040 3450 93150 3460
rect 93040 3360 93050 3450
rect 93140 3360 93150 3450
rect 93040 3350 93150 3360
rect 93060 3000 93130 3350
rect 93500 3000 93570 3550
rect 94020 3000 94090 4040
rect 96480 3650 96590 3660
rect 96480 3560 96490 3650
rect 96580 3560 96590 3650
rect 96480 3550 96590 3560
rect 96040 3450 96150 3460
rect 96040 3360 96050 3450
rect 96140 3360 96150 3450
rect 96040 3350 96150 3360
rect 96060 3000 96130 3350
rect 96500 3000 96570 3550
rect 97020 3000 97090 4040
rect 99480 3650 99590 3660
rect 99480 3560 99490 3650
rect 99580 3560 99590 3650
rect 99480 3550 99590 3560
rect 99040 3450 99150 3460
rect 99040 3360 99050 3450
rect 99140 3360 99150 3450
rect 99040 3350 99150 3360
rect 99060 3000 99130 3350
rect 99500 3000 99570 3550
rect 100020 3000 100090 4040
rect 102480 3650 102590 3660
rect 102480 3560 102490 3650
rect 102580 3560 102590 3650
rect 102480 3550 102590 3560
rect 102040 3450 102150 3460
rect 102040 3360 102050 3450
rect 102140 3360 102150 3450
rect 102040 3350 102150 3360
rect 102060 3000 102130 3350
rect 102500 3000 102570 3550
rect 103020 3000 103090 4040
rect 105480 3650 105590 3660
rect 105480 3560 105490 3650
rect 105580 3560 105590 3650
rect 105480 3550 105590 3560
rect 105040 3450 105150 3460
rect 105040 3360 105050 3450
rect 105140 3360 105150 3450
rect 105040 3350 105150 3360
rect 105060 3000 105130 3350
rect 105500 3000 105570 3550
rect 106020 3000 106090 4040
rect 108480 3650 108590 3660
rect 108480 3560 108490 3650
rect 108580 3560 108590 3650
rect 108480 3550 108590 3560
rect 108040 3450 108150 3460
rect 108040 3360 108050 3450
rect 108140 3360 108150 3450
rect 108040 3350 108150 3360
rect 108060 3000 108130 3350
rect 108500 3000 108570 3550
rect 109020 3000 109090 4040
rect 111480 3650 111590 3660
rect 111480 3560 111490 3650
rect 111580 3560 111590 3650
rect 111480 3550 111590 3560
rect 111040 3450 111150 3460
rect 111040 3360 111050 3450
rect 111140 3360 111150 3450
rect 111040 3350 111150 3360
rect 111060 3000 111130 3350
rect 111500 3000 111570 3550
rect 112020 3000 112090 4040
rect 114480 3650 114590 3660
rect 114480 3560 114490 3650
rect 114580 3560 114590 3650
rect 114480 3550 114590 3560
rect 114040 3450 114150 3460
rect 114040 3360 114050 3450
rect 114140 3360 114150 3450
rect 114040 3350 114150 3360
rect 114060 3000 114130 3350
rect 114500 3000 114570 3550
rect 115020 3000 115090 4040
rect 117480 3650 117590 3660
rect 117480 3560 117490 3650
rect 117580 3560 117590 3650
rect 117480 3550 117590 3560
rect 117040 3450 117150 3460
rect 117040 3360 117050 3450
rect 117140 3360 117150 3450
rect 117040 3350 117150 3360
rect 117060 3000 117130 3350
rect 117500 3000 117570 3550
rect 118020 3000 118090 4040
rect 120480 3650 120590 3660
rect 120480 3560 120490 3650
rect 120580 3560 120590 3650
rect 120480 3550 120590 3560
rect 120040 3450 120150 3460
rect 120040 3360 120050 3450
rect 120140 3360 120150 3450
rect 120040 3350 120150 3360
rect 120060 3000 120130 3350
rect 120500 3000 120570 3550
rect 121020 3000 121090 4040
rect 123480 3650 123590 3660
rect 123480 3560 123490 3650
rect 123580 3560 123590 3650
rect 123480 3550 123590 3560
rect 123040 3450 123150 3460
rect 123040 3360 123050 3450
rect 123140 3360 123150 3450
rect 123040 3350 123150 3360
rect 123060 3000 123130 3350
rect 123500 3000 123570 3550
rect 124020 3000 124090 4040
rect 126480 3650 126590 3660
rect 126480 3560 126490 3650
rect 126580 3560 126590 3650
rect 126480 3550 126590 3560
rect 126040 3450 126150 3460
rect 126040 3360 126050 3450
rect 126140 3360 126150 3450
rect 126040 3350 126150 3360
rect 126060 3000 126130 3350
rect 126500 3000 126570 3550
rect 127020 3000 127090 4040
rect 129480 3650 129590 3660
rect 129480 3560 129490 3650
rect 129580 3560 129590 3650
rect 129480 3550 129590 3560
rect 129040 3450 129150 3460
rect 129040 3360 129050 3450
rect 129140 3360 129150 3450
rect 129040 3350 129150 3360
rect 129060 3000 129130 3350
rect 129500 3000 129570 3550
rect 130020 3000 130090 4040
rect 132480 3650 132590 3660
rect 132480 3560 132490 3650
rect 132580 3560 132590 3650
rect 132480 3550 132590 3560
rect 132040 3450 132150 3460
rect 132040 3360 132050 3450
rect 132140 3360 132150 3450
rect 132040 3350 132150 3360
rect 132060 3000 132130 3350
rect 132500 3000 132570 3550
rect 133020 3000 133090 4040
rect 135480 3650 135590 3660
rect 135480 3560 135490 3650
rect 135580 3560 135590 3650
rect 135480 3550 135590 3560
rect 135040 3450 135150 3460
rect 135040 3360 135050 3450
rect 135140 3360 135150 3450
rect 135040 3350 135150 3360
rect 135060 3000 135130 3350
rect 135500 3000 135570 3550
rect 136020 3000 136090 4040
rect 138480 3650 138590 3660
rect 138480 3560 138490 3650
rect 138580 3560 138590 3650
rect 138480 3550 138590 3560
rect 138040 3450 138150 3460
rect 138040 3360 138050 3450
rect 138140 3360 138150 3450
rect 138040 3350 138150 3360
rect 138060 3000 138130 3350
rect 138500 3000 138570 3550
rect 139020 3000 139090 4040
rect 141480 3650 141590 3660
rect 141480 3560 141490 3650
rect 141580 3560 141590 3650
rect 141480 3550 141590 3560
rect 141040 3450 141150 3460
rect 141040 3360 141050 3450
rect 141140 3360 141150 3450
rect 141040 3350 141150 3360
rect 141060 3000 141130 3350
rect 141500 3000 141570 3550
rect 142020 3000 142090 4040
rect 144480 3650 144590 3660
rect 144480 3560 144490 3650
rect 144580 3560 144590 3650
rect 144480 3550 144590 3560
rect 144040 3450 144150 3460
rect 144040 3360 144050 3450
rect 144140 3360 144150 3450
rect 144040 3350 144150 3360
rect 144060 3000 144130 3350
rect 144500 3000 144570 3550
rect 145020 3000 145090 4040
rect 147480 3650 147590 3660
rect 147480 3560 147490 3650
rect 147580 3560 147590 3650
rect 147480 3550 147590 3560
rect 147040 3450 147150 3460
rect 147040 3360 147050 3450
rect 147140 3360 147150 3450
rect 147040 3350 147150 3360
rect 147060 3000 147130 3350
rect 147500 3000 147570 3550
rect 148020 3000 148090 4040
rect -560 1560 -260 1570
rect -560 1490 -540 1560
rect -560 1480 -260 1490
rect -750 160 -740 230
rect -650 160 -640 230
rect -3000 -1440 -1000 -1430
rect -3000 -1510 -1580 -1440
rect -1180 -1510 -1000 -1440
rect -3000 -1520 -1000 -1510
rect -750 -2770 -640 160
rect -560 -1440 -260 -1430
rect -560 -1510 -540 -1440
rect -560 -1520 -260 -1510
rect -750 -2840 -740 -2770
rect -650 -2840 -640 -2770
rect -3000 -4440 -1000 -4430
rect -3000 -4510 -1580 -4440
rect -1180 -4510 -1000 -4440
rect -3000 -4520 -1000 -4510
rect -750 -5770 -640 -2840
rect -560 -4440 -260 -4430
rect -560 -4510 -540 -4440
rect -560 -4520 -260 -4510
rect -750 -5840 -740 -5770
rect -650 -5840 -640 -5770
rect -3000 -7440 -1000 -7430
rect -3000 -7510 -1580 -7440
rect -1180 -7510 -1000 -7440
rect -3000 -7520 -1000 -7510
rect -750 -8770 -640 -5840
rect -560 -7440 -260 -7430
rect -560 -7510 -540 -7440
rect -560 -7520 -260 -7510
rect -750 -8840 -740 -8770
rect -650 -8840 -640 -8770
rect -3000 -10440 -1000 -10430
rect -3000 -10510 -1580 -10440
rect -1180 -10510 -1000 -10440
rect -3000 -10520 -1000 -10510
rect -750 -11770 -640 -8840
rect -560 -10440 -260 -10430
rect -560 -10510 -540 -10440
rect -560 -10520 -260 -10510
rect -750 -11840 -740 -11770
rect -650 -11840 -640 -11770
rect -3000 -13440 -1000 -13430
rect -3000 -13510 -1580 -13440
rect -1180 -13510 -1000 -13440
rect -3000 -13520 -1000 -13510
rect -750 -14770 -640 -11840
rect -560 -13440 -260 -13430
rect -560 -13510 -540 -13440
rect -560 -13520 -260 -13510
rect -750 -14840 -740 -14770
rect -650 -14840 -640 -14770
rect -3000 -16440 -1000 -16430
rect -3000 -16510 -1580 -16440
rect -1180 -16510 -1000 -16440
rect -3000 -16520 -1000 -16510
rect -750 -17770 -640 -14840
rect -560 -16440 -260 -16430
rect -560 -16510 -540 -16440
rect -560 -16520 -260 -16510
rect -750 -17840 -740 -17770
rect -650 -17840 -640 -17770
rect -3000 -19440 -1000 -19430
rect -3000 -19510 -1580 -19440
rect -1180 -19510 -1000 -19440
rect -3000 -19520 -1000 -19510
rect -750 -20770 -640 -17840
rect -560 -19440 -260 -19430
rect -560 -19510 -540 -19440
rect -560 -19520 -260 -19510
rect -750 -20840 -740 -20770
rect -650 -20840 -640 -20770
rect -3000 -22440 -1000 -22430
rect -3000 -22510 -1580 -22440
rect -1180 -22510 -1000 -22440
rect -3000 -22520 -1000 -22510
rect -750 -23770 -640 -20840
rect -560 -22440 -260 -22430
rect -560 -22510 -540 -22440
rect -560 -22520 -260 -22510
rect -750 -23840 -740 -23770
rect -650 -23840 -640 -23770
rect -3000 -25440 -1000 -25430
rect -3000 -25510 -1580 -25440
rect -1180 -25510 -1000 -25440
rect -3000 -25520 -1000 -25510
rect -750 -26770 -640 -23840
rect -560 -25440 -260 -25430
rect -560 -25510 -540 -25440
rect -560 -25520 -260 -25510
rect -750 -26840 -740 -26770
rect -650 -26840 -640 -26770
rect -3000 -28440 -1000 -28430
rect -3000 -28510 -1580 -28440
rect -1180 -28510 -1000 -28440
rect -3000 -28520 -1000 -28510
rect -750 -29770 -640 -26840
rect -560 -28440 -260 -28430
rect -560 -28510 -540 -28440
rect -560 -28520 -260 -28510
rect -750 -29840 -740 -29770
rect -650 -29840 -640 -29770
rect -3000 -31440 -1000 -31430
rect -3000 -31510 -1580 -31440
rect -1180 -31510 -1000 -31440
rect -3000 -31520 -1000 -31510
rect -750 -32770 -640 -29840
rect -560 -31440 -260 -31430
rect -560 -31510 -540 -31440
rect -560 -31520 -260 -31510
rect -750 -32840 -740 -32770
rect -650 -32840 -640 -32770
rect -3000 -34440 -1000 -34430
rect -3000 -34510 -1580 -34440
rect -1180 -34510 -1000 -34440
rect -3000 -34520 -1000 -34510
rect -750 -35770 -640 -32840
rect -560 -34440 -260 -34430
rect -560 -34510 -540 -34440
rect -560 -34520 -260 -34510
rect -750 -35840 -740 -35770
rect -650 -35840 -640 -35770
rect -3000 -37440 -1000 -37430
rect -3000 -37510 -1580 -37440
rect -1180 -37510 -1000 -37440
rect -3000 -37520 -1000 -37510
rect -750 -38770 -640 -35840
rect -560 -37440 -260 -37430
rect -560 -37510 -540 -37440
rect -560 -37520 -260 -37510
rect -750 -38840 -740 -38770
rect -650 -38840 -640 -38770
rect -3000 -40440 -1000 -40430
rect -3000 -40510 -1580 -40440
rect -1180 -40510 -1000 -40440
rect -3000 -40520 -1000 -40510
rect -750 -41770 -640 -38840
rect -560 -40440 -260 -40430
rect -560 -40510 -540 -40440
rect -560 -40520 -260 -40510
rect -750 -41840 -740 -41770
rect -650 -41840 -640 -41770
rect -3000 -43440 -1000 -43430
rect -3000 -43510 -1580 -43440
rect -1180 -43510 -1000 -43440
rect -3000 -43520 -1000 -43510
rect -750 -44770 -640 -41840
rect -560 -43440 -260 -43430
rect -560 -43510 -540 -43440
rect -560 -43520 -260 -43510
rect -750 -44840 -740 -44770
rect -650 -44840 -640 -44770
rect -3000 -46440 -1000 -46430
rect -3000 -46510 -1580 -46440
rect -1180 -46510 -1000 -46440
rect -3000 -46520 -1000 -46510
rect -750 -47770 -640 -44840
rect -560 -46440 -260 -46430
rect -560 -46510 -540 -46440
rect -560 -46520 -260 -46510
rect -750 -47840 -740 -47770
rect -650 -47840 -640 -47770
rect -3000 -49440 -1000 -49430
rect -3000 -49510 -1580 -49440
rect -1180 -49510 -1000 -49440
rect -3000 -49520 -1000 -49510
rect -750 -50770 -640 -47840
rect -560 -49440 -260 -49430
rect -560 -49510 -540 -49440
rect -560 -49520 -260 -49510
rect -750 -50840 -740 -50770
rect -650 -50840 -640 -50770
rect -3000 -52440 -1000 -52430
rect -3000 -52510 -1580 -52440
rect -1180 -52510 -1000 -52440
rect -3000 -52520 -1000 -52510
rect -750 -53770 -640 -50840
rect -560 -52440 -260 -52430
rect -560 -52510 -540 -52440
rect -560 -52520 -260 -52510
rect -750 -53840 -740 -53770
rect -650 -53840 -640 -53770
rect -3000 -55440 -1000 -55430
rect -3000 -55510 -1580 -55440
rect -1180 -55510 -1000 -55440
rect -3000 -55520 -1000 -55510
rect -750 -56770 -640 -53840
rect -560 -55440 -260 -55430
rect -560 -55510 -540 -55440
rect -560 -55520 -260 -55510
rect -750 -56840 -740 -56770
rect -650 -56840 -640 -56770
rect -3000 -58440 -1000 -58430
rect -3000 -58510 -1580 -58440
rect -1180 -58510 -1000 -58440
rect -3000 -58520 -1000 -58510
rect -750 -59770 -640 -56840
rect -560 -58440 -260 -58430
rect -560 -58510 -540 -58440
rect -560 -58520 -260 -58510
rect -750 -59840 -740 -59770
rect -650 -59840 -640 -59770
rect -3000 -61440 -1000 -61430
rect -3000 -61510 -1580 -61440
rect -1180 -61510 -1000 -61440
rect -3000 -61520 -1000 -61510
rect -750 -62770 -640 -59840
rect -560 -61440 -260 -61430
rect -560 -61510 -540 -61440
rect -560 -61520 -260 -61510
rect -750 -62840 -740 -62770
rect -650 -62840 -640 -62770
rect -3000 -64440 -1000 -64430
rect -3000 -64510 -1580 -64440
rect -1180 -64510 -1000 -64440
rect -3000 -64520 -1000 -64510
rect -750 -65770 -640 -62840
rect -560 -64440 -260 -64430
rect -560 -64510 -540 -64440
rect -560 -64520 -260 -64510
rect -750 -65840 -740 -65770
rect -650 -65840 -640 -65770
rect -3000 -67440 -1000 -67430
rect -3000 -67510 -1580 -67440
rect -1180 -67510 -1000 -67440
rect -3000 -67520 -1000 -67510
rect -750 -68770 -640 -65840
rect -560 -67440 -260 -67430
rect -560 -67510 -540 -67440
rect -560 -67520 -260 -67510
rect -750 -68840 -740 -68770
rect -650 -68840 -640 -68770
rect -3000 -70440 -1000 -70430
rect -3000 -70510 -1580 -70440
rect -1180 -70510 -1000 -70440
rect -3000 -70520 -1000 -70510
rect -750 -71770 -640 -68840
rect -560 -70440 -260 -70430
rect -560 -70510 -540 -70440
rect -560 -70520 -260 -70510
rect -750 -71840 -740 -71770
rect -650 -71840 -640 -71770
rect -3000 -73440 -1000 -73430
rect -3000 -73510 -1580 -73440
rect -1180 -73510 -1000 -73440
rect -3000 -73520 -1000 -73510
rect -750 -74770 -640 -71840
rect -560 -73440 -260 -73430
rect -560 -73510 -540 -73440
rect -560 -73520 -260 -73510
rect -750 -74840 -740 -74770
rect -650 -74840 -640 -74770
rect -3000 -76440 -1000 -76430
rect -3000 -76510 -1580 -76440
rect -1180 -76510 -1000 -76440
rect -3000 -76520 -1000 -76510
rect -750 -77770 -640 -74840
rect -560 -76440 -260 -76430
rect -560 -76510 -540 -76440
rect -560 -76520 -260 -76510
rect -750 -77840 -740 -77770
rect -650 -77840 -640 -77770
rect -3000 -79440 -1000 -79430
rect -3000 -79510 -1580 -79440
rect -1180 -79510 -1000 -79440
rect -3000 -79520 -1000 -79510
rect -750 -80770 -640 -77840
rect -560 -79440 -260 -79430
rect -560 -79510 -540 -79440
rect -560 -79520 -260 -79510
rect -750 -80840 -740 -80770
rect -650 -80840 -640 -80770
rect -3000 -82440 -1000 -82430
rect -3000 -82510 -1580 -82440
rect -1180 -82510 -1000 -82440
rect -3000 -82520 -1000 -82510
rect -750 -83770 -640 -80840
rect -560 -82440 -260 -82430
rect -560 -82510 -540 -82440
rect -560 -82520 -260 -82510
rect -750 -83840 -740 -83770
rect -650 -83840 -640 -83770
rect -3000 -85440 -1000 -85430
rect -3000 -85510 -1580 -85440
rect -1180 -85510 -1000 -85440
rect -3000 -85520 -1000 -85510
rect -750 -86770 -640 -83840
rect -560 -85440 -260 -85430
rect -560 -85510 -540 -85440
rect -560 -85520 -260 -85510
rect -750 -86840 -740 -86770
rect -650 -86840 -640 -86770
rect -3000 -88440 -1000 -88430
rect -3000 -88510 -1580 -88440
rect -1180 -88510 -1000 -88440
rect -3000 -88520 -1000 -88510
rect -750 -89770 -640 -86840
rect -560 -88440 -260 -88430
rect -560 -88510 -540 -88440
rect -560 -88520 -260 -88510
rect -750 -89840 -740 -89770
rect -650 -89840 -640 -89770
rect -3000 -91440 -1000 -91430
rect -3000 -91510 -1580 -91440
rect -1180 -91510 -1000 -91440
rect -3000 -91520 -1000 -91510
rect -750 -92770 -640 -89840
rect -560 -91440 -260 -91430
rect -560 -91510 -540 -91440
rect -560 -91520 -260 -91510
rect -750 -92840 -740 -92770
rect -650 -92840 -640 -92770
rect -3000 -94440 -1000 -94430
rect -3000 -94510 -1580 -94440
rect -1180 -94510 -1000 -94440
rect -3000 -94520 -1000 -94510
rect -750 -95770 -640 -92840
rect -560 -94440 -260 -94430
rect -560 -94510 -540 -94440
rect -560 -94520 -260 -94510
rect -750 -95840 -740 -95770
rect -650 -95840 -640 -95770
rect -3000 -97440 -1000 -97430
rect -3000 -97510 -1580 -97440
rect -1180 -97510 -1000 -97440
rect -3000 -97520 -1000 -97510
rect -750 -98770 -640 -95840
rect -560 -97440 -260 -97430
rect -560 -97510 -540 -97440
rect -560 -97520 -260 -97510
rect -750 -98840 -740 -98770
rect -650 -98840 -640 -98770
rect -3000 -100440 -1000 -100430
rect -3000 -100510 -1580 -100440
rect -1180 -100510 -1000 -100440
rect -3000 -100520 -1000 -100510
rect -750 -101770 -640 -98840
rect -560 -100440 -260 -100430
rect -560 -100510 -540 -100440
rect -560 -100520 -260 -100510
rect -750 -101840 -740 -101770
rect -650 -101840 -640 -101770
rect -3000 -103440 -1000 -103430
rect -3000 -103510 -1580 -103440
rect -1180 -103510 -1000 -103440
rect -3000 -103520 -1000 -103510
rect -750 -104770 -640 -101840
rect -560 -103440 -260 -103430
rect -560 -103510 -540 -103440
rect -560 -103520 -260 -103510
rect -750 -104840 -740 -104770
rect -650 -104840 -640 -104770
rect -3000 -106440 -1000 -106430
rect -3000 -106510 -1580 -106440
rect -1180 -106510 -1000 -106440
rect -3000 -106520 -1000 -106510
rect -750 -107770 -640 -104840
rect -560 -106440 -260 -106430
rect -560 -106510 -540 -106440
rect -560 -106520 -260 -106510
rect -750 -107840 -740 -107770
rect -650 -107840 -640 -107770
rect -3000 -109440 -1000 -109430
rect -3000 -109510 -1580 -109440
rect -1180 -109510 -1000 -109440
rect -3000 -109520 -1000 -109510
rect -750 -110770 -640 -107840
rect -560 -109440 -260 -109430
rect -560 -109510 -540 -109440
rect -560 -109520 -260 -109510
rect -750 -110840 -740 -110770
rect -650 -110840 -640 -110770
rect -3000 -112440 -1000 -112430
rect -3000 -112510 -1580 -112440
rect -1180 -112510 -1000 -112440
rect -3000 -112520 -1000 -112510
rect -750 -113770 -640 -110840
rect -560 -112440 -260 -112430
rect -560 -112510 -540 -112440
rect -560 -112520 -260 -112510
rect -750 -113840 -740 -113770
rect -650 -113840 -640 -113770
rect -3000 -115440 -1000 -115430
rect -3000 -115510 -1580 -115440
rect -1180 -115510 -1000 -115440
rect -3000 -115520 -1000 -115510
rect -750 -116770 -640 -113840
rect -560 -115440 -260 -115430
rect -560 -115510 -540 -115440
rect -560 -115520 -260 -115510
rect -750 -116840 -740 -116770
rect -650 -116840 -640 -116770
rect -3000 -118440 -1000 -118430
rect -3000 -118510 -1580 -118440
rect -1180 -118510 -1000 -118440
rect -3000 -118520 -1000 -118510
rect -750 -119770 -640 -116840
rect -560 -118440 -260 -118430
rect -560 -118510 -540 -118440
rect -560 -118520 -260 -118510
rect -750 -119840 -740 -119770
rect -650 -119840 -640 -119770
rect -3000 -121440 -1000 -121430
rect -3000 -121510 -1580 -121440
rect -1180 -121510 -1000 -121440
rect -3000 -121520 -1000 -121510
rect -750 -122770 -640 -119840
rect -560 -121440 -260 -121430
rect -560 -121510 -540 -121440
rect -560 -121520 -260 -121510
rect -750 -122840 -740 -122770
rect -650 -122840 -640 -122770
rect -3000 -124440 -1000 -124430
rect -3000 -124510 -1580 -124440
rect -1180 -124510 -1000 -124440
rect -3000 -124520 -1000 -124510
rect -750 -125770 -640 -122840
rect -560 -124440 -260 -124430
rect -560 -124510 -540 -124440
rect -560 -124520 -260 -124510
rect -750 -125840 -740 -125770
rect -650 -125840 -640 -125770
rect -3000 -127440 -1000 -127430
rect -3000 -127510 -1580 -127440
rect -1180 -127510 -1000 -127440
rect -3000 -127520 -1000 -127510
rect -750 -128770 -640 -125840
rect -560 -127440 -260 -127430
rect -560 -127510 -540 -127440
rect -560 -127520 -260 -127510
rect -750 -128840 -740 -128770
rect -650 -128840 -640 -128770
rect -3000 -130440 -1000 -130430
rect -3000 -130510 -1580 -130440
rect -1180 -130510 -1000 -130440
rect -3000 -130520 -1000 -130510
rect -750 -131770 -640 -128840
rect -560 -130440 -260 -130430
rect -560 -130510 -540 -130440
rect -560 -130520 -260 -130510
rect -750 -131840 -740 -131770
rect -650 -131840 -640 -131770
rect -3000 -133440 -1000 -133430
rect -3000 -133510 -1580 -133440
rect -1180 -133510 -1000 -133440
rect -3000 -133520 -1000 -133510
rect -750 -134770 -640 -131840
rect -560 -133440 -260 -133430
rect -560 -133510 -540 -133440
rect -560 -133520 -260 -133510
rect -750 -134840 -740 -134770
rect -650 -134840 -640 -134770
rect -3000 -136440 -1000 -136430
rect -3000 -136510 -1580 -136440
rect -1180 -136510 -1000 -136440
rect -3000 -136520 -1000 -136510
rect -750 -137770 -640 -134840
rect -560 -136440 -260 -136430
rect -560 -136510 -540 -136440
rect -560 -136520 -260 -136510
rect -750 -137840 -740 -137770
rect -650 -137840 -640 -137770
rect -3000 -139440 -1000 -139430
rect -3000 -139510 -1580 -139440
rect -1180 -139510 -1000 -139440
rect -3000 -139520 -1000 -139510
rect -750 -140770 -640 -137840
rect -560 -139440 -260 -139430
rect -560 -139510 -540 -139440
rect -560 -139520 -260 -139510
rect -750 -140840 -740 -140770
rect -650 -140840 -640 -140770
rect -3000 -142440 -1000 -142430
rect -3000 -142510 -1580 -142440
rect -1180 -142510 -1000 -142440
rect -3000 -142520 -1000 -142510
rect -750 -143770 -640 -140840
rect -560 -142440 -260 -142430
rect -560 -142510 -540 -142440
rect -560 -142520 -260 -142510
rect -750 -143840 -740 -143770
rect -650 -143840 -640 -143770
rect -3000 -145440 -1000 -145430
rect -3000 -145510 -1580 -145440
rect -1180 -145510 -1000 -145440
rect -3000 -145520 -1000 -145510
rect -750 -146770 -640 -143840
rect -560 -145440 -260 -145430
rect -560 -145510 -540 -145440
rect -560 -145520 -260 -145510
rect -750 -146840 -740 -146770
rect -650 -146840 -640 -146770
rect -750 -147000 -640 -146840
rect 540 -147080 2780 -147060
rect 540 -147200 560 -147080
rect 2760 -147180 2780 -147080
rect 2120 -147200 2780 -147180
rect 3540 -147080 5780 -147060
rect 3540 -147200 3560 -147080
rect 5760 -147180 5780 -147080
rect 5120 -147200 5780 -147180
rect 6540 -147080 8780 -147060
rect 6540 -147200 6560 -147080
rect 8760 -147180 8780 -147080
rect 8120 -147200 8780 -147180
rect 9540 -147080 11780 -147060
rect 9540 -147200 9560 -147080
rect 11760 -147180 11780 -147080
rect 11120 -147200 11780 -147180
rect 12540 -147080 14780 -147060
rect 12540 -147200 12560 -147080
rect 14760 -147180 14780 -147080
rect 14120 -147200 14780 -147180
rect 15540 -147080 17780 -147060
rect 15540 -147200 15560 -147080
rect 17760 -147180 17780 -147080
rect 17120 -147200 17780 -147180
rect 18540 -147080 20780 -147060
rect 18540 -147200 18560 -147080
rect 20760 -147180 20780 -147080
rect 20120 -147200 20780 -147180
rect 21540 -147080 23780 -147060
rect 21540 -147200 21560 -147080
rect 23760 -147180 23780 -147080
rect 23120 -147200 23780 -147180
rect 24540 -147080 26780 -147060
rect 24540 -147200 24560 -147080
rect 26760 -147180 26780 -147080
rect 26120 -147200 26780 -147180
rect 27540 -147080 29780 -147060
rect 27540 -147200 27560 -147080
rect 29760 -147180 29780 -147080
rect 29120 -147200 29780 -147180
rect 30540 -147080 32780 -147060
rect 30540 -147200 30560 -147080
rect 32760 -147180 32780 -147080
rect 32120 -147200 32780 -147180
rect 33540 -147080 35780 -147060
rect 33540 -147200 33560 -147080
rect 35760 -147180 35780 -147080
rect 35120 -147200 35780 -147180
rect 36540 -147080 38780 -147060
rect 36540 -147200 36560 -147080
rect 38760 -147180 38780 -147080
rect 38120 -147200 38780 -147180
rect 39540 -147080 41780 -147060
rect 39540 -147200 39560 -147080
rect 41760 -147180 41780 -147080
rect 41120 -147200 41780 -147180
rect 42540 -147080 44780 -147060
rect 42540 -147200 42560 -147080
rect 44760 -147180 44780 -147080
rect 44120 -147200 44780 -147180
rect 45540 -147080 47780 -147060
rect 45540 -147200 45560 -147080
rect 47760 -147180 47780 -147080
rect 47120 -147200 47780 -147180
rect 48540 -147080 50780 -147060
rect 48540 -147200 48560 -147080
rect 50760 -147180 50780 -147080
rect 50120 -147200 50780 -147180
rect 51540 -147080 53780 -147060
rect 51540 -147200 51560 -147080
rect 53760 -147180 53780 -147080
rect 53120 -147200 53780 -147180
rect 54540 -147080 56780 -147060
rect 54540 -147200 54560 -147080
rect 56760 -147180 56780 -147080
rect 56120 -147200 56780 -147180
rect 57540 -147080 59780 -147060
rect 57540 -147200 57560 -147080
rect 59760 -147180 59780 -147080
rect 59120 -147200 59780 -147180
rect 60540 -147080 62780 -147060
rect 60540 -147200 60560 -147080
rect 62760 -147180 62780 -147080
rect 62120 -147200 62780 -147180
rect 63540 -147080 65780 -147060
rect 63540 -147200 63560 -147080
rect 65760 -147180 65780 -147080
rect 65120 -147200 65780 -147180
rect 66540 -147080 68780 -147060
rect 66540 -147200 66560 -147080
rect 68760 -147180 68780 -147080
rect 68120 -147200 68780 -147180
rect 69540 -147080 71780 -147060
rect 69540 -147200 69560 -147080
rect 71760 -147180 71780 -147080
rect 71120 -147200 71780 -147180
rect 72540 -147080 74780 -147060
rect 72540 -147200 72560 -147080
rect 74760 -147180 74780 -147080
rect 74120 -147200 74780 -147180
rect 75540 -147080 77780 -147060
rect 75540 -147200 75560 -147080
rect 77760 -147180 77780 -147080
rect 77120 -147200 77780 -147180
rect 78540 -147080 80780 -147060
rect 78540 -147200 78560 -147080
rect 80760 -147180 80780 -147080
rect 80120 -147200 80780 -147180
rect 81540 -147080 83780 -147060
rect 81540 -147200 81560 -147080
rect 83760 -147180 83780 -147080
rect 83120 -147200 83780 -147180
rect 84540 -147080 86780 -147060
rect 84540 -147200 84560 -147080
rect 86760 -147180 86780 -147080
rect 86120 -147200 86780 -147180
rect 87540 -147080 89780 -147060
rect 87540 -147200 87560 -147080
rect 89760 -147180 89780 -147080
rect 89120 -147200 89780 -147180
rect 90540 -147080 92780 -147060
rect 90540 -147200 90560 -147080
rect 92760 -147180 92780 -147080
rect 92120 -147200 92780 -147180
rect 93540 -147080 95780 -147060
rect 93540 -147200 93560 -147080
rect 95760 -147180 95780 -147080
rect 95120 -147200 95780 -147180
rect 96540 -147080 98780 -147060
rect 96540 -147200 96560 -147080
rect 98760 -147180 98780 -147080
rect 98120 -147200 98780 -147180
rect 99540 -147080 101780 -147060
rect 99540 -147200 99560 -147080
rect 101760 -147180 101780 -147080
rect 101120 -147200 101780 -147180
rect 102540 -147080 104780 -147060
rect 102540 -147200 102560 -147080
rect 104760 -147180 104780 -147080
rect 104120 -147200 104780 -147180
rect 105540 -147080 107780 -147060
rect 105540 -147200 105560 -147080
rect 107760 -147180 107780 -147080
rect 107120 -147200 107780 -147180
rect 108540 -147080 110780 -147060
rect 108540 -147200 108560 -147080
rect 110760 -147180 110780 -147080
rect 110120 -147200 110780 -147180
rect 111540 -147080 113780 -147060
rect 111540 -147200 111560 -147080
rect 113760 -147180 113780 -147080
rect 113120 -147200 113780 -147180
rect 114540 -147080 116780 -147060
rect 114540 -147200 114560 -147080
rect 116760 -147180 116780 -147080
rect 116120 -147200 116780 -147180
rect 117540 -147080 119780 -147060
rect 117540 -147200 117560 -147080
rect 119760 -147180 119780 -147080
rect 119120 -147200 119780 -147180
rect 120540 -147080 122780 -147060
rect 120540 -147200 120560 -147080
rect 122760 -147180 122780 -147080
rect 122120 -147200 122780 -147180
rect 123540 -147080 125780 -147060
rect 123540 -147200 123560 -147080
rect 125760 -147180 125780 -147080
rect 125120 -147200 125780 -147180
rect 126540 -147080 128780 -147060
rect 126540 -147200 126560 -147080
rect 128760 -147180 128780 -147080
rect 128120 -147200 128780 -147180
rect 129540 -147080 131780 -147060
rect 129540 -147200 129560 -147080
rect 131760 -147180 131780 -147080
rect 131120 -147200 131780 -147180
rect 132540 -147080 134780 -147060
rect 132540 -147200 132560 -147080
rect 134760 -147180 134780 -147080
rect 134120 -147200 134780 -147180
rect 135540 -147080 137780 -147060
rect 135540 -147200 135560 -147080
rect 137760 -147180 137780 -147080
rect 137120 -147200 137780 -147180
rect 138540 -147080 140780 -147060
rect 138540 -147200 138560 -147080
rect 140760 -147180 140780 -147080
rect 140120 -147200 140780 -147180
rect 141540 -147080 143780 -147060
rect 141540 -147200 141560 -147080
rect 143760 -147180 143780 -147080
rect 143120 -147200 143780 -147180
rect 144540 -147080 146780 -147060
rect 144540 -147200 144560 -147080
rect 146760 -147180 146780 -147080
rect 146120 -147200 146780 -147180
rect 147540 -147080 149780 -147060
rect 147540 -147200 147560 -147080
rect 149760 -147180 149780 -147080
rect 149120 -147200 149780 -147180
rect 220 -147500 440 -147490
rect 220 -147700 240 -147500
rect 420 -147700 440 -147500
rect 220 -147710 440 -147700
rect 3220 -147500 3440 -147490
rect 3220 -147700 3240 -147500
rect 3420 -147700 3440 -147500
rect 3220 -147710 3440 -147700
rect 6220 -147500 6440 -147490
rect 6220 -147700 6240 -147500
rect 6420 -147700 6440 -147500
rect 6220 -147710 6440 -147700
rect 9220 -147500 9440 -147490
rect 9220 -147700 9240 -147500
rect 9420 -147700 9440 -147500
rect 9220 -147710 9440 -147700
rect 12220 -147500 12440 -147490
rect 12220 -147700 12240 -147500
rect 12420 -147700 12440 -147500
rect 12220 -147710 12440 -147700
rect 15220 -147500 15440 -147490
rect 15220 -147700 15240 -147500
rect 15420 -147700 15440 -147500
rect 15220 -147710 15440 -147700
rect 18220 -147500 18440 -147490
rect 18220 -147700 18240 -147500
rect 18420 -147700 18440 -147500
rect 18220 -147710 18440 -147700
rect 21220 -147500 21440 -147490
rect 21220 -147700 21240 -147500
rect 21420 -147700 21440 -147500
rect 21220 -147710 21440 -147700
rect 24220 -147500 24440 -147490
rect 24220 -147700 24240 -147500
rect 24420 -147700 24440 -147500
rect 24220 -147710 24440 -147700
rect 27220 -147500 27440 -147490
rect 27220 -147700 27240 -147500
rect 27420 -147700 27440 -147500
rect 27220 -147710 27440 -147700
rect 30220 -147500 30440 -147490
rect 30220 -147700 30240 -147500
rect 30420 -147700 30440 -147500
rect 30220 -147710 30440 -147700
rect 33220 -147500 33440 -147490
rect 33220 -147700 33240 -147500
rect 33420 -147700 33440 -147500
rect 33220 -147710 33440 -147700
rect 36220 -147500 36440 -147490
rect 36220 -147700 36240 -147500
rect 36420 -147700 36440 -147500
rect 36220 -147710 36440 -147700
rect 39220 -147500 39440 -147490
rect 39220 -147700 39240 -147500
rect 39420 -147700 39440 -147500
rect 39220 -147710 39440 -147700
rect 42220 -147500 42440 -147490
rect 42220 -147700 42240 -147500
rect 42420 -147700 42440 -147500
rect 42220 -147710 42440 -147700
rect 45220 -147500 45440 -147490
rect 45220 -147700 45240 -147500
rect 45420 -147700 45440 -147500
rect 45220 -147710 45440 -147700
rect 48220 -147500 48440 -147490
rect 48220 -147700 48240 -147500
rect 48420 -147700 48440 -147500
rect 48220 -147710 48440 -147700
rect 51220 -147500 51440 -147490
rect 51220 -147700 51240 -147500
rect 51420 -147700 51440 -147500
rect 51220 -147710 51440 -147700
rect 54220 -147500 54440 -147490
rect 54220 -147700 54240 -147500
rect 54420 -147700 54440 -147500
rect 54220 -147710 54440 -147700
rect 57220 -147500 57440 -147490
rect 57220 -147700 57240 -147500
rect 57420 -147700 57440 -147500
rect 57220 -147710 57440 -147700
rect 60220 -147500 60440 -147490
rect 60220 -147700 60240 -147500
rect 60420 -147700 60440 -147500
rect 60220 -147710 60440 -147700
rect 63220 -147500 63440 -147490
rect 63220 -147700 63240 -147500
rect 63420 -147700 63440 -147500
rect 63220 -147710 63440 -147700
rect 66220 -147500 66440 -147490
rect 66220 -147700 66240 -147500
rect 66420 -147700 66440 -147500
rect 66220 -147710 66440 -147700
rect 69220 -147500 69440 -147490
rect 69220 -147700 69240 -147500
rect 69420 -147700 69440 -147500
rect 69220 -147710 69440 -147700
rect 72220 -147500 72440 -147490
rect 72220 -147700 72240 -147500
rect 72420 -147700 72440 -147500
rect 72220 -147710 72440 -147700
rect 75220 -147500 75440 -147490
rect 75220 -147700 75240 -147500
rect 75420 -147700 75440 -147500
rect 75220 -147710 75440 -147700
rect 78220 -147500 78440 -147490
rect 78220 -147700 78240 -147500
rect 78420 -147700 78440 -147500
rect 78220 -147710 78440 -147700
rect 81220 -147500 81440 -147490
rect 81220 -147700 81240 -147500
rect 81420 -147700 81440 -147500
rect 81220 -147710 81440 -147700
rect 84220 -147500 84440 -147490
rect 84220 -147700 84240 -147500
rect 84420 -147700 84440 -147500
rect 84220 -147710 84440 -147700
rect 87220 -147500 87440 -147490
rect 87220 -147700 87240 -147500
rect 87420 -147700 87440 -147500
rect 87220 -147710 87440 -147700
rect 90220 -147500 90440 -147490
rect 90220 -147700 90240 -147500
rect 90420 -147700 90440 -147500
rect 90220 -147710 90440 -147700
rect 93220 -147500 93440 -147490
rect 93220 -147700 93240 -147500
rect 93420 -147700 93440 -147500
rect 93220 -147710 93440 -147700
rect 96220 -147500 96440 -147490
rect 96220 -147700 96240 -147500
rect 96420 -147700 96440 -147500
rect 96220 -147710 96440 -147700
rect 99220 -147500 99440 -147490
rect 99220 -147700 99240 -147500
rect 99420 -147700 99440 -147500
rect 99220 -147710 99440 -147700
rect 102220 -147500 102440 -147490
rect 102220 -147700 102240 -147500
rect 102420 -147700 102440 -147500
rect 102220 -147710 102440 -147700
rect 105220 -147500 105440 -147490
rect 105220 -147700 105240 -147500
rect 105420 -147700 105440 -147500
rect 105220 -147710 105440 -147700
rect 108220 -147500 108440 -147490
rect 108220 -147700 108240 -147500
rect 108420 -147700 108440 -147500
rect 108220 -147710 108440 -147700
rect 111220 -147500 111440 -147490
rect 111220 -147700 111240 -147500
rect 111420 -147700 111440 -147500
rect 111220 -147710 111440 -147700
rect 114220 -147500 114440 -147490
rect 114220 -147700 114240 -147500
rect 114420 -147700 114440 -147500
rect 114220 -147710 114440 -147700
rect 117220 -147500 117440 -147490
rect 117220 -147700 117240 -147500
rect 117420 -147700 117440 -147500
rect 117220 -147710 117440 -147700
rect 120220 -147500 120440 -147490
rect 120220 -147700 120240 -147500
rect 120420 -147700 120440 -147500
rect 120220 -147710 120440 -147700
rect 123220 -147500 123440 -147490
rect 123220 -147700 123240 -147500
rect 123420 -147700 123440 -147500
rect 123220 -147710 123440 -147700
rect 126220 -147500 126440 -147490
rect 126220 -147700 126240 -147500
rect 126420 -147700 126440 -147500
rect 126220 -147710 126440 -147700
rect 129220 -147500 129440 -147490
rect 129220 -147700 129240 -147500
rect 129420 -147700 129440 -147500
rect 129220 -147710 129440 -147700
rect 132220 -147500 132440 -147490
rect 132220 -147700 132240 -147500
rect 132420 -147700 132440 -147500
rect 132220 -147710 132440 -147700
rect 135220 -147500 135440 -147490
rect 135220 -147700 135240 -147500
rect 135420 -147700 135440 -147500
rect 135220 -147710 135440 -147700
rect 138220 -147500 138440 -147490
rect 138220 -147700 138240 -147500
rect 138420 -147700 138440 -147500
rect 138220 -147710 138440 -147700
rect 141220 -147500 141440 -147490
rect 141220 -147700 141240 -147500
rect 141420 -147700 141440 -147500
rect 141220 -147710 141440 -147700
rect 144220 -147500 144440 -147490
rect 144220 -147700 144240 -147500
rect 144420 -147700 144440 -147500
rect 144220 -147710 144440 -147700
rect 147220 -147500 147440 -147490
rect 147220 -147700 147240 -147500
rect 147420 -147700 147440 -147500
rect 147220 -147710 147440 -147700
rect 540 -147920 150740 -147900
rect 540 -148080 560 -147920
rect 540 -148100 150740 -148080
<< via2 >>
rect 490 3560 580 3650
rect 3490 3560 3580 3650
rect 6490 3560 6580 3650
rect 9490 3560 9580 3650
rect 12490 3560 12580 3650
rect 15490 3560 15580 3650
rect 18490 3560 18580 3650
rect 21490 3560 21580 3650
rect 24490 3560 24580 3650
rect 27490 3560 27580 3650
rect 30490 3560 30580 3650
rect 33490 3560 33580 3650
rect 36490 3560 36580 3650
rect 39490 3560 39580 3650
rect 42490 3560 42580 3650
rect 45490 3560 45580 3650
rect 48490 3560 48580 3650
rect 51490 3560 51580 3650
rect 54490 3560 54580 3650
rect 57490 3560 57580 3650
rect 60490 3560 60580 3650
rect 63490 3560 63580 3650
rect 66490 3560 66580 3650
rect 69490 3560 69580 3650
rect 72490 3560 72580 3650
rect 75490 3560 75580 3650
rect 78490 3560 78580 3650
rect 81490 3560 81580 3650
rect 84490 3560 84580 3650
rect 87490 3560 87580 3650
rect 90490 3560 90580 3650
rect 93490 3560 93580 3650
rect 96490 3560 96580 3650
rect 99490 3560 99580 3650
rect 102490 3560 102580 3650
rect 105490 3560 105580 3650
rect 108490 3560 108580 3650
rect 111490 3560 111580 3650
rect 114490 3560 114580 3650
rect 117490 3560 117580 3650
rect 120490 3560 120580 3650
rect 123490 3560 123580 3650
rect 126490 3560 126580 3650
rect 129490 3560 129580 3650
rect 132490 3560 132580 3650
rect 135490 3560 135580 3650
rect 138490 3560 138580 3650
rect 141490 3560 141580 3650
rect 144490 3560 144580 3650
rect 147490 3560 147580 3650
rect -540 1490 -260 1560
rect -740 160 -650 230
rect -540 -1510 -260 -1440
rect -740 -2840 -650 -2770
rect -540 -4510 -260 -4440
rect -740 -5840 -650 -5770
rect -540 -7510 -260 -7440
rect -740 -8840 -650 -8770
rect -540 -10510 -260 -10440
rect -740 -11840 -650 -11770
rect -540 -13510 -260 -13440
rect -740 -14840 -650 -14770
rect -540 -16510 -260 -16440
rect -740 -17840 -650 -17770
rect -540 -19510 -260 -19440
rect -740 -20840 -650 -20770
rect -540 -22510 -260 -22440
rect -740 -23840 -650 -23770
rect -540 -25510 -260 -25440
rect -740 -26840 -650 -26770
rect -540 -28510 -260 -28440
rect -740 -29840 -650 -29770
rect -540 -31510 -260 -31440
rect -740 -32840 -650 -32770
rect -540 -34510 -260 -34440
rect -740 -35840 -650 -35770
rect -540 -37510 -260 -37440
rect -740 -38840 -650 -38770
rect -540 -40510 -260 -40440
rect -740 -41840 -650 -41770
rect -540 -43510 -260 -43440
rect -740 -44840 -650 -44770
rect -540 -46510 -260 -46440
rect -740 -47840 -650 -47770
rect -540 -49510 -260 -49440
rect -740 -50840 -650 -50770
rect -540 -52510 -260 -52440
rect -740 -53840 -650 -53770
rect -540 -55510 -260 -55440
rect -740 -56840 -650 -56770
rect -540 -58510 -260 -58440
rect -740 -59840 -650 -59770
rect -540 -61510 -260 -61440
rect -740 -62840 -650 -62770
rect -540 -64510 -260 -64440
rect -740 -65840 -650 -65770
rect -540 -67510 -260 -67440
rect -740 -68840 -650 -68770
rect -540 -70510 -260 -70440
rect -740 -71840 -650 -71770
rect -540 -73510 -260 -73440
rect -740 -74840 -650 -74770
rect -540 -76510 -260 -76440
rect -740 -77840 -650 -77770
rect -540 -79510 -260 -79440
rect -740 -80840 -650 -80770
rect -540 -82510 -260 -82440
rect -740 -83840 -650 -83770
rect -540 -85510 -260 -85440
rect -740 -86840 -650 -86770
rect -540 -88510 -260 -88440
rect -740 -89840 -650 -89770
rect -540 -91510 -260 -91440
rect -740 -92840 -650 -92770
rect -540 -94510 -260 -94440
rect -740 -95840 -650 -95770
rect -540 -97510 -260 -97440
rect -740 -98840 -650 -98770
rect -540 -100510 -260 -100440
rect -740 -101840 -650 -101770
rect -540 -103510 -260 -103440
rect -740 -104840 -650 -104770
rect -540 -106510 -260 -106440
rect -740 -107840 -650 -107770
rect -540 -109510 -260 -109440
rect -740 -110840 -650 -110770
rect -540 -112510 -260 -112440
rect -740 -113840 -650 -113770
rect -540 -115510 -260 -115440
rect -740 -116840 -650 -116770
rect -540 -118510 -260 -118440
rect -740 -119840 -650 -119770
rect -540 -121510 -260 -121440
rect -740 -122840 -650 -122770
rect -540 -124510 -260 -124440
rect -740 -125840 -650 -125770
rect -540 -127510 -260 -127440
rect -740 -128840 -650 -128770
rect -540 -130510 -260 -130440
rect -740 -131840 -650 -131770
rect -540 -133510 -260 -133440
rect -740 -134840 -650 -134770
rect -540 -136510 -260 -136440
rect -740 -137840 -650 -137770
rect -540 -139510 -260 -139440
rect -740 -140840 -650 -140770
rect -540 -142510 -260 -142440
rect -740 -143840 -650 -143770
rect -540 -145510 -260 -145440
rect -740 -146840 -650 -146770
rect 560 -147130 2760 -147080
rect 560 -147180 2120 -147130
rect 2120 -147180 2760 -147130
rect 3560 -147130 5760 -147080
rect 3560 -147180 5120 -147130
rect 5120 -147180 5760 -147130
rect 6560 -147130 8760 -147080
rect 6560 -147180 8120 -147130
rect 8120 -147180 8760 -147130
rect 9560 -147130 11760 -147080
rect 9560 -147180 11120 -147130
rect 11120 -147180 11760 -147130
rect 12560 -147130 14760 -147080
rect 12560 -147180 14120 -147130
rect 14120 -147180 14760 -147130
rect 15560 -147130 17760 -147080
rect 15560 -147180 17120 -147130
rect 17120 -147180 17760 -147130
rect 18560 -147130 20760 -147080
rect 18560 -147180 20120 -147130
rect 20120 -147180 20760 -147130
rect 21560 -147130 23760 -147080
rect 21560 -147180 23120 -147130
rect 23120 -147180 23760 -147130
rect 24560 -147130 26760 -147080
rect 24560 -147180 26120 -147130
rect 26120 -147180 26760 -147130
rect 27560 -147130 29760 -147080
rect 27560 -147180 29120 -147130
rect 29120 -147180 29760 -147130
rect 30560 -147130 32760 -147080
rect 30560 -147180 32120 -147130
rect 32120 -147180 32760 -147130
rect 33560 -147130 35760 -147080
rect 33560 -147180 35120 -147130
rect 35120 -147180 35760 -147130
rect 36560 -147130 38760 -147080
rect 36560 -147180 38120 -147130
rect 38120 -147180 38760 -147130
rect 39560 -147130 41760 -147080
rect 39560 -147180 41120 -147130
rect 41120 -147180 41760 -147130
rect 42560 -147130 44760 -147080
rect 42560 -147180 44120 -147130
rect 44120 -147180 44760 -147130
rect 45560 -147130 47760 -147080
rect 45560 -147180 47120 -147130
rect 47120 -147180 47760 -147130
rect 48560 -147130 50760 -147080
rect 48560 -147180 50120 -147130
rect 50120 -147180 50760 -147130
rect 51560 -147130 53760 -147080
rect 51560 -147180 53120 -147130
rect 53120 -147180 53760 -147130
rect 54560 -147130 56760 -147080
rect 54560 -147180 56120 -147130
rect 56120 -147180 56760 -147130
rect 57560 -147130 59760 -147080
rect 57560 -147180 59120 -147130
rect 59120 -147180 59760 -147130
rect 60560 -147130 62760 -147080
rect 60560 -147180 62120 -147130
rect 62120 -147180 62760 -147130
rect 63560 -147130 65760 -147080
rect 63560 -147180 65120 -147130
rect 65120 -147180 65760 -147130
rect 66560 -147130 68760 -147080
rect 66560 -147180 68120 -147130
rect 68120 -147180 68760 -147130
rect 69560 -147130 71760 -147080
rect 69560 -147180 71120 -147130
rect 71120 -147180 71760 -147130
rect 72560 -147130 74760 -147080
rect 72560 -147180 74120 -147130
rect 74120 -147180 74760 -147130
rect 75560 -147130 77760 -147080
rect 75560 -147180 77120 -147130
rect 77120 -147180 77760 -147130
rect 78560 -147130 80760 -147080
rect 78560 -147180 80120 -147130
rect 80120 -147180 80760 -147130
rect 81560 -147130 83760 -147080
rect 81560 -147180 83120 -147130
rect 83120 -147180 83760 -147130
rect 84560 -147130 86760 -147080
rect 84560 -147180 86120 -147130
rect 86120 -147180 86760 -147130
rect 87560 -147130 89760 -147080
rect 87560 -147180 89120 -147130
rect 89120 -147180 89760 -147130
rect 90560 -147130 92760 -147080
rect 90560 -147180 92120 -147130
rect 92120 -147180 92760 -147130
rect 93560 -147130 95760 -147080
rect 93560 -147180 95120 -147130
rect 95120 -147180 95760 -147130
rect 96560 -147130 98760 -147080
rect 96560 -147180 98120 -147130
rect 98120 -147180 98760 -147130
rect 99560 -147130 101760 -147080
rect 99560 -147180 101120 -147130
rect 101120 -147180 101760 -147130
rect 102560 -147130 104760 -147080
rect 102560 -147180 104120 -147130
rect 104120 -147180 104760 -147130
rect 105560 -147130 107760 -147080
rect 105560 -147180 107120 -147130
rect 107120 -147180 107760 -147130
rect 108560 -147130 110760 -147080
rect 108560 -147180 110120 -147130
rect 110120 -147180 110760 -147130
rect 111560 -147130 113760 -147080
rect 111560 -147180 113120 -147130
rect 113120 -147180 113760 -147130
rect 114560 -147130 116760 -147080
rect 114560 -147180 116120 -147130
rect 116120 -147180 116760 -147130
rect 117560 -147130 119760 -147080
rect 117560 -147180 119120 -147130
rect 119120 -147180 119760 -147130
rect 120560 -147130 122760 -147080
rect 120560 -147180 122120 -147130
rect 122120 -147180 122760 -147130
rect 123560 -147130 125760 -147080
rect 123560 -147180 125120 -147130
rect 125120 -147180 125760 -147130
rect 126560 -147130 128760 -147080
rect 126560 -147180 128120 -147130
rect 128120 -147180 128760 -147130
rect 129560 -147130 131760 -147080
rect 129560 -147180 131120 -147130
rect 131120 -147180 131760 -147130
rect 132560 -147130 134760 -147080
rect 132560 -147180 134120 -147130
rect 134120 -147180 134760 -147130
rect 135560 -147130 137760 -147080
rect 135560 -147180 137120 -147130
rect 137120 -147180 137760 -147130
rect 138560 -147130 140760 -147080
rect 138560 -147180 140120 -147130
rect 140120 -147180 140760 -147130
rect 141560 -147130 143760 -147080
rect 141560 -147180 143120 -147130
rect 143120 -147180 143760 -147130
rect 144560 -147130 146760 -147080
rect 144560 -147180 146120 -147130
rect 146120 -147180 146760 -147130
rect 147560 -147130 149760 -147080
rect 147560 -147180 149120 -147130
rect 149120 -147180 149760 -147130
rect 240 -147700 420 -147500
rect 3240 -147700 3420 -147500
rect 6240 -147700 6420 -147500
rect 9240 -147700 9420 -147500
rect 12240 -147700 12420 -147500
rect 15240 -147700 15420 -147500
rect 18240 -147700 18420 -147500
rect 21240 -147700 21420 -147500
rect 24240 -147700 24420 -147500
rect 27240 -147700 27420 -147500
rect 30240 -147700 30420 -147500
rect 33240 -147700 33420 -147500
rect 36240 -147700 36420 -147500
rect 39240 -147700 39420 -147500
rect 42240 -147700 42420 -147500
rect 45240 -147700 45420 -147500
rect 48240 -147700 48420 -147500
rect 51240 -147700 51420 -147500
rect 54240 -147700 54420 -147500
rect 57240 -147700 57420 -147500
rect 60240 -147700 60420 -147500
rect 63240 -147700 63420 -147500
rect 66240 -147700 66420 -147500
rect 69240 -147700 69420 -147500
rect 72240 -147700 72420 -147500
rect 75240 -147700 75420 -147500
rect 78240 -147700 78420 -147500
rect 81240 -147700 81420 -147500
rect 84240 -147700 84420 -147500
rect 87240 -147700 87420 -147500
rect 90240 -147700 90420 -147500
rect 93240 -147700 93420 -147500
rect 96240 -147700 96420 -147500
rect 99240 -147700 99420 -147500
rect 102240 -147700 102420 -147500
rect 105240 -147700 105420 -147500
rect 108240 -147700 108420 -147500
rect 111240 -147700 111420 -147500
rect 114240 -147700 114420 -147500
rect 117240 -147700 117420 -147500
rect 120240 -147700 120420 -147500
rect 123240 -147700 123420 -147500
rect 126240 -147700 126420 -147500
rect 129240 -147700 129420 -147500
rect 132240 -147700 132420 -147500
rect 135240 -147700 135420 -147500
rect 138240 -147700 138420 -147500
rect 141240 -147700 141420 -147500
rect 144240 -147700 144420 -147500
rect 147240 -147700 147420 -147500
<< metal3 >>
rect -1200 2840 -1110 5000
rect 480 3650 590 3660
rect 480 3560 490 3650
rect 580 3560 590 3650
rect 480 3550 590 3560
rect 3480 3650 3590 3660
rect 3480 3560 3490 3650
rect 3580 3560 3590 3650
rect 3480 3550 3590 3560
rect 6480 3650 6590 3660
rect 6480 3560 6490 3650
rect 6580 3560 6590 3650
rect 6480 3550 6590 3560
rect 9480 3650 9590 3660
rect 9480 3560 9490 3650
rect 9580 3560 9590 3650
rect 9480 3550 9590 3560
rect 12480 3650 12590 3660
rect 12480 3560 12490 3650
rect 12580 3560 12590 3650
rect 12480 3550 12590 3560
rect 15480 3650 15590 3660
rect 15480 3560 15490 3650
rect 15580 3560 15590 3650
rect 15480 3550 15590 3560
rect 18480 3650 18590 3660
rect 18480 3560 18490 3650
rect 18580 3560 18590 3650
rect 18480 3550 18590 3560
rect 21480 3650 21590 3660
rect 21480 3560 21490 3650
rect 21580 3560 21590 3650
rect 21480 3550 21590 3560
rect 24480 3650 24590 3660
rect 24480 3560 24490 3650
rect 24580 3560 24590 3650
rect 24480 3550 24590 3560
rect 27480 3650 27590 3660
rect 27480 3560 27490 3650
rect 27580 3560 27590 3650
rect 27480 3550 27590 3560
rect 30480 3650 30590 3660
rect 30480 3560 30490 3650
rect 30580 3560 30590 3650
rect 30480 3550 30590 3560
rect 33480 3650 33590 3660
rect 33480 3560 33490 3650
rect 33580 3560 33590 3650
rect 33480 3550 33590 3560
rect 36480 3650 36590 3660
rect 36480 3560 36490 3650
rect 36580 3560 36590 3650
rect 36480 3550 36590 3560
rect 39480 3650 39590 3660
rect 39480 3560 39490 3650
rect 39580 3560 39590 3650
rect 39480 3550 39590 3560
rect 42480 3650 42590 3660
rect 42480 3560 42490 3650
rect 42580 3560 42590 3650
rect 42480 3550 42590 3560
rect 45480 3650 45590 3660
rect 45480 3560 45490 3650
rect 45580 3560 45590 3650
rect 45480 3550 45590 3560
rect 48480 3650 48590 3660
rect 48480 3560 48490 3650
rect 48580 3560 48590 3650
rect 48480 3550 48590 3560
rect 51480 3650 51590 3660
rect 51480 3560 51490 3650
rect 51580 3560 51590 3650
rect 51480 3550 51590 3560
rect 54480 3650 54590 3660
rect 54480 3560 54490 3650
rect 54580 3560 54590 3650
rect 54480 3550 54590 3560
rect 57480 3650 57590 3660
rect 57480 3560 57490 3650
rect 57580 3560 57590 3650
rect 57480 3550 57590 3560
rect 60480 3650 60590 3660
rect 60480 3560 60490 3650
rect 60580 3560 60590 3650
rect 60480 3550 60590 3560
rect 63480 3650 63590 3660
rect 63480 3560 63490 3650
rect 63580 3560 63590 3650
rect 63480 3550 63590 3560
rect 66480 3650 66590 3660
rect 66480 3560 66490 3650
rect 66580 3560 66590 3650
rect 66480 3550 66590 3560
rect 69480 3650 69590 3660
rect 69480 3560 69490 3650
rect 69580 3560 69590 3650
rect 69480 3550 69590 3560
rect 72480 3650 72590 3660
rect 72480 3560 72490 3650
rect 72580 3560 72590 3650
rect 72480 3550 72590 3560
rect 75480 3650 75590 3660
rect 75480 3560 75490 3650
rect 75580 3560 75590 3650
rect 75480 3550 75590 3560
rect 78480 3650 78590 3660
rect 78480 3560 78490 3650
rect 78580 3560 78590 3650
rect 78480 3550 78590 3560
rect 81480 3650 81590 3660
rect 81480 3560 81490 3650
rect 81580 3560 81590 3650
rect 81480 3550 81590 3560
rect 84480 3650 84590 3660
rect 84480 3560 84490 3650
rect 84580 3560 84590 3650
rect 84480 3550 84590 3560
rect 87480 3650 87590 3660
rect 87480 3560 87490 3650
rect 87580 3560 87590 3650
rect 87480 3550 87590 3560
rect 90480 3650 90590 3660
rect 90480 3560 90490 3650
rect 90580 3560 90590 3650
rect 90480 3550 90590 3560
rect 93480 3650 93590 3660
rect 93480 3560 93490 3650
rect 93580 3560 93590 3650
rect 93480 3550 93590 3560
rect 96480 3650 96590 3660
rect 96480 3560 96490 3650
rect 96580 3560 96590 3650
rect 96480 3550 96590 3560
rect 99480 3650 99590 3660
rect 99480 3560 99490 3650
rect 99580 3560 99590 3650
rect 99480 3550 99590 3560
rect 102480 3650 102590 3660
rect 102480 3560 102490 3650
rect 102580 3560 102590 3650
rect 102480 3550 102590 3560
rect 105480 3650 105590 3660
rect 105480 3560 105490 3650
rect 105580 3560 105590 3650
rect 105480 3550 105590 3560
rect 108480 3650 108590 3660
rect 108480 3560 108490 3650
rect 108580 3560 108590 3650
rect 108480 3550 108590 3560
rect 111480 3650 111590 3660
rect 111480 3560 111490 3650
rect 111580 3560 111590 3650
rect 111480 3550 111590 3560
rect 114480 3650 114590 3660
rect 114480 3560 114490 3650
rect 114580 3560 114590 3650
rect 114480 3550 114590 3560
rect 117480 3650 117590 3660
rect 117480 3560 117490 3650
rect 117580 3560 117590 3650
rect 117480 3550 117590 3560
rect 120480 3650 120590 3660
rect 120480 3560 120490 3650
rect 120580 3560 120590 3650
rect 120480 3550 120590 3560
rect 123480 3650 123590 3660
rect 123480 3560 123490 3650
rect 123580 3560 123590 3650
rect 123480 3550 123590 3560
rect 126480 3650 126590 3660
rect 126480 3560 126490 3650
rect 126580 3560 126590 3650
rect 126480 3550 126590 3560
rect 129480 3650 129590 3660
rect 129480 3560 129490 3650
rect 129580 3560 129590 3650
rect 129480 3550 129590 3560
rect 132480 3650 132590 3660
rect 132480 3560 132490 3650
rect 132580 3560 132590 3650
rect 132480 3550 132590 3560
rect 135480 3650 135590 3660
rect 135480 3560 135490 3650
rect 135580 3560 135590 3650
rect 135480 3550 135590 3560
rect 138480 3650 138590 3660
rect 138480 3560 138490 3650
rect 138580 3560 138590 3650
rect 138480 3550 138590 3560
rect 141480 3650 141590 3660
rect 141480 3560 141490 3650
rect 141580 3560 141590 3650
rect 141480 3550 141590 3560
rect 144480 3650 144590 3660
rect 144480 3560 144490 3650
rect 144580 3560 144590 3650
rect 144480 3550 144590 3560
rect 147480 3650 147590 3660
rect 147480 3560 147490 3650
rect 147580 3560 147590 3650
rect 147480 3550 147590 3560
rect -1200 2750 200 2840
rect -1200 -160 -1110 2750
rect -480 2550 -370 2560
rect -480 2540 520 2550
rect -480 2470 -470 2540
rect -380 2470 520 2540
rect -480 2460 520 2470
rect -480 2450 -370 2460
rect -560 1560 440 1570
rect -560 1490 -540 1560
rect -260 1490 440 1560
rect -560 1480 440 1490
rect -760 230 40 250
rect -760 160 -740 230
rect -650 160 40 230
rect -750 140 -640 160
rect -1200 -250 200 -160
rect -1200 -3160 -1110 -250
rect -480 -450 -370 -440
rect -480 -460 520 -450
rect -480 -530 -470 -460
rect -380 -530 520 -460
rect -480 -540 520 -530
rect -480 -550 -370 -540
rect -560 -1440 440 -1430
rect -560 -1510 -540 -1440
rect -260 -1510 440 -1440
rect -560 -1520 440 -1510
rect -760 -2770 40 -2750
rect -760 -2840 -740 -2770
rect -650 -2840 40 -2770
rect -750 -2860 -640 -2840
rect -1200 -3250 200 -3160
rect -1200 -6160 -1110 -3250
rect -480 -3450 -370 -3440
rect -480 -3460 520 -3450
rect -480 -3530 -470 -3460
rect -380 -3530 520 -3460
rect -480 -3540 520 -3530
rect -480 -3550 -370 -3540
rect -560 -4440 440 -4430
rect -560 -4510 -540 -4440
rect -260 -4510 440 -4440
rect -560 -4520 440 -4510
rect -760 -5770 40 -5750
rect -760 -5840 -740 -5770
rect -650 -5840 40 -5770
rect -750 -5860 -640 -5840
rect -1200 -6250 200 -6160
rect -1200 -9160 -1110 -6250
rect -480 -6450 -370 -6440
rect -480 -6460 520 -6450
rect -480 -6530 -470 -6460
rect -380 -6530 520 -6460
rect -480 -6540 520 -6530
rect -480 -6550 -370 -6540
rect -560 -7440 440 -7430
rect -560 -7510 -540 -7440
rect -260 -7510 440 -7440
rect -560 -7520 440 -7510
rect -760 -8770 40 -8750
rect -760 -8840 -740 -8770
rect -650 -8840 40 -8770
rect -750 -8860 -640 -8840
rect -1200 -9250 200 -9160
rect -1200 -12160 -1110 -9250
rect -480 -9450 -370 -9440
rect -480 -9460 520 -9450
rect -480 -9530 -470 -9460
rect -380 -9530 520 -9460
rect -480 -9540 520 -9530
rect -480 -9550 -370 -9540
rect -560 -10440 440 -10430
rect -560 -10510 -540 -10440
rect -260 -10510 440 -10440
rect -560 -10520 440 -10510
rect -760 -11770 40 -11750
rect -760 -11840 -740 -11770
rect -650 -11840 40 -11770
rect -750 -11860 -640 -11840
rect -1200 -12250 200 -12160
rect -1200 -15160 -1110 -12250
rect -480 -12450 -370 -12440
rect -480 -12460 520 -12450
rect -480 -12530 -470 -12460
rect -380 -12530 520 -12460
rect -480 -12540 520 -12530
rect -480 -12550 -370 -12540
rect -560 -13440 440 -13430
rect -560 -13510 -540 -13440
rect -260 -13510 440 -13440
rect -560 -13520 440 -13510
rect -760 -14770 40 -14750
rect -760 -14840 -740 -14770
rect -650 -14840 40 -14770
rect -750 -14860 -640 -14840
rect -1200 -15250 200 -15160
rect -1200 -18160 -1110 -15250
rect -480 -15450 -370 -15440
rect -480 -15460 520 -15450
rect -480 -15530 -470 -15460
rect -380 -15530 520 -15460
rect -480 -15540 520 -15530
rect -480 -15550 -370 -15540
rect -560 -16440 440 -16430
rect -560 -16510 -540 -16440
rect -260 -16510 440 -16440
rect -560 -16520 440 -16510
rect -760 -17770 40 -17750
rect -760 -17840 -740 -17770
rect -650 -17840 40 -17770
rect -750 -17860 -640 -17840
rect -1200 -18250 200 -18160
rect -1200 -21160 -1110 -18250
rect -480 -18450 -370 -18440
rect -480 -18460 520 -18450
rect -480 -18530 -470 -18460
rect -380 -18530 520 -18460
rect -480 -18540 520 -18530
rect -480 -18550 -370 -18540
rect -560 -19440 440 -19430
rect -560 -19510 -540 -19440
rect -260 -19510 440 -19440
rect -560 -19520 440 -19510
rect -760 -20770 40 -20750
rect -760 -20840 -740 -20770
rect -650 -20840 40 -20770
rect -750 -20860 -640 -20840
rect -1200 -21250 200 -21160
rect -1200 -24160 -1110 -21250
rect -480 -21450 -370 -21440
rect -480 -21460 520 -21450
rect -480 -21530 -470 -21460
rect -380 -21530 520 -21460
rect -480 -21540 520 -21530
rect -480 -21550 -370 -21540
rect -560 -22440 440 -22430
rect -560 -22510 -540 -22440
rect -260 -22510 440 -22440
rect -560 -22520 440 -22510
rect -760 -23770 40 -23750
rect -760 -23840 -740 -23770
rect -650 -23840 40 -23770
rect -750 -23860 -640 -23840
rect -1200 -24250 200 -24160
rect -1200 -27160 -1110 -24250
rect -480 -24450 -370 -24440
rect -480 -24460 520 -24450
rect -480 -24530 -470 -24460
rect -380 -24530 520 -24460
rect -480 -24540 520 -24530
rect -480 -24550 -370 -24540
rect -560 -25440 440 -25430
rect -560 -25510 -540 -25440
rect -260 -25510 440 -25440
rect -560 -25520 440 -25510
rect -760 -26770 40 -26750
rect -760 -26840 -740 -26770
rect -650 -26840 40 -26770
rect -750 -26860 -640 -26840
rect -1200 -27250 200 -27160
rect -1200 -30160 -1110 -27250
rect -480 -27450 -370 -27440
rect -480 -27460 520 -27450
rect -480 -27530 -470 -27460
rect -380 -27530 520 -27460
rect -480 -27540 520 -27530
rect -480 -27550 -370 -27540
rect -560 -28440 440 -28430
rect -560 -28510 -540 -28440
rect -260 -28510 440 -28440
rect -560 -28520 440 -28510
rect -760 -29770 40 -29750
rect -760 -29840 -740 -29770
rect -650 -29840 40 -29770
rect -750 -29860 -640 -29840
rect -1200 -30250 200 -30160
rect -1200 -33160 -1110 -30250
rect -480 -30450 -370 -30440
rect -480 -30460 520 -30450
rect -480 -30530 -470 -30460
rect -380 -30530 520 -30460
rect -480 -30540 520 -30530
rect -480 -30550 -370 -30540
rect -560 -31440 440 -31430
rect -560 -31510 -540 -31440
rect -260 -31510 440 -31440
rect -560 -31520 440 -31510
rect -760 -32770 40 -32750
rect -760 -32840 -740 -32770
rect -650 -32840 40 -32770
rect -750 -32860 -640 -32840
rect -1200 -33250 200 -33160
rect -1200 -36160 -1110 -33250
rect -480 -33450 -370 -33440
rect -480 -33460 520 -33450
rect -480 -33530 -470 -33460
rect -380 -33530 520 -33460
rect -480 -33540 520 -33530
rect -480 -33550 -370 -33540
rect -560 -34440 440 -34430
rect -560 -34510 -540 -34440
rect -260 -34510 440 -34440
rect -560 -34520 440 -34510
rect -760 -35770 40 -35750
rect -760 -35840 -740 -35770
rect -650 -35840 40 -35770
rect -750 -35860 -640 -35840
rect -1200 -36250 200 -36160
rect -1200 -39160 -1110 -36250
rect -480 -36450 -370 -36440
rect -480 -36460 520 -36450
rect -480 -36530 -470 -36460
rect -380 -36530 520 -36460
rect -480 -36540 520 -36530
rect -480 -36550 -370 -36540
rect -560 -37440 440 -37430
rect -560 -37510 -540 -37440
rect -260 -37510 440 -37440
rect -560 -37520 440 -37510
rect -760 -38770 40 -38750
rect -760 -38840 -740 -38770
rect -650 -38840 40 -38770
rect -750 -38860 -640 -38840
rect -1200 -39250 200 -39160
rect -1200 -42160 -1110 -39250
rect -480 -39450 -370 -39440
rect -480 -39460 520 -39450
rect -480 -39530 -470 -39460
rect -380 -39530 520 -39460
rect -480 -39540 520 -39530
rect -480 -39550 -370 -39540
rect -560 -40440 440 -40430
rect -560 -40510 -540 -40440
rect -260 -40510 440 -40440
rect -560 -40520 440 -40510
rect -760 -41770 40 -41750
rect -760 -41840 -740 -41770
rect -650 -41840 40 -41770
rect -750 -41860 -640 -41840
rect -1200 -42250 200 -42160
rect -1200 -45160 -1110 -42250
rect -480 -42450 -370 -42440
rect -480 -42460 520 -42450
rect -480 -42530 -470 -42460
rect -380 -42530 520 -42460
rect -480 -42540 520 -42530
rect -480 -42550 -370 -42540
rect -560 -43440 440 -43430
rect -560 -43510 -540 -43440
rect -260 -43510 440 -43440
rect -560 -43520 440 -43510
rect -760 -44770 40 -44750
rect -760 -44840 -740 -44770
rect -650 -44840 40 -44770
rect -750 -44860 -640 -44840
rect -1200 -45250 200 -45160
rect -1200 -48160 -1110 -45250
rect -480 -45450 -370 -45440
rect -480 -45460 520 -45450
rect -480 -45530 -470 -45460
rect -380 -45530 520 -45460
rect -480 -45540 520 -45530
rect -480 -45550 -370 -45540
rect -560 -46440 440 -46430
rect -560 -46510 -540 -46440
rect -260 -46510 440 -46440
rect -560 -46520 440 -46510
rect -760 -47770 40 -47750
rect -760 -47840 -740 -47770
rect -650 -47840 40 -47770
rect -750 -47860 -640 -47840
rect -1200 -48250 200 -48160
rect -1200 -51160 -1110 -48250
rect -480 -48450 -370 -48440
rect -480 -48460 520 -48450
rect -480 -48530 -470 -48460
rect -380 -48530 520 -48460
rect -480 -48540 520 -48530
rect -480 -48550 -370 -48540
rect -560 -49440 440 -49430
rect -560 -49510 -540 -49440
rect -260 -49510 440 -49440
rect -560 -49520 440 -49510
rect -760 -50770 40 -50750
rect -760 -50840 -740 -50770
rect -650 -50840 40 -50770
rect -750 -50860 -640 -50840
rect -1200 -51250 200 -51160
rect -1200 -54160 -1110 -51250
rect -480 -51450 -370 -51440
rect -480 -51460 520 -51450
rect -480 -51530 -470 -51460
rect -380 -51530 520 -51460
rect -480 -51540 520 -51530
rect -480 -51550 -370 -51540
rect -560 -52440 440 -52430
rect -560 -52510 -540 -52440
rect -260 -52510 440 -52440
rect -560 -52520 440 -52510
rect -760 -53770 40 -53750
rect -760 -53840 -740 -53770
rect -650 -53840 40 -53770
rect -750 -53860 -640 -53840
rect -1200 -54250 200 -54160
rect -1200 -57160 -1110 -54250
rect -480 -54450 -370 -54440
rect -480 -54460 520 -54450
rect -480 -54530 -470 -54460
rect -380 -54530 520 -54460
rect -480 -54540 520 -54530
rect -480 -54550 -370 -54540
rect -560 -55440 440 -55430
rect -560 -55510 -540 -55440
rect -260 -55510 440 -55440
rect -560 -55520 440 -55510
rect -760 -56770 40 -56750
rect -760 -56840 -740 -56770
rect -650 -56840 40 -56770
rect -750 -56860 -640 -56840
rect -1200 -57250 200 -57160
rect -1200 -60160 -1110 -57250
rect -480 -57450 -370 -57440
rect -480 -57460 520 -57450
rect -480 -57530 -470 -57460
rect -380 -57530 520 -57460
rect -480 -57540 520 -57530
rect -480 -57550 -370 -57540
rect -560 -58440 440 -58430
rect -560 -58510 -540 -58440
rect -260 -58510 440 -58440
rect -560 -58520 440 -58510
rect -760 -59770 40 -59750
rect -760 -59840 -740 -59770
rect -650 -59840 40 -59770
rect -750 -59860 -640 -59840
rect -1200 -60250 200 -60160
rect -1200 -63160 -1110 -60250
rect -480 -60450 -370 -60440
rect -480 -60460 520 -60450
rect -480 -60530 -470 -60460
rect -380 -60530 520 -60460
rect -480 -60540 520 -60530
rect -480 -60550 -370 -60540
rect -560 -61440 440 -61430
rect -560 -61510 -540 -61440
rect -260 -61510 440 -61440
rect -560 -61520 440 -61510
rect -760 -62770 40 -62750
rect -760 -62840 -740 -62770
rect -650 -62840 40 -62770
rect -750 -62860 -640 -62840
rect -1200 -63250 200 -63160
rect -1200 -66160 -1110 -63250
rect -480 -63450 -370 -63440
rect -480 -63460 520 -63450
rect -480 -63530 -470 -63460
rect -380 -63530 520 -63460
rect -480 -63540 520 -63530
rect -480 -63550 -370 -63540
rect -560 -64440 440 -64430
rect -560 -64510 -540 -64440
rect -260 -64510 440 -64440
rect -560 -64520 440 -64510
rect -760 -65770 40 -65750
rect -760 -65840 -740 -65770
rect -650 -65840 40 -65770
rect -750 -65860 -640 -65840
rect -1200 -66250 200 -66160
rect -1200 -69160 -1110 -66250
rect -480 -66450 -370 -66440
rect -480 -66460 520 -66450
rect -480 -66530 -470 -66460
rect -380 -66530 520 -66460
rect -480 -66540 520 -66530
rect -480 -66550 -370 -66540
rect -560 -67440 440 -67430
rect -560 -67510 -540 -67440
rect -260 -67510 440 -67440
rect -560 -67520 440 -67510
rect -760 -68770 40 -68750
rect -760 -68840 -740 -68770
rect -650 -68840 40 -68770
rect -750 -68860 -640 -68840
rect -1200 -69250 200 -69160
rect -1200 -72160 -1110 -69250
rect -480 -69450 -370 -69440
rect -480 -69460 520 -69450
rect -480 -69530 -470 -69460
rect -380 -69530 520 -69460
rect -480 -69540 520 -69530
rect -480 -69550 -370 -69540
rect -560 -70440 440 -70430
rect -560 -70510 -540 -70440
rect -260 -70510 440 -70440
rect -560 -70520 440 -70510
rect -760 -71770 40 -71750
rect -760 -71840 -740 -71770
rect -650 -71840 40 -71770
rect -750 -71860 -640 -71840
rect -1200 -72250 200 -72160
rect -1200 -75160 -1110 -72250
rect -480 -72450 -370 -72440
rect -480 -72460 520 -72450
rect -480 -72530 -470 -72460
rect -380 -72530 520 -72460
rect -480 -72540 520 -72530
rect -480 -72550 -370 -72540
rect -560 -73440 440 -73430
rect -560 -73510 -540 -73440
rect -260 -73510 440 -73440
rect -560 -73520 440 -73510
rect -760 -74770 40 -74750
rect -760 -74840 -740 -74770
rect -650 -74840 40 -74770
rect -750 -74860 -640 -74840
rect -1200 -75250 200 -75160
rect -1200 -78160 -1110 -75250
rect -480 -75450 -370 -75440
rect -480 -75460 520 -75450
rect -480 -75530 -470 -75460
rect -380 -75530 520 -75460
rect -480 -75540 520 -75530
rect -480 -75550 -370 -75540
rect -560 -76440 440 -76430
rect -560 -76510 -540 -76440
rect -260 -76510 440 -76440
rect -560 -76520 440 -76510
rect -760 -77770 40 -77750
rect -760 -77840 -740 -77770
rect -650 -77840 40 -77770
rect -750 -77860 -640 -77840
rect -1200 -78250 200 -78160
rect -1200 -81160 -1110 -78250
rect -480 -78450 -370 -78440
rect -480 -78460 520 -78450
rect -480 -78530 -470 -78460
rect -380 -78530 520 -78460
rect -480 -78540 520 -78530
rect -480 -78550 -370 -78540
rect -560 -79440 440 -79430
rect -560 -79510 -540 -79440
rect -260 -79510 440 -79440
rect -560 -79520 440 -79510
rect -760 -80770 40 -80750
rect -760 -80840 -740 -80770
rect -650 -80840 40 -80770
rect -750 -80860 -640 -80840
rect -1200 -81250 200 -81160
rect -1200 -84160 -1110 -81250
rect -480 -81450 -370 -81440
rect -480 -81460 520 -81450
rect -480 -81530 -470 -81460
rect -380 -81530 520 -81460
rect -480 -81540 520 -81530
rect -480 -81550 -370 -81540
rect -560 -82440 440 -82430
rect -560 -82510 -540 -82440
rect -260 -82510 440 -82440
rect -560 -82520 440 -82510
rect -760 -83770 40 -83750
rect -760 -83840 -740 -83770
rect -650 -83840 40 -83770
rect -750 -83860 -640 -83840
rect -1200 -84250 200 -84160
rect -1200 -87160 -1110 -84250
rect -480 -84450 -370 -84440
rect -480 -84460 520 -84450
rect -480 -84530 -470 -84460
rect -380 -84530 520 -84460
rect -480 -84540 520 -84530
rect -480 -84550 -370 -84540
rect -560 -85440 440 -85430
rect -560 -85510 -540 -85440
rect -260 -85510 440 -85440
rect -560 -85520 440 -85510
rect -760 -86770 40 -86750
rect -760 -86840 -740 -86770
rect -650 -86840 40 -86770
rect -750 -86860 -640 -86840
rect -1200 -87250 200 -87160
rect -1200 -90160 -1110 -87250
rect -480 -87450 -370 -87440
rect -480 -87460 520 -87450
rect -480 -87530 -470 -87460
rect -380 -87530 520 -87460
rect -480 -87540 520 -87530
rect -480 -87550 -370 -87540
rect -560 -88440 440 -88430
rect -560 -88510 -540 -88440
rect -260 -88510 440 -88440
rect -560 -88520 440 -88510
rect -760 -89770 40 -89750
rect -760 -89840 -740 -89770
rect -650 -89840 40 -89770
rect -750 -89860 -640 -89840
rect -1200 -90250 200 -90160
rect -1200 -93160 -1110 -90250
rect -480 -90450 -370 -90440
rect -480 -90460 520 -90450
rect -480 -90530 -470 -90460
rect -380 -90530 520 -90460
rect -480 -90540 520 -90530
rect -480 -90550 -370 -90540
rect -560 -91440 440 -91430
rect -560 -91510 -540 -91440
rect -260 -91510 440 -91440
rect -560 -91520 440 -91510
rect -760 -92770 40 -92750
rect -760 -92840 -740 -92770
rect -650 -92840 40 -92770
rect -750 -92860 -640 -92840
rect -1200 -93250 200 -93160
rect -1200 -96160 -1110 -93250
rect -480 -93450 -370 -93440
rect -480 -93460 520 -93450
rect -480 -93530 -470 -93460
rect -380 -93530 520 -93460
rect -480 -93540 520 -93530
rect -480 -93550 -370 -93540
rect -560 -94440 440 -94430
rect -560 -94510 -540 -94440
rect -260 -94510 440 -94440
rect -560 -94520 440 -94510
rect -760 -95770 40 -95750
rect -760 -95840 -740 -95770
rect -650 -95840 40 -95770
rect -750 -95860 -640 -95840
rect -1200 -96250 200 -96160
rect -1200 -99160 -1110 -96250
rect -480 -96450 -370 -96440
rect -480 -96460 520 -96450
rect -480 -96530 -470 -96460
rect -380 -96530 520 -96460
rect -480 -96540 520 -96530
rect -480 -96550 -370 -96540
rect -560 -97440 440 -97430
rect -560 -97510 -540 -97440
rect -260 -97510 440 -97440
rect -560 -97520 440 -97510
rect -760 -98770 40 -98750
rect -760 -98840 -740 -98770
rect -650 -98840 40 -98770
rect -750 -98860 -640 -98840
rect -1200 -99250 200 -99160
rect -1200 -102160 -1110 -99250
rect -480 -99450 -370 -99440
rect -480 -99460 520 -99450
rect -480 -99530 -470 -99460
rect -380 -99530 520 -99460
rect -480 -99540 520 -99530
rect -480 -99550 -370 -99540
rect -560 -100440 440 -100430
rect -560 -100510 -540 -100440
rect -260 -100510 440 -100440
rect -560 -100520 440 -100510
rect -760 -101770 40 -101750
rect -760 -101840 -740 -101770
rect -650 -101840 40 -101770
rect -750 -101860 -640 -101840
rect -1200 -102250 200 -102160
rect -1200 -105160 -1110 -102250
rect -480 -102450 -370 -102440
rect -480 -102460 520 -102450
rect -480 -102530 -470 -102460
rect -380 -102530 520 -102460
rect -480 -102540 520 -102530
rect -480 -102550 -370 -102540
rect -560 -103440 440 -103430
rect -560 -103510 -540 -103440
rect -260 -103510 440 -103440
rect -560 -103520 440 -103510
rect -760 -104770 40 -104750
rect -760 -104840 -740 -104770
rect -650 -104840 40 -104770
rect -750 -104860 -640 -104840
rect -1200 -105250 200 -105160
rect -1200 -108160 -1110 -105250
rect -480 -105450 -370 -105440
rect -480 -105460 520 -105450
rect -480 -105530 -470 -105460
rect -380 -105530 520 -105460
rect -480 -105540 520 -105530
rect -480 -105550 -370 -105540
rect -560 -106440 440 -106430
rect -560 -106510 -540 -106440
rect -260 -106510 440 -106440
rect -560 -106520 440 -106510
rect -760 -107770 40 -107750
rect -760 -107840 -740 -107770
rect -650 -107840 40 -107770
rect -750 -107860 -640 -107840
rect -1200 -108250 200 -108160
rect -1200 -111160 -1110 -108250
rect -480 -108450 -370 -108440
rect -480 -108460 520 -108450
rect -480 -108530 -470 -108460
rect -380 -108530 520 -108460
rect -480 -108540 520 -108530
rect -480 -108550 -370 -108540
rect -560 -109440 440 -109430
rect -560 -109510 -540 -109440
rect -260 -109510 440 -109440
rect -560 -109520 440 -109510
rect -760 -110770 40 -110750
rect -760 -110840 -740 -110770
rect -650 -110840 40 -110770
rect -750 -110860 -640 -110840
rect -1200 -111250 200 -111160
rect -1200 -114160 -1110 -111250
rect -480 -111450 -370 -111440
rect -480 -111460 520 -111450
rect -480 -111530 -470 -111460
rect -380 -111530 520 -111460
rect -480 -111540 520 -111530
rect -480 -111550 -370 -111540
rect -560 -112440 440 -112430
rect -560 -112510 -540 -112440
rect -260 -112510 440 -112440
rect -560 -112520 440 -112510
rect -760 -113770 40 -113750
rect -760 -113840 -740 -113770
rect -650 -113840 40 -113770
rect -750 -113860 -640 -113840
rect -1200 -114250 200 -114160
rect -1200 -117160 -1110 -114250
rect -480 -114450 -370 -114440
rect -480 -114460 520 -114450
rect -480 -114530 -470 -114460
rect -380 -114530 520 -114460
rect -480 -114540 520 -114530
rect -480 -114550 -370 -114540
rect -560 -115440 440 -115430
rect -560 -115510 -540 -115440
rect -260 -115510 440 -115440
rect -560 -115520 440 -115510
rect -760 -116770 40 -116750
rect -760 -116840 -740 -116770
rect -650 -116840 40 -116770
rect -750 -116860 -640 -116840
rect -1200 -117250 200 -117160
rect -1200 -120160 -1110 -117250
rect -480 -117450 -370 -117440
rect -480 -117460 520 -117450
rect -480 -117530 -470 -117460
rect -380 -117530 520 -117460
rect -480 -117540 520 -117530
rect -480 -117550 -370 -117540
rect -560 -118440 440 -118430
rect -560 -118510 -540 -118440
rect -260 -118510 440 -118440
rect -560 -118520 440 -118510
rect -760 -119770 40 -119750
rect -760 -119840 -740 -119770
rect -650 -119840 40 -119770
rect -750 -119860 -640 -119840
rect -1200 -120250 200 -120160
rect -1200 -123160 -1110 -120250
rect -480 -120450 -370 -120440
rect -480 -120460 520 -120450
rect -480 -120530 -470 -120460
rect -380 -120530 520 -120460
rect -480 -120540 520 -120530
rect -480 -120550 -370 -120540
rect -560 -121440 440 -121430
rect -560 -121510 -540 -121440
rect -260 -121510 440 -121440
rect -560 -121520 440 -121510
rect -760 -122770 40 -122750
rect -760 -122840 -740 -122770
rect -650 -122840 40 -122770
rect -750 -122860 -640 -122840
rect -1200 -123250 200 -123160
rect -1200 -126160 -1110 -123250
rect -480 -123450 -370 -123440
rect -480 -123460 520 -123450
rect -480 -123530 -470 -123460
rect -380 -123530 520 -123460
rect -480 -123540 520 -123530
rect -480 -123550 -370 -123540
rect -560 -124440 440 -124430
rect -560 -124510 -540 -124440
rect -260 -124510 440 -124440
rect -560 -124520 440 -124510
rect -760 -125770 40 -125750
rect -760 -125840 -740 -125770
rect -650 -125840 40 -125770
rect -750 -125860 -640 -125840
rect -1200 -126250 200 -126160
rect -1200 -129160 -1110 -126250
rect -480 -126450 -370 -126440
rect -480 -126460 520 -126450
rect -480 -126530 -470 -126460
rect -380 -126530 520 -126460
rect -480 -126540 520 -126530
rect -480 -126550 -370 -126540
rect -560 -127440 440 -127430
rect -560 -127510 -540 -127440
rect -260 -127510 440 -127440
rect -560 -127520 440 -127510
rect -760 -128770 40 -128750
rect -760 -128840 -740 -128770
rect -650 -128840 40 -128770
rect -750 -128860 -640 -128840
rect -1200 -129250 200 -129160
rect -1200 -132160 -1110 -129250
rect -480 -129450 -370 -129440
rect -480 -129460 520 -129450
rect -480 -129530 -470 -129460
rect -380 -129530 520 -129460
rect -480 -129540 520 -129530
rect -480 -129550 -370 -129540
rect -560 -130440 440 -130430
rect -560 -130510 -540 -130440
rect -260 -130510 440 -130440
rect -560 -130520 440 -130510
rect -760 -131770 40 -131750
rect -760 -131840 -740 -131770
rect -650 -131840 40 -131770
rect -750 -131860 -640 -131840
rect -1200 -132250 200 -132160
rect -1200 -135160 -1110 -132250
rect -480 -132450 -370 -132440
rect -480 -132460 520 -132450
rect -480 -132530 -470 -132460
rect -380 -132530 520 -132460
rect -480 -132540 520 -132530
rect -480 -132550 -370 -132540
rect -560 -133440 440 -133430
rect -560 -133510 -540 -133440
rect -260 -133510 440 -133440
rect -560 -133520 440 -133510
rect -760 -134770 40 -134750
rect -760 -134840 -740 -134770
rect -650 -134840 40 -134770
rect -750 -134860 -640 -134840
rect -1200 -135250 200 -135160
rect -1200 -138160 -1110 -135250
rect -480 -135450 -370 -135440
rect -480 -135460 520 -135450
rect -480 -135530 -470 -135460
rect -380 -135530 520 -135460
rect -480 -135540 520 -135530
rect -480 -135550 -370 -135540
rect -560 -136440 440 -136430
rect -560 -136510 -540 -136440
rect -260 -136510 440 -136440
rect -560 -136520 440 -136510
rect -760 -137770 40 -137750
rect -760 -137840 -740 -137770
rect -650 -137840 40 -137770
rect -750 -137860 -640 -137840
rect -1200 -138250 200 -138160
rect -1200 -141160 -1110 -138250
rect -480 -138450 -370 -138440
rect -480 -138460 520 -138450
rect -480 -138530 -470 -138460
rect -380 -138530 520 -138460
rect -480 -138540 520 -138530
rect -480 -138550 -370 -138540
rect -560 -139440 440 -139430
rect -560 -139510 -540 -139440
rect -260 -139510 440 -139440
rect -560 -139520 440 -139510
rect -760 -140770 40 -140750
rect -760 -140840 -740 -140770
rect -650 -140840 40 -140770
rect -750 -140860 -640 -140840
rect -1200 -141250 200 -141160
rect -1200 -144160 -1110 -141250
rect -480 -141450 -370 -141440
rect -480 -141460 520 -141450
rect -480 -141530 -470 -141460
rect -380 -141530 520 -141460
rect -480 -141540 520 -141530
rect -480 -141550 -370 -141540
rect -560 -142440 440 -142430
rect -560 -142510 -540 -142440
rect -260 -142510 440 -142440
rect -560 -142520 440 -142510
rect -760 -143770 40 -143750
rect -760 -143840 -740 -143770
rect -650 -143840 40 -143770
rect -750 -143860 -640 -143840
rect -1200 -144250 200 -144160
rect -1200 -145000 -1110 -144250
rect -480 -144450 -370 -144440
rect -480 -144460 520 -144450
rect -480 -144530 -470 -144460
rect -380 -144530 520 -144460
rect -480 -144540 520 -144530
rect -480 -144550 -370 -144540
rect -560 -145440 440 -145430
rect -560 -145510 -540 -145440
rect -260 -145510 440 -145440
rect -560 -145520 440 -145510
rect -760 -146770 40 -146750
rect -760 -146840 -740 -146770
rect -650 -146840 40 -146770
rect -750 -146860 -640 -146840
rect 540 -147080 2780 -147060
rect 540 -147180 560 -147080
rect 2760 -147180 2780 -147080
rect 540 -147200 2780 -147180
rect 3540 -147080 5780 -147060
rect 3540 -147180 3560 -147080
rect 5760 -147180 5780 -147080
rect 3540 -147200 5780 -147180
rect 6540 -147080 8780 -147060
rect 6540 -147180 6560 -147080
rect 8760 -147180 8780 -147080
rect 6540 -147200 8780 -147180
rect 9540 -147080 11780 -147060
rect 9540 -147180 9560 -147080
rect 11760 -147180 11780 -147080
rect 9540 -147200 11780 -147180
rect 12540 -147080 14780 -147060
rect 12540 -147180 12560 -147080
rect 14760 -147180 14780 -147080
rect 12540 -147200 14780 -147180
rect 15540 -147080 17780 -147060
rect 15540 -147180 15560 -147080
rect 17760 -147180 17780 -147080
rect 15540 -147200 17780 -147180
rect 18540 -147080 20780 -147060
rect 18540 -147180 18560 -147080
rect 20760 -147180 20780 -147080
rect 18540 -147200 20780 -147180
rect 21540 -147080 23780 -147060
rect 21540 -147180 21560 -147080
rect 23760 -147180 23780 -147080
rect 21540 -147200 23780 -147180
rect 24540 -147080 26780 -147060
rect 24540 -147180 24560 -147080
rect 26760 -147180 26780 -147080
rect 24540 -147200 26780 -147180
rect 27540 -147080 29780 -147060
rect 27540 -147180 27560 -147080
rect 29760 -147180 29780 -147080
rect 27540 -147200 29780 -147180
rect 30540 -147080 32780 -147060
rect 30540 -147180 30560 -147080
rect 32760 -147180 32780 -147080
rect 30540 -147200 32780 -147180
rect 33540 -147080 35780 -147060
rect 33540 -147180 33560 -147080
rect 35760 -147180 35780 -147080
rect 33540 -147200 35780 -147180
rect 36540 -147080 38780 -147060
rect 36540 -147180 36560 -147080
rect 38760 -147180 38780 -147080
rect 36540 -147200 38780 -147180
rect 39540 -147080 41780 -147060
rect 39540 -147180 39560 -147080
rect 41760 -147180 41780 -147080
rect 39540 -147200 41780 -147180
rect 42540 -147080 44780 -147060
rect 42540 -147180 42560 -147080
rect 44760 -147180 44780 -147080
rect 42540 -147200 44780 -147180
rect 45540 -147080 47780 -147060
rect 45540 -147180 45560 -147080
rect 47760 -147180 47780 -147080
rect 45540 -147200 47780 -147180
rect 48540 -147080 50780 -147060
rect 48540 -147180 48560 -147080
rect 50760 -147180 50780 -147080
rect 48540 -147200 50780 -147180
rect 51540 -147080 53780 -147060
rect 51540 -147180 51560 -147080
rect 53760 -147180 53780 -147080
rect 51540 -147200 53780 -147180
rect 54540 -147080 56780 -147060
rect 54540 -147180 54560 -147080
rect 56760 -147180 56780 -147080
rect 54540 -147200 56780 -147180
rect 57540 -147080 59780 -147060
rect 57540 -147180 57560 -147080
rect 59760 -147180 59780 -147080
rect 57540 -147200 59780 -147180
rect 60540 -147080 62780 -147060
rect 60540 -147180 60560 -147080
rect 62760 -147180 62780 -147080
rect 60540 -147200 62780 -147180
rect 63540 -147080 65780 -147060
rect 63540 -147180 63560 -147080
rect 65760 -147180 65780 -147080
rect 63540 -147200 65780 -147180
rect 66540 -147080 68780 -147060
rect 66540 -147180 66560 -147080
rect 68760 -147180 68780 -147080
rect 66540 -147200 68780 -147180
rect 69540 -147080 71780 -147060
rect 69540 -147180 69560 -147080
rect 71760 -147180 71780 -147080
rect 69540 -147200 71780 -147180
rect 72540 -147080 74780 -147060
rect 72540 -147180 72560 -147080
rect 74760 -147180 74780 -147080
rect 72540 -147200 74780 -147180
rect 75540 -147080 77780 -147060
rect 75540 -147180 75560 -147080
rect 77760 -147180 77780 -147080
rect 75540 -147200 77780 -147180
rect 78540 -147080 80780 -147060
rect 78540 -147180 78560 -147080
rect 80760 -147180 80780 -147080
rect 78540 -147200 80780 -147180
rect 81540 -147080 83780 -147060
rect 81540 -147180 81560 -147080
rect 83760 -147180 83780 -147080
rect 81540 -147200 83780 -147180
rect 84540 -147080 86780 -147060
rect 84540 -147180 84560 -147080
rect 86760 -147180 86780 -147080
rect 84540 -147200 86780 -147180
rect 87540 -147080 89780 -147060
rect 87540 -147180 87560 -147080
rect 89760 -147180 89780 -147080
rect 87540 -147200 89780 -147180
rect 90540 -147080 92780 -147060
rect 90540 -147180 90560 -147080
rect 92760 -147180 92780 -147080
rect 90540 -147200 92780 -147180
rect 93540 -147080 95780 -147060
rect 93540 -147180 93560 -147080
rect 95760 -147180 95780 -147080
rect 93540 -147200 95780 -147180
rect 96540 -147080 98780 -147060
rect 96540 -147180 96560 -147080
rect 98760 -147180 98780 -147080
rect 96540 -147200 98780 -147180
rect 99540 -147080 101780 -147060
rect 99540 -147180 99560 -147080
rect 101760 -147180 101780 -147080
rect 99540 -147200 101780 -147180
rect 102540 -147080 104780 -147060
rect 102540 -147180 102560 -147080
rect 104760 -147180 104780 -147080
rect 102540 -147200 104780 -147180
rect 105540 -147080 107780 -147060
rect 105540 -147180 105560 -147080
rect 107760 -147180 107780 -147080
rect 105540 -147200 107780 -147180
rect 108540 -147080 110780 -147060
rect 108540 -147180 108560 -147080
rect 110760 -147180 110780 -147080
rect 108540 -147200 110780 -147180
rect 111540 -147080 113780 -147060
rect 111540 -147180 111560 -147080
rect 113760 -147180 113780 -147080
rect 111540 -147200 113780 -147180
rect 114540 -147080 116780 -147060
rect 114540 -147180 114560 -147080
rect 116760 -147180 116780 -147080
rect 114540 -147200 116780 -147180
rect 117540 -147080 119780 -147060
rect 117540 -147180 117560 -147080
rect 119760 -147180 119780 -147080
rect 117540 -147200 119780 -147180
rect 120540 -147080 122780 -147060
rect 120540 -147180 120560 -147080
rect 122760 -147180 122780 -147080
rect 120540 -147200 122780 -147180
rect 123540 -147080 125780 -147060
rect 123540 -147180 123560 -147080
rect 125760 -147180 125780 -147080
rect 123540 -147200 125780 -147180
rect 126540 -147080 128780 -147060
rect 126540 -147180 126560 -147080
rect 128760 -147180 128780 -147080
rect 126540 -147200 128780 -147180
rect 129540 -147080 131780 -147060
rect 129540 -147180 129560 -147080
rect 131760 -147180 131780 -147080
rect 129540 -147200 131780 -147180
rect 132540 -147080 134780 -147060
rect 132540 -147180 132560 -147080
rect 134760 -147180 134780 -147080
rect 132540 -147200 134780 -147180
rect 135540 -147080 137780 -147060
rect 135540 -147180 135560 -147080
rect 137760 -147180 137780 -147080
rect 135540 -147200 137780 -147180
rect 138540 -147080 140780 -147060
rect 138540 -147180 138560 -147080
rect 140760 -147180 140780 -147080
rect 138540 -147200 140780 -147180
rect 141540 -147080 143780 -147060
rect 141540 -147180 141560 -147080
rect 143760 -147180 143780 -147080
rect 141540 -147200 143780 -147180
rect 144540 -147080 146780 -147060
rect 144540 -147180 144560 -147080
rect 146760 -147180 146780 -147080
rect 144540 -147200 146780 -147180
rect 147540 -147080 149780 -147060
rect 147540 -147180 147560 -147080
rect 149760 -147180 149780 -147080
rect 147540 -147200 149780 -147180
rect 220 -147500 440 -147490
rect 220 -147700 240 -147500
rect 420 -147700 440 -147500
rect 220 -147710 440 -147700
rect 3220 -147500 3440 -147490
rect 3220 -147700 3240 -147500
rect 3420 -147700 3440 -147500
rect 3220 -147710 3440 -147700
rect 6220 -147500 6440 -147490
rect 6220 -147700 6240 -147500
rect 6420 -147700 6440 -147500
rect 6220 -147710 6440 -147700
rect 9220 -147500 9440 -147490
rect 9220 -147700 9240 -147500
rect 9420 -147700 9440 -147500
rect 9220 -147710 9440 -147700
rect 12220 -147500 12440 -147490
rect 12220 -147700 12240 -147500
rect 12420 -147700 12440 -147500
rect 12220 -147710 12440 -147700
rect 15220 -147500 15440 -147490
rect 15220 -147700 15240 -147500
rect 15420 -147700 15440 -147500
rect 15220 -147710 15440 -147700
rect 18220 -147500 18440 -147490
rect 18220 -147700 18240 -147500
rect 18420 -147700 18440 -147500
rect 18220 -147710 18440 -147700
rect 21220 -147500 21440 -147490
rect 21220 -147700 21240 -147500
rect 21420 -147700 21440 -147500
rect 21220 -147710 21440 -147700
rect 24220 -147500 24440 -147490
rect 24220 -147700 24240 -147500
rect 24420 -147700 24440 -147500
rect 24220 -147710 24440 -147700
rect 27220 -147500 27440 -147490
rect 27220 -147700 27240 -147500
rect 27420 -147700 27440 -147500
rect 27220 -147710 27440 -147700
rect 30220 -147500 30440 -147490
rect 30220 -147700 30240 -147500
rect 30420 -147700 30440 -147500
rect 30220 -147710 30440 -147700
rect 33220 -147500 33440 -147490
rect 33220 -147700 33240 -147500
rect 33420 -147700 33440 -147500
rect 33220 -147710 33440 -147700
rect 36220 -147500 36440 -147490
rect 36220 -147700 36240 -147500
rect 36420 -147700 36440 -147500
rect 36220 -147710 36440 -147700
rect 39220 -147500 39440 -147490
rect 39220 -147700 39240 -147500
rect 39420 -147700 39440 -147500
rect 39220 -147710 39440 -147700
rect 42220 -147500 42440 -147490
rect 42220 -147700 42240 -147500
rect 42420 -147700 42440 -147500
rect 42220 -147710 42440 -147700
rect 45220 -147500 45440 -147490
rect 45220 -147700 45240 -147500
rect 45420 -147700 45440 -147500
rect 45220 -147710 45440 -147700
rect 48220 -147500 48440 -147490
rect 48220 -147700 48240 -147500
rect 48420 -147700 48440 -147500
rect 48220 -147710 48440 -147700
rect 51220 -147500 51440 -147490
rect 51220 -147700 51240 -147500
rect 51420 -147700 51440 -147500
rect 51220 -147710 51440 -147700
rect 54220 -147500 54440 -147490
rect 54220 -147700 54240 -147500
rect 54420 -147700 54440 -147500
rect 54220 -147710 54440 -147700
rect 57220 -147500 57440 -147490
rect 57220 -147700 57240 -147500
rect 57420 -147700 57440 -147500
rect 57220 -147710 57440 -147700
rect 60220 -147500 60440 -147490
rect 60220 -147700 60240 -147500
rect 60420 -147700 60440 -147500
rect 60220 -147710 60440 -147700
rect 63220 -147500 63440 -147490
rect 63220 -147700 63240 -147500
rect 63420 -147700 63440 -147500
rect 63220 -147710 63440 -147700
rect 66220 -147500 66440 -147490
rect 66220 -147700 66240 -147500
rect 66420 -147700 66440 -147500
rect 66220 -147710 66440 -147700
rect 69220 -147500 69440 -147490
rect 69220 -147700 69240 -147500
rect 69420 -147700 69440 -147500
rect 69220 -147710 69440 -147700
rect 72220 -147500 72440 -147490
rect 72220 -147700 72240 -147500
rect 72420 -147700 72440 -147500
rect 72220 -147710 72440 -147700
rect 75220 -147500 75440 -147490
rect 75220 -147700 75240 -147500
rect 75420 -147700 75440 -147500
rect 75220 -147710 75440 -147700
rect 78220 -147500 78440 -147490
rect 78220 -147700 78240 -147500
rect 78420 -147700 78440 -147500
rect 78220 -147710 78440 -147700
rect 81220 -147500 81440 -147490
rect 81220 -147700 81240 -147500
rect 81420 -147700 81440 -147500
rect 81220 -147710 81440 -147700
rect 84220 -147500 84440 -147490
rect 84220 -147700 84240 -147500
rect 84420 -147700 84440 -147500
rect 84220 -147710 84440 -147700
rect 87220 -147500 87440 -147490
rect 87220 -147700 87240 -147500
rect 87420 -147700 87440 -147500
rect 87220 -147710 87440 -147700
rect 90220 -147500 90440 -147490
rect 90220 -147700 90240 -147500
rect 90420 -147700 90440 -147500
rect 90220 -147710 90440 -147700
rect 93220 -147500 93440 -147490
rect 93220 -147700 93240 -147500
rect 93420 -147700 93440 -147500
rect 93220 -147710 93440 -147700
rect 96220 -147500 96440 -147490
rect 96220 -147700 96240 -147500
rect 96420 -147700 96440 -147500
rect 96220 -147710 96440 -147700
rect 99220 -147500 99440 -147490
rect 99220 -147700 99240 -147500
rect 99420 -147700 99440 -147500
rect 99220 -147710 99440 -147700
rect 102220 -147500 102440 -147490
rect 102220 -147700 102240 -147500
rect 102420 -147700 102440 -147500
rect 102220 -147710 102440 -147700
rect 105220 -147500 105440 -147490
rect 105220 -147700 105240 -147500
rect 105420 -147700 105440 -147500
rect 105220 -147710 105440 -147700
rect 108220 -147500 108440 -147490
rect 108220 -147700 108240 -147500
rect 108420 -147700 108440 -147500
rect 108220 -147710 108440 -147700
rect 111220 -147500 111440 -147490
rect 111220 -147700 111240 -147500
rect 111420 -147700 111440 -147500
rect 111220 -147710 111440 -147700
rect 114220 -147500 114440 -147490
rect 114220 -147700 114240 -147500
rect 114420 -147700 114440 -147500
rect 114220 -147710 114440 -147700
rect 117220 -147500 117440 -147490
rect 117220 -147700 117240 -147500
rect 117420 -147700 117440 -147500
rect 117220 -147710 117440 -147700
rect 120220 -147500 120440 -147490
rect 120220 -147700 120240 -147500
rect 120420 -147700 120440 -147500
rect 120220 -147710 120440 -147700
rect 123220 -147500 123440 -147490
rect 123220 -147700 123240 -147500
rect 123420 -147700 123440 -147500
rect 123220 -147710 123440 -147700
rect 126220 -147500 126440 -147490
rect 126220 -147700 126240 -147500
rect 126420 -147700 126440 -147500
rect 126220 -147710 126440 -147700
rect 129220 -147500 129440 -147490
rect 129220 -147700 129240 -147500
rect 129420 -147700 129440 -147500
rect 129220 -147710 129440 -147700
rect 132220 -147500 132440 -147490
rect 132220 -147700 132240 -147500
rect 132420 -147700 132440 -147500
rect 132220 -147710 132440 -147700
rect 135220 -147500 135440 -147490
rect 135220 -147700 135240 -147500
rect 135420 -147700 135440 -147500
rect 135220 -147710 135440 -147700
rect 138220 -147500 138440 -147490
rect 138220 -147700 138240 -147500
rect 138420 -147700 138440 -147500
rect 138220 -147710 138440 -147700
rect 141220 -147500 141440 -147490
rect 141220 -147700 141240 -147500
rect 141420 -147700 141440 -147500
rect 141220 -147710 141440 -147700
rect 144220 -147500 144440 -147490
rect 144220 -147700 144240 -147500
rect 144420 -147700 144440 -147500
rect 144220 -147710 144440 -147700
rect 147220 -147500 147440 -147490
rect 147220 -147700 147240 -147500
rect 147420 -147700 147440 -147500
rect 147220 -147710 147440 -147700
<< via3 >>
rect 490 3560 580 3650
rect 3490 3560 3580 3650
rect 6490 3560 6580 3650
rect 9490 3560 9580 3650
rect 12490 3560 12580 3650
rect 15490 3560 15580 3650
rect 18490 3560 18580 3650
rect 21490 3560 21580 3650
rect 24490 3560 24580 3650
rect 27490 3560 27580 3650
rect 30490 3560 30580 3650
rect 33490 3560 33580 3650
rect 36490 3560 36580 3650
rect 39490 3560 39580 3650
rect 42490 3560 42580 3650
rect 45490 3560 45580 3650
rect 48490 3560 48580 3650
rect 51490 3560 51580 3650
rect 54490 3560 54580 3650
rect 57490 3560 57580 3650
rect 60490 3560 60580 3650
rect 63490 3560 63580 3650
rect 66490 3560 66580 3650
rect 69490 3560 69580 3650
rect 72490 3560 72580 3650
rect 75490 3560 75580 3650
rect 78490 3560 78580 3650
rect 81490 3560 81580 3650
rect 84490 3560 84580 3650
rect 87490 3560 87580 3650
rect 90490 3560 90580 3650
rect 93490 3560 93580 3650
rect 96490 3560 96580 3650
rect 99490 3560 99580 3650
rect 102490 3560 102580 3650
rect 105490 3560 105580 3650
rect 108490 3560 108580 3650
rect 111490 3560 111580 3650
rect 114490 3560 114580 3650
rect 117490 3560 117580 3650
rect 120490 3560 120580 3650
rect 123490 3560 123580 3650
rect 126490 3560 126580 3650
rect 129490 3560 129580 3650
rect 132490 3560 132580 3650
rect 135490 3560 135580 3650
rect 138490 3560 138580 3650
rect 141490 3560 141580 3650
rect 144490 3560 144580 3650
rect 147490 3560 147580 3650
rect -470 2470 -380 2540
rect -470 -530 -380 -460
rect -470 -3530 -380 -3460
rect -470 -6530 -380 -6460
rect -470 -9530 -380 -9460
rect -470 -12530 -380 -12460
rect -470 -15530 -380 -15460
rect -470 -18530 -380 -18460
rect -470 -21530 -380 -21460
rect -470 -24530 -380 -24460
rect -470 -27530 -380 -27460
rect -470 -30530 -380 -30460
rect -470 -33530 -380 -33460
rect -470 -36530 -380 -36460
rect -470 -39530 -380 -39460
rect -470 -42530 -380 -42460
rect -470 -45530 -380 -45460
rect -470 -48530 -380 -48460
rect -470 -51530 -380 -51460
rect -470 -54530 -380 -54460
rect -470 -57530 -380 -57460
rect -470 -60530 -380 -60460
rect -470 -63530 -380 -63460
rect -470 -66530 -380 -66460
rect -470 -69530 -380 -69460
rect -470 -72530 -380 -72460
rect -470 -75530 -380 -75460
rect -470 -78530 -380 -78460
rect -470 -81530 -380 -81460
rect -470 -84530 -380 -84460
rect -470 -87530 -380 -87460
rect -470 -90530 -380 -90460
rect -470 -93530 -380 -93460
rect -470 -96530 -380 -96460
rect -470 -99530 -380 -99460
rect -470 -102530 -380 -102460
rect -470 -105530 -380 -105460
rect -470 -108530 -380 -108460
rect -470 -111530 -380 -111460
rect -470 -114530 -380 -114460
rect -470 -117530 -380 -117460
rect -470 -120530 -380 -120460
rect -470 -123530 -380 -123460
rect -470 -126530 -380 -126460
rect -470 -129530 -380 -129460
rect -470 -132530 -380 -132460
rect -470 -135530 -380 -135460
rect -470 -138530 -380 -138460
rect -470 -141530 -380 -141460
rect -470 -144530 -380 -144460
rect 560 -147180 2760 -147080
rect 3560 -147180 5760 -147080
rect 6560 -147180 8760 -147080
rect 9560 -147180 11760 -147080
rect 12560 -147180 14760 -147080
rect 15560 -147180 17760 -147080
rect 18560 -147180 20760 -147080
rect 21560 -147180 23760 -147080
rect 24560 -147180 26760 -147080
rect 27560 -147180 29760 -147080
rect 30560 -147180 32760 -147080
rect 33560 -147180 35760 -147080
rect 36560 -147180 38760 -147080
rect 39560 -147180 41760 -147080
rect 42560 -147180 44760 -147080
rect 45560 -147180 47760 -147080
rect 48560 -147180 50760 -147080
rect 51560 -147180 53760 -147080
rect 54560 -147180 56760 -147080
rect 57560 -147180 59760 -147080
rect 60560 -147180 62760 -147080
rect 63560 -147180 65760 -147080
rect 66560 -147180 68760 -147080
rect 69560 -147180 71760 -147080
rect 72560 -147180 74760 -147080
rect 75560 -147180 77760 -147080
rect 78560 -147180 80760 -147080
rect 81560 -147180 83760 -147080
rect 84560 -147180 86760 -147080
rect 87560 -147180 89760 -147080
rect 90560 -147180 92760 -147080
rect 93560 -147180 95760 -147080
rect 96560 -147180 98760 -147080
rect 99560 -147180 101760 -147080
rect 102560 -147180 104760 -147080
rect 105560 -147180 107760 -147080
rect 108560 -147180 110760 -147080
rect 111560 -147180 113760 -147080
rect 114560 -147180 116760 -147080
rect 117560 -147180 119760 -147080
rect 120560 -147180 122760 -147080
rect 123560 -147180 125760 -147080
rect 126560 -147180 128760 -147080
rect 129560 -147180 131760 -147080
rect 132560 -147180 134760 -147080
rect 135560 -147180 137760 -147080
rect 138560 -147180 140760 -147080
rect 141560 -147180 143760 -147080
rect 144560 -147180 146760 -147080
rect 147560 -147180 149760 -147080
rect 240 -147700 420 -147500
rect 3240 -147700 3420 -147500
rect 6240 -147700 6420 -147500
rect 9240 -147700 9420 -147500
rect 12240 -147700 12420 -147500
rect 15240 -147700 15420 -147500
rect 18240 -147700 18420 -147500
rect 21240 -147700 21420 -147500
rect 24240 -147700 24420 -147500
rect 27240 -147700 27420 -147500
rect 30240 -147700 30420 -147500
rect 33240 -147700 33420 -147500
rect 36240 -147700 36420 -147500
rect 39240 -147700 39420 -147500
rect 42240 -147700 42420 -147500
rect 45240 -147700 45420 -147500
rect 48240 -147700 48420 -147500
rect 51240 -147700 51420 -147500
rect 54240 -147700 54420 -147500
rect 57240 -147700 57420 -147500
rect 60240 -147700 60420 -147500
rect 63240 -147700 63420 -147500
rect 66240 -147700 66420 -147500
rect 69240 -147700 69420 -147500
rect 72240 -147700 72420 -147500
rect 75240 -147700 75420 -147500
rect 78240 -147700 78420 -147500
rect 81240 -147700 81420 -147500
rect 84240 -147700 84420 -147500
rect 87240 -147700 87420 -147500
rect 90240 -147700 90420 -147500
rect 93240 -147700 93420 -147500
rect 96240 -147700 96420 -147500
rect 99240 -147700 99420 -147500
rect 102240 -147700 102420 -147500
rect 105240 -147700 105420 -147500
rect 108240 -147700 108420 -147500
rect 111240 -147700 111420 -147500
rect 114240 -147700 114420 -147500
rect 117240 -147700 117420 -147500
rect 120240 -147700 120420 -147500
rect 123240 -147700 123420 -147500
rect 126240 -147700 126420 -147500
rect 129240 -147700 129420 -147500
rect 132240 -147700 132420 -147500
rect 135240 -147700 135420 -147500
rect 138240 -147700 138420 -147500
rect 141240 -147700 141420 -147500
rect 144240 -147700 144420 -147500
rect 147240 -147700 147420 -147500
<< metal4 >>
rect -3000 3650 149200 3660
rect -3000 3560 490 3650
rect 580 3560 3490 3650
rect 3580 3560 6490 3650
rect 6580 3560 9490 3650
rect 9580 3560 12490 3650
rect 12580 3560 15490 3650
rect 15580 3560 18490 3650
rect 18580 3560 21490 3650
rect 21580 3560 24490 3650
rect 24580 3560 27490 3650
rect 27580 3560 30490 3650
rect 30580 3560 33490 3650
rect 33580 3560 36490 3650
rect 36580 3560 39490 3650
rect 39580 3560 42490 3650
rect 42580 3560 45490 3650
rect 45580 3560 48490 3650
rect 48580 3560 51490 3650
rect 51580 3560 54490 3650
rect 54580 3560 57490 3650
rect 57580 3560 60490 3650
rect 60580 3560 63490 3650
rect 63580 3560 66490 3650
rect 66580 3560 69490 3650
rect 69580 3560 72490 3650
rect 72580 3560 75490 3650
rect 75580 3560 78490 3650
rect 78580 3560 81490 3650
rect 81580 3560 84490 3650
rect 84580 3560 87490 3650
rect 87580 3560 90490 3650
rect 90580 3560 93490 3650
rect 93580 3560 96490 3650
rect 96580 3560 99490 3650
rect 99580 3560 102490 3650
rect 102580 3560 105490 3650
rect 105580 3560 108490 3650
rect 108580 3560 111490 3650
rect 111580 3560 114490 3650
rect 114580 3560 117490 3650
rect 117580 3560 120490 3650
rect 120580 3560 123490 3650
rect 123580 3560 126490 3650
rect 126580 3560 129490 3650
rect 129580 3560 132490 3650
rect 132580 3560 135490 3650
rect 135580 3560 138490 3650
rect 138580 3560 141490 3650
rect 141580 3560 144490 3650
rect 144580 3560 147490 3650
rect 147580 3560 149200 3650
rect -3000 3550 149200 3560
rect -480 2540 -370 2600
rect -480 2470 -470 2540
rect -380 2470 -370 2540
rect -480 -460 -370 2470
rect -480 -530 -470 -460
rect -380 -530 -370 -460
rect -480 -3460 -370 -530
rect -480 -3530 -470 -3460
rect -380 -3530 -370 -3460
rect -480 -6460 -370 -3530
rect -480 -6530 -470 -6460
rect -380 -6530 -370 -6460
rect -480 -9460 -370 -6530
rect -480 -9530 -470 -9460
rect -380 -9530 -370 -9460
rect -480 -12460 -370 -9530
rect -480 -12530 -470 -12460
rect -380 -12530 -370 -12460
rect -480 -15460 -370 -12530
rect -480 -15530 -470 -15460
rect -380 -15530 -370 -15460
rect -480 -18460 -370 -15530
rect -480 -18530 -470 -18460
rect -380 -18530 -370 -18460
rect -480 -21460 -370 -18530
rect -480 -21530 -470 -21460
rect -380 -21530 -370 -21460
rect -480 -24460 -370 -21530
rect -480 -24530 -470 -24460
rect -380 -24530 -370 -24460
rect -480 -27460 -370 -24530
rect -480 -27530 -470 -27460
rect -380 -27530 -370 -27460
rect -480 -30460 -370 -27530
rect -480 -30530 -470 -30460
rect -380 -30530 -370 -30460
rect -480 -33460 -370 -30530
rect -480 -33530 -470 -33460
rect -380 -33530 -370 -33460
rect -480 -36460 -370 -33530
rect -480 -36530 -470 -36460
rect -380 -36530 -370 -36460
rect -480 -39460 -370 -36530
rect -480 -39530 -470 -39460
rect -380 -39530 -370 -39460
rect -480 -42460 -370 -39530
rect -480 -42530 -470 -42460
rect -380 -42530 -370 -42460
rect -480 -45460 -370 -42530
rect -480 -45530 -470 -45460
rect -380 -45530 -370 -45460
rect -480 -48460 -370 -45530
rect -480 -48530 -470 -48460
rect -380 -48530 -370 -48460
rect -480 -51460 -370 -48530
rect -480 -51530 -470 -51460
rect -380 -51530 -370 -51460
rect -480 -54460 -370 -51530
rect -480 -54530 -470 -54460
rect -380 -54530 -370 -54460
rect -480 -57460 -370 -54530
rect -480 -57530 -470 -57460
rect -380 -57530 -370 -57460
rect -480 -60460 -370 -57530
rect -480 -60530 -470 -60460
rect -380 -60530 -370 -60460
rect -480 -63460 -370 -60530
rect -480 -63530 -470 -63460
rect -380 -63530 -370 -63460
rect -480 -66460 -370 -63530
rect -480 -66530 -470 -66460
rect -380 -66530 -370 -66460
rect -480 -69460 -370 -66530
rect -480 -69530 -470 -69460
rect -380 -69530 -370 -69460
rect -480 -72460 -370 -69530
rect -480 -72530 -470 -72460
rect -380 -72530 -370 -72460
rect -480 -75460 -370 -72530
rect -480 -75530 -470 -75460
rect -380 -75530 -370 -75460
rect -480 -78460 -370 -75530
rect -480 -78530 -470 -78460
rect -380 -78530 -370 -78460
rect -480 -81460 -370 -78530
rect -480 -81530 -470 -81460
rect -380 -81530 -370 -81460
rect -480 -84460 -370 -81530
rect -480 -84530 -470 -84460
rect -380 -84530 -370 -84460
rect -480 -87460 -370 -84530
rect -480 -87530 -470 -87460
rect -380 -87530 -370 -87460
rect -480 -90460 -370 -87530
rect -480 -90530 -470 -90460
rect -380 -90530 -370 -90460
rect -480 -93460 -370 -90530
rect -480 -93530 -470 -93460
rect -380 -93530 -370 -93460
rect -480 -96460 -370 -93530
rect -480 -96530 -470 -96460
rect -380 -96530 -370 -96460
rect -480 -99460 -370 -96530
rect -480 -99530 -470 -99460
rect -380 -99530 -370 -99460
rect -480 -102460 -370 -99530
rect -480 -102530 -470 -102460
rect -380 -102530 -370 -102460
rect -480 -105460 -370 -102530
rect -480 -105530 -470 -105460
rect -380 -105530 -370 -105460
rect -480 -108460 -370 -105530
rect -480 -108530 -470 -108460
rect -380 -108530 -370 -108460
rect -480 -111460 -370 -108530
rect -480 -111530 -470 -111460
rect -380 -111530 -370 -111460
rect -480 -114460 -370 -111530
rect -480 -114530 -470 -114460
rect -380 -114530 -370 -114460
rect -480 -117460 -370 -114530
rect -480 -117530 -470 -117460
rect -380 -117530 -370 -117460
rect -480 -120460 -370 -117530
rect -480 -120530 -470 -120460
rect -380 -120530 -370 -120460
rect -480 -123460 -370 -120530
rect -480 -123530 -470 -123460
rect -380 -123530 -370 -123460
rect -480 -126460 -370 -123530
rect -480 -126530 -470 -126460
rect -380 -126530 -370 -126460
rect -480 -129460 -370 -126530
rect -480 -129530 -470 -129460
rect -380 -129530 -370 -129460
rect -480 -132460 -370 -129530
rect -480 -132530 -470 -132460
rect -380 -132530 -370 -132460
rect -480 -135460 -370 -132530
rect -480 -135530 -470 -135460
rect -380 -135530 -370 -135460
rect -480 -138460 -370 -135530
rect -480 -138530 -470 -138460
rect -380 -138530 -370 -138460
rect -480 -141460 -370 -138530
rect -480 -141530 -470 -141460
rect -380 -141530 -370 -141460
rect -480 -144460 -370 -141530
rect -480 -144530 -470 -144460
rect -380 -144530 -370 -144460
rect -480 -148600 -370 -144530
rect 2630 -147060 2780 -147000
rect 5630 -147060 5780 -147000
rect 8630 -147060 8780 -147000
rect 11630 -147060 11780 -147000
rect 14630 -147060 14780 -147000
rect 17630 -147060 17780 -147000
rect 20630 -147060 20780 -147000
rect 23630 -147060 23780 -147000
rect 26630 -147060 26780 -147000
rect 29630 -147060 29780 -147000
rect 32630 -147060 32780 -147000
rect 35630 -147060 35780 -147000
rect 38630 -147060 38780 -147000
rect 41630 -147060 41780 -147000
rect 44630 -147060 44780 -147000
rect 47630 -147060 47780 -147000
rect 50630 -147060 50780 -147000
rect 53630 -147060 53780 -147000
rect 56630 -147060 56780 -147000
rect 59630 -147060 59780 -147000
rect 62630 -147060 62780 -147000
rect 65630 -147060 65780 -147000
rect 68630 -147060 68780 -147000
rect 71630 -147060 71780 -147000
rect 74630 -147060 74780 -147000
rect 77630 -147060 77780 -147000
rect 80630 -147060 80780 -147000
rect 83630 -147060 83780 -147000
rect 86630 -147060 86780 -147000
rect 89630 -147060 89780 -147000
rect 92630 -147060 92780 -147000
rect 95630 -147060 95780 -147000
rect 98630 -147060 98780 -147000
rect 101630 -147060 101780 -147000
rect 104630 -147060 104780 -147000
rect 107630 -147060 107780 -147000
rect 110630 -147060 110780 -147000
rect 113630 -147060 113780 -147000
rect 116630 -147060 116780 -147000
rect 119630 -147060 119780 -147000
rect 122630 -147060 122780 -147000
rect 125630 -147060 125780 -147000
rect 128630 -147060 128780 -147000
rect 131630 -147060 131780 -147000
rect 134630 -147060 134780 -147000
rect 137630 -147060 137780 -147000
rect 140630 -147060 140780 -147000
rect 143630 -147060 143780 -147000
rect 146630 -147060 146780 -147000
rect 149630 -147060 149780 -147000
rect 540 -147080 2780 -147060
rect 540 -147180 560 -147080
rect 2760 -147180 2780 -147080
rect 540 -147200 2780 -147180
rect 3540 -147080 5780 -147060
rect 3540 -147180 3560 -147080
rect 5760 -147180 5780 -147080
rect 3540 -147200 5780 -147180
rect 6540 -147080 8780 -147060
rect 6540 -147180 6560 -147080
rect 8760 -147180 8780 -147080
rect 6540 -147200 8780 -147180
rect 9540 -147080 11780 -147060
rect 9540 -147180 9560 -147080
rect 11760 -147180 11780 -147080
rect 9540 -147200 11780 -147180
rect 12540 -147080 14780 -147060
rect 12540 -147180 12560 -147080
rect 14760 -147180 14780 -147080
rect 12540 -147200 14780 -147180
rect 15540 -147080 17780 -147060
rect 15540 -147180 15560 -147080
rect 17760 -147180 17780 -147080
rect 15540 -147200 17780 -147180
rect 18540 -147080 20780 -147060
rect 18540 -147180 18560 -147080
rect 20760 -147180 20780 -147080
rect 18540 -147200 20780 -147180
rect 21540 -147080 23780 -147060
rect 21540 -147180 21560 -147080
rect 23760 -147180 23780 -147080
rect 21540 -147200 23780 -147180
rect 24540 -147080 26780 -147060
rect 24540 -147180 24560 -147080
rect 26760 -147180 26780 -147080
rect 24540 -147200 26780 -147180
rect 27540 -147080 29780 -147060
rect 27540 -147180 27560 -147080
rect 29760 -147180 29780 -147080
rect 27540 -147200 29780 -147180
rect 30540 -147080 32780 -147060
rect 30540 -147180 30560 -147080
rect 32760 -147180 32780 -147080
rect 30540 -147200 32780 -147180
rect 33540 -147080 35780 -147060
rect 33540 -147180 33560 -147080
rect 35760 -147180 35780 -147080
rect 33540 -147200 35780 -147180
rect 36540 -147080 38780 -147060
rect 36540 -147180 36560 -147080
rect 38760 -147180 38780 -147080
rect 36540 -147200 38780 -147180
rect 39540 -147080 41780 -147060
rect 39540 -147180 39560 -147080
rect 41760 -147180 41780 -147080
rect 39540 -147200 41780 -147180
rect 42540 -147080 44780 -147060
rect 42540 -147180 42560 -147080
rect 44760 -147180 44780 -147080
rect 42540 -147200 44780 -147180
rect 45540 -147080 47780 -147060
rect 45540 -147180 45560 -147080
rect 47760 -147180 47780 -147080
rect 45540 -147200 47780 -147180
rect 48540 -147080 50780 -147060
rect 48540 -147180 48560 -147080
rect 50760 -147180 50780 -147080
rect 48540 -147200 50780 -147180
rect 51540 -147080 53780 -147060
rect 51540 -147180 51560 -147080
rect 53760 -147180 53780 -147080
rect 51540 -147200 53780 -147180
rect 54540 -147080 56780 -147060
rect 54540 -147180 54560 -147080
rect 56760 -147180 56780 -147080
rect 54540 -147200 56780 -147180
rect 57540 -147080 59780 -147060
rect 57540 -147180 57560 -147080
rect 59760 -147180 59780 -147080
rect 57540 -147200 59780 -147180
rect 60540 -147080 62780 -147060
rect 60540 -147180 60560 -147080
rect 62760 -147180 62780 -147080
rect 60540 -147200 62780 -147180
rect 63540 -147080 65780 -147060
rect 63540 -147180 63560 -147080
rect 65760 -147180 65780 -147080
rect 63540 -147200 65780 -147180
rect 66540 -147080 68780 -147060
rect 66540 -147180 66560 -147080
rect 68760 -147180 68780 -147080
rect 66540 -147200 68780 -147180
rect 69540 -147080 71780 -147060
rect 69540 -147180 69560 -147080
rect 71760 -147180 71780 -147080
rect 69540 -147200 71780 -147180
rect 72540 -147080 74780 -147060
rect 72540 -147180 72560 -147080
rect 74760 -147180 74780 -147080
rect 72540 -147200 74780 -147180
rect 75540 -147080 77780 -147060
rect 75540 -147180 75560 -147080
rect 77760 -147180 77780 -147080
rect 75540 -147200 77780 -147180
rect 78540 -147080 80780 -147060
rect 78540 -147180 78560 -147080
rect 80760 -147180 80780 -147080
rect 78540 -147200 80780 -147180
rect 81540 -147080 83780 -147060
rect 81540 -147180 81560 -147080
rect 83760 -147180 83780 -147080
rect 81540 -147200 83780 -147180
rect 84540 -147080 86780 -147060
rect 84540 -147180 84560 -147080
rect 86760 -147180 86780 -147080
rect 84540 -147200 86780 -147180
rect 87540 -147080 89780 -147060
rect 87540 -147180 87560 -147080
rect 89760 -147180 89780 -147080
rect 87540 -147200 89780 -147180
rect 90540 -147080 92780 -147060
rect 90540 -147180 90560 -147080
rect 92760 -147180 92780 -147080
rect 90540 -147200 92780 -147180
rect 93540 -147080 95780 -147060
rect 93540 -147180 93560 -147080
rect 95760 -147180 95780 -147080
rect 93540 -147200 95780 -147180
rect 96540 -147080 98780 -147060
rect 96540 -147180 96560 -147080
rect 98760 -147180 98780 -147080
rect 96540 -147200 98780 -147180
rect 99540 -147080 101780 -147060
rect 99540 -147180 99560 -147080
rect 101760 -147180 101780 -147080
rect 99540 -147200 101780 -147180
rect 102540 -147080 104780 -147060
rect 102540 -147180 102560 -147080
rect 104760 -147180 104780 -147080
rect 102540 -147200 104780 -147180
rect 105540 -147080 107780 -147060
rect 105540 -147180 105560 -147080
rect 107760 -147180 107780 -147080
rect 105540 -147200 107780 -147180
rect 108540 -147080 110780 -147060
rect 108540 -147180 108560 -147080
rect 110760 -147180 110780 -147080
rect 108540 -147200 110780 -147180
rect 111540 -147080 113780 -147060
rect 111540 -147180 111560 -147080
rect 113760 -147180 113780 -147080
rect 111540 -147200 113780 -147180
rect 114540 -147080 116780 -147060
rect 114540 -147180 114560 -147080
rect 116760 -147180 116780 -147080
rect 114540 -147200 116780 -147180
rect 117540 -147080 119780 -147060
rect 117540 -147180 117560 -147080
rect 119760 -147180 119780 -147080
rect 117540 -147200 119780 -147180
rect 120540 -147080 122780 -147060
rect 120540 -147180 120560 -147080
rect 122760 -147180 122780 -147080
rect 120540 -147200 122780 -147180
rect 123540 -147080 125780 -147060
rect 123540 -147180 123560 -147080
rect 125760 -147180 125780 -147080
rect 123540 -147200 125780 -147180
rect 126540 -147080 128780 -147060
rect 126540 -147180 126560 -147080
rect 128760 -147180 128780 -147080
rect 126540 -147200 128780 -147180
rect 129540 -147080 131780 -147060
rect 129540 -147180 129560 -147080
rect 131760 -147180 131780 -147080
rect 129540 -147200 131780 -147180
rect 132540 -147080 134780 -147060
rect 132540 -147180 132560 -147080
rect 134760 -147180 134780 -147080
rect 132540 -147200 134780 -147180
rect 135540 -147080 137780 -147060
rect 135540 -147180 135560 -147080
rect 137760 -147180 137780 -147080
rect 135540 -147200 137780 -147180
rect 138540 -147080 140780 -147060
rect 138540 -147180 138560 -147080
rect 140760 -147180 140780 -147080
rect 138540 -147200 140780 -147180
rect 141540 -147080 143780 -147060
rect 141540 -147180 141560 -147080
rect 143760 -147180 143780 -147080
rect 141540 -147200 143780 -147180
rect 144540 -147080 146780 -147060
rect 144540 -147180 144560 -147080
rect 146760 -147180 146780 -147080
rect 144540 -147200 146780 -147180
rect 147540 -147080 149780 -147060
rect 147540 -147180 147560 -147080
rect 149760 -147180 149780 -147080
rect 147540 -147200 149780 -147180
rect 220 -147500 440 -147490
rect 220 -147700 240 -147500
rect 420 -147700 440 -147500
rect 220 -148100 440 -147700
rect 3220 -147500 3440 -147490
rect 3220 -147700 3240 -147500
rect 3420 -147700 3440 -147500
rect 3220 -148100 3440 -147700
rect 6220 -147500 6440 -147490
rect 6220 -147700 6240 -147500
rect 6420 -147700 6440 -147500
rect 6220 -148100 6440 -147700
rect 9220 -147500 9440 -147490
rect 9220 -147700 9240 -147500
rect 9420 -147700 9440 -147500
rect 9220 -148100 9440 -147700
rect 12220 -147500 12440 -147490
rect 12220 -147700 12240 -147500
rect 12420 -147700 12440 -147500
rect 12220 -148100 12440 -147700
rect 15220 -147500 15440 -147490
rect 15220 -147700 15240 -147500
rect 15420 -147700 15440 -147500
rect 15220 -148100 15440 -147700
rect 18220 -147500 18440 -147490
rect 18220 -147700 18240 -147500
rect 18420 -147700 18440 -147500
rect 18220 -148100 18440 -147700
rect 21220 -147500 21440 -147490
rect 21220 -147700 21240 -147500
rect 21420 -147700 21440 -147500
rect 21220 -148100 21440 -147700
rect 24220 -147500 24440 -147490
rect 24220 -147700 24240 -147500
rect 24420 -147700 24440 -147500
rect 24220 -148100 24440 -147700
rect 27220 -147500 27440 -147490
rect 27220 -147700 27240 -147500
rect 27420 -147700 27440 -147500
rect 27220 -148100 27440 -147700
rect 30220 -147500 30440 -147490
rect 30220 -147700 30240 -147500
rect 30420 -147700 30440 -147500
rect 30220 -148100 30440 -147700
rect 33220 -147500 33440 -147490
rect 33220 -147700 33240 -147500
rect 33420 -147700 33440 -147500
rect 33220 -148100 33440 -147700
rect 36220 -147500 36440 -147490
rect 36220 -147700 36240 -147500
rect 36420 -147700 36440 -147500
rect 36220 -148100 36440 -147700
rect 39220 -147500 39440 -147490
rect 39220 -147700 39240 -147500
rect 39420 -147700 39440 -147500
rect 39220 -148100 39440 -147700
rect 42220 -147500 42440 -147490
rect 42220 -147700 42240 -147500
rect 42420 -147700 42440 -147500
rect 42220 -148100 42440 -147700
rect 45220 -147500 45440 -147490
rect 45220 -147700 45240 -147500
rect 45420 -147700 45440 -147500
rect 45220 -148100 45440 -147700
rect 48220 -147500 48440 -147490
rect 48220 -147700 48240 -147500
rect 48420 -147700 48440 -147500
rect 48220 -148100 48440 -147700
rect 51220 -147500 51440 -147490
rect 51220 -147700 51240 -147500
rect 51420 -147700 51440 -147500
rect 51220 -148100 51440 -147700
rect 54220 -147500 54440 -147490
rect 54220 -147700 54240 -147500
rect 54420 -147700 54440 -147500
rect 54220 -148100 54440 -147700
rect 57220 -147500 57440 -147490
rect 57220 -147700 57240 -147500
rect 57420 -147700 57440 -147500
rect 57220 -148100 57440 -147700
rect 60220 -147500 60440 -147490
rect 60220 -147700 60240 -147500
rect 60420 -147700 60440 -147500
rect 60220 -148100 60440 -147700
rect 63220 -147500 63440 -147490
rect 63220 -147700 63240 -147500
rect 63420 -147700 63440 -147500
rect 63220 -148100 63440 -147700
rect 66220 -147500 66440 -147490
rect 66220 -147700 66240 -147500
rect 66420 -147700 66440 -147500
rect 66220 -148100 66440 -147700
rect 69220 -147500 69440 -147490
rect 69220 -147700 69240 -147500
rect 69420 -147700 69440 -147500
rect 69220 -148100 69440 -147700
rect 72220 -147500 72440 -147490
rect 72220 -147700 72240 -147500
rect 72420 -147700 72440 -147500
rect 72220 -148100 72440 -147700
rect 75220 -147500 75440 -147490
rect 75220 -147700 75240 -147500
rect 75420 -147700 75440 -147500
rect 75220 -148100 75440 -147700
rect 78220 -147500 78440 -147490
rect 78220 -147700 78240 -147500
rect 78420 -147700 78440 -147500
rect 78220 -148100 78440 -147700
rect 81220 -147500 81440 -147490
rect 81220 -147700 81240 -147500
rect 81420 -147700 81440 -147500
rect 81220 -148100 81440 -147700
rect 84220 -147500 84440 -147490
rect 84220 -147700 84240 -147500
rect 84420 -147700 84440 -147500
rect 84220 -148100 84440 -147700
rect 87220 -147500 87440 -147490
rect 87220 -147700 87240 -147500
rect 87420 -147700 87440 -147500
rect 87220 -148100 87440 -147700
rect 90220 -147500 90440 -147490
rect 90220 -147700 90240 -147500
rect 90420 -147700 90440 -147500
rect 90220 -148100 90440 -147700
rect 93220 -147500 93440 -147490
rect 93220 -147700 93240 -147500
rect 93420 -147700 93440 -147500
rect 93220 -148100 93440 -147700
rect 96220 -147500 96440 -147490
rect 96220 -147700 96240 -147500
rect 96420 -147700 96440 -147500
rect 96220 -148100 96440 -147700
rect 99220 -147500 99440 -147490
rect 99220 -147700 99240 -147500
rect 99420 -147700 99440 -147500
rect 99220 -148100 99440 -147700
rect 102220 -147500 102440 -147490
rect 102220 -147700 102240 -147500
rect 102420 -147700 102440 -147500
rect 102220 -148100 102440 -147700
rect 105220 -147500 105440 -147490
rect 105220 -147700 105240 -147500
rect 105420 -147700 105440 -147500
rect 105220 -148100 105440 -147700
rect 108220 -147500 108440 -147490
rect 108220 -147700 108240 -147500
rect 108420 -147700 108440 -147500
rect 108220 -148100 108440 -147700
rect 111220 -147500 111440 -147490
rect 111220 -147700 111240 -147500
rect 111420 -147700 111440 -147500
rect 111220 -148100 111440 -147700
rect 114220 -147500 114440 -147490
rect 114220 -147700 114240 -147500
rect 114420 -147700 114440 -147500
rect 114220 -148100 114440 -147700
rect 117220 -147500 117440 -147490
rect 117220 -147700 117240 -147500
rect 117420 -147700 117440 -147500
rect 117220 -148100 117440 -147700
rect 120220 -147500 120440 -147490
rect 120220 -147700 120240 -147500
rect 120420 -147700 120440 -147500
rect 120220 -148100 120440 -147700
rect 123220 -147500 123440 -147490
rect 123220 -147700 123240 -147500
rect 123420 -147700 123440 -147500
rect 123220 -148100 123440 -147700
rect 126220 -147500 126440 -147490
rect 126220 -147700 126240 -147500
rect 126420 -147700 126440 -147500
rect 126220 -148100 126440 -147700
rect 129220 -147500 129440 -147490
rect 129220 -147700 129240 -147500
rect 129420 -147700 129440 -147500
rect 129220 -148100 129440 -147700
rect 132220 -147500 132440 -147490
rect 132220 -147700 132240 -147500
rect 132420 -147700 132440 -147500
rect 132220 -148100 132440 -147700
rect 135220 -147500 135440 -147490
rect 135220 -147700 135240 -147500
rect 135420 -147700 135440 -147500
rect 135220 -148100 135440 -147700
rect 138220 -147500 138440 -147490
rect 138220 -147700 138240 -147500
rect 138420 -147700 138440 -147500
rect 138220 -148100 138440 -147700
rect 141220 -147500 141440 -147490
rect 141220 -147700 141240 -147500
rect 141420 -147700 141440 -147500
rect 141220 -148100 141440 -147700
rect 144220 -147500 144440 -147490
rect 144220 -147700 144240 -147500
rect 144420 -147700 144440 -147500
rect 144220 -148100 144440 -147700
rect 147220 -147500 147440 -147490
rect 147220 -147700 147240 -147500
rect 147420 -147700 147440 -147500
rect 147220 -148100 147440 -147700
<< metal5 >>
rect -2000 2840 0 3160
rect 1040 1040 1240 1240
rect 4040 1040 4240 1240
rect 7040 1040 7240 1240
rect 10040 1040 10240 1240
rect 13040 1040 13240 1240
rect 16040 1040 16240 1240
rect 19040 1040 19240 1240
rect 22040 1040 22240 1240
rect 25040 1040 25240 1240
rect 28040 1040 28240 1240
rect 31040 1040 31240 1240
rect 34040 1040 34240 1240
rect 37040 1040 37240 1240
rect 40040 1040 40240 1240
rect 43040 1040 43240 1240
rect 46040 1040 46240 1240
rect 49040 1040 49240 1240
rect 52040 1040 52240 1240
rect 55040 1040 55240 1240
rect 58040 1040 58240 1240
rect 61040 1040 61240 1240
rect 64040 1040 64240 1240
rect 67040 1040 67240 1240
rect 70040 1040 70240 1240
rect 73040 1040 73240 1240
rect 76040 1040 76240 1240
rect 79040 1040 79240 1240
rect 82040 1040 82240 1240
rect 85040 1040 85240 1240
rect 88040 1040 88240 1240
rect 91040 1040 91240 1240
rect 94040 1040 94240 1240
rect 97040 1040 97240 1240
rect 100040 1040 100240 1240
rect 103040 1040 103240 1240
rect 106040 1040 106240 1240
rect 109040 1040 109240 1240
rect 112040 1040 112240 1240
rect 115040 1040 115240 1240
rect 118040 1040 118240 1240
rect 121040 1040 121240 1240
rect 124040 1040 124240 1240
rect 127040 1040 127240 1240
rect 130040 1040 130240 1240
rect 133040 1040 133240 1240
rect 136040 1040 136240 1240
rect 139040 1040 139240 1240
rect 142040 1040 142240 1240
rect 145040 1040 145240 1240
rect 148040 1040 148240 1240
rect 1040 -1960 1240 -1760
rect 4040 -1960 4240 -1760
rect 7040 -1960 7240 -1760
rect 10040 -1960 10240 -1760
rect 13040 -1960 13240 -1760
rect 16040 -1960 16240 -1760
rect 19040 -1960 19240 -1760
rect 22040 -1960 22240 -1760
rect 25040 -1960 25240 -1760
rect 28040 -1960 28240 -1760
rect 31040 -1960 31240 -1760
rect 34040 -1960 34240 -1760
rect 37040 -1960 37240 -1760
rect 40040 -1960 40240 -1760
rect 43040 -1960 43240 -1760
rect 46040 -1960 46240 -1760
rect 49040 -1960 49240 -1760
rect 52040 -1960 52240 -1760
rect 55040 -1960 55240 -1760
rect 58040 -1960 58240 -1760
rect 61040 -1960 61240 -1760
rect 64040 -1960 64240 -1760
rect 67040 -1960 67240 -1760
rect 70040 -1960 70240 -1760
rect 73040 -1960 73240 -1760
rect 76040 -1960 76240 -1760
rect 79040 -1960 79240 -1760
rect 82040 -1960 82240 -1760
rect 85040 -1960 85240 -1760
rect 88040 -1960 88240 -1760
rect 91040 -1960 91240 -1760
rect 94040 -1960 94240 -1760
rect 97040 -1960 97240 -1760
rect 100040 -1960 100240 -1760
rect 103040 -1960 103240 -1760
rect 106040 -1960 106240 -1760
rect 109040 -1960 109240 -1760
rect 112040 -1960 112240 -1760
rect 115040 -1960 115240 -1760
rect 118040 -1960 118240 -1760
rect 121040 -1960 121240 -1760
rect 124040 -1960 124240 -1760
rect 127040 -1960 127240 -1760
rect 130040 -1960 130240 -1760
rect 133040 -1960 133240 -1760
rect 136040 -1960 136240 -1760
rect 139040 -1960 139240 -1760
rect 142040 -1960 142240 -1760
rect 145040 -1960 145240 -1760
rect 148040 -1960 148240 -1760
rect 1040 -4960 1240 -4760
rect 4040 -4960 4240 -4760
rect 7040 -4960 7240 -4760
rect 10040 -4960 10240 -4760
rect 13040 -4960 13240 -4760
rect 16040 -4960 16240 -4760
rect 19040 -4960 19240 -4760
rect 22040 -4960 22240 -4760
rect 25040 -4960 25240 -4760
rect 28040 -4960 28240 -4760
rect 31040 -4960 31240 -4760
rect 34040 -4960 34240 -4760
rect 37040 -4960 37240 -4760
rect 40040 -4960 40240 -4760
rect 43040 -4960 43240 -4760
rect 46040 -4960 46240 -4760
rect 49040 -4960 49240 -4760
rect 52040 -4960 52240 -4760
rect 55040 -4960 55240 -4760
rect 58040 -4960 58240 -4760
rect 61040 -4960 61240 -4760
rect 64040 -4960 64240 -4760
rect 67040 -4960 67240 -4760
rect 70040 -4960 70240 -4760
rect 73040 -4960 73240 -4760
rect 76040 -4960 76240 -4760
rect 79040 -4960 79240 -4760
rect 82040 -4960 82240 -4760
rect 85040 -4960 85240 -4760
rect 88040 -4960 88240 -4760
rect 91040 -4960 91240 -4760
rect 94040 -4960 94240 -4760
rect 97040 -4960 97240 -4760
rect 100040 -4960 100240 -4760
rect 103040 -4960 103240 -4760
rect 106040 -4960 106240 -4760
rect 109040 -4960 109240 -4760
rect 112040 -4960 112240 -4760
rect 115040 -4960 115240 -4760
rect 118040 -4960 118240 -4760
rect 121040 -4960 121240 -4760
rect 124040 -4960 124240 -4760
rect 127040 -4960 127240 -4760
rect 130040 -4960 130240 -4760
rect 133040 -4960 133240 -4760
rect 136040 -4960 136240 -4760
rect 139040 -4960 139240 -4760
rect 142040 -4960 142240 -4760
rect 145040 -4960 145240 -4760
rect 148040 -4960 148240 -4760
rect 1040 -7960 1240 -7760
rect 4040 -7960 4240 -7760
rect 7040 -7960 7240 -7760
rect 10040 -7960 10240 -7760
rect 13040 -7960 13240 -7760
rect 16040 -7960 16240 -7760
rect 19040 -7960 19240 -7760
rect 22040 -7960 22240 -7760
rect 25040 -7960 25240 -7760
rect 28040 -7960 28240 -7760
rect 31040 -7960 31240 -7760
rect 34040 -7960 34240 -7760
rect 37040 -7960 37240 -7760
rect 40040 -7960 40240 -7760
rect 43040 -7960 43240 -7760
rect 46040 -7960 46240 -7760
rect 49040 -7960 49240 -7760
rect 52040 -7960 52240 -7760
rect 55040 -7960 55240 -7760
rect 58040 -7960 58240 -7760
rect 61040 -7960 61240 -7760
rect 64040 -7960 64240 -7760
rect 67040 -7960 67240 -7760
rect 70040 -7960 70240 -7760
rect 73040 -7960 73240 -7760
rect 76040 -7960 76240 -7760
rect 79040 -7960 79240 -7760
rect 82040 -7960 82240 -7760
rect 85040 -7960 85240 -7760
rect 88040 -7960 88240 -7760
rect 91040 -7960 91240 -7760
rect 94040 -7960 94240 -7760
rect 97040 -7960 97240 -7760
rect 100040 -7960 100240 -7760
rect 103040 -7960 103240 -7760
rect 106040 -7960 106240 -7760
rect 109040 -7960 109240 -7760
rect 112040 -7960 112240 -7760
rect 115040 -7960 115240 -7760
rect 118040 -7960 118240 -7760
rect 121040 -7960 121240 -7760
rect 124040 -7960 124240 -7760
rect 127040 -7960 127240 -7760
rect 130040 -7960 130240 -7760
rect 133040 -7960 133240 -7760
rect 136040 -7960 136240 -7760
rect 139040 -7960 139240 -7760
rect 142040 -7960 142240 -7760
rect 145040 -7960 145240 -7760
rect 148040 -7960 148240 -7760
rect 1040 -10960 1240 -10760
rect 4040 -10960 4240 -10760
rect 7040 -10960 7240 -10760
rect 10040 -10960 10240 -10760
rect 13040 -10960 13240 -10760
rect 16040 -10960 16240 -10760
rect 19040 -10960 19240 -10760
rect 22040 -10960 22240 -10760
rect 25040 -10960 25240 -10760
rect 28040 -10960 28240 -10760
rect 31040 -10960 31240 -10760
rect 34040 -10960 34240 -10760
rect 37040 -10960 37240 -10760
rect 40040 -10960 40240 -10760
rect 43040 -10960 43240 -10760
rect 46040 -10960 46240 -10760
rect 49040 -10960 49240 -10760
rect 52040 -10960 52240 -10760
rect 55040 -10960 55240 -10760
rect 58040 -10960 58240 -10760
rect 61040 -10960 61240 -10760
rect 64040 -10960 64240 -10760
rect 67040 -10960 67240 -10760
rect 70040 -10960 70240 -10760
rect 73040 -10960 73240 -10760
rect 76040 -10960 76240 -10760
rect 79040 -10960 79240 -10760
rect 82040 -10960 82240 -10760
rect 85040 -10960 85240 -10760
rect 88040 -10960 88240 -10760
rect 91040 -10960 91240 -10760
rect 94040 -10960 94240 -10760
rect 97040 -10960 97240 -10760
rect 100040 -10960 100240 -10760
rect 103040 -10960 103240 -10760
rect 106040 -10960 106240 -10760
rect 109040 -10960 109240 -10760
rect 112040 -10960 112240 -10760
rect 115040 -10960 115240 -10760
rect 118040 -10960 118240 -10760
rect 121040 -10960 121240 -10760
rect 124040 -10960 124240 -10760
rect 127040 -10960 127240 -10760
rect 130040 -10960 130240 -10760
rect 133040 -10960 133240 -10760
rect 136040 -10960 136240 -10760
rect 139040 -10960 139240 -10760
rect 142040 -10960 142240 -10760
rect 145040 -10960 145240 -10760
rect 148040 -10960 148240 -10760
rect 1040 -13960 1240 -13760
rect 4040 -13960 4240 -13760
rect 7040 -13960 7240 -13760
rect 10040 -13960 10240 -13760
rect 13040 -13960 13240 -13760
rect 16040 -13960 16240 -13760
rect 19040 -13960 19240 -13760
rect 22040 -13960 22240 -13760
rect 25040 -13960 25240 -13760
rect 28040 -13960 28240 -13760
rect 31040 -13960 31240 -13760
rect 34040 -13960 34240 -13760
rect 37040 -13960 37240 -13760
rect 40040 -13960 40240 -13760
rect 43040 -13960 43240 -13760
rect 46040 -13960 46240 -13760
rect 49040 -13960 49240 -13760
rect 52040 -13960 52240 -13760
rect 55040 -13960 55240 -13760
rect 58040 -13960 58240 -13760
rect 61040 -13960 61240 -13760
rect 64040 -13960 64240 -13760
rect 67040 -13960 67240 -13760
rect 70040 -13960 70240 -13760
rect 73040 -13960 73240 -13760
rect 76040 -13960 76240 -13760
rect 79040 -13960 79240 -13760
rect 82040 -13960 82240 -13760
rect 85040 -13960 85240 -13760
rect 88040 -13960 88240 -13760
rect 91040 -13960 91240 -13760
rect 94040 -13960 94240 -13760
rect 97040 -13960 97240 -13760
rect 100040 -13960 100240 -13760
rect 103040 -13960 103240 -13760
rect 106040 -13960 106240 -13760
rect 109040 -13960 109240 -13760
rect 112040 -13960 112240 -13760
rect 115040 -13960 115240 -13760
rect 118040 -13960 118240 -13760
rect 121040 -13960 121240 -13760
rect 124040 -13960 124240 -13760
rect 127040 -13960 127240 -13760
rect 130040 -13960 130240 -13760
rect 133040 -13960 133240 -13760
rect 136040 -13960 136240 -13760
rect 139040 -13960 139240 -13760
rect 142040 -13960 142240 -13760
rect 145040 -13960 145240 -13760
rect 148040 -13960 148240 -13760
rect 1040 -16960 1240 -16760
rect 4040 -16960 4240 -16760
rect 7040 -16960 7240 -16760
rect 10040 -16960 10240 -16760
rect 13040 -16960 13240 -16760
rect 16040 -16960 16240 -16760
rect 19040 -16960 19240 -16760
rect 22040 -16960 22240 -16760
rect 25040 -16960 25240 -16760
rect 28040 -16960 28240 -16760
rect 31040 -16960 31240 -16760
rect 34040 -16960 34240 -16760
rect 37040 -16960 37240 -16760
rect 40040 -16960 40240 -16760
rect 43040 -16960 43240 -16760
rect 46040 -16960 46240 -16760
rect 49040 -16960 49240 -16760
rect 52040 -16960 52240 -16760
rect 55040 -16960 55240 -16760
rect 58040 -16960 58240 -16760
rect 61040 -16960 61240 -16760
rect 64040 -16960 64240 -16760
rect 67040 -16960 67240 -16760
rect 70040 -16960 70240 -16760
rect 73040 -16960 73240 -16760
rect 76040 -16960 76240 -16760
rect 79040 -16960 79240 -16760
rect 82040 -16960 82240 -16760
rect 85040 -16960 85240 -16760
rect 88040 -16960 88240 -16760
rect 91040 -16960 91240 -16760
rect 94040 -16960 94240 -16760
rect 97040 -16960 97240 -16760
rect 100040 -16960 100240 -16760
rect 103040 -16960 103240 -16760
rect 106040 -16960 106240 -16760
rect 109040 -16960 109240 -16760
rect 112040 -16960 112240 -16760
rect 115040 -16960 115240 -16760
rect 118040 -16960 118240 -16760
rect 121040 -16960 121240 -16760
rect 124040 -16960 124240 -16760
rect 127040 -16960 127240 -16760
rect 130040 -16960 130240 -16760
rect 133040 -16960 133240 -16760
rect 136040 -16960 136240 -16760
rect 139040 -16960 139240 -16760
rect 142040 -16960 142240 -16760
rect 145040 -16960 145240 -16760
rect 148040 -16960 148240 -16760
rect 1040 -19960 1240 -19760
rect 4040 -19960 4240 -19760
rect 7040 -19960 7240 -19760
rect 10040 -19960 10240 -19760
rect 13040 -19960 13240 -19760
rect 16040 -19960 16240 -19760
rect 19040 -19960 19240 -19760
rect 22040 -19960 22240 -19760
rect 25040 -19960 25240 -19760
rect 28040 -19960 28240 -19760
rect 31040 -19960 31240 -19760
rect 34040 -19960 34240 -19760
rect 37040 -19960 37240 -19760
rect 40040 -19960 40240 -19760
rect 43040 -19960 43240 -19760
rect 46040 -19960 46240 -19760
rect 49040 -19960 49240 -19760
rect 52040 -19960 52240 -19760
rect 55040 -19960 55240 -19760
rect 58040 -19960 58240 -19760
rect 61040 -19960 61240 -19760
rect 64040 -19960 64240 -19760
rect 67040 -19960 67240 -19760
rect 70040 -19960 70240 -19760
rect 73040 -19960 73240 -19760
rect 76040 -19960 76240 -19760
rect 79040 -19960 79240 -19760
rect 82040 -19960 82240 -19760
rect 85040 -19960 85240 -19760
rect 88040 -19960 88240 -19760
rect 91040 -19960 91240 -19760
rect 94040 -19960 94240 -19760
rect 97040 -19960 97240 -19760
rect 100040 -19960 100240 -19760
rect 103040 -19960 103240 -19760
rect 106040 -19960 106240 -19760
rect 109040 -19960 109240 -19760
rect 112040 -19960 112240 -19760
rect 115040 -19960 115240 -19760
rect 118040 -19960 118240 -19760
rect 121040 -19960 121240 -19760
rect 124040 -19960 124240 -19760
rect 127040 -19960 127240 -19760
rect 130040 -19960 130240 -19760
rect 133040 -19960 133240 -19760
rect 136040 -19960 136240 -19760
rect 139040 -19960 139240 -19760
rect 142040 -19960 142240 -19760
rect 145040 -19960 145240 -19760
rect 148040 -19960 148240 -19760
rect 1040 -22960 1240 -22760
rect 4040 -22960 4240 -22760
rect 7040 -22960 7240 -22760
rect 10040 -22960 10240 -22760
rect 13040 -22960 13240 -22760
rect 16040 -22960 16240 -22760
rect 19040 -22960 19240 -22760
rect 22040 -22960 22240 -22760
rect 25040 -22960 25240 -22760
rect 28040 -22960 28240 -22760
rect 31040 -22960 31240 -22760
rect 34040 -22960 34240 -22760
rect 37040 -22960 37240 -22760
rect 40040 -22960 40240 -22760
rect 43040 -22960 43240 -22760
rect 46040 -22960 46240 -22760
rect 49040 -22960 49240 -22760
rect 52040 -22960 52240 -22760
rect 55040 -22960 55240 -22760
rect 58040 -22960 58240 -22760
rect 61040 -22960 61240 -22760
rect 64040 -22960 64240 -22760
rect 67040 -22960 67240 -22760
rect 70040 -22960 70240 -22760
rect 73040 -22960 73240 -22760
rect 76040 -22960 76240 -22760
rect 79040 -22960 79240 -22760
rect 82040 -22960 82240 -22760
rect 85040 -22960 85240 -22760
rect 88040 -22960 88240 -22760
rect 91040 -22960 91240 -22760
rect 94040 -22960 94240 -22760
rect 97040 -22960 97240 -22760
rect 100040 -22960 100240 -22760
rect 103040 -22960 103240 -22760
rect 106040 -22960 106240 -22760
rect 109040 -22960 109240 -22760
rect 112040 -22960 112240 -22760
rect 115040 -22960 115240 -22760
rect 118040 -22960 118240 -22760
rect 121040 -22960 121240 -22760
rect 124040 -22960 124240 -22760
rect 127040 -22960 127240 -22760
rect 130040 -22960 130240 -22760
rect 133040 -22960 133240 -22760
rect 136040 -22960 136240 -22760
rect 139040 -22960 139240 -22760
rect 142040 -22960 142240 -22760
rect 145040 -22960 145240 -22760
rect 148040 -22960 148240 -22760
rect 1040 -25960 1240 -25760
rect 4040 -25960 4240 -25760
rect 7040 -25960 7240 -25760
rect 10040 -25960 10240 -25760
rect 13040 -25960 13240 -25760
rect 16040 -25960 16240 -25760
rect 19040 -25960 19240 -25760
rect 22040 -25960 22240 -25760
rect 25040 -25960 25240 -25760
rect 28040 -25960 28240 -25760
rect 31040 -25960 31240 -25760
rect 34040 -25960 34240 -25760
rect 37040 -25960 37240 -25760
rect 40040 -25960 40240 -25760
rect 43040 -25960 43240 -25760
rect 46040 -25960 46240 -25760
rect 49040 -25960 49240 -25760
rect 52040 -25960 52240 -25760
rect 55040 -25960 55240 -25760
rect 58040 -25960 58240 -25760
rect 61040 -25960 61240 -25760
rect 64040 -25960 64240 -25760
rect 67040 -25960 67240 -25760
rect 70040 -25960 70240 -25760
rect 73040 -25960 73240 -25760
rect 76040 -25960 76240 -25760
rect 79040 -25960 79240 -25760
rect 82040 -25960 82240 -25760
rect 85040 -25960 85240 -25760
rect 88040 -25960 88240 -25760
rect 91040 -25960 91240 -25760
rect 94040 -25960 94240 -25760
rect 97040 -25960 97240 -25760
rect 100040 -25960 100240 -25760
rect 103040 -25960 103240 -25760
rect 106040 -25960 106240 -25760
rect 109040 -25960 109240 -25760
rect 112040 -25960 112240 -25760
rect 115040 -25960 115240 -25760
rect 118040 -25960 118240 -25760
rect 121040 -25960 121240 -25760
rect 124040 -25960 124240 -25760
rect 127040 -25960 127240 -25760
rect 130040 -25960 130240 -25760
rect 133040 -25960 133240 -25760
rect 136040 -25960 136240 -25760
rect 139040 -25960 139240 -25760
rect 142040 -25960 142240 -25760
rect 145040 -25960 145240 -25760
rect 148040 -25960 148240 -25760
rect 1040 -28960 1240 -28760
rect 4040 -28960 4240 -28760
rect 7040 -28960 7240 -28760
rect 10040 -28960 10240 -28760
rect 13040 -28960 13240 -28760
rect 16040 -28960 16240 -28760
rect 19040 -28960 19240 -28760
rect 22040 -28960 22240 -28760
rect 25040 -28960 25240 -28760
rect 28040 -28960 28240 -28760
rect 31040 -28960 31240 -28760
rect 34040 -28960 34240 -28760
rect 37040 -28960 37240 -28760
rect 40040 -28960 40240 -28760
rect 43040 -28960 43240 -28760
rect 46040 -28960 46240 -28760
rect 49040 -28960 49240 -28760
rect 52040 -28960 52240 -28760
rect 55040 -28960 55240 -28760
rect 58040 -28960 58240 -28760
rect 61040 -28960 61240 -28760
rect 64040 -28960 64240 -28760
rect 67040 -28960 67240 -28760
rect 70040 -28960 70240 -28760
rect 73040 -28960 73240 -28760
rect 76040 -28960 76240 -28760
rect 79040 -28960 79240 -28760
rect 82040 -28960 82240 -28760
rect 85040 -28960 85240 -28760
rect 88040 -28960 88240 -28760
rect 91040 -28960 91240 -28760
rect 94040 -28960 94240 -28760
rect 97040 -28960 97240 -28760
rect 100040 -28960 100240 -28760
rect 103040 -28960 103240 -28760
rect 106040 -28960 106240 -28760
rect 109040 -28960 109240 -28760
rect 112040 -28960 112240 -28760
rect 115040 -28960 115240 -28760
rect 118040 -28960 118240 -28760
rect 121040 -28960 121240 -28760
rect 124040 -28960 124240 -28760
rect 127040 -28960 127240 -28760
rect 130040 -28960 130240 -28760
rect 133040 -28960 133240 -28760
rect 136040 -28960 136240 -28760
rect 139040 -28960 139240 -28760
rect 142040 -28960 142240 -28760
rect 145040 -28960 145240 -28760
rect 148040 -28960 148240 -28760
rect 1040 -31960 1240 -31760
rect 4040 -31960 4240 -31760
rect 7040 -31960 7240 -31760
rect 10040 -31960 10240 -31760
rect 13040 -31960 13240 -31760
rect 16040 -31960 16240 -31760
rect 19040 -31960 19240 -31760
rect 22040 -31960 22240 -31760
rect 25040 -31960 25240 -31760
rect 28040 -31960 28240 -31760
rect 31040 -31960 31240 -31760
rect 34040 -31960 34240 -31760
rect 37040 -31960 37240 -31760
rect 40040 -31960 40240 -31760
rect 43040 -31960 43240 -31760
rect 46040 -31960 46240 -31760
rect 49040 -31960 49240 -31760
rect 52040 -31960 52240 -31760
rect 55040 -31960 55240 -31760
rect 58040 -31960 58240 -31760
rect 61040 -31960 61240 -31760
rect 64040 -31960 64240 -31760
rect 67040 -31960 67240 -31760
rect 70040 -31960 70240 -31760
rect 73040 -31960 73240 -31760
rect 76040 -31960 76240 -31760
rect 79040 -31960 79240 -31760
rect 82040 -31960 82240 -31760
rect 85040 -31960 85240 -31760
rect 88040 -31960 88240 -31760
rect 91040 -31960 91240 -31760
rect 94040 -31960 94240 -31760
rect 97040 -31960 97240 -31760
rect 100040 -31960 100240 -31760
rect 103040 -31960 103240 -31760
rect 106040 -31960 106240 -31760
rect 109040 -31960 109240 -31760
rect 112040 -31960 112240 -31760
rect 115040 -31960 115240 -31760
rect 118040 -31960 118240 -31760
rect 121040 -31960 121240 -31760
rect 124040 -31960 124240 -31760
rect 127040 -31960 127240 -31760
rect 130040 -31960 130240 -31760
rect 133040 -31960 133240 -31760
rect 136040 -31960 136240 -31760
rect 139040 -31960 139240 -31760
rect 142040 -31960 142240 -31760
rect 145040 -31960 145240 -31760
rect 148040 -31960 148240 -31760
rect 1040 -34960 1240 -34760
rect 4040 -34960 4240 -34760
rect 7040 -34960 7240 -34760
rect 10040 -34960 10240 -34760
rect 13040 -34960 13240 -34760
rect 16040 -34960 16240 -34760
rect 19040 -34960 19240 -34760
rect 22040 -34960 22240 -34760
rect 25040 -34960 25240 -34760
rect 28040 -34960 28240 -34760
rect 31040 -34960 31240 -34760
rect 34040 -34960 34240 -34760
rect 37040 -34960 37240 -34760
rect 40040 -34960 40240 -34760
rect 43040 -34960 43240 -34760
rect 46040 -34960 46240 -34760
rect 49040 -34960 49240 -34760
rect 52040 -34960 52240 -34760
rect 55040 -34960 55240 -34760
rect 58040 -34960 58240 -34760
rect 61040 -34960 61240 -34760
rect 64040 -34960 64240 -34760
rect 67040 -34960 67240 -34760
rect 70040 -34960 70240 -34760
rect 73040 -34960 73240 -34760
rect 76040 -34960 76240 -34760
rect 79040 -34960 79240 -34760
rect 82040 -34960 82240 -34760
rect 85040 -34960 85240 -34760
rect 88040 -34960 88240 -34760
rect 91040 -34960 91240 -34760
rect 94040 -34960 94240 -34760
rect 97040 -34960 97240 -34760
rect 100040 -34960 100240 -34760
rect 103040 -34960 103240 -34760
rect 106040 -34960 106240 -34760
rect 109040 -34960 109240 -34760
rect 112040 -34960 112240 -34760
rect 115040 -34960 115240 -34760
rect 118040 -34960 118240 -34760
rect 121040 -34960 121240 -34760
rect 124040 -34960 124240 -34760
rect 127040 -34960 127240 -34760
rect 130040 -34960 130240 -34760
rect 133040 -34960 133240 -34760
rect 136040 -34960 136240 -34760
rect 139040 -34960 139240 -34760
rect 142040 -34960 142240 -34760
rect 145040 -34960 145240 -34760
rect 148040 -34960 148240 -34760
rect 1040 -37960 1240 -37760
rect 4040 -37960 4240 -37760
rect 7040 -37960 7240 -37760
rect 10040 -37960 10240 -37760
rect 13040 -37960 13240 -37760
rect 16040 -37960 16240 -37760
rect 19040 -37960 19240 -37760
rect 22040 -37960 22240 -37760
rect 25040 -37960 25240 -37760
rect 28040 -37960 28240 -37760
rect 31040 -37960 31240 -37760
rect 34040 -37960 34240 -37760
rect 37040 -37960 37240 -37760
rect 40040 -37960 40240 -37760
rect 43040 -37960 43240 -37760
rect 46040 -37960 46240 -37760
rect 49040 -37960 49240 -37760
rect 52040 -37960 52240 -37760
rect 55040 -37960 55240 -37760
rect 58040 -37960 58240 -37760
rect 61040 -37960 61240 -37760
rect 64040 -37960 64240 -37760
rect 67040 -37960 67240 -37760
rect 70040 -37960 70240 -37760
rect 73040 -37960 73240 -37760
rect 76040 -37960 76240 -37760
rect 79040 -37960 79240 -37760
rect 82040 -37960 82240 -37760
rect 85040 -37960 85240 -37760
rect 88040 -37960 88240 -37760
rect 91040 -37960 91240 -37760
rect 94040 -37960 94240 -37760
rect 97040 -37960 97240 -37760
rect 100040 -37960 100240 -37760
rect 103040 -37960 103240 -37760
rect 106040 -37960 106240 -37760
rect 109040 -37960 109240 -37760
rect 112040 -37960 112240 -37760
rect 115040 -37960 115240 -37760
rect 118040 -37960 118240 -37760
rect 121040 -37960 121240 -37760
rect 124040 -37960 124240 -37760
rect 127040 -37960 127240 -37760
rect 130040 -37960 130240 -37760
rect 133040 -37960 133240 -37760
rect 136040 -37960 136240 -37760
rect 139040 -37960 139240 -37760
rect 142040 -37960 142240 -37760
rect 145040 -37960 145240 -37760
rect 148040 -37960 148240 -37760
rect 1040 -40960 1240 -40760
rect 4040 -40960 4240 -40760
rect 7040 -40960 7240 -40760
rect 10040 -40960 10240 -40760
rect 13040 -40960 13240 -40760
rect 16040 -40960 16240 -40760
rect 19040 -40960 19240 -40760
rect 22040 -40960 22240 -40760
rect 25040 -40960 25240 -40760
rect 28040 -40960 28240 -40760
rect 31040 -40960 31240 -40760
rect 34040 -40960 34240 -40760
rect 37040 -40960 37240 -40760
rect 40040 -40960 40240 -40760
rect 43040 -40960 43240 -40760
rect 46040 -40960 46240 -40760
rect 49040 -40960 49240 -40760
rect 52040 -40960 52240 -40760
rect 55040 -40960 55240 -40760
rect 58040 -40960 58240 -40760
rect 61040 -40960 61240 -40760
rect 64040 -40960 64240 -40760
rect 67040 -40960 67240 -40760
rect 70040 -40960 70240 -40760
rect 73040 -40960 73240 -40760
rect 76040 -40960 76240 -40760
rect 79040 -40960 79240 -40760
rect 82040 -40960 82240 -40760
rect 85040 -40960 85240 -40760
rect 88040 -40960 88240 -40760
rect 91040 -40960 91240 -40760
rect 94040 -40960 94240 -40760
rect 97040 -40960 97240 -40760
rect 100040 -40960 100240 -40760
rect 103040 -40960 103240 -40760
rect 106040 -40960 106240 -40760
rect 109040 -40960 109240 -40760
rect 112040 -40960 112240 -40760
rect 115040 -40960 115240 -40760
rect 118040 -40960 118240 -40760
rect 121040 -40960 121240 -40760
rect 124040 -40960 124240 -40760
rect 127040 -40960 127240 -40760
rect 130040 -40960 130240 -40760
rect 133040 -40960 133240 -40760
rect 136040 -40960 136240 -40760
rect 139040 -40960 139240 -40760
rect 142040 -40960 142240 -40760
rect 145040 -40960 145240 -40760
rect 148040 -40960 148240 -40760
rect 1040 -43960 1240 -43760
rect 4040 -43960 4240 -43760
rect 7040 -43960 7240 -43760
rect 10040 -43960 10240 -43760
rect 13040 -43960 13240 -43760
rect 16040 -43960 16240 -43760
rect 19040 -43960 19240 -43760
rect 22040 -43960 22240 -43760
rect 25040 -43960 25240 -43760
rect 28040 -43960 28240 -43760
rect 31040 -43960 31240 -43760
rect 34040 -43960 34240 -43760
rect 37040 -43960 37240 -43760
rect 40040 -43960 40240 -43760
rect 43040 -43960 43240 -43760
rect 46040 -43960 46240 -43760
rect 49040 -43960 49240 -43760
rect 52040 -43960 52240 -43760
rect 55040 -43960 55240 -43760
rect 58040 -43960 58240 -43760
rect 61040 -43960 61240 -43760
rect 64040 -43960 64240 -43760
rect 67040 -43960 67240 -43760
rect 70040 -43960 70240 -43760
rect 73040 -43960 73240 -43760
rect 76040 -43960 76240 -43760
rect 79040 -43960 79240 -43760
rect 82040 -43960 82240 -43760
rect 85040 -43960 85240 -43760
rect 88040 -43960 88240 -43760
rect 91040 -43960 91240 -43760
rect 94040 -43960 94240 -43760
rect 97040 -43960 97240 -43760
rect 100040 -43960 100240 -43760
rect 103040 -43960 103240 -43760
rect 106040 -43960 106240 -43760
rect 109040 -43960 109240 -43760
rect 112040 -43960 112240 -43760
rect 115040 -43960 115240 -43760
rect 118040 -43960 118240 -43760
rect 121040 -43960 121240 -43760
rect 124040 -43960 124240 -43760
rect 127040 -43960 127240 -43760
rect 130040 -43960 130240 -43760
rect 133040 -43960 133240 -43760
rect 136040 -43960 136240 -43760
rect 139040 -43960 139240 -43760
rect 142040 -43960 142240 -43760
rect 145040 -43960 145240 -43760
rect 148040 -43960 148240 -43760
rect 1040 -46960 1240 -46760
rect 4040 -46960 4240 -46760
rect 7040 -46960 7240 -46760
rect 10040 -46960 10240 -46760
rect 13040 -46960 13240 -46760
rect 16040 -46960 16240 -46760
rect 19040 -46960 19240 -46760
rect 22040 -46960 22240 -46760
rect 25040 -46960 25240 -46760
rect 28040 -46960 28240 -46760
rect 31040 -46960 31240 -46760
rect 34040 -46960 34240 -46760
rect 37040 -46960 37240 -46760
rect 40040 -46960 40240 -46760
rect 43040 -46960 43240 -46760
rect 46040 -46960 46240 -46760
rect 49040 -46960 49240 -46760
rect 52040 -46960 52240 -46760
rect 55040 -46960 55240 -46760
rect 58040 -46960 58240 -46760
rect 61040 -46960 61240 -46760
rect 64040 -46960 64240 -46760
rect 67040 -46960 67240 -46760
rect 70040 -46960 70240 -46760
rect 73040 -46960 73240 -46760
rect 76040 -46960 76240 -46760
rect 79040 -46960 79240 -46760
rect 82040 -46960 82240 -46760
rect 85040 -46960 85240 -46760
rect 88040 -46960 88240 -46760
rect 91040 -46960 91240 -46760
rect 94040 -46960 94240 -46760
rect 97040 -46960 97240 -46760
rect 100040 -46960 100240 -46760
rect 103040 -46960 103240 -46760
rect 106040 -46960 106240 -46760
rect 109040 -46960 109240 -46760
rect 112040 -46960 112240 -46760
rect 115040 -46960 115240 -46760
rect 118040 -46960 118240 -46760
rect 121040 -46960 121240 -46760
rect 124040 -46960 124240 -46760
rect 127040 -46960 127240 -46760
rect 130040 -46960 130240 -46760
rect 133040 -46960 133240 -46760
rect 136040 -46960 136240 -46760
rect 139040 -46960 139240 -46760
rect 142040 -46960 142240 -46760
rect 145040 -46960 145240 -46760
rect 148040 -46960 148240 -46760
rect 1040 -49960 1240 -49760
rect 4040 -49960 4240 -49760
rect 7040 -49960 7240 -49760
rect 10040 -49960 10240 -49760
rect 13040 -49960 13240 -49760
rect 16040 -49960 16240 -49760
rect 19040 -49960 19240 -49760
rect 22040 -49960 22240 -49760
rect 25040 -49960 25240 -49760
rect 28040 -49960 28240 -49760
rect 31040 -49960 31240 -49760
rect 34040 -49960 34240 -49760
rect 37040 -49960 37240 -49760
rect 40040 -49960 40240 -49760
rect 43040 -49960 43240 -49760
rect 46040 -49960 46240 -49760
rect 49040 -49960 49240 -49760
rect 52040 -49960 52240 -49760
rect 55040 -49960 55240 -49760
rect 58040 -49960 58240 -49760
rect 61040 -49960 61240 -49760
rect 64040 -49960 64240 -49760
rect 67040 -49960 67240 -49760
rect 70040 -49960 70240 -49760
rect 73040 -49960 73240 -49760
rect 76040 -49960 76240 -49760
rect 79040 -49960 79240 -49760
rect 82040 -49960 82240 -49760
rect 85040 -49960 85240 -49760
rect 88040 -49960 88240 -49760
rect 91040 -49960 91240 -49760
rect 94040 -49960 94240 -49760
rect 97040 -49960 97240 -49760
rect 100040 -49960 100240 -49760
rect 103040 -49960 103240 -49760
rect 106040 -49960 106240 -49760
rect 109040 -49960 109240 -49760
rect 112040 -49960 112240 -49760
rect 115040 -49960 115240 -49760
rect 118040 -49960 118240 -49760
rect 121040 -49960 121240 -49760
rect 124040 -49960 124240 -49760
rect 127040 -49960 127240 -49760
rect 130040 -49960 130240 -49760
rect 133040 -49960 133240 -49760
rect 136040 -49960 136240 -49760
rect 139040 -49960 139240 -49760
rect 142040 -49960 142240 -49760
rect 145040 -49960 145240 -49760
rect 148040 -49960 148240 -49760
rect 1040 -52960 1240 -52760
rect 4040 -52960 4240 -52760
rect 7040 -52960 7240 -52760
rect 10040 -52960 10240 -52760
rect 13040 -52960 13240 -52760
rect 16040 -52960 16240 -52760
rect 19040 -52960 19240 -52760
rect 22040 -52960 22240 -52760
rect 25040 -52960 25240 -52760
rect 28040 -52960 28240 -52760
rect 31040 -52960 31240 -52760
rect 34040 -52960 34240 -52760
rect 37040 -52960 37240 -52760
rect 40040 -52960 40240 -52760
rect 43040 -52960 43240 -52760
rect 46040 -52960 46240 -52760
rect 49040 -52960 49240 -52760
rect 52040 -52960 52240 -52760
rect 55040 -52960 55240 -52760
rect 58040 -52960 58240 -52760
rect 61040 -52960 61240 -52760
rect 64040 -52960 64240 -52760
rect 67040 -52960 67240 -52760
rect 70040 -52960 70240 -52760
rect 73040 -52960 73240 -52760
rect 76040 -52960 76240 -52760
rect 79040 -52960 79240 -52760
rect 82040 -52960 82240 -52760
rect 85040 -52960 85240 -52760
rect 88040 -52960 88240 -52760
rect 91040 -52960 91240 -52760
rect 94040 -52960 94240 -52760
rect 97040 -52960 97240 -52760
rect 100040 -52960 100240 -52760
rect 103040 -52960 103240 -52760
rect 106040 -52960 106240 -52760
rect 109040 -52960 109240 -52760
rect 112040 -52960 112240 -52760
rect 115040 -52960 115240 -52760
rect 118040 -52960 118240 -52760
rect 121040 -52960 121240 -52760
rect 124040 -52960 124240 -52760
rect 127040 -52960 127240 -52760
rect 130040 -52960 130240 -52760
rect 133040 -52960 133240 -52760
rect 136040 -52960 136240 -52760
rect 139040 -52960 139240 -52760
rect 142040 -52960 142240 -52760
rect 145040 -52960 145240 -52760
rect 148040 -52960 148240 -52760
rect 1040 -55960 1240 -55760
rect 4040 -55960 4240 -55760
rect 7040 -55960 7240 -55760
rect 10040 -55960 10240 -55760
rect 13040 -55960 13240 -55760
rect 16040 -55960 16240 -55760
rect 19040 -55960 19240 -55760
rect 22040 -55960 22240 -55760
rect 25040 -55960 25240 -55760
rect 28040 -55960 28240 -55760
rect 31040 -55960 31240 -55760
rect 34040 -55960 34240 -55760
rect 37040 -55960 37240 -55760
rect 40040 -55960 40240 -55760
rect 43040 -55960 43240 -55760
rect 46040 -55960 46240 -55760
rect 49040 -55960 49240 -55760
rect 52040 -55960 52240 -55760
rect 55040 -55960 55240 -55760
rect 58040 -55960 58240 -55760
rect 61040 -55960 61240 -55760
rect 64040 -55960 64240 -55760
rect 67040 -55960 67240 -55760
rect 70040 -55960 70240 -55760
rect 73040 -55960 73240 -55760
rect 76040 -55960 76240 -55760
rect 79040 -55960 79240 -55760
rect 82040 -55960 82240 -55760
rect 85040 -55960 85240 -55760
rect 88040 -55960 88240 -55760
rect 91040 -55960 91240 -55760
rect 94040 -55960 94240 -55760
rect 97040 -55960 97240 -55760
rect 100040 -55960 100240 -55760
rect 103040 -55960 103240 -55760
rect 106040 -55960 106240 -55760
rect 109040 -55960 109240 -55760
rect 112040 -55960 112240 -55760
rect 115040 -55960 115240 -55760
rect 118040 -55960 118240 -55760
rect 121040 -55960 121240 -55760
rect 124040 -55960 124240 -55760
rect 127040 -55960 127240 -55760
rect 130040 -55960 130240 -55760
rect 133040 -55960 133240 -55760
rect 136040 -55960 136240 -55760
rect 139040 -55960 139240 -55760
rect 142040 -55960 142240 -55760
rect 145040 -55960 145240 -55760
rect 148040 -55960 148240 -55760
rect 1040 -58960 1240 -58760
rect 4040 -58960 4240 -58760
rect 7040 -58960 7240 -58760
rect 10040 -58960 10240 -58760
rect 13040 -58960 13240 -58760
rect 16040 -58960 16240 -58760
rect 19040 -58960 19240 -58760
rect 22040 -58960 22240 -58760
rect 25040 -58960 25240 -58760
rect 28040 -58960 28240 -58760
rect 31040 -58960 31240 -58760
rect 34040 -58960 34240 -58760
rect 37040 -58960 37240 -58760
rect 40040 -58960 40240 -58760
rect 43040 -58960 43240 -58760
rect 46040 -58960 46240 -58760
rect 49040 -58960 49240 -58760
rect 52040 -58960 52240 -58760
rect 55040 -58960 55240 -58760
rect 58040 -58960 58240 -58760
rect 61040 -58960 61240 -58760
rect 64040 -58960 64240 -58760
rect 67040 -58960 67240 -58760
rect 70040 -58960 70240 -58760
rect 73040 -58960 73240 -58760
rect 76040 -58960 76240 -58760
rect 79040 -58960 79240 -58760
rect 82040 -58960 82240 -58760
rect 85040 -58960 85240 -58760
rect 88040 -58960 88240 -58760
rect 91040 -58960 91240 -58760
rect 94040 -58960 94240 -58760
rect 97040 -58960 97240 -58760
rect 100040 -58960 100240 -58760
rect 103040 -58960 103240 -58760
rect 106040 -58960 106240 -58760
rect 109040 -58960 109240 -58760
rect 112040 -58960 112240 -58760
rect 115040 -58960 115240 -58760
rect 118040 -58960 118240 -58760
rect 121040 -58960 121240 -58760
rect 124040 -58960 124240 -58760
rect 127040 -58960 127240 -58760
rect 130040 -58960 130240 -58760
rect 133040 -58960 133240 -58760
rect 136040 -58960 136240 -58760
rect 139040 -58960 139240 -58760
rect 142040 -58960 142240 -58760
rect 145040 -58960 145240 -58760
rect 148040 -58960 148240 -58760
rect 1040 -61960 1240 -61760
rect 4040 -61960 4240 -61760
rect 7040 -61960 7240 -61760
rect 10040 -61960 10240 -61760
rect 13040 -61960 13240 -61760
rect 16040 -61960 16240 -61760
rect 19040 -61960 19240 -61760
rect 22040 -61960 22240 -61760
rect 25040 -61960 25240 -61760
rect 28040 -61960 28240 -61760
rect 31040 -61960 31240 -61760
rect 34040 -61960 34240 -61760
rect 37040 -61960 37240 -61760
rect 40040 -61960 40240 -61760
rect 43040 -61960 43240 -61760
rect 46040 -61960 46240 -61760
rect 49040 -61960 49240 -61760
rect 52040 -61960 52240 -61760
rect 55040 -61960 55240 -61760
rect 58040 -61960 58240 -61760
rect 61040 -61960 61240 -61760
rect 64040 -61960 64240 -61760
rect 67040 -61960 67240 -61760
rect 70040 -61960 70240 -61760
rect 73040 -61960 73240 -61760
rect 76040 -61960 76240 -61760
rect 79040 -61960 79240 -61760
rect 82040 -61960 82240 -61760
rect 85040 -61960 85240 -61760
rect 88040 -61960 88240 -61760
rect 91040 -61960 91240 -61760
rect 94040 -61960 94240 -61760
rect 97040 -61960 97240 -61760
rect 100040 -61960 100240 -61760
rect 103040 -61960 103240 -61760
rect 106040 -61960 106240 -61760
rect 109040 -61960 109240 -61760
rect 112040 -61960 112240 -61760
rect 115040 -61960 115240 -61760
rect 118040 -61960 118240 -61760
rect 121040 -61960 121240 -61760
rect 124040 -61960 124240 -61760
rect 127040 -61960 127240 -61760
rect 130040 -61960 130240 -61760
rect 133040 -61960 133240 -61760
rect 136040 -61960 136240 -61760
rect 139040 -61960 139240 -61760
rect 142040 -61960 142240 -61760
rect 145040 -61960 145240 -61760
rect 148040 -61960 148240 -61760
rect 1040 -64960 1240 -64760
rect 4040 -64960 4240 -64760
rect 7040 -64960 7240 -64760
rect 10040 -64960 10240 -64760
rect 13040 -64960 13240 -64760
rect 16040 -64960 16240 -64760
rect 19040 -64960 19240 -64760
rect 22040 -64960 22240 -64760
rect 25040 -64960 25240 -64760
rect 28040 -64960 28240 -64760
rect 31040 -64960 31240 -64760
rect 34040 -64960 34240 -64760
rect 37040 -64960 37240 -64760
rect 40040 -64960 40240 -64760
rect 43040 -64960 43240 -64760
rect 46040 -64960 46240 -64760
rect 49040 -64960 49240 -64760
rect 52040 -64960 52240 -64760
rect 55040 -64960 55240 -64760
rect 58040 -64960 58240 -64760
rect 61040 -64960 61240 -64760
rect 64040 -64960 64240 -64760
rect 67040 -64960 67240 -64760
rect 70040 -64960 70240 -64760
rect 73040 -64960 73240 -64760
rect 76040 -64960 76240 -64760
rect 79040 -64960 79240 -64760
rect 82040 -64960 82240 -64760
rect 85040 -64960 85240 -64760
rect 88040 -64960 88240 -64760
rect 91040 -64960 91240 -64760
rect 94040 -64960 94240 -64760
rect 97040 -64960 97240 -64760
rect 100040 -64960 100240 -64760
rect 103040 -64960 103240 -64760
rect 106040 -64960 106240 -64760
rect 109040 -64960 109240 -64760
rect 112040 -64960 112240 -64760
rect 115040 -64960 115240 -64760
rect 118040 -64960 118240 -64760
rect 121040 -64960 121240 -64760
rect 124040 -64960 124240 -64760
rect 127040 -64960 127240 -64760
rect 130040 -64960 130240 -64760
rect 133040 -64960 133240 -64760
rect 136040 -64960 136240 -64760
rect 139040 -64960 139240 -64760
rect 142040 -64960 142240 -64760
rect 145040 -64960 145240 -64760
rect 148040 -64960 148240 -64760
rect 1040 -67960 1240 -67760
rect 4040 -67960 4240 -67760
rect 7040 -67960 7240 -67760
rect 10040 -67960 10240 -67760
rect 13040 -67960 13240 -67760
rect 16040 -67960 16240 -67760
rect 19040 -67960 19240 -67760
rect 22040 -67960 22240 -67760
rect 25040 -67960 25240 -67760
rect 28040 -67960 28240 -67760
rect 31040 -67960 31240 -67760
rect 34040 -67960 34240 -67760
rect 37040 -67960 37240 -67760
rect 40040 -67960 40240 -67760
rect 43040 -67960 43240 -67760
rect 46040 -67960 46240 -67760
rect 49040 -67960 49240 -67760
rect 52040 -67960 52240 -67760
rect 55040 -67960 55240 -67760
rect 58040 -67960 58240 -67760
rect 61040 -67960 61240 -67760
rect 64040 -67960 64240 -67760
rect 67040 -67960 67240 -67760
rect 70040 -67960 70240 -67760
rect 73040 -67960 73240 -67760
rect 76040 -67960 76240 -67760
rect 79040 -67960 79240 -67760
rect 82040 -67960 82240 -67760
rect 85040 -67960 85240 -67760
rect 88040 -67960 88240 -67760
rect 91040 -67960 91240 -67760
rect 94040 -67960 94240 -67760
rect 97040 -67960 97240 -67760
rect 100040 -67960 100240 -67760
rect 103040 -67960 103240 -67760
rect 106040 -67960 106240 -67760
rect 109040 -67960 109240 -67760
rect 112040 -67960 112240 -67760
rect 115040 -67960 115240 -67760
rect 118040 -67960 118240 -67760
rect 121040 -67960 121240 -67760
rect 124040 -67960 124240 -67760
rect 127040 -67960 127240 -67760
rect 130040 -67960 130240 -67760
rect 133040 -67960 133240 -67760
rect 136040 -67960 136240 -67760
rect 139040 -67960 139240 -67760
rect 142040 -67960 142240 -67760
rect 145040 -67960 145240 -67760
rect 148040 -67960 148240 -67760
rect 1040 -70960 1240 -70760
rect 4040 -70960 4240 -70760
rect 7040 -70960 7240 -70760
rect 10040 -70960 10240 -70760
rect 13040 -70960 13240 -70760
rect 16040 -70960 16240 -70760
rect 19040 -70960 19240 -70760
rect 22040 -70960 22240 -70760
rect 25040 -70960 25240 -70760
rect 28040 -70960 28240 -70760
rect 31040 -70960 31240 -70760
rect 34040 -70960 34240 -70760
rect 37040 -70960 37240 -70760
rect 40040 -70960 40240 -70760
rect 43040 -70960 43240 -70760
rect 46040 -70960 46240 -70760
rect 49040 -70960 49240 -70760
rect 52040 -70960 52240 -70760
rect 55040 -70960 55240 -70760
rect 58040 -70960 58240 -70760
rect 61040 -70960 61240 -70760
rect 64040 -70960 64240 -70760
rect 67040 -70960 67240 -70760
rect 70040 -70960 70240 -70760
rect 73040 -70960 73240 -70760
rect 76040 -70960 76240 -70760
rect 79040 -70960 79240 -70760
rect 82040 -70960 82240 -70760
rect 85040 -70960 85240 -70760
rect 88040 -70960 88240 -70760
rect 91040 -70960 91240 -70760
rect 94040 -70960 94240 -70760
rect 97040 -70960 97240 -70760
rect 100040 -70960 100240 -70760
rect 103040 -70960 103240 -70760
rect 106040 -70960 106240 -70760
rect 109040 -70960 109240 -70760
rect 112040 -70960 112240 -70760
rect 115040 -70960 115240 -70760
rect 118040 -70960 118240 -70760
rect 121040 -70960 121240 -70760
rect 124040 -70960 124240 -70760
rect 127040 -70960 127240 -70760
rect 130040 -70960 130240 -70760
rect 133040 -70960 133240 -70760
rect 136040 -70960 136240 -70760
rect 139040 -70960 139240 -70760
rect 142040 -70960 142240 -70760
rect 145040 -70960 145240 -70760
rect 148040 -70960 148240 -70760
rect 1040 -73960 1240 -73760
rect 4040 -73960 4240 -73760
rect 7040 -73960 7240 -73760
rect 10040 -73960 10240 -73760
rect 13040 -73960 13240 -73760
rect 16040 -73960 16240 -73760
rect 19040 -73960 19240 -73760
rect 22040 -73960 22240 -73760
rect 25040 -73960 25240 -73760
rect 28040 -73960 28240 -73760
rect 31040 -73960 31240 -73760
rect 34040 -73960 34240 -73760
rect 37040 -73960 37240 -73760
rect 40040 -73960 40240 -73760
rect 43040 -73960 43240 -73760
rect 46040 -73960 46240 -73760
rect 49040 -73960 49240 -73760
rect 52040 -73960 52240 -73760
rect 55040 -73960 55240 -73760
rect 58040 -73960 58240 -73760
rect 61040 -73960 61240 -73760
rect 64040 -73960 64240 -73760
rect 67040 -73960 67240 -73760
rect 70040 -73960 70240 -73760
rect 73040 -73960 73240 -73760
rect 76040 -73960 76240 -73760
rect 79040 -73960 79240 -73760
rect 82040 -73960 82240 -73760
rect 85040 -73960 85240 -73760
rect 88040 -73960 88240 -73760
rect 91040 -73960 91240 -73760
rect 94040 -73960 94240 -73760
rect 97040 -73960 97240 -73760
rect 100040 -73960 100240 -73760
rect 103040 -73960 103240 -73760
rect 106040 -73960 106240 -73760
rect 109040 -73960 109240 -73760
rect 112040 -73960 112240 -73760
rect 115040 -73960 115240 -73760
rect 118040 -73960 118240 -73760
rect 121040 -73960 121240 -73760
rect 124040 -73960 124240 -73760
rect 127040 -73960 127240 -73760
rect 130040 -73960 130240 -73760
rect 133040 -73960 133240 -73760
rect 136040 -73960 136240 -73760
rect 139040 -73960 139240 -73760
rect 142040 -73960 142240 -73760
rect 145040 -73960 145240 -73760
rect 148040 -73960 148240 -73760
rect 1040 -76960 1240 -76760
rect 4040 -76960 4240 -76760
rect 7040 -76960 7240 -76760
rect 10040 -76960 10240 -76760
rect 13040 -76960 13240 -76760
rect 16040 -76960 16240 -76760
rect 19040 -76960 19240 -76760
rect 22040 -76960 22240 -76760
rect 25040 -76960 25240 -76760
rect 28040 -76960 28240 -76760
rect 31040 -76960 31240 -76760
rect 34040 -76960 34240 -76760
rect 37040 -76960 37240 -76760
rect 40040 -76960 40240 -76760
rect 43040 -76960 43240 -76760
rect 46040 -76960 46240 -76760
rect 49040 -76960 49240 -76760
rect 52040 -76960 52240 -76760
rect 55040 -76960 55240 -76760
rect 58040 -76960 58240 -76760
rect 61040 -76960 61240 -76760
rect 64040 -76960 64240 -76760
rect 67040 -76960 67240 -76760
rect 70040 -76960 70240 -76760
rect 73040 -76960 73240 -76760
rect 76040 -76960 76240 -76760
rect 79040 -76960 79240 -76760
rect 82040 -76960 82240 -76760
rect 85040 -76960 85240 -76760
rect 88040 -76960 88240 -76760
rect 91040 -76960 91240 -76760
rect 94040 -76960 94240 -76760
rect 97040 -76960 97240 -76760
rect 100040 -76960 100240 -76760
rect 103040 -76960 103240 -76760
rect 106040 -76960 106240 -76760
rect 109040 -76960 109240 -76760
rect 112040 -76960 112240 -76760
rect 115040 -76960 115240 -76760
rect 118040 -76960 118240 -76760
rect 121040 -76960 121240 -76760
rect 124040 -76960 124240 -76760
rect 127040 -76960 127240 -76760
rect 130040 -76960 130240 -76760
rect 133040 -76960 133240 -76760
rect 136040 -76960 136240 -76760
rect 139040 -76960 139240 -76760
rect 142040 -76960 142240 -76760
rect 145040 -76960 145240 -76760
rect 148040 -76960 148240 -76760
rect 1040 -79960 1240 -79760
rect 4040 -79960 4240 -79760
rect 7040 -79960 7240 -79760
rect 10040 -79960 10240 -79760
rect 13040 -79960 13240 -79760
rect 16040 -79960 16240 -79760
rect 19040 -79960 19240 -79760
rect 22040 -79960 22240 -79760
rect 25040 -79960 25240 -79760
rect 28040 -79960 28240 -79760
rect 31040 -79960 31240 -79760
rect 34040 -79960 34240 -79760
rect 37040 -79960 37240 -79760
rect 40040 -79960 40240 -79760
rect 43040 -79960 43240 -79760
rect 46040 -79960 46240 -79760
rect 49040 -79960 49240 -79760
rect 52040 -79960 52240 -79760
rect 55040 -79960 55240 -79760
rect 58040 -79960 58240 -79760
rect 61040 -79960 61240 -79760
rect 64040 -79960 64240 -79760
rect 67040 -79960 67240 -79760
rect 70040 -79960 70240 -79760
rect 73040 -79960 73240 -79760
rect 76040 -79960 76240 -79760
rect 79040 -79960 79240 -79760
rect 82040 -79960 82240 -79760
rect 85040 -79960 85240 -79760
rect 88040 -79960 88240 -79760
rect 91040 -79960 91240 -79760
rect 94040 -79960 94240 -79760
rect 97040 -79960 97240 -79760
rect 100040 -79960 100240 -79760
rect 103040 -79960 103240 -79760
rect 106040 -79960 106240 -79760
rect 109040 -79960 109240 -79760
rect 112040 -79960 112240 -79760
rect 115040 -79960 115240 -79760
rect 118040 -79960 118240 -79760
rect 121040 -79960 121240 -79760
rect 124040 -79960 124240 -79760
rect 127040 -79960 127240 -79760
rect 130040 -79960 130240 -79760
rect 133040 -79960 133240 -79760
rect 136040 -79960 136240 -79760
rect 139040 -79960 139240 -79760
rect 142040 -79960 142240 -79760
rect 145040 -79960 145240 -79760
rect 148040 -79960 148240 -79760
rect 1040 -82960 1240 -82760
rect 4040 -82960 4240 -82760
rect 7040 -82960 7240 -82760
rect 10040 -82960 10240 -82760
rect 13040 -82960 13240 -82760
rect 16040 -82960 16240 -82760
rect 19040 -82960 19240 -82760
rect 22040 -82960 22240 -82760
rect 25040 -82960 25240 -82760
rect 28040 -82960 28240 -82760
rect 31040 -82960 31240 -82760
rect 34040 -82960 34240 -82760
rect 37040 -82960 37240 -82760
rect 40040 -82960 40240 -82760
rect 43040 -82960 43240 -82760
rect 46040 -82960 46240 -82760
rect 49040 -82960 49240 -82760
rect 52040 -82960 52240 -82760
rect 55040 -82960 55240 -82760
rect 58040 -82960 58240 -82760
rect 61040 -82960 61240 -82760
rect 64040 -82960 64240 -82760
rect 67040 -82960 67240 -82760
rect 70040 -82960 70240 -82760
rect 73040 -82960 73240 -82760
rect 76040 -82960 76240 -82760
rect 79040 -82960 79240 -82760
rect 82040 -82960 82240 -82760
rect 85040 -82960 85240 -82760
rect 88040 -82960 88240 -82760
rect 91040 -82960 91240 -82760
rect 94040 -82960 94240 -82760
rect 97040 -82960 97240 -82760
rect 100040 -82960 100240 -82760
rect 103040 -82960 103240 -82760
rect 106040 -82960 106240 -82760
rect 109040 -82960 109240 -82760
rect 112040 -82960 112240 -82760
rect 115040 -82960 115240 -82760
rect 118040 -82960 118240 -82760
rect 121040 -82960 121240 -82760
rect 124040 -82960 124240 -82760
rect 127040 -82960 127240 -82760
rect 130040 -82960 130240 -82760
rect 133040 -82960 133240 -82760
rect 136040 -82960 136240 -82760
rect 139040 -82960 139240 -82760
rect 142040 -82960 142240 -82760
rect 145040 -82960 145240 -82760
rect 148040 -82960 148240 -82760
rect 1040 -85960 1240 -85760
rect 4040 -85960 4240 -85760
rect 7040 -85960 7240 -85760
rect 10040 -85960 10240 -85760
rect 13040 -85960 13240 -85760
rect 16040 -85960 16240 -85760
rect 19040 -85960 19240 -85760
rect 22040 -85960 22240 -85760
rect 25040 -85960 25240 -85760
rect 28040 -85960 28240 -85760
rect 31040 -85960 31240 -85760
rect 34040 -85960 34240 -85760
rect 37040 -85960 37240 -85760
rect 40040 -85960 40240 -85760
rect 43040 -85960 43240 -85760
rect 46040 -85960 46240 -85760
rect 49040 -85960 49240 -85760
rect 52040 -85960 52240 -85760
rect 55040 -85960 55240 -85760
rect 58040 -85960 58240 -85760
rect 61040 -85960 61240 -85760
rect 64040 -85960 64240 -85760
rect 67040 -85960 67240 -85760
rect 70040 -85960 70240 -85760
rect 73040 -85960 73240 -85760
rect 76040 -85960 76240 -85760
rect 79040 -85960 79240 -85760
rect 82040 -85960 82240 -85760
rect 85040 -85960 85240 -85760
rect 88040 -85960 88240 -85760
rect 91040 -85960 91240 -85760
rect 94040 -85960 94240 -85760
rect 97040 -85960 97240 -85760
rect 100040 -85960 100240 -85760
rect 103040 -85960 103240 -85760
rect 106040 -85960 106240 -85760
rect 109040 -85960 109240 -85760
rect 112040 -85960 112240 -85760
rect 115040 -85960 115240 -85760
rect 118040 -85960 118240 -85760
rect 121040 -85960 121240 -85760
rect 124040 -85960 124240 -85760
rect 127040 -85960 127240 -85760
rect 130040 -85960 130240 -85760
rect 133040 -85960 133240 -85760
rect 136040 -85960 136240 -85760
rect 139040 -85960 139240 -85760
rect 142040 -85960 142240 -85760
rect 145040 -85960 145240 -85760
rect 148040 -85960 148240 -85760
rect 1040 -88960 1240 -88760
rect 4040 -88960 4240 -88760
rect 7040 -88960 7240 -88760
rect 10040 -88960 10240 -88760
rect 13040 -88960 13240 -88760
rect 16040 -88960 16240 -88760
rect 19040 -88960 19240 -88760
rect 22040 -88960 22240 -88760
rect 25040 -88960 25240 -88760
rect 28040 -88960 28240 -88760
rect 31040 -88960 31240 -88760
rect 34040 -88960 34240 -88760
rect 37040 -88960 37240 -88760
rect 40040 -88960 40240 -88760
rect 43040 -88960 43240 -88760
rect 46040 -88960 46240 -88760
rect 49040 -88960 49240 -88760
rect 52040 -88960 52240 -88760
rect 55040 -88960 55240 -88760
rect 58040 -88960 58240 -88760
rect 61040 -88960 61240 -88760
rect 64040 -88960 64240 -88760
rect 67040 -88960 67240 -88760
rect 70040 -88960 70240 -88760
rect 73040 -88960 73240 -88760
rect 76040 -88960 76240 -88760
rect 79040 -88960 79240 -88760
rect 82040 -88960 82240 -88760
rect 85040 -88960 85240 -88760
rect 88040 -88960 88240 -88760
rect 91040 -88960 91240 -88760
rect 94040 -88960 94240 -88760
rect 97040 -88960 97240 -88760
rect 100040 -88960 100240 -88760
rect 103040 -88960 103240 -88760
rect 106040 -88960 106240 -88760
rect 109040 -88960 109240 -88760
rect 112040 -88960 112240 -88760
rect 115040 -88960 115240 -88760
rect 118040 -88960 118240 -88760
rect 121040 -88960 121240 -88760
rect 124040 -88960 124240 -88760
rect 127040 -88960 127240 -88760
rect 130040 -88960 130240 -88760
rect 133040 -88960 133240 -88760
rect 136040 -88960 136240 -88760
rect 139040 -88960 139240 -88760
rect 142040 -88960 142240 -88760
rect 145040 -88960 145240 -88760
rect 148040 -88960 148240 -88760
rect 1040 -91960 1240 -91760
rect 4040 -91960 4240 -91760
rect 7040 -91960 7240 -91760
rect 10040 -91960 10240 -91760
rect 13040 -91960 13240 -91760
rect 16040 -91960 16240 -91760
rect 19040 -91960 19240 -91760
rect 22040 -91960 22240 -91760
rect 25040 -91960 25240 -91760
rect 28040 -91960 28240 -91760
rect 31040 -91960 31240 -91760
rect 34040 -91960 34240 -91760
rect 37040 -91960 37240 -91760
rect 40040 -91960 40240 -91760
rect 43040 -91960 43240 -91760
rect 46040 -91960 46240 -91760
rect 49040 -91960 49240 -91760
rect 52040 -91960 52240 -91760
rect 55040 -91960 55240 -91760
rect 58040 -91960 58240 -91760
rect 61040 -91960 61240 -91760
rect 64040 -91960 64240 -91760
rect 67040 -91960 67240 -91760
rect 70040 -91960 70240 -91760
rect 73040 -91960 73240 -91760
rect 76040 -91960 76240 -91760
rect 79040 -91960 79240 -91760
rect 82040 -91960 82240 -91760
rect 85040 -91960 85240 -91760
rect 88040 -91960 88240 -91760
rect 91040 -91960 91240 -91760
rect 94040 -91960 94240 -91760
rect 97040 -91960 97240 -91760
rect 100040 -91960 100240 -91760
rect 103040 -91960 103240 -91760
rect 106040 -91960 106240 -91760
rect 109040 -91960 109240 -91760
rect 112040 -91960 112240 -91760
rect 115040 -91960 115240 -91760
rect 118040 -91960 118240 -91760
rect 121040 -91960 121240 -91760
rect 124040 -91960 124240 -91760
rect 127040 -91960 127240 -91760
rect 130040 -91960 130240 -91760
rect 133040 -91960 133240 -91760
rect 136040 -91960 136240 -91760
rect 139040 -91960 139240 -91760
rect 142040 -91960 142240 -91760
rect 145040 -91960 145240 -91760
rect 148040 -91960 148240 -91760
rect 1040 -94960 1240 -94760
rect 4040 -94960 4240 -94760
rect 7040 -94960 7240 -94760
rect 10040 -94960 10240 -94760
rect 13040 -94960 13240 -94760
rect 16040 -94960 16240 -94760
rect 19040 -94960 19240 -94760
rect 22040 -94960 22240 -94760
rect 25040 -94960 25240 -94760
rect 28040 -94960 28240 -94760
rect 31040 -94960 31240 -94760
rect 34040 -94960 34240 -94760
rect 37040 -94960 37240 -94760
rect 40040 -94960 40240 -94760
rect 43040 -94960 43240 -94760
rect 46040 -94960 46240 -94760
rect 49040 -94960 49240 -94760
rect 52040 -94960 52240 -94760
rect 55040 -94960 55240 -94760
rect 58040 -94960 58240 -94760
rect 61040 -94960 61240 -94760
rect 64040 -94960 64240 -94760
rect 67040 -94960 67240 -94760
rect 70040 -94960 70240 -94760
rect 73040 -94960 73240 -94760
rect 76040 -94960 76240 -94760
rect 79040 -94960 79240 -94760
rect 82040 -94960 82240 -94760
rect 85040 -94960 85240 -94760
rect 88040 -94960 88240 -94760
rect 91040 -94960 91240 -94760
rect 94040 -94960 94240 -94760
rect 97040 -94960 97240 -94760
rect 100040 -94960 100240 -94760
rect 103040 -94960 103240 -94760
rect 106040 -94960 106240 -94760
rect 109040 -94960 109240 -94760
rect 112040 -94960 112240 -94760
rect 115040 -94960 115240 -94760
rect 118040 -94960 118240 -94760
rect 121040 -94960 121240 -94760
rect 124040 -94960 124240 -94760
rect 127040 -94960 127240 -94760
rect 130040 -94960 130240 -94760
rect 133040 -94960 133240 -94760
rect 136040 -94960 136240 -94760
rect 139040 -94960 139240 -94760
rect 142040 -94960 142240 -94760
rect 145040 -94960 145240 -94760
rect 148040 -94960 148240 -94760
rect 1040 -97960 1240 -97760
rect 4040 -97960 4240 -97760
rect 7040 -97960 7240 -97760
rect 10040 -97960 10240 -97760
rect 13040 -97960 13240 -97760
rect 16040 -97960 16240 -97760
rect 19040 -97960 19240 -97760
rect 22040 -97960 22240 -97760
rect 25040 -97960 25240 -97760
rect 28040 -97960 28240 -97760
rect 31040 -97960 31240 -97760
rect 34040 -97960 34240 -97760
rect 37040 -97960 37240 -97760
rect 40040 -97960 40240 -97760
rect 43040 -97960 43240 -97760
rect 46040 -97960 46240 -97760
rect 49040 -97960 49240 -97760
rect 52040 -97960 52240 -97760
rect 55040 -97960 55240 -97760
rect 58040 -97960 58240 -97760
rect 61040 -97960 61240 -97760
rect 64040 -97960 64240 -97760
rect 67040 -97960 67240 -97760
rect 70040 -97960 70240 -97760
rect 73040 -97960 73240 -97760
rect 76040 -97960 76240 -97760
rect 79040 -97960 79240 -97760
rect 82040 -97960 82240 -97760
rect 85040 -97960 85240 -97760
rect 88040 -97960 88240 -97760
rect 91040 -97960 91240 -97760
rect 94040 -97960 94240 -97760
rect 97040 -97960 97240 -97760
rect 100040 -97960 100240 -97760
rect 103040 -97960 103240 -97760
rect 106040 -97960 106240 -97760
rect 109040 -97960 109240 -97760
rect 112040 -97960 112240 -97760
rect 115040 -97960 115240 -97760
rect 118040 -97960 118240 -97760
rect 121040 -97960 121240 -97760
rect 124040 -97960 124240 -97760
rect 127040 -97960 127240 -97760
rect 130040 -97960 130240 -97760
rect 133040 -97960 133240 -97760
rect 136040 -97960 136240 -97760
rect 139040 -97960 139240 -97760
rect 142040 -97960 142240 -97760
rect 145040 -97960 145240 -97760
rect 148040 -97960 148240 -97760
rect 1040 -100960 1240 -100760
rect 4040 -100960 4240 -100760
rect 7040 -100960 7240 -100760
rect 10040 -100960 10240 -100760
rect 13040 -100960 13240 -100760
rect 16040 -100960 16240 -100760
rect 19040 -100960 19240 -100760
rect 22040 -100960 22240 -100760
rect 25040 -100960 25240 -100760
rect 28040 -100960 28240 -100760
rect 31040 -100960 31240 -100760
rect 34040 -100960 34240 -100760
rect 37040 -100960 37240 -100760
rect 40040 -100960 40240 -100760
rect 43040 -100960 43240 -100760
rect 46040 -100960 46240 -100760
rect 49040 -100960 49240 -100760
rect 52040 -100960 52240 -100760
rect 55040 -100960 55240 -100760
rect 58040 -100960 58240 -100760
rect 61040 -100960 61240 -100760
rect 64040 -100960 64240 -100760
rect 67040 -100960 67240 -100760
rect 70040 -100960 70240 -100760
rect 73040 -100960 73240 -100760
rect 76040 -100960 76240 -100760
rect 79040 -100960 79240 -100760
rect 82040 -100960 82240 -100760
rect 85040 -100960 85240 -100760
rect 88040 -100960 88240 -100760
rect 91040 -100960 91240 -100760
rect 94040 -100960 94240 -100760
rect 97040 -100960 97240 -100760
rect 100040 -100960 100240 -100760
rect 103040 -100960 103240 -100760
rect 106040 -100960 106240 -100760
rect 109040 -100960 109240 -100760
rect 112040 -100960 112240 -100760
rect 115040 -100960 115240 -100760
rect 118040 -100960 118240 -100760
rect 121040 -100960 121240 -100760
rect 124040 -100960 124240 -100760
rect 127040 -100960 127240 -100760
rect 130040 -100960 130240 -100760
rect 133040 -100960 133240 -100760
rect 136040 -100960 136240 -100760
rect 139040 -100960 139240 -100760
rect 142040 -100960 142240 -100760
rect 145040 -100960 145240 -100760
rect 148040 -100960 148240 -100760
rect 1040 -103960 1240 -103760
rect 4040 -103960 4240 -103760
rect 7040 -103960 7240 -103760
rect 10040 -103960 10240 -103760
rect 13040 -103960 13240 -103760
rect 16040 -103960 16240 -103760
rect 19040 -103960 19240 -103760
rect 22040 -103960 22240 -103760
rect 25040 -103960 25240 -103760
rect 28040 -103960 28240 -103760
rect 31040 -103960 31240 -103760
rect 34040 -103960 34240 -103760
rect 37040 -103960 37240 -103760
rect 40040 -103960 40240 -103760
rect 43040 -103960 43240 -103760
rect 46040 -103960 46240 -103760
rect 49040 -103960 49240 -103760
rect 52040 -103960 52240 -103760
rect 55040 -103960 55240 -103760
rect 58040 -103960 58240 -103760
rect 61040 -103960 61240 -103760
rect 64040 -103960 64240 -103760
rect 67040 -103960 67240 -103760
rect 70040 -103960 70240 -103760
rect 73040 -103960 73240 -103760
rect 76040 -103960 76240 -103760
rect 79040 -103960 79240 -103760
rect 82040 -103960 82240 -103760
rect 85040 -103960 85240 -103760
rect 88040 -103960 88240 -103760
rect 91040 -103960 91240 -103760
rect 94040 -103960 94240 -103760
rect 97040 -103960 97240 -103760
rect 100040 -103960 100240 -103760
rect 103040 -103960 103240 -103760
rect 106040 -103960 106240 -103760
rect 109040 -103960 109240 -103760
rect 112040 -103960 112240 -103760
rect 115040 -103960 115240 -103760
rect 118040 -103960 118240 -103760
rect 121040 -103960 121240 -103760
rect 124040 -103960 124240 -103760
rect 127040 -103960 127240 -103760
rect 130040 -103960 130240 -103760
rect 133040 -103960 133240 -103760
rect 136040 -103960 136240 -103760
rect 139040 -103960 139240 -103760
rect 142040 -103960 142240 -103760
rect 145040 -103960 145240 -103760
rect 148040 -103960 148240 -103760
rect 1040 -106960 1240 -106760
rect 4040 -106960 4240 -106760
rect 7040 -106960 7240 -106760
rect 10040 -106960 10240 -106760
rect 13040 -106960 13240 -106760
rect 16040 -106960 16240 -106760
rect 19040 -106960 19240 -106760
rect 22040 -106960 22240 -106760
rect 25040 -106960 25240 -106760
rect 28040 -106960 28240 -106760
rect 31040 -106960 31240 -106760
rect 34040 -106960 34240 -106760
rect 37040 -106960 37240 -106760
rect 40040 -106960 40240 -106760
rect 43040 -106960 43240 -106760
rect 46040 -106960 46240 -106760
rect 49040 -106960 49240 -106760
rect 52040 -106960 52240 -106760
rect 55040 -106960 55240 -106760
rect 58040 -106960 58240 -106760
rect 61040 -106960 61240 -106760
rect 64040 -106960 64240 -106760
rect 67040 -106960 67240 -106760
rect 70040 -106960 70240 -106760
rect 73040 -106960 73240 -106760
rect 76040 -106960 76240 -106760
rect 79040 -106960 79240 -106760
rect 82040 -106960 82240 -106760
rect 85040 -106960 85240 -106760
rect 88040 -106960 88240 -106760
rect 91040 -106960 91240 -106760
rect 94040 -106960 94240 -106760
rect 97040 -106960 97240 -106760
rect 100040 -106960 100240 -106760
rect 103040 -106960 103240 -106760
rect 106040 -106960 106240 -106760
rect 109040 -106960 109240 -106760
rect 112040 -106960 112240 -106760
rect 115040 -106960 115240 -106760
rect 118040 -106960 118240 -106760
rect 121040 -106960 121240 -106760
rect 124040 -106960 124240 -106760
rect 127040 -106960 127240 -106760
rect 130040 -106960 130240 -106760
rect 133040 -106960 133240 -106760
rect 136040 -106960 136240 -106760
rect 139040 -106960 139240 -106760
rect 142040 -106960 142240 -106760
rect 145040 -106960 145240 -106760
rect 148040 -106960 148240 -106760
rect 1040 -109960 1240 -109760
rect 4040 -109960 4240 -109760
rect 7040 -109960 7240 -109760
rect 10040 -109960 10240 -109760
rect 13040 -109960 13240 -109760
rect 16040 -109960 16240 -109760
rect 19040 -109960 19240 -109760
rect 22040 -109960 22240 -109760
rect 25040 -109960 25240 -109760
rect 28040 -109960 28240 -109760
rect 31040 -109960 31240 -109760
rect 34040 -109960 34240 -109760
rect 37040 -109960 37240 -109760
rect 40040 -109960 40240 -109760
rect 43040 -109960 43240 -109760
rect 46040 -109960 46240 -109760
rect 49040 -109960 49240 -109760
rect 52040 -109960 52240 -109760
rect 55040 -109960 55240 -109760
rect 58040 -109960 58240 -109760
rect 61040 -109960 61240 -109760
rect 64040 -109960 64240 -109760
rect 67040 -109960 67240 -109760
rect 70040 -109960 70240 -109760
rect 73040 -109960 73240 -109760
rect 76040 -109960 76240 -109760
rect 79040 -109960 79240 -109760
rect 82040 -109960 82240 -109760
rect 85040 -109960 85240 -109760
rect 88040 -109960 88240 -109760
rect 91040 -109960 91240 -109760
rect 94040 -109960 94240 -109760
rect 97040 -109960 97240 -109760
rect 100040 -109960 100240 -109760
rect 103040 -109960 103240 -109760
rect 106040 -109960 106240 -109760
rect 109040 -109960 109240 -109760
rect 112040 -109960 112240 -109760
rect 115040 -109960 115240 -109760
rect 118040 -109960 118240 -109760
rect 121040 -109960 121240 -109760
rect 124040 -109960 124240 -109760
rect 127040 -109960 127240 -109760
rect 130040 -109960 130240 -109760
rect 133040 -109960 133240 -109760
rect 136040 -109960 136240 -109760
rect 139040 -109960 139240 -109760
rect 142040 -109960 142240 -109760
rect 145040 -109960 145240 -109760
rect 148040 -109960 148240 -109760
rect 1040 -112960 1240 -112760
rect 4040 -112960 4240 -112760
rect 7040 -112960 7240 -112760
rect 10040 -112960 10240 -112760
rect 13040 -112960 13240 -112760
rect 16040 -112960 16240 -112760
rect 19040 -112960 19240 -112760
rect 22040 -112960 22240 -112760
rect 25040 -112960 25240 -112760
rect 28040 -112960 28240 -112760
rect 31040 -112960 31240 -112760
rect 34040 -112960 34240 -112760
rect 37040 -112960 37240 -112760
rect 40040 -112960 40240 -112760
rect 43040 -112960 43240 -112760
rect 46040 -112960 46240 -112760
rect 49040 -112960 49240 -112760
rect 52040 -112960 52240 -112760
rect 55040 -112960 55240 -112760
rect 58040 -112960 58240 -112760
rect 61040 -112960 61240 -112760
rect 64040 -112960 64240 -112760
rect 67040 -112960 67240 -112760
rect 70040 -112960 70240 -112760
rect 73040 -112960 73240 -112760
rect 76040 -112960 76240 -112760
rect 79040 -112960 79240 -112760
rect 82040 -112960 82240 -112760
rect 85040 -112960 85240 -112760
rect 88040 -112960 88240 -112760
rect 91040 -112960 91240 -112760
rect 94040 -112960 94240 -112760
rect 97040 -112960 97240 -112760
rect 100040 -112960 100240 -112760
rect 103040 -112960 103240 -112760
rect 106040 -112960 106240 -112760
rect 109040 -112960 109240 -112760
rect 112040 -112960 112240 -112760
rect 115040 -112960 115240 -112760
rect 118040 -112960 118240 -112760
rect 121040 -112960 121240 -112760
rect 124040 -112960 124240 -112760
rect 127040 -112960 127240 -112760
rect 130040 -112960 130240 -112760
rect 133040 -112960 133240 -112760
rect 136040 -112960 136240 -112760
rect 139040 -112960 139240 -112760
rect 142040 -112960 142240 -112760
rect 145040 -112960 145240 -112760
rect 148040 -112960 148240 -112760
rect 1040 -115960 1240 -115760
rect 4040 -115960 4240 -115760
rect 7040 -115960 7240 -115760
rect 10040 -115960 10240 -115760
rect 13040 -115960 13240 -115760
rect 16040 -115960 16240 -115760
rect 19040 -115960 19240 -115760
rect 22040 -115960 22240 -115760
rect 25040 -115960 25240 -115760
rect 28040 -115960 28240 -115760
rect 31040 -115960 31240 -115760
rect 34040 -115960 34240 -115760
rect 37040 -115960 37240 -115760
rect 40040 -115960 40240 -115760
rect 43040 -115960 43240 -115760
rect 46040 -115960 46240 -115760
rect 49040 -115960 49240 -115760
rect 52040 -115960 52240 -115760
rect 55040 -115960 55240 -115760
rect 58040 -115960 58240 -115760
rect 61040 -115960 61240 -115760
rect 64040 -115960 64240 -115760
rect 67040 -115960 67240 -115760
rect 70040 -115960 70240 -115760
rect 73040 -115960 73240 -115760
rect 76040 -115960 76240 -115760
rect 79040 -115960 79240 -115760
rect 82040 -115960 82240 -115760
rect 85040 -115960 85240 -115760
rect 88040 -115960 88240 -115760
rect 91040 -115960 91240 -115760
rect 94040 -115960 94240 -115760
rect 97040 -115960 97240 -115760
rect 100040 -115960 100240 -115760
rect 103040 -115960 103240 -115760
rect 106040 -115960 106240 -115760
rect 109040 -115960 109240 -115760
rect 112040 -115960 112240 -115760
rect 115040 -115960 115240 -115760
rect 118040 -115960 118240 -115760
rect 121040 -115960 121240 -115760
rect 124040 -115960 124240 -115760
rect 127040 -115960 127240 -115760
rect 130040 -115960 130240 -115760
rect 133040 -115960 133240 -115760
rect 136040 -115960 136240 -115760
rect 139040 -115960 139240 -115760
rect 142040 -115960 142240 -115760
rect 145040 -115960 145240 -115760
rect 148040 -115960 148240 -115760
rect 1040 -118960 1240 -118760
rect 4040 -118960 4240 -118760
rect 7040 -118960 7240 -118760
rect 10040 -118960 10240 -118760
rect 13040 -118960 13240 -118760
rect 16040 -118960 16240 -118760
rect 19040 -118960 19240 -118760
rect 22040 -118960 22240 -118760
rect 25040 -118960 25240 -118760
rect 28040 -118960 28240 -118760
rect 31040 -118960 31240 -118760
rect 34040 -118960 34240 -118760
rect 37040 -118960 37240 -118760
rect 40040 -118960 40240 -118760
rect 43040 -118960 43240 -118760
rect 46040 -118960 46240 -118760
rect 49040 -118960 49240 -118760
rect 52040 -118960 52240 -118760
rect 55040 -118960 55240 -118760
rect 58040 -118960 58240 -118760
rect 61040 -118960 61240 -118760
rect 64040 -118960 64240 -118760
rect 67040 -118960 67240 -118760
rect 70040 -118960 70240 -118760
rect 73040 -118960 73240 -118760
rect 76040 -118960 76240 -118760
rect 79040 -118960 79240 -118760
rect 82040 -118960 82240 -118760
rect 85040 -118960 85240 -118760
rect 88040 -118960 88240 -118760
rect 91040 -118960 91240 -118760
rect 94040 -118960 94240 -118760
rect 97040 -118960 97240 -118760
rect 100040 -118960 100240 -118760
rect 103040 -118960 103240 -118760
rect 106040 -118960 106240 -118760
rect 109040 -118960 109240 -118760
rect 112040 -118960 112240 -118760
rect 115040 -118960 115240 -118760
rect 118040 -118960 118240 -118760
rect 121040 -118960 121240 -118760
rect 124040 -118960 124240 -118760
rect 127040 -118960 127240 -118760
rect 130040 -118960 130240 -118760
rect 133040 -118960 133240 -118760
rect 136040 -118960 136240 -118760
rect 139040 -118960 139240 -118760
rect 142040 -118960 142240 -118760
rect 145040 -118960 145240 -118760
rect 148040 -118960 148240 -118760
rect 1040 -121960 1240 -121760
rect 4040 -121960 4240 -121760
rect 7040 -121960 7240 -121760
rect 10040 -121960 10240 -121760
rect 13040 -121960 13240 -121760
rect 16040 -121960 16240 -121760
rect 19040 -121960 19240 -121760
rect 22040 -121960 22240 -121760
rect 25040 -121960 25240 -121760
rect 28040 -121960 28240 -121760
rect 31040 -121960 31240 -121760
rect 34040 -121960 34240 -121760
rect 37040 -121960 37240 -121760
rect 40040 -121960 40240 -121760
rect 43040 -121960 43240 -121760
rect 46040 -121960 46240 -121760
rect 49040 -121960 49240 -121760
rect 52040 -121960 52240 -121760
rect 55040 -121960 55240 -121760
rect 58040 -121960 58240 -121760
rect 61040 -121960 61240 -121760
rect 64040 -121960 64240 -121760
rect 67040 -121960 67240 -121760
rect 70040 -121960 70240 -121760
rect 73040 -121960 73240 -121760
rect 76040 -121960 76240 -121760
rect 79040 -121960 79240 -121760
rect 82040 -121960 82240 -121760
rect 85040 -121960 85240 -121760
rect 88040 -121960 88240 -121760
rect 91040 -121960 91240 -121760
rect 94040 -121960 94240 -121760
rect 97040 -121960 97240 -121760
rect 100040 -121960 100240 -121760
rect 103040 -121960 103240 -121760
rect 106040 -121960 106240 -121760
rect 109040 -121960 109240 -121760
rect 112040 -121960 112240 -121760
rect 115040 -121960 115240 -121760
rect 118040 -121960 118240 -121760
rect 121040 -121960 121240 -121760
rect 124040 -121960 124240 -121760
rect 127040 -121960 127240 -121760
rect 130040 -121960 130240 -121760
rect 133040 -121960 133240 -121760
rect 136040 -121960 136240 -121760
rect 139040 -121960 139240 -121760
rect 142040 -121960 142240 -121760
rect 145040 -121960 145240 -121760
rect 148040 -121960 148240 -121760
rect 1040 -124960 1240 -124760
rect 4040 -124960 4240 -124760
rect 7040 -124960 7240 -124760
rect 10040 -124960 10240 -124760
rect 13040 -124960 13240 -124760
rect 16040 -124960 16240 -124760
rect 19040 -124960 19240 -124760
rect 22040 -124960 22240 -124760
rect 25040 -124960 25240 -124760
rect 28040 -124960 28240 -124760
rect 31040 -124960 31240 -124760
rect 34040 -124960 34240 -124760
rect 37040 -124960 37240 -124760
rect 40040 -124960 40240 -124760
rect 43040 -124960 43240 -124760
rect 46040 -124960 46240 -124760
rect 49040 -124960 49240 -124760
rect 52040 -124960 52240 -124760
rect 55040 -124960 55240 -124760
rect 58040 -124960 58240 -124760
rect 61040 -124960 61240 -124760
rect 64040 -124960 64240 -124760
rect 67040 -124960 67240 -124760
rect 70040 -124960 70240 -124760
rect 73040 -124960 73240 -124760
rect 76040 -124960 76240 -124760
rect 79040 -124960 79240 -124760
rect 82040 -124960 82240 -124760
rect 85040 -124960 85240 -124760
rect 88040 -124960 88240 -124760
rect 91040 -124960 91240 -124760
rect 94040 -124960 94240 -124760
rect 97040 -124960 97240 -124760
rect 100040 -124960 100240 -124760
rect 103040 -124960 103240 -124760
rect 106040 -124960 106240 -124760
rect 109040 -124960 109240 -124760
rect 112040 -124960 112240 -124760
rect 115040 -124960 115240 -124760
rect 118040 -124960 118240 -124760
rect 121040 -124960 121240 -124760
rect 124040 -124960 124240 -124760
rect 127040 -124960 127240 -124760
rect 130040 -124960 130240 -124760
rect 133040 -124960 133240 -124760
rect 136040 -124960 136240 -124760
rect 139040 -124960 139240 -124760
rect 142040 -124960 142240 -124760
rect 145040 -124960 145240 -124760
rect 148040 -124960 148240 -124760
rect 1040 -127960 1240 -127760
rect 4040 -127960 4240 -127760
rect 7040 -127960 7240 -127760
rect 10040 -127960 10240 -127760
rect 13040 -127960 13240 -127760
rect 16040 -127960 16240 -127760
rect 19040 -127960 19240 -127760
rect 22040 -127960 22240 -127760
rect 25040 -127960 25240 -127760
rect 28040 -127960 28240 -127760
rect 31040 -127960 31240 -127760
rect 34040 -127960 34240 -127760
rect 37040 -127960 37240 -127760
rect 40040 -127960 40240 -127760
rect 43040 -127960 43240 -127760
rect 46040 -127960 46240 -127760
rect 49040 -127960 49240 -127760
rect 52040 -127960 52240 -127760
rect 55040 -127960 55240 -127760
rect 58040 -127960 58240 -127760
rect 61040 -127960 61240 -127760
rect 64040 -127960 64240 -127760
rect 67040 -127960 67240 -127760
rect 70040 -127960 70240 -127760
rect 73040 -127960 73240 -127760
rect 76040 -127960 76240 -127760
rect 79040 -127960 79240 -127760
rect 82040 -127960 82240 -127760
rect 85040 -127960 85240 -127760
rect 88040 -127960 88240 -127760
rect 91040 -127960 91240 -127760
rect 94040 -127960 94240 -127760
rect 97040 -127960 97240 -127760
rect 100040 -127960 100240 -127760
rect 103040 -127960 103240 -127760
rect 106040 -127960 106240 -127760
rect 109040 -127960 109240 -127760
rect 112040 -127960 112240 -127760
rect 115040 -127960 115240 -127760
rect 118040 -127960 118240 -127760
rect 121040 -127960 121240 -127760
rect 124040 -127960 124240 -127760
rect 127040 -127960 127240 -127760
rect 130040 -127960 130240 -127760
rect 133040 -127960 133240 -127760
rect 136040 -127960 136240 -127760
rect 139040 -127960 139240 -127760
rect 142040 -127960 142240 -127760
rect 145040 -127960 145240 -127760
rect 148040 -127960 148240 -127760
rect 1040 -130960 1240 -130760
rect 4040 -130960 4240 -130760
rect 7040 -130960 7240 -130760
rect 10040 -130960 10240 -130760
rect 13040 -130960 13240 -130760
rect 16040 -130960 16240 -130760
rect 19040 -130960 19240 -130760
rect 22040 -130960 22240 -130760
rect 25040 -130960 25240 -130760
rect 28040 -130960 28240 -130760
rect 31040 -130960 31240 -130760
rect 34040 -130960 34240 -130760
rect 37040 -130960 37240 -130760
rect 40040 -130960 40240 -130760
rect 43040 -130960 43240 -130760
rect 46040 -130960 46240 -130760
rect 49040 -130960 49240 -130760
rect 52040 -130960 52240 -130760
rect 55040 -130960 55240 -130760
rect 58040 -130960 58240 -130760
rect 61040 -130960 61240 -130760
rect 64040 -130960 64240 -130760
rect 67040 -130960 67240 -130760
rect 70040 -130960 70240 -130760
rect 73040 -130960 73240 -130760
rect 76040 -130960 76240 -130760
rect 79040 -130960 79240 -130760
rect 82040 -130960 82240 -130760
rect 85040 -130960 85240 -130760
rect 88040 -130960 88240 -130760
rect 91040 -130960 91240 -130760
rect 94040 -130960 94240 -130760
rect 97040 -130960 97240 -130760
rect 100040 -130960 100240 -130760
rect 103040 -130960 103240 -130760
rect 106040 -130960 106240 -130760
rect 109040 -130960 109240 -130760
rect 112040 -130960 112240 -130760
rect 115040 -130960 115240 -130760
rect 118040 -130960 118240 -130760
rect 121040 -130960 121240 -130760
rect 124040 -130960 124240 -130760
rect 127040 -130960 127240 -130760
rect 130040 -130960 130240 -130760
rect 133040 -130960 133240 -130760
rect 136040 -130960 136240 -130760
rect 139040 -130960 139240 -130760
rect 142040 -130960 142240 -130760
rect 145040 -130960 145240 -130760
rect 148040 -130960 148240 -130760
rect 1040 -133960 1240 -133760
rect 4040 -133960 4240 -133760
rect 7040 -133960 7240 -133760
rect 10040 -133960 10240 -133760
rect 13040 -133960 13240 -133760
rect 16040 -133960 16240 -133760
rect 19040 -133960 19240 -133760
rect 22040 -133960 22240 -133760
rect 25040 -133960 25240 -133760
rect 28040 -133960 28240 -133760
rect 31040 -133960 31240 -133760
rect 34040 -133960 34240 -133760
rect 37040 -133960 37240 -133760
rect 40040 -133960 40240 -133760
rect 43040 -133960 43240 -133760
rect 46040 -133960 46240 -133760
rect 49040 -133960 49240 -133760
rect 52040 -133960 52240 -133760
rect 55040 -133960 55240 -133760
rect 58040 -133960 58240 -133760
rect 61040 -133960 61240 -133760
rect 64040 -133960 64240 -133760
rect 67040 -133960 67240 -133760
rect 70040 -133960 70240 -133760
rect 73040 -133960 73240 -133760
rect 76040 -133960 76240 -133760
rect 79040 -133960 79240 -133760
rect 82040 -133960 82240 -133760
rect 85040 -133960 85240 -133760
rect 88040 -133960 88240 -133760
rect 91040 -133960 91240 -133760
rect 94040 -133960 94240 -133760
rect 97040 -133960 97240 -133760
rect 100040 -133960 100240 -133760
rect 103040 -133960 103240 -133760
rect 106040 -133960 106240 -133760
rect 109040 -133960 109240 -133760
rect 112040 -133960 112240 -133760
rect 115040 -133960 115240 -133760
rect 118040 -133960 118240 -133760
rect 121040 -133960 121240 -133760
rect 124040 -133960 124240 -133760
rect 127040 -133960 127240 -133760
rect 130040 -133960 130240 -133760
rect 133040 -133960 133240 -133760
rect 136040 -133960 136240 -133760
rect 139040 -133960 139240 -133760
rect 142040 -133960 142240 -133760
rect 145040 -133960 145240 -133760
rect 148040 -133960 148240 -133760
rect 1040 -136960 1240 -136760
rect 4040 -136960 4240 -136760
rect 7040 -136960 7240 -136760
rect 10040 -136960 10240 -136760
rect 13040 -136960 13240 -136760
rect 16040 -136960 16240 -136760
rect 19040 -136960 19240 -136760
rect 22040 -136960 22240 -136760
rect 25040 -136960 25240 -136760
rect 28040 -136960 28240 -136760
rect 31040 -136960 31240 -136760
rect 34040 -136960 34240 -136760
rect 37040 -136960 37240 -136760
rect 40040 -136960 40240 -136760
rect 43040 -136960 43240 -136760
rect 46040 -136960 46240 -136760
rect 49040 -136960 49240 -136760
rect 52040 -136960 52240 -136760
rect 55040 -136960 55240 -136760
rect 58040 -136960 58240 -136760
rect 61040 -136960 61240 -136760
rect 64040 -136960 64240 -136760
rect 67040 -136960 67240 -136760
rect 70040 -136960 70240 -136760
rect 73040 -136960 73240 -136760
rect 76040 -136960 76240 -136760
rect 79040 -136960 79240 -136760
rect 82040 -136960 82240 -136760
rect 85040 -136960 85240 -136760
rect 88040 -136960 88240 -136760
rect 91040 -136960 91240 -136760
rect 94040 -136960 94240 -136760
rect 97040 -136960 97240 -136760
rect 100040 -136960 100240 -136760
rect 103040 -136960 103240 -136760
rect 106040 -136960 106240 -136760
rect 109040 -136960 109240 -136760
rect 112040 -136960 112240 -136760
rect 115040 -136960 115240 -136760
rect 118040 -136960 118240 -136760
rect 121040 -136960 121240 -136760
rect 124040 -136960 124240 -136760
rect 127040 -136960 127240 -136760
rect 130040 -136960 130240 -136760
rect 133040 -136960 133240 -136760
rect 136040 -136960 136240 -136760
rect 139040 -136960 139240 -136760
rect 142040 -136960 142240 -136760
rect 145040 -136960 145240 -136760
rect 148040 -136960 148240 -136760
rect 1040 -139960 1240 -139760
rect 4040 -139960 4240 -139760
rect 7040 -139960 7240 -139760
rect 10040 -139960 10240 -139760
rect 13040 -139960 13240 -139760
rect 16040 -139960 16240 -139760
rect 19040 -139960 19240 -139760
rect 22040 -139960 22240 -139760
rect 25040 -139960 25240 -139760
rect 28040 -139960 28240 -139760
rect 31040 -139960 31240 -139760
rect 34040 -139960 34240 -139760
rect 37040 -139960 37240 -139760
rect 40040 -139960 40240 -139760
rect 43040 -139960 43240 -139760
rect 46040 -139960 46240 -139760
rect 49040 -139960 49240 -139760
rect 52040 -139960 52240 -139760
rect 55040 -139960 55240 -139760
rect 58040 -139960 58240 -139760
rect 61040 -139960 61240 -139760
rect 64040 -139960 64240 -139760
rect 67040 -139960 67240 -139760
rect 70040 -139960 70240 -139760
rect 73040 -139960 73240 -139760
rect 76040 -139960 76240 -139760
rect 79040 -139960 79240 -139760
rect 82040 -139960 82240 -139760
rect 85040 -139960 85240 -139760
rect 88040 -139960 88240 -139760
rect 91040 -139960 91240 -139760
rect 94040 -139960 94240 -139760
rect 97040 -139960 97240 -139760
rect 100040 -139960 100240 -139760
rect 103040 -139960 103240 -139760
rect 106040 -139960 106240 -139760
rect 109040 -139960 109240 -139760
rect 112040 -139960 112240 -139760
rect 115040 -139960 115240 -139760
rect 118040 -139960 118240 -139760
rect 121040 -139960 121240 -139760
rect 124040 -139960 124240 -139760
rect 127040 -139960 127240 -139760
rect 130040 -139960 130240 -139760
rect 133040 -139960 133240 -139760
rect 136040 -139960 136240 -139760
rect 139040 -139960 139240 -139760
rect 142040 -139960 142240 -139760
rect 145040 -139960 145240 -139760
rect 148040 -139960 148240 -139760
rect 1040 -142960 1240 -142760
rect 4040 -142960 4240 -142760
rect 7040 -142960 7240 -142760
rect 10040 -142960 10240 -142760
rect 13040 -142960 13240 -142760
rect 16040 -142960 16240 -142760
rect 19040 -142960 19240 -142760
rect 22040 -142960 22240 -142760
rect 25040 -142960 25240 -142760
rect 28040 -142960 28240 -142760
rect 31040 -142960 31240 -142760
rect 34040 -142960 34240 -142760
rect 37040 -142960 37240 -142760
rect 40040 -142960 40240 -142760
rect 43040 -142960 43240 -142760
rect 46040 -142960 46240 -142760
rect 49040 -142960 49240 -142760
rect 52040 -142960 52240 -142760
rect 55040 -142960 55240 -142760
rect 58040 -142960 58240 -142760
rect 61040 -142960 61240 -142760
rect 64040 -142960 64240 -142760
rect 67040 -142960 67240 -142760
rect 70040 -142960 70240 -142760
rect 73040 -142960 73240 -142760
rect 76040 -142960 76240 -142760
rect 79040 -142960 79240 -142760
rect 82040 -142960 82240 -142760
rect 85040 -142960 85240 -142760
rect 88040 -142960 88240 -142760
rect 91040 -142960 91240 -142760
rect 94040 -142960 94240 -142760
rect 97040 -142960 97240 -142760
rect 100040 -142960 100240 -142760
rect 103040 -142960 103240 -142760
rect 106040 -142960 106240 -142760
rect 109040 -142960 109240 -142760
rect 112040 -142960 112240 -142760
rect 115040 -142960 115240 -142760
rect 118040 -142960 118240 -142760
rect 121040 -142960 121240 -142760
rect 124040 -142960 124240 -142760
rect 127040 -142960 127240 -142760
rect 130040 -142960 130240 -142760
rect 133040 -142960 133240 -142760
rect 136040 -142960 136240 -142760
rect 139040 -142960 139240 -142760
rect 142040 -142960 142240 -142760
rect 145040 -142960 145240 -142760
rect 148040 -142960 148240 -142760
rect 1040 -145960 1240 -145760
rect 4040 -145960 4240 -145760
rect 7040 -145960 7240 -145760
rect 10040 -145960 10240 -145760
rect 13040 -145960 13240 -145760
rect 16040 -145960 16240 -145760
rect 19040 -145960 19240 -145760
rect 22040 -145960 22240 -145760
rect 25040 -145960 25240 -145760
rect 28040 -145960 28240 -145760
rect 31040 -145960 31240 -145760
rect 34040 -145960 34240 -145760
rect 37040 -145960 37240 -145760
rect 40040 -145960 40240 -145760
rect 43040 -145960 43240 -145760
rect 46040 -145960 46240 -145760
rect 49040 -145960 49240 -145760
rect 52040 -145960 52240 -145760
rect 55040 -145960 55240 -145760
rect 58040 -145960 58240 -145760
rect 61040 -145960 61240 -145760
rect 64040 -145960 64240 -145760
rect 67040 -145960 67240 -145760
rect 70040 -145960 70240 -145760
rect 73040 -145960 73240 -145760
rect 76040 -145960 76240 -145760
rect 79040 -145960 79240 -145760
rect 82040 -145960 82240 -145760
rect 85040 -145960 85240 -145760
rect 88040 -145960 88240 -145760
rect 91040 -145960 91240 -145760
rect 94040 -145960 94240 -145760
rect 97040 -145960 97240 -145760
rect 100040 -145960 100240 -145760
rect 103040 -145960 103240 -145760
rect 106040 -145960 106240 -145760
rect 109040 -145960 109240 -145760
rect 112040 -145960 112240 -145760
rect 115040 -145960 115240 -145760
rect 118040 -145960 118240 -145760
rect 121040 -145960 121240 -145760
rect 124040 -145960 124240 -145760
rect 127040 -145960 127240 -145760
rect 130040 -145960 130240 -145760
rect 133040 -145960 133240 -145760
rect 136040 -145960 136240 -145760
rect 139040 -145960 139240 -145760
rect 142040 -145960 142240 -145760
rect 145040 -145960 145240 -145760
rect 148040 -145960 148240 -145760
use pixel  pixel_2451
timestamp 1654648307
transform 1 0 -800 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2450
timestamp 1654648307
transform 1 0 -3800 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2453
timestamp 1654648307
transform 1 0 5200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2452
timestamp 1654648307
transform 1 0 2200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2455
timestamp 1654648307
transform 1 0 11200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2454
timestamp 1654648307
transform 1 0 8200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2457
timestamp 1654648307
transform 1 0 17200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2456
timestamp 1654648307
transform 1 0 14200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2459
timestamp 1654648307
transform 1 0 23200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2458
timestamp 1654648307
transform 1 0 20200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2461
timestamp 1654648307
transform 1 0 29200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2460
timestamp 1654648307
transform 1 0 26200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2463
timestamp 1654648307
transform 1 0 35200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2462
timestamp 1654648307
transform 1 0 32200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2465
timestamp 1654648307
transform 1 0 41200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2464
timestamp 1654648307
transform 1 0 38200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2467
timestamp 1654648307
transform 1 0 47200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2466
timestamp 1654648307
transform 1 0 44200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2469
timestamp 1654648307
transform 1 0 53200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2468
timestamp 1654648307
transform 1 0 50200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2471
timestamp 1654648307
transform 1 0 59200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2470
timestamp 1654648307
transform 1 0 56200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2473
timestamp 1654648307
transform 1 0 65200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2472
timestamp 1654648307
transform 1 0 62200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2475
timestamp 1654648307
transform 1 0 71200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2474
timestamp 1654648307
transform 1 0 68200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2477
timestamp 1654648307
transform 1 0 77200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2476
timestamp 1654648307
transform 1 0 74200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2479
timestamp 1654648307
transform 1 0 83200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2478
timestamp 1654648307
transform 1 0 80200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2481
timestamp 1654648307
transform 1 0 89200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2480
timestamp 1654648307
transform 1 0 86200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2483
timestamp 1654648307
transform 1 0 95200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2482
timestamp 1654648307
transform 1 0 92200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2485
timestamp 1654648307
transform 1 0 101200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2484
timestamp 1654648307
transform 1 0 98200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2487
timestamp 1654648307
transform 1 0 107200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2486
timestamp 1654648307
transform 1 0 104200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2489
timestamp 1654648307
transform 1 0 113200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2488
timestamp 1654648307
transform 1 0 110200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2491
timestamp 1654648307
transform 1 0 119200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2490
timestamp 1654648307
transform 1 0 116200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2493
timestamp 1654648307
transform 1 0 125200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2492
timestamp 1654648307
transform 1 0 122200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2495
timestamp 1654648307
transform 1 0 131200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2494
timestamp 1654648307
transform 1 0 128200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2497
timestamp 1654648307
transform 1 0 137200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2496
timestamp 1654648307
transform 1 0 134200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2499
timestamp 1654648307
transform 1 0 143200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2498
timestamp 1654648307
transform 1 0 140200 0 1 -144300
box 3640 -2860 6960 460
use pixel  pixel_2401
timestamp 1654648307
transform 1 0 -800 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2400
timestamp 1654648307
transform 1 0 -3800 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2351
timestamp 1654648307
transform 1 0 -800 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2350
timestamp 1654648307
transform 1 0 -3800 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2403
timestamp 1654648307
transform 1 0 5200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2402
timestamp 1654648307
transform 1 0 2200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2353
timestamp 1654648307
transform 1 0 5200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2352
timestamp 1654648307
transform 1 0 2200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2405
timestamp 1654648307
transform 1 0 11200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2404
timestamp 1654648307
transform 1 0 8200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2355
timestamp 1654648307
transform 1 0 11200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2354
timestamp 1654648307
transform 1 0 8200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2407
timestamp 1654648307
transform 1 0 17200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2406
timestamp 1654648307
transform 1 0 14200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2357
timestamp 1654648307
transform 1 0 17200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2356
timestamp 1654648307
transform 1 0 14200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2409
timestamp 1654648307
transform 1 0 23200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2408
timestamp 1654648307
transform 1 0 20200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2359
timestamp 1654648307
transform 1 0 23200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2358
timestamp 1654648307
transform 1 0 20200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2411
timestamp 1654648307
transform 1 0 29200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2410
timestamp 1654648307
transform 1 0 26200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2361
timestamp 1654648307
transform 1 0 29200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2360
timestamp 1654648307
transform 1 0 26200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2413
timestamp 1654648307
transform 1 0 35200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2412
timestamp 1654648307
transform 1 0 32200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2363
timestamp 1654648307
transform 1 0 35200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2362
timestamp 1654648307
transform 1 0 32200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2415
timestamp 1654648307
transform 1 0 41200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2414
timestamp 1654648307
transform 1 0 38200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2365
timestamp 1654648307
transform 1 0 41200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2364
timestamp 1654648307
transform 1 0 38200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2417
timestamp 1654648307
transform 1 0 47200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2416
timestamp 1654648307
transform 1 0 44200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2367
timestamp 1654648307
transform 1 0 47200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2366
timestamp 1654648307
transform 1 0 44200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2419
timestamp 1654648307
transform 1 0 53200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2418
timestamp 1654648307
transform 1 0 50200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2369
timestamp 1654648307
transform 1 0 53200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2368
timestamp 1654648307
transform 1 0 50200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2421
timestamp 1654648307
transform 1 0 59200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2420
timestamp 1654648307
transform 1 0 56200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2371
timestamp 1654648307
transform 1 0 59200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2370
timestamp 1654648307
transform 1 0 56200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2423
timestamp 1654648307
transform 1 0 65200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2422
timestamp 1654648307
transform 1 0 62200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2373
timestamp 1654648307
transform 1 0 65200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2372
timestamp 1654648307
transform 1 0 62200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2425
timestamp 1654648307
transform 1 0 71200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2424
timestamp 1654648307
transform 1 0 68200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2375
timestamp 1654648307
transform 1 0 71200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2374
timestamp 1654648307
transform 1 0 68200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2427
timestamp 1654648307
transform 1 0 77200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2426
timestamp 1654648307
transform 1 0 74200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2377
timestamp 1654648307
transform 1 0 77200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2376
timestamp 1654648307
transform 1 0 74200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2429
timestamp 1654648307
transform 1 0 83200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2428
timestamp 1654648307
transform 1 0 80200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2379
timestamp 1654648307
transform 1 0 83200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2378
timestamp 1654648307
transform 1 0 80200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2431
timestamp 1654648307
transform 1 0 89200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2430
timestamp 1654648307
transform 1 0 86200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2381
timestamp 1654648307
transform 1 0 89200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2380
timestamp 1654648307
transform 1 0 86200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2433
timestamp 1654648307
transform 1 0 95200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2432
timestamp 1654648307
transform 1 0 92200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2383
timestamp 1654648307
transform 1 0 95200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2382
timestamp 1654648307
transform 1 0 92200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2435
timestamp 1654648307
transform 1 0 101200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2434
timestamp 1654648307
transform 1 0 98200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2385
timestamp 1654648307
transform 1 0 101200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2384
timestamp 1654648307
transform 1 0 98200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2437
timestamp 1654648307
transform 1 0 107200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2436
timestamp 1654648307
transform 1 0 104200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2387
timestamp 1654648307
transform 1 0 107200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2386
timestamp 1654648307
transform 1 0 104200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2439
timestamp 1654648307
transform 1 0 113200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2438
timestamp 1654648307
transform 1 0 110200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2389
timestamp 1654648307
transform 1 0 113200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2388
timestamp 1654648307
transform 1 0 110200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2441
timestamp 1654648307
transform 1 0 119200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2440
timestamp 1654648307
transform 1 0 116200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2391
timestamp 1654648307
transform 1 0 119200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2390
timestamp 1654648307
transform 1 0 116200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2443
timestamp 1654648307
transform 1 0 125200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2442
timestamp 1654648307
transform 1 0 122200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2393
timestamp 1654648307
transform 1 0 125200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2392
timestamp 1654648307
transform 1 0 122200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2445
timestamp 1654648307
transform 1 0 131200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2444
timestamp 1654648307
transform 1 0 128200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2395
timestamp 1654648307
transform 1 0 131200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2394
timestamp 1654648307
transform 1 0 128200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2447
timestamp 1654648307
transform 1 0 137200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2446
timestamp 1654648307
transform 1 0 134200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2397
timestamp 1654648307
transform 1 0 137200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2396
timestamp 1654648307
transform 1 0 134200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2449
timestamp 1654648307
transform 1 0 143200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2448
timestamp 1654648307
transform 1 0 140200 0 1 -141300
box 3640 -2860 6960 460
use pixel  pixel_2399
timestamp 1654648307
transform 1 0 143200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2398
timestamp 1654648307
transform 1 0 140200 0 1 -138300
box 3640 -2860 6960 460
use pixel  pixel_2301
timestamp 1654648307
transform 1 0 -800 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2300
timestamp 1654648307
transform 1 0 -3800 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2251
timestamp 1654648307
transform 1 0 -800 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2250
timestamp 1654648307
transform 1 0 -3800 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2303
timestamp 1654648307
transform 1 0 5200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2302
timestamp 1654648307
transform 1 0 2200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2253
timestamp 1654648307
transform 1 0 5200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2252
timestamp 1654648307
transform 1 0 2200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2305
timestamp 1654648307
transform 1 0 11200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2304
timestamp 1654648307
transform 1 0 8200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2255
timestamp 1654648307
transform 1 0 11200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2254
timestamp 1654648307
transform 1 0 8200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2307
timestamp 1654648307
transform 1 0 17200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2306
timestamp 1654648307
transform 1 0 14200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2257
timestamp 1654648307
transform 1 0 17200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2256
timestamp 1654648307
transform 1 0 14200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2309
timestamp 1654648307
transform 1 0 23200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2308
timestamp 1654648307
transform 1 0 20200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2259
timestamp 1654648307
transform 1 0 23200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2258
timestamp 1654648307
transform 1 0 20200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2311
timestamp 1654648307
transform 1 0 29200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2310
timestamp 1654648307
transform 1 0 26200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2261
timestamp 1654648307
transform 1 0 29200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2260
timestamp 1654648307
transform 1 0 26200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2313
timestamp 1654648307
transform 1 0 35200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2312
timestamp 1654648307
transform 1 0 32200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2263
timestamp 1654648307
transform 1 0 35200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2262
timestamp 1654648307
transform 1 0 32200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2315
timestamp 1654648307
transform 1 0 41200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2314
timestamp 1654648307
transform 1 0 38200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2265
timestamp 1654648307
transform 1 0 41200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2264
timestamp 1654648307
transform 1 0 38200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2317
timestamp 1654648307
transform 1 0 47200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2316
timestamp 1654648307
transform 1 0 44200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2267
timestamp 1654648307
transform 1 0 47200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2266
timestamp 1654648307
transform 1 0 44200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2319
timestamp 1654648307
transform 1 0 53200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2318
timestamp 1654648307
transform 1 0 50200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2269
timestamp 1654648307
transform 1 0 53200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2268
timestamp 1654648307
transform 1 0 50200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2321
timestamp 1654648307
transform 1 0 59200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2320
timestamp 1654648307
transform 1 0 56200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2271
timestamp 1654648307
transform 1 0 59200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2270
timestamp 1654648307
transform 1 0 56200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2323
timestamp 1654648307
transform 1 0 65200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2322
timestamp 1654648307
transform 1 0 62200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2273
timestamp 1654648307
transform 1 0 65200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2272
timestamp 1654648307
transform 1 0 62200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2325
timestamp 1654648307
transform 1 0 71200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2324
timestamp 1654648307
transform 1 0 68200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2275
timestamp 1654648307
transform 1 0 71200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2274
timestamp 1654648307
transform 1 0 68200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2327
timestamp 1654648307
transform 1 0 77200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2326
timestamp 1654648307
transform 1 0 74200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2277
timestamp 1654648307
transform 1 0 77200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2276
timestamp 1654648307
transform 1 0 74200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2329
timestamp 1654648307
transform 1 0 83200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2328
timestamp 1654648307
transform 1 0 80200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2279
timestamp 1654648307
transform 1 0 83200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2278
timestamp 1654648307
transform 1 0 80200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2331
timestamp 1654648307
transform 1 0 89200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2330
timestamp 1654648307
transform 1 0 86200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2281
timestamp 1654648307
transform 1 0 89200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2280
timestamp 1654648307
transform 1 0 86200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2333
timestamp 1654648307
transform 1 0 95200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2332
timestamp 1654648307
transform 1 0 92200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2283
timestamp 1654648307
transform 1 0 95200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2282
timestamp 1654648307
transform 1 0 92200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2335
timestamp 1654648307
transform 1 0 101200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2334
timestamp 1654648307
transform 1 0 98200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2285
timestamp 1654648307
transform 1 0 101200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2284
timestamp 1654648307
transform 1 0 98200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2337
timestamp 1654648307
transform 1 0 107200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2336
timestamp 1654648307
transform 1 0 104200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2287
timestamp 1654648307
transform 1 0 107200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2286
timestamp 1654648307
transform 1 0 104200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2339
timestamp 1654648307
transform 1 0 113200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2338
timestamp 1654648307
transform 1 0 110200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2289
timestamp 1654648307
transform 1 0 113200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2288
timestamp 1654648307
transform 1 0 110200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2341
timestamp 1654648307
transform 1 0 119200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2340
timestamp 1654648307
transform 1 0 116200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2291
timestamp 1654648307
transform 1 0 119200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2290
timestamp 1654648307
transform 1 0 116200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2343
timestamp 1654648307
transform 1 0 125200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2342
timestamp 1654648307
transform 1 0 122200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2293
timestamp 1654648307
transform 1 0 125200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2292
timestamp 1654648307
transform 1 0 122200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2345
timestamp 1654648307
transform 1 0 131200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2344
timestamp 1654648307
transform 1 0 128200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2295
timestamp 1654648307
transform 1 0 131200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2294
timestamp 1654648307
transform 1 0 128200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2347
timestamp 1654648307
transform 1 0 137200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2346
timestamp 1654648307
transform 1 0 134200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2297
timestamp 1654648307
transform 1 0 137200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2296
timestamp 1654648307
transform 1 0 134200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2349
timestamp 1654648307
transform 1 0 143200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2348
timestamp 1654648307
transform 1 0 140200 0 1 -135300
box 3640 -2860 6960 460
use pixel  pixel_2299
timestamp 1654648307
transform 1 0 143200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2298
timestamp 1654648307
transform 1 0 140200 0 1 -132300
box 3640 -2860 6960 460
use pixel  pixel_2201
timestamp 1654648307
transform 1 0 -800 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2200
timestamp 1654648307
transform 1 0 -3800 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2151
timestamp 1654648307
transform 1 0 -800 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2150
timestamp 1654648307
transform 1 0 -3800 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2203
timestamp 1654648307
transform 1 0 5200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2202
timestamp 1654648307
transform 1 0 2200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2153
timestamp 1654648307
transform 1 0 5200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2152
timestamp 1654648307
transform 1 0 2200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2205
timestamp 1654648307
transform 1 0 11200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2204
timestamp 1654648307
transform 1 0 8200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2155
timestamp 1654648307
transform 1 0 11200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2154
timestamp 1654648307
transform 1 0 8200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2207
timestamp 1654648307
transform 1 0 17200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2206
timestamp 1654648307
transform 1 0 14200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2157
timestamp 1654648307
transform 1 0 17200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2156
timestamp 1654648307
transform 1 0 14200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2209
timestamp 1654648307
transform 1 0 23200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2208
timestamp 1654648307
transform 1 0 20200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2159
timestamp 1654648307
transform 1 0 23200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2158
timestamp 1654648307
transform 1 0 20200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2211
timestamp 1654648307
transform 1 0 29200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2210
timestamp 1654648307
transform 1 0 26200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2161
timestamp 1654648307
transform 1 0 29200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2160
timestamp 1654648307
transform 1 0 26200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2213
timestamp 1654648307
transform 1 0 35200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2212
timestamp 1654648307
transform 1 0 32200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2163
timestamp 1654648307
transform 1 0 35200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2162
timestamp 1654648307
transform 1 0 32200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2215
timestamp 1654648307
transform 1 0 41200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2214
timestamp 1654648307
transform 1 0 38200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2165
timestamp 1654648307
transform 1 0 41200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2164
timestamp 1654648307
transform 1 0 38200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2217
timestamp 1654648307
transform 1 0 47200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2216
timestamp 1654648307
transform 1 0 44200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2167
timestamp 1654648307
transform 1 0 47200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2166
timestamp 1654648307
transform 1 0 44200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2219
timestamp 1654648307
transform 1 0 53200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2218
timestamp 1654648307
transform 1 0 50200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2169
timestamp 1654648307
transform 1 0 53200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2168
timestamp 1654648307
transform 1 0 50200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2221
timestamp 1654648307
transform 1 0 59200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2220
timestamp 1654648307
transform 1 0 56200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2171
timestamp 1654648307
transform 1 0 59200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2170
timestamp 1654648307
transform 1 0 56200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2223
timestamp 1654648307
transform 1 0 65200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2222
timestamp 1654648307
transform 1 0 62200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2173
timestamp 1654648307
transform 1 0 65200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2172
timestamp 1654648307
transform 1 0 62200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2225
timestamp 1654648307
transform 1 0 71200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2224
timestamp 1654648307
transform 1 0 68200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2175
timestamp 1654648307
transform 1 0 71200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2174
timestamp 1654648307
transform 1 0 68200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2227
timestamp 1654648307
transform 1 0 77200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2226
timestamp 1654648307
transform 1 0 74200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2177
timestamp 1654648307
transform 1 0 77200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2176
timestamp 1654648307
transform 1 0 74200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2229
timestamp 1654648307
transform 1 0 83200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2228
timestamp 1654648307
transform 1 0 80200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2179
timestamp 1654648307
transform 1 0 83200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2178
timestamp 1654648307
transform 1 0 80200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2231
timestamp 1654648307
transform 1 0 89200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2230
timestamp 1654648307
transform 1 0 86200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2181
timestamp 1654648307
transform 1 0 89200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2180
timestamp 1654648307
transform 1 0 86200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2233
timestamp 1654648307
transform 1 0 95200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2232
timestamp 1654648307
transform 1 0 92200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2183
timestamp 1654648307
transform 1 0 95200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2182
timestamp 1654648307
transform 1 0 92200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2235
timestamp 1654648307
transform 1 0 101200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2234
timestamp 1654648307
transform 1 0 98200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2185
timestamp 1654648307
transform 1 0 101200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2184
timestamp 1654648307
transform 1 0 98200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2237
timestamp 1654648307
transform 1 0 107200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2236
timestamp 1654648307
transform 1 0 104200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2187
timestamp 1654648307
transform 1 0 107200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2186
timestamp 1654648307
transform 1 0 104200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2239
timestamp 1654648307
transform 1 0 113200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2238
timestamp 1654648307
transform 1 0 110200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2189
timestamp 1654648307
transform 1 0 113200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2188
timestamp 1654648307
transform 1 0 110200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2241
timestamp 1654648307
transform 1 0 119200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2240
timestamp 1654648307
transform 1 0 116200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2191
timestamp 1654648307
transform 1 0 119200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2190
timestamp 1654648307
transform 1 0 116200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2243
timestamp 1654648307
transform 1 0 125200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2242
timestamp 1654648307
transform 1 0 122200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2193
timestamp 1654648307
transform 1 0 125200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2192
timestamp 1654648307
transform 1 0 122200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2245
timestamp 1654648307
transform 1 0 131200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2244
timestamp 1654648307
transform 1 0 128200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2195
timestamp 1654648307
transform 1 0 131200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2194
timestamp 1654648307
transform 1 0 128200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2247
timestamp 1654648307
transform 1 0 137200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2246
timestamp 1654648307
transform 1 0 134200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2197
timestamp 1654648307
transform 1 0 137200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2196
timestamp 1654648307
transform 1 0 134200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2249
timestamp 1654648307
transform 1 0 143200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2248
timestamp 1654648307
transform 1 0 140200 0 1 -129300
box 3640 -2860 6960 460
use pixel  pixel_2199
timestamp 1654648307
transform 1 0 143200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2198
timestamp 1654648307
transform 1 0 140200 0 1 -126300
box 3640 -2860 6960 460
use pixel  pixel_2101
timestamp 1654648307
transform 1 0 -800 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2100
timestamp 1654648307
transform 1 0 -3800 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2051
timestamp 1654648307
transform 1 0 -800 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2050
timestamp 1654648307
transform 1 0 -3800 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2103
timestamp 1654648307
transform 1 0 5200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2102
timestamp 1654648307
transform 1 0 2200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2053
timestamp 1654648307
transform 1 0 5200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2052
timestamp 1654648307
transform 1 0 2200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2105
timestamp 1654648307
transform 1 0 11200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2104
timestamp 1654648307
transform 1 0 8200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2055
timestamp 1654648307
transform 1 0 11200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2054
timestamp 1654648307
transform 1 0 8200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2107
timestamp 1654648307
transform 1 0 17200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2106
timestamp 1654648307
transform 1 0 14200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2057
timestamp 1654648307
transform 1 0 17200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2056
timestamp 1654648307
transform 1 0 14200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2109
timestamp 1654648307
transform 1 0 23200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2108
timestamp 1654648307
transform 1 0 20200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2059
timestamp 1654648307
transform 1 0 23200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2058
timestamp 1654648307
transform 1 0 20200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2111
timestamp 1654648307
transform 1 0 29200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2110
timestamp 1654648307
transform 1 0 26200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2061
timestamp 1654648307
transform 1 0 29200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2060
timestamp 1654648307
transform 1 0 26200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2113
timestamp 1654648307
transform 1 0 35200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2112
timestamp 1654648307
transform 1 0 32200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2063
timestamp 1654648307
transform 1 0 35200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2062
timestamp 1654648307
transform 1 0 32200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2115
timestamp 1654648307
transform 1 0 41200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2114
timestamp 1654648307
transform 1 0 38200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2065
timestamp 1654648307
transform 1 0 41200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2064
timestamp 1654648307
transform 1 0 38200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2117
timestamp 1654648307
transform 1 0 47200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2116
timestamp 1654648307
transform 1 0 44200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2067
timestamp 1654648307
transform 1 0 47200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2066
timestamp 1654648307
transform 1 0 44200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2119
timestamp 1654648307
transform 1 0 53200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2118
timestamp 1654648307
transform 1 0 50200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2069
timestamp 1654648307
transform 1 0 53200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2068
timestamp 1654648307
transform 1 0 50200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2121
timestamp 1654648307
transform 1 0 59200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2120
timestamp 1654648307
transform 1 0 56200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2071
timestamp 1654648307
transform 1 0 59200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2070
timestamp 1654648307
transform 1 0 56200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2123
timestamp 1654648307
transform 1 0 65200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2122
timestamp 1654648307
transform 1 0 62200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2073
timestamp 1654648307
transform 1 0 65200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2072
timestamp 1654648307
transform 1 0 62200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2125
timestamp 1654648307
transform 1 0 71200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2124
timestamp 1654648307
transform 1 0 68200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2075
timestamp 1654648307
transform 1 0 71200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2074
timestamp 1654648307
transform 1 0 68200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2127
timestamp 1654648307
transform 1 0 77200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2126
timestamp 1654648307
transform 1 0 74200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2077
timestamp 1654648307
transform 1 0 77200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2076
timestamp 1654648307
transform 1 0 74200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2129
timestamp 1654648307
transform 1 0 83200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2128
timestamp 1654648307
transform 1 0 80200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2079
timestamp 1654648307
transform 1 0 83200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2078
timestamp 1654648307
transform 1 0 80200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2131
timestamp 1654648307
transform 1 0 89200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2130
timestamp 1654648307
transform 1 0 86200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2081
timestamp 1654648307
transform 1 0 89200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2080
timestamp 1654648307
transform 1 0 86200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2133
timestamp 1654648307
transform 1 0 95200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2132
timestamp 1654648307
transform 1 0 92200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2083
timestamp 1654648307
transform 1 0 95200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2082
timestamp 1654648307
transform 1 0 92200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2135
timestamp 1654648307
transform 1 0 101200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2134
timestamp 1654648307
transform 1 0 98200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2085
timestamp 1654648307
transform 1 0 101200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2084
timestamp 1654648307
transform 1 0 98200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2137
timestamp 1654648307
transform 1 0 107200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2136
timestamp 1654648307
transform 1 0 104200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2087
timestamp 1654648307
transform 1 0 107200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2086
timestamp 1654648307
transform 1 0 104200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2139
timestamp 1654648307
transform 1 0 113200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2138
timestamp 1654648307
transform 1 0 110200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2089
timestamp 1654648307
transform 1 0 113200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2088
timestamp 1654648307
transform 1 0 110200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2141
timestamp 1654648307
transform 1 0 119200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2140
timestamp 1654648307
transform 1 0 116200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2091
timestamp 1654648307
transform 1 0 119200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2090
timestamp 1654648307
transform 1 0 116200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2143
timestamp 1654648307
transform 1 0 125200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2142
timestamp 1654648307
transform 1 0 122200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2093
timestamp 1654648307
transform 1 0 125200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2092
timestamp 1654648307
transform 1 0 122200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2145
timestamp 1654648307
transform 1 0 131200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2144
timestamp 1654648307
transform 1 0 128200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2095
timestamp 1654648307
transform 1 0 131200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2094
timestamp 1654648307
transform 1 0 128200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2147
timestamp 1654648307
transform 1 0 137200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2146
timestamp 1654648307
transform 1 0 134200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2097
timestamp 1654648307
transform 1 0 137200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2096
timestamp 1654648307
transform 1 0 134200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2149
timestamp 1654648307
transform 1 0 143200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2148
timestamp 1654648307
transform 1 0 140200 0 1 -123300
box 3640 -2860 6960 460
use pixel  pixel_2099
timestamp 1654648307
transform 1 0 143200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2098
timestamp 1654648307
transform 1 0 140200 0 1 -120300
box 3640 -2860 6960 460
use pixel  pixel_2001
timestamp 1654648307
transform 1 0 -800 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_2000
timestamp 1654648307
transform 1 0 -3800 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_1951
timestamp 1654648307
transform 1 0 -800 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_1950
timestamp 1654648307
transform 1 0 -3800 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_2003
timestamp 1654648307
transform 1 0 5200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_2002
timestamp 1654648307
transform 1 0 2200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_1953
timestamp 1654648307
transform 1 0 5200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_1952
timestamp 1654648307
transform 1 0 2200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_2005
timestamp 1654648307
transform 1 0 11200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_2004
timestamp 1654648307
transform 1 0 8200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_1955
timestamp 1654648307
transform 1 0 11200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_1954
timestamp 1654648307
transform 1 0 8200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_2007
timestamp 1654648307
transform 1 0 17200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_2006
timestamp 1654648307
transform 1 0 14200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_1957
timestamp 1654648307
transform 1 0 17200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_1956
timestamp 1654648307
transform 1 0 14200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_2009
timestamp 1654648307
transform 1 0 23200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_2008
timestamp 1654648307
transform 1 0 20200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_1959
timestamp 1654648307
transform 1 0 23200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_1958
timestamp 1654648307
transform 1 0 20200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_2011
timestamp 1654648307
transform 1 0 29200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_2010
timestamp 1654648307
transform 1 0 26200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_1961
timestamp 1654648307
transform 1 0 29200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_1960
timestamp 1654648307
transform 1 0 26200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_2013
timestamp 1654648307
transform 1 0 35200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_2012
timestamp 1654648307
transform 1 0 32200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_1963
timestamp 1654648307
transform 1 0 35200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_1962
timestamp 1654648307
transform 1 0 32200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_2015
timestamp 1654648307
transform 1 0 41200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_2014
timestamp 1654648307
transform 1 0 38200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_1965
timestamp 1654648307
transform 1 0 41200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_1964
timestamp 1654648307
transform 1 0 38200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_2017
timestamp 1654648307
transform 1 0 47200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_2016
timestamp 1654648307
transform 1 0 44200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_1967
timestamp 1654648307
transform 1 0 47200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_1966
timestamp 1654648307
transform 1 0 44200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_2019
timestamp 1654648307
transform 1 0 53200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_2018
timestamp 1654648307
transform 1 0 50200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_1969
timestamp 1654648307
transform 1 0 53200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_1968
timestamp 1654648307
transform 1 0 50200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_2021
timestamp 1654648307
transform 1 0 59200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_2020
timestamp 1654648307
transform 1 0 56200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_1971
timestamp 1654648307
transform 1 0 59200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_1970
timestamp 1654648307
transform 1 0 56200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_2023
timestamp 1654648307
transform 1 0 65200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_2022
timestamp 1654648307
transform 1 0 62200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_1973
timestamp 1654648307
transform 1 0 65200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_1972
timestamp 1654648307
transform 1 0 62200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_2025
timestamp 1654648307
transform 1 0 71200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_2024
timestamp 1654648307
transform 1 0 68200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_1975
timestamp 1654648307
transform 1 0 71200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_1974
timestamp 1654648307
transform 1 0 68200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_2027
timestamp 1654648307
transform 1 0 77200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_2026
timestamp 1654648307
transform 1 0 74200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_1977
timestamp 1654648307
transform 1 0 77200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_1976
timestamp 1654648307
transform 1 0 74200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_2029
timestamp 1654648307
transform 1 0 83200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_2028
timestamp 1654648307
transform 1 0 80200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_1979
timestamp 1654648307
transform 1 0 83200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_1978
timestamp 1654648307
transform 1 0 80200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_2031
timestamp 1654648307
transform 1 0 89200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_2030
timestamp 1654648307
transform 1 0 86200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_1981
timestamp 1654648307
transform 1 0 89200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_1980
timestamp 1654648307
transform 1 0 86200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_2033
timestamp 1654648307
transform 1 0 95200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_2032
timestamp 1654648307
transform 1 0 92200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_1983
timestamp 1654648307
transform 1 0 95200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_1982
timestamp 1654648307
transform 1 0 92200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_2035
timestamp 1654648307
transform 1 0 101200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_2034
timestamp 1654648307
transform 1 0 98200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_1985
timestamp 1654648307
transform 1 0 101200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_1984
timestamp 1654648307
transform 1 0 98200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_2037
timestamp 1654648307
transform 1 0 107200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_2036
timestamp 1654648307
transform 1 0 104200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_1987
timestamp 1654648307
transform 1 0 107200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_1986
timestamp 1654648307
transform 1 0 104200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_2039
timestamp 1654648307
transform 1 0 113200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_2038
timestamp 1654648307
transform 1 0 110200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_1989
timestamp 1654648307
transform 1 0 113200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_1988
timestamp 1654648307
transform 1 0 110200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_2041
timestamp 1654648307
transform 1 0 119200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_2040
timestamp 1654648307
transform 1 0 116200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_1991
timestamp 1654648307
transform 1 0 119200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_1990
timestamp 1654648307
transform 1 0 116200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_2043
timestamp 1654648307
transform 1 0 125200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_2042
timestamp 1654648307
transform 1 0 122200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_1993
timestamp 1654648307
transform 1 0 125200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_1992
timestamp 1654648307
transform 1 0 122200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_2045
timestamp 1654648307
transform 1 0 131200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_2044
timestamp 1654648307
transform 1 0 128200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_1995
timestamp 1654648307
transform 1 0 131200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_1994
timestamp 1654648307
transform 1 0 128200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_2047
timestamp 1654648307
transform 1 0 137200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_2046
timestamp 1654648307
transform 1 0 134200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_1997
timestamp 1654648307
transform 1 0 137200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_1996
timestamp 1654648307
transform 1 0 134200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_2049
timestamp 1654648307
transform 1 0 143200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_2048
timestamp 1654648307
transform 1 0 140200 0 1 -117300
box 3640 -2860 6960 460
use pixel  pixel_1999
timestamp 1654648307
transform 1 0 143200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_1998
timestamp 1654648307
transform 1 0 140200 0 1 -114300
box 3640 -2860 6960 460
use pixel  pixel_1901
timestamp 1654648307
transform 1 0 -800 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1900
timestamp 1654648307
transform 1 0 -3800 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1851
timestamp 1654648307
transform 1 0 -800 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1850
timestamp 1654648307
transform 1 0 -3800 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1903
timestamp 1654648307
transform 1 0 5200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1902
timestamp 1654648307
transform 1 0 2200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1853
timestamp 1654648307
transform 1 0 5200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1852
timestamp 1654648307
transform 1 0 2200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1905
timestamp 1654648307
transform 1 0 11200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1904
timestamp 1654648307
transform 1 0 8200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1855
timestamp 1654648307
transform 1 0 11200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1854
timestamp 1654648307
transform 1 0 8200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1907
timestamp 1654648307
transform 1 0 17200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1906
timestamp 1654648307
transform 1 0 14200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1857
timestamp 1654648307
transform 1 0 17200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1856
timestamp 1654648307
transform 1 0 14200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1909
timestamp 1654648307
transform 1 0 23200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1908
timestamp 1654648307
transform 1 0 20200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1859
timestamp 1654648307
transform 1 0 23200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1858
timestamp 1654648307
transform 1 0 20200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1911
timestamp 1654648307
transform 1 0 29200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1910
timestamp 1654648307
transform 1 0 26200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1861
timestamp 1654648307
transform 1 0 29200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1860
timestamp 1654648307
transform 1 0 26200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1913
timestamp 1654648307
transform 1 0 35200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1912
timestamp 1654648307
transform 1 0 32200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1863
timestamp 1654648307
transform 1 0 35200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1862
timestamp 1654648307
transform 1 0 32200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1915
timestamp 1654648307
transform 1 0 41200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1914
timestamp 1654648307
transform 1 0 38200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1865
timestamp 1654648307
transform 1 0 41200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1864
timestamp 1654648307
transform 1 0 38200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1917
timestamp 1654648307
transform 1 0 47200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1916
timestamp 1654648307
transform 1 0 44200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1867
timestamp 1654648307
transform 1 0 47200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1866
timestamp 1654648307
transform 1 0 44200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1919
timestamp 1654648307
transform 1 0 53200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1918
timestamp 1654648307
transform 1 0 50200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1869
timestamp 1654648307
transform 1 0 53200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1868
timestamp 1654648307
transform 1 0 50200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1921
timestamp 1654648307
transform 1 0 59200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1920
timestamp 1654648307
transform 1 0 56200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1871
timestamp 1654648307
transform 1 0 59200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1870
timestamp 1654648307
transform 1 0 56200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1923
timestamp 1654648307
transform 1 0 65200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1922
timestamp 1654648307
transform 1 0 62200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1873
timestamp 1654648307
transform 1 0 65200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1872
timestamp 1654648307
transform 1 0 62200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1925
timestamp 1654648307
transform 1 0 71200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1924
timestamp 1654648307
transform 1 0 68200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1875
timestamp 1654648307
transform 1 0 71200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1874
timestamp 1654648307
transform 1 0 68200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1927
timestamp 1654648307
transform 1 0 77200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1926
timestamp 1654648307
transform 1 0 74200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1877
timestamp 1654648307
transform 1 0 77200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1876
timestamp 1654648307
transform 1 0 74200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1929
timestamp 1654648307
transform 1 0 83200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1928
timestamp 1654648307
transform 1 0 80200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1879
timestamp 1654648307
transform 1 0 83200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1878
timestamp 1654648307
transform 1 0 80200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1931
timestamp 1654648307
transform 1 0 89200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1930
timestamp 1654648307
transform 1 0 86200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1881
timestamp 1654648307
transform 1 0 89200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1880
timestamp 1654648307
transform 1 0 86200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1932
timestamp 1654648307
transform 1 0 92200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1882
timestamp 1654648307
transform 1 0 92200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1933
timestamp 1654648307
transform 1 0 95200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1883
timestamp 1654648307
transform 1 0 95200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1934
timestamp 1654648307
transform 1 0 98200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1884
timestamp 1654648307
transform 1 0 98200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1935
timestamp 1654648307
transform 1 0 101200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1885
timestamp 1654648307
transform 1 0 101200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1936
timestamp 1654648307
transform 1 0 104200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1886
timestamp 1654648307
transform 1 0 104200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1937
timestamp 1654648307
transform 1 0 107200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1887
timestamp 1654648307
transform 1 0 107200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1938
timestamp 1654648307
transform 1 0 110200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1888
timestamp 1654648307
transform 1 0 110200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1939
timestamp 1654648307
transform 1 0 113200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1889
timestamp 1654648307
transform 1 0 113200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1940
timestamp 1654648307
transform 1 0 116200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1890
timestamp 1654648307
transform 1 0 116200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1941
timestamp 1654648307
transform 1 0 119200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1891
timestamp 1654648307
transform 1 0 119200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1942
timestamp 1654648307
transform 1 0 122200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1892
timestamp 1654648307
transform 1 0 122200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1943
timestamp 1654648307
transform 1 0 125200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1893
timestamp 1654648307
transform 1 0 125200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1944
timestamp 1654648307
transform 1 0 128200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1894
timestamp 1654648307
transform 1 0 128200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1945
timestamp 1654648307
transform 1 0 131200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1895
timestamp 1654648307
transform 1 0 131200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1946
timestamp 1654648307
transform 1 0 134200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1896
timestamp 1654648307
transform 1 0 134200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1947
timestamp 1654648307
transform 1 0 137200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1897
timestamp 1654648307
transform 1 0 137200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1948
timestamp 1654648307
transform 1 0 140200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1898
timestamp 1654648307
transform 1 0 140200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1949
timestamp 1654648307
transform 1 0 143200 0 1 -111300
box 3640 -2860 6960 460
use pixel  pixel_1899
timestamp 1654648307
transform 1 0 143200 0 1 -108300
box 3640 -2860 6960 460
use pixel  pixel_1801
timestamp 1654648307
transform 1 0 -800 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1800
timestamp 1654648307
transform 1 0 -3800 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1751
timestamp 1654648307
transform 1 0 -800 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1750
timestamp 1654648307
transform 1 0 -3800 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1803
timestamp 1654648307
transform 1 0 5200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1802
timestamp 1654648307
transform 1 0 2200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1753
timestamp 1654648307
transform 1 0 5200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1752
timestamp 1654648307
transform 1 0 2200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1805
timestamp 1654648307
transform 1 0 11200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1804
timestamp 1654648307
transform 1 0 8200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1755
timestamp 1654648307
transform 1 0 11200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1754
timestamp 1654648307
transform 1 0 8200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1807
timestamp 1654648307
transform 1 0 17200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1806
timestamp 1654648307
transform 1 0 14200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1757
timestamp 1654648307
transform 1 0 17200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1756
timestamp 1654648307
transform 1 0 14200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1809
timestamp 1654648307
transform 1 0 23200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1808
timestamp 1654648307
transform 1 0 20200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1759
timestamp 1654648307
transform 1 0 23200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1758
timestamp 1654648307
transform 1 0 20200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1811
timestamp 1654648307
transform 1 0 29200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1810
timestamp 1654648307
transform 1 0 26200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1761
timestamp 1654648307
transform 1 0 29200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1760
timestamp 1654648307
transform 1 0 26200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1813
timestamp 1654648307
transform 1 0 35200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1812
timestamp 1654648307
transform 1 0 32200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1763
timestamp 1654648307
transform 1 0 35200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1762
timestamp 1654648307
transform 1 0 32200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1815
timestamp 1654648307
transform 1 0 41200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1814
timestamp 1654648307
transform 1 0 38200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1765
timestamp 1654648307
transform 1 0 41200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1764
timestamp 1654648307
transform 1 0 38200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1817
timestamp 1654648307
transform 1 0 47200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1816
timestamp 1654648307
transform 1 0 44200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1767
timestamp 1654648307
transform 1 0 47200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1766
timestamp 1654648307
transform 1 0 44200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1819
timestamp 1654648307
transform 1 0 53200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1818
timestamp 1654648307
transform 1 0 50200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1769
timestamp 1654648307
transform 1 0 53200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1768
timestamp 1654648307
transform 1 0 50200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1821
timestamp 1654648307
transform 1 0 59200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1820
timestamp 1654648307
transform 1 0 56200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1771
timestamp 1654648307
transform 1 0 59200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1770
timestamp 1654648307
transform 1 0 56200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1823
timestamp 1654648307
transform 1 0 65200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1822
timestamp 1654648307
transform 1 0 62200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1773
timestamp 1654648307
transform 1 0 65200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1772
timestamp 1654648307
transform 1 0 62200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1825
timestamp 1654648307
transform 1 0 71200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1824
timestamp 1654648307
transform 1 0 68200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1775
timestamp 1654648307
transform 1 0 71200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1774
timestamp 1654648307
transform 1 0 68200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1827
timestamp 1654648307
transform 1 0 77200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1826
timestamp 1654648307
transform 1 0 74200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1777
timestamp 1654648307
transform 1 0 77200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1776
timestamp 1654648307
transform 1 0 74200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1829
timestamp 1654648307
transform 1 0 83200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1828
timestamp 1654648307
transform 1 0 80200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1779
timestamp 1654648307
transform 1 0 83200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1778
timestamp 1654648307
transform 1 0 80200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1831
timestamp 1654648307
transform 1 0 89200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1830
timestamp 1654648307
transform 1 0 86200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1781
timestamp 1654648307
transform 1 0 89200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1780
timestamp 1654648307
transform 1 0 86200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1832
timestamp 1654648307
transform 1 0 92200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1782
timestamp 1654648307
transform 1 0 92200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1833
timestamp 1654648307
transform 1 0 95200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1783
timestamp 1654648307
transform 1 0 95200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1834
timestamp 1654648307
transform 1 0 98200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1784
timestamp 1654648307
transform 1 0 98200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1835
timestamp 1654648307
transform 1 0 101200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1785
timestamp 1654648307
transform 1 0 101200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1836
timestamp 1654648307
transform 1 0 104200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1786
timestamp 1654648307
transform 1 0 104200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1837
timestamp 1654648307
transform 1 0 107200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1787
timestamp 1654648307
transform 1 0 107200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1838
timestamp 1654648307
transform 1 0 110200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1788
timestamp 1654648307
transform 1 0 110200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1839
timestamp 1654648307
transform 1 0 113200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1789
timestamp 1654648307
transform 1 0 113200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1840
timestamp 1654648307
transform 1 0 116200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1790
timestamp 1654648307
transform 1 0 116200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1841
timestamp 1654648307
transform 1 0 119200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1791
timestamp 1654648307
transform 1 0 119200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1842
timestamp 1654648307
transform 1 0 122200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1792
timestamp 1654648307
transform 1 0 122200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1843
timestamp 1654648307
transform 1 0 125200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1793
timestamp 1654648307
transform 1 0 125200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1844
timestamp 1654648307
transform 1 0 128200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1794
timestamp 1654648307
transform 1 0 128200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1845
timestamp 1654648307
transform 1 0 131200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1795
timestamp 1654648307
transform 1 0 131200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1846
timestamp 1654648307
transform 1 0 134200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1796
timestamp 1654648307
transform 1 0 134200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1847
timestamp 1654648307
transform 1 0 137200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1797
timestamp 1654648307
transform 1 0 137200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1848
timestamp 1654648307
transform 1 0 140200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1798
timestamp 1654648307
transform 1 0 140200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1849
timestamp 1654648307
transform 1 0 143200 0 1 -105300
box 3640 -2860 6960 460
use pixel  pixel_1799
timestamp 1654648307
transform 1 0 143200 0 1 -102300
box 3640 -2860 6960 460
use pixel  pixel_1701
timestamp 1654648307
transform 1 0 -800 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1700
timestamp 1654648307
transform 1 0 -3800 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1651
timestamp 1654648307
transform 1 0 -800 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1650
timestamp 1654648307
transform 1 0 -3800 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1703
timestamp 1654648307
transform 1 0 5200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1702
timestamp 1654648307
transform 1 0 2200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1653
timestamp 1654648307
transform 1 0 5200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1652
timestamp 1654648307
transform 1 0 2200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1705
timestamp 1654648307
transform 1 0 11200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1704
timestamp 1654648307
transform 1 0 8200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1655
timestamp 1654648307
transform 1 0 11200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1654
timestamp 1654648307
transform 1 0 8200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1707
timestamp 1654648307
transform 1 0 17200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1706
timestamp 1654648307
transform 1 0 14200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1657
timestamp 1654648307
transform 1 0 17200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1656
timestamp 1654648307
transform 1 0 14200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1709
timestamp 1654648307
transform 1 0 23200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1708
timestamp 1654648307
transform 1 0 20200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1659
timestamp 1654648307
transform 1 0 23200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1658
timestamp 1654648307
transform 1 0 20200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1711
timestamp 1654648307
transform 1 0 29200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1710
timestamp 1654648307
transform 1 0 26200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1661
timestamp 1654648307
transform 1 0 29200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1660
timestamp 1654648307
transform 1 0 26200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1713
timestamp 1654648307
transform 1 0 35200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1712
timestamp 1654648307
transform 1 0 32200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1663
timestamp 1654648307
transform 1 0 35200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1662
timestamp 1654648307
transform 1 0 32200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1715
timestamp 1654648307
transform 1 0 41200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1714
timestamp 1654648307
transform 1 0 38200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1665
timestamp 1654648307
transform 1 0 41200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1664
timestamp 1654648307
transform 1 0 38200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1717
timestamp 1654648307
transform 1 0 47200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1716
timestamp 1654648307
transform 1 0 44200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1667
timestamp 1654648307
transform 1 0 47200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1666
timestamp 1654648307
transform 1 0 44200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1719
timestamp 1654648307
transform 1 0 53200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1718
timestamp 1654648307
transform 1 0 50200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1669
timestamp 1654648307
transform 1 0 53200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1668
timestamp 1654648307
transform 1 0 50200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1721
timestamp 1654648307
transform 1 0 59200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1720
timestamp 1654648307
transform 1 0 56200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1671
timestamp 1654648307
transform 1 0 59200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1670
timestamp 1654648307
transform 1 0 56200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1723
timestamp 1654648307
transform 1 0 65200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1722
timestamp 1654648307
transform 1 0 62200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1673
timestamp 1654648307
transform 1 0 65200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1672
timestamp 1654648307
transform 1 0 62200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1725
timestamp 1654648307
transform 1 0 71200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1724
timestamp 1654648307
transform 1 0 68200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1675
timestamp 1654648307
transform 1 0 71200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1674
timestamp 1654648307
transform 1 0 68200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1727
timestamp 1654648307
transform 1 0 77200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1726
timestamp 1654648307
transform 1 0 74200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1677
timestamp 1654648307
transform 1 0 77200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1676
timestamp 1654648307
transform 1 0 74200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1729
timestamp 1654648307
transform 1 0 83200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1728
timestamp 1654648307
transform 1 0 80200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1679
timestamp 1654648307
transform 1 0 83200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1678
timestamp 1654648307
transform 1 0 80200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1731
timestamp 1654648307
transform 1 0 89200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1730
timestamp 1654648307
transform 1 0 86200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1681
timestamp 1654648307
transform 1 0 89200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1680
timestamp 1654648307
transform 1 0 86200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1732
timestamp 1654648307
transform 1 0 92200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1733
timestamp 1654648307
transform 1 0 95200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1682
timestamp 1654648307
transform 1 0 92200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1683
timestamp 1654648307
transform 1 0 95200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1734
timestamp 1654648307
transform 1 0 98200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1735
timestamp 1654648307
transform 1 0 101200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1684
timestamp 1654648307
transform 1 0 98200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1685
timestamp 1654648307
transform 1 0 101200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1736
timestamp 1654648307
transform 1 0 104200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1737
timestamp 1654648307
transform 1 0 107200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1686
timestamp 1654648307
transform 1 0 104200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1687
timestamp 1654648307
transform 1 0 107200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1738
timestamp 1654648307
transform 1 0 110200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1739
timestamp 1654648307
transform 1 0 113200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1688
timestamp 1654648307
transform 1 0 110200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1689
timestamp 1654648307
transform 1 0 113200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1740
timestamp 1654648307
transform 1 0 116200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1741
timestamp 1654648307
transform 1 0 119200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1690
timestamp 1654648307
transform 1 0 116200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1691
timestamp 1654648307
transform 1 0 119200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1742
timestamp 1654648307
transform 1 0 122200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1743
timestamp 1654648307
transform 1 0 125200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1692
timestamp 1654648307
transform 1 0 122200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1693
timestamp 1654648307
transform 1 0 125200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1744
timestamp 1654648307
transform 1 0 128200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1745
timestamp 1654648307
transform 1 0 131200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1694
timestamp 1654648307
transform 1 0 128200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1695
timestamp 1654648307
transform 1 0 131200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1746
timestamp 1654648307
transform 1 0 134200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1747
timestamp 1654648307
transform 1 0 137200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1696
timestamp 1654648307
transform 1 0 134200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1697
timestamp 1654648307
transform 1 0 137200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1748
timestamp 1654648307
transform 1 0 140200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1749
timestamp 1654648307
transform 1 0 143200 0 1 -99300
box 3640 -2860 6960 460
use pixel  pixel_1698
timestamp 1654648307
transform 1 0 140200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1699
timestamp 1654648307
transform 1 0 143200 0 1 -96300
box 3640 -2860 6960 460
use pixel  pixel_1601
timestamp 1654648307
transform 1 0 -800 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1600
timestamp 1654648307
transform 1 0 -3800 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1551
timestamp 1654648307
transform 1 0 -800 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1550
timestamp 1654648307
transform 1 0 -3800 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1603
timestamp 1654648307
transform 1 0 5200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1602
timestamp 1654648307
transform 1 0 2200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1553
timestamp 1654648307
transform 1 0 5200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1552
timestamp 1654648307
transform 1 0 2200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1605
timestamp 1654648307
transform 1 0 11200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1604
timestamp 1654648307
transform 1 0 8200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1555
timestamp 1654648307
transform 1 0 11200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1554
timestamp 1654648307
transform 1 0 8200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1607
timestamp 1654648307
transform 1 0 17200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1606
timestamp 1654648307
transform 1 0 14200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1557
timestamp 1654648307
transform 1 0 17200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1556
timestamp 1654648307
transform 1 0 14200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1609
timestamp 1654648307
transform 1 0 23200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1608
timestamp 1654648307
transform 1 0 20200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1559
timestamp 1654648307
transform 1 0 23200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1558
timestamp 1654648307
transform 1 0 20200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1611
timestamp 1654648307
transform 1 0 29200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1610
timestamp 1654648307
transform 1 0 26200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1561
timestamp 1654648307
transform 1 0 29200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1560
timestamp 1654648307
transform 1 0 26200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1613
timestamp 1654648307
transform 1 0 35200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1612
timestamp 1654648307
transform 1 0 32200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1563
timestamp 1654648307
transform 1 0 35200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1562
timestamp 1654648307
transform 1 0 32200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1615
timestamp 1654648307
transform 1 0 41200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1614
timestamp 1654648307
transform 1 0 38200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1565
timestamp 1654648307
transform 1 0 41200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1564
timestamp 1654648307
transform 1 0 38200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1617
timestamp 1654648307
transform 1 0 47200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1616
timestamp 1654648307
transform 1 0 44200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1567
timestamp 1654648307
transform 1 0 47200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1566
timestamp 1654648307
transform 1 0 44200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1619
timestamp 1654648307
transform 1 0 53200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1618
timestamp 1654648307
transform 1 0 50200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1569
timestamp 1654648307
transform 1 0 53200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1568
timestamp 1654648307
transform 1 0 50200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1621
timestamp 1654648307
transform 1 0 59200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1620
timestamp 1654648307
transform 1 0 56200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1571
timestamp 1654648307
transform 1 0 59200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1570
timestamp 1654648307
transform 1 0 56200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1623
timestamp 1654648307
transform 1 0 65200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1622
timestamp 1654648307
transform 1 0 62200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1573
timestamp 1654648307
transform 1 0 65200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1572
timestamp 1654648307
transform 1 0 62200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1625
timestamp 1654648307
transform 1 0 71200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1624
timestamp 1654648307
transform 1 0 68200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1575
timestamp 1654648307
transform 1 0 71200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1574
timestamp 1654648307
transform 1 0 68200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1627
timestamp 1654648307
transform 1 0 77200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1626
timestamp 1654648307
transform 1 0 74200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1577
timestamp 1654648307
transform 1 0 77200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1576
timestamp 1654648307
transform 1 0 74200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1629
timestamp 1654648307
transform 1 0 83200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1628
timestamp 1654648307
transform 1 0 80200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1579
timestamp 1654648307
transform 1 0 83200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1578
timestamp 1654648307
transform 1 0 80200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1631
timestamp 1654648307
transform 1 0 89200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1630
timestamp 1654648307
transform 1 0 86200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1581
timestamp 1654648307
transform 1 0 89200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1580
timestamp 1654648307
transform 1 0 86200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1632
timestamp 1654648307
transform 1 0 92200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1633
timestamp 1654648307
transform 1 0 95200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1582
timestamp 1654648307
transform 1 0 92200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1583
timestamp 1654648307
transform 1 0 95200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1634
timestamp 1654648307
transform 1 0 98200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1635
timestamp 1654648307
transform 1 0 101200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1584
timestamp 1654648307
transform 1 0 98200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1585
timestamp 1654648307
transform 1 0 101200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1636
timestamp 1654648307
transform 1 0 104200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1637
timestamp 1654648307
transform 1 0 107200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1586
timestamp 1654648307
transform 1 0 104200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1587
timestamp 1654648307
transform 1 0 107200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1638
timestamp 1654648307
transform 1 0 110200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1639
timestamp 1654648307
transform 1 0 113200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1588
timestamp 1654648307
transform 1 0 110200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1589
timestamp 1654648307
transform 1 0 113200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1640
timestamp 1654648307
transform 1 0 116200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1641
timestamp 1654648307
transform 1 0 119200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1590
timestamp 1654648307
transform 1 0 116200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1591
timestamp 1654648307
transform 1 0 119200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1642
timestamp 1654648307
transform 1 0 122200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1643
timestamp 1654648307
transform 1 0 125200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1592
timestamp 1654648307
transform 1 0 122200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1593
timestamp 1654648307
transform 1 0 125200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1644
timestamp 1654648307
transform 1 0 128200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1645
timestamp 1654648307
transform 1 0 131200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1594
timestamp 1654648307
transform 1 0 128200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1595
timestamp 1654648307
transform 1 0 131200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1646
timestamp 1654648307
transform 1 0 134200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1647
timestamp 1654648307
transform 1 0 137200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1596
timestamp 1654648307
transform 1 0 134200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1597
timestamp 1654648307
transform 1 0 137200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1648
timestamp 1654648307
transform 1 0 140200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1649
timestamp 1654648307
transform 1 0 143200 0 1 -93300
box 3640 -2860 6960 460
use pixel  pixel_1598
timestamp 1654648307
transform 1 0 140200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1599
timestamp 1654648307
transform 1 0 143200 0 1 -90300
box 3640 -2860 6960 460
use pixel  pixel_1501
timestamp 1654648307
transform 1 0 -800 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1500
timestamp 1654648307
transform 1 0 -3800 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1451
timestamp 1654648307
transform 1 0 -800 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1450
timestamp 1654648307
transform 1 0 -3800 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1503
timestamp 1654648307
transform 1 0 5200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1502
timestamp 1654648307
transform 1 0 2200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1453
timestamp 1654648307
transform 1 0 5200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1452
timestamp 1654648307
transform 1 0 2200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1505
timestamp 1654648307
transform 1 0 11200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1504
timestamp 1654648307
transform 1 0 8200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1455
timestamp 1654648307
transform 1 0 11200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1454
timestamp 1654648307
transform 1 0 8200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1507
timestamp 1654648307
transform 1 0 17200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1506
timestamp 1654648307
transform 1 0 14200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1457
timestamp 1654648307
transform 1 0 17200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1456
timestamp 1654648307
transform 1 0 14200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1509
timestamp 1654648307
transform 1 0 23200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1508
timestamp 1654648307
transform 1 0 20200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1459
timestamp 1654648307
transform 1 0 23200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1458
timestamp 1654648307
transform 1 0 20200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1511
timestamp 1654648307
transform 1 0 29200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1510
timestamp 1654648307
transform 1 0 26200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1461
timestamp 1654648307
transform 1 0 29200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1460
timestamp 1654648307
transform 1 0 26200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1513
timestamp 1654648307
transform 1 0 35200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1512
timestamp 1654648307
transform 1 0 32200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1463
timestamp 1654648307
transform 1 0 35200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1462
timestamp 1654648307
transform 1 0 32200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1515
timestamp 1654648307
transform 1 0 41200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1514
timestamp 1654648307
transform 1 0 38200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1465
timestamp 1654648307
transform 1 0 41200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1464
timestamp 1654648307
transform 1 0 38200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1517
timestamp 1654648307
transform 1 0 47200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1516
timestamp 1654648307
transform 1 0 44200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1467
timestamp 1654648307
transform 1 0 47200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1466
timestamp 1654648307
transform 1 0 44200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1519
timestamp 1654648307
transform 1 0 53200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1518
timestamp 1654648307
transform 1 0 50200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1469
timestamp 1654648307
transform 1 0 53200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1468
timestamp 1654648307
transform 1 0 50200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1521
timestamp 1654648307
transform 1 0 59200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1520
timestamp 1654648307
transform 1 0 56200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1471
timestamp 1654648307
transform 1 0 59200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1470
timestamp 1654648307
transform 1 0 56200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1523
timestamp 1654648307
transform 1 0 65200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1522
timestamp 1654648307
transform 1 0 62200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1473
timestamp 1654648307
transform 1 0 65200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1472
timestamp 1654648307
transform 1 0 62200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1525
timestamp 1654648307
transform 1 0 71200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1524
timestamp 1654648307
transform 1 0 68200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1475
timestamp 1654648307
transform 1 0 71200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1474
timestamp 1654648307
transform 1 0 68200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1527
timestamp 1654648307
transform 1 0 77200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1526
timestamp 1654648307
transform 1 0 74200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1477
timestamp 1654648307
transform 1 0 77200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1476
timestamp 1654648307
transform 1 0 74200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1529
timestamp 1654648307
transform 1 0 83200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1528
timestamp 1654648307
transform 1 0 80200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1479
timestamp 1654648307
transform 1 0 83200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1478
timestamp 1654648307
transform 1 0 80200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1531
timestamp 1654648307
transform 1 0 89200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1530
timestamp 1654648307
transform 1 0 86200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1481
timestamp 1654648307
transform 1 0 89200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1480
timestamp 1654648307
transform 1 0 86200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1532
timestamp 1654648307
transform 1 0 92200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1533
timestamp 1654648307
transform 1 0 95200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1482
timestamp 1654648307
transform 1 0 92200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1483
timestamp 1654648307
transform 1 0 95200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1534
timestamp 1654648307
transform 1 0 98200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1535
timestamp 1654648307
transform 1 0 101200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1484
timestamp 1654648307
transform 1 0 98200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1485
timestamp 1654648307
transform 1 0 101200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1536
timestamp 1654648307
transform 1 0 104200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1537
timestamp 1654648307
transform 1 0 107200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1486
timestamp 1654648307
transform 1 0 104200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1487
timestamp 1654648307
transform 1 0 107200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1538
timestamp 1654648307
transform 1 0 110200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1539
timestamp 1654648307
transform 1 0 113200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1488
timestamp 1654648307
transform 1 0 110200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1489
timestamp 1654648307
transform 1 0 113200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1540
timestamp 1654648307
transform 1 0 116200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1541
timestamp 1654648307
transform 1 0 119200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1490
timestamp 1654648307
transform 1 0 116200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1491
timestamp 1654648307
transform 1 0 119200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1542
timestamp 1654648307
transform 1 0 122200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1543
timestamp 1654648307
transform 1 0 125200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1492
timestamp 1654648307
transform 1 0 122200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1493
timestamp 1654648307
transform 1 0 125200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1544
timestamp 1654648307
transform 1 0 128200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1545
timestamp 1654648307
transform 1 0 131200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1494
timestamp 1654648307
transform 1 0 128200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1495
timestamp 1654648307
transform 1 0 131200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1546
timestamp 1654648307
transform 1 0 134200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1547
timestamp 1654648307
transform 1 0 137200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1496
timestamp 1654648307
transform 1 0 134200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1497
timestamp 1654648307
transform 1 0 137200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1548
timestamp 1654648307
transform 1 0 140200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1549
timestamp 1654648307
transform 1 0 143200 0 1 -87300
box 3640 -2860 6960 460
use pixel  pixel_1498
timestamp 1654648307
transform 1 0 140200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1499
timestamp 1654648307
transform 1 0 143200 0 1 -84300
box 3640 -2860 6960 460
use pixel  pixel_1401
timestamp 1654648307
transform 1 0 -800 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1400
timestamp 1654648307
transform 1 0 -3800 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1351
timestamp 1654648307
transform 1 0 -800 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1350
timestamp 1654648307
transform 1 0 -3800 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1403
timestamp 1654648307
transform 1 0 5200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1402
timestamp 1654648307
transform 1 0 2200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1353
timestamp 1654648307
transform 1 0 5200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1352
timestamp 1654648307
transform 1 0 2200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1405
timestamp 1654648307
transform 1 0 11200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1404
timestamp 1654648307
transform 1 0 8200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1355
timestamp 1654648307
transform 1 0 11200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1354
timestamp 1654648307
transform 1 0 8200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1407
timestamp 1654648307
transform 1 0 17200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1406
timestamp 1654648307
transform 1 0 14200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1357
timestamp 1654648307
transform 1 0 17200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1356
timestamp 1654648307
transform 1 0 14200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1409
timestamp 1654648307
transform 1 0 23200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1408
timestamp 1654648307
transform 1 0 20200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1359
timestamp 1654648307
transform 1 0 23200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1358
timestamp 1654648307
transform 1 0 20200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1411
timestamp 1654648307
transform 1 0 29200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1410
timestamp 1654648307
transform 1 0 26200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1361
timestamp 1654648307
transform 1 0 29200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1360
timestamp 1654648307
transform 1 0 26200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1413
timestamp 1654648307
transform 1 0 35200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1412
timestamp 1654648307
transform 1 0 32200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1363
timestamp 1654648307
transform 1 0 35200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1362
timestamp 1654648307
transform 1 0 32200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1415
timestamp 1654648307
transform 1 0 41200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1414
timestamp 1654648307
transform 1 0 38200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1365
timestamp 1654648307
transform 1 0 41200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1364
timestamp 1654648307
transform 1 0 38200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1417
timestamp 1654648307
transform 1 0 47200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1416
timestamp 1654648307
transform 1 0 44200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1367
timestamp 1654648307
transform 1 0 47200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1366
timestamp 1654648307
transform 1 0 44200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1419
timestamp 1654648307
transform 1 0 53200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1418
timestamp 1654648307
transform 1 0 50200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1369
timestamp 1654648307
transform 1 0 53200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1368
timestamp 1654648307
transform 1 0 50200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1421
timestamp 1654648307
transform 1 0 59200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1420
timestamp 1654648307
transform 1 0 56200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1371
timestamp 1654648307
transform 1 0 59200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1370
timestamp 1654648307
transform 1 0 56200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1423
timestamp 1654648307
transform 1 0 65200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1422
timestamp 1654648307
transform 1 0 62200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1373
timestamp 1654648307
transform 1 0 65200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1372
timestamp 1654648307
transform 1 0 62200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1425
timestamp 1654648307
transform 1 0 71200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1424
timestamp 1654648307
transform 1 0 68200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1375
timestamp 1654648307
transform 1 0 71200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1374
timestamp 1654648307
transform 1 0 68200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1427
timestamp 1654648307
transform 1 0 77200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1426
timestamp 1654648307
transform 1 0 74200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1377
timestamp 1654648307
transform 1 0 77200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1376
timestamp 1654648307
transform 1 0 74200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1429
timestamp 1654648307
transform 1 0 83200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1428
timestamp 1654648307
transform 1 0 80200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1379
timestamp 1654648307
transform 1 0 83200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1378
timestamp 1654648307
transform 1 0 80200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1431
timestamp 1654648307
transform 1 0 89200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1430
timestamp 1654648307
transform 1 0 86200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1381
timestamp 1654648307
transform 1 0 89200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1380
timestamp 1654648307
transform 1 0 86200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1432
timestamp 1654648307
transform 1 0 92200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1433
timestamp 1654648307
transform 1 0 95200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1382
timestamp 1654648307
transform 1 0 92200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1383
timestamp 1654648307
transform 1 0 95200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1434
timestamp 1654648307
transform 1 0 98200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1435
timestamp 1654648307
transform 1 0 101200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1384
timestamp 1654648307
transform 1 0 98200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1385
timestamp 1654648307
transform 1 0 101200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1436
timestamp 1654648307
transform 1 0 104200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1437
timestamp 1654648307
transform 1 0 107200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1386
timestamp 1654648307
transform 1 0 104200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1387
timestamp 1654648307
transform 1 0 107200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1438
timestamp 1654648307
transform 1 0 110200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1439
timestamp 1654648307
transform 1 0 113200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1388
timestamp 1654648307
transform 1 0 110200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1389
timestamp 1654648307
transform 1 0 113200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1440
timestamp 1654648307
transform 1 0 116200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1441
timestamp 1654648307
transform 1 0 119200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1390
timestamp 1654648307
transform 1 0 116200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1391
timestamp 1654648307
transform 1 0 119200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1442
timestamp 1654648307
transform 1 0 122200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1443
timestamp 1654648307
transform 1 0 125200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1392
timestamp 1654648307
transform 1 0 122200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1393
timestamp 1654648307
transform 1 0 125200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1444
timestamp 1654648307
transform 1 0 128200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1445
timestamp 1654648307
transform 1 0 131200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1394
timestamp 1654648307
transform 1 0 128200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1395
timestamp 1654648307
transform 1 0 131200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1446
timestamp 1654648307
transform 1 0 134200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1447
timestamp 1654648307
transform 1 0 137200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1396
timestamp 1654648307
transform 1 0 134200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1397
timestamp 1654648307
transform 1 0 137200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1448
timestamp 1654648307
transform 1 0 140200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1449
timestamp 1654648307
transform 1 0 143200 0 1 -81300
box 3640 -2860 6960 460
use pixel  pixel_1398
timestamp 1654648307
transform 1 0 140200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1399
timestamp 1654648307
transform 1 0 143200 0 1 -78300
box 3640 -2860 6960 460
use pixel  pixel_1301
timestamp 1654648307
transform 1 0 -800 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1300
timestamp 1654648307
transform 1 0 -3800 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1251
timestamp 1654648307
transform 1 0 -800 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1250
timestamp 1654648307
transform 1 0 -3800 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1303
timestamp 1654648307
transform 1 0 5200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1302
timestamp 1654648307
transform 1 0 2200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1253
timestamp 1654648307
transform 1 0 5200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1252
timestamp 1654648307
transform 1 0 2200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1305
timestamp 1654648307
transform 1 0 11200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1304
timestamp 1654648307
transform 1 0 8200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1255
timestamp 1654648307
transform 1 0 11200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1254
timestamp 1654648307
transform 1 0 8200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1307
timestamp 1654648307
transform 1 0 17200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1306
timestamp 1654648307
transform 1 0 14200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1257
timestamp 1654648307
transform 1 0 17200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1256
timestamp 1654648307
transform 1 0 14200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1309
timestamp 1654648307
transform 1 0 23200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1308
timestamp 1654648307
transform 1 0 20200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1259
timestamp 1654648307
transform 1 0 23200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1258
timestamp 1654648307
transform 1 0 20200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1311
timestamp 1654648307
transform 1 0 29200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1310
timestamp 1654648307
transform 1 0 26200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1261
timestamp 1654648307
transform 1 0 29200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1260
timestamp 1654648307
transform 1 0 26200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1313
timestamp 1654648307
transform 1 0 35200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1312
timestamp 1654648307
transform 1 0 32200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1263
timestamp 1654648307
transform 1 0 35200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1262
timestamp 1654648307
transform 1 0 32200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1315
timestamp 1654648307
transform 1 0 41200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1314
timestamp 1654648307
transform 1 0 38200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1265
timestamp 1654648307
transform 1 0 41200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1264
timestamp 1654648307
transform 1 0 38200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1317
timestamp 1654648307
transform 1 0 47200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1316
timestamp 1654648307
transform 1 0 44200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1267
timestamp 1654648307
transform 1 0 47200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1266
timestamp 1654648307
transform 1 0 44200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1319
timestamp 1654648307
transform 1 0 53200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1318
timestamp 1654648307
transform 1 0 50200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1269
timestamp 1654648307
transform 1 0 53200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1268
timestamp 1654648307
transform 1 0 50200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1321
timestamp 1654648307
transform 1 0 59200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1320
timestamp 1654648307
transform 1 0 56200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1271
timestamp 1654648307
transform 1 0 59200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1270
timestamp 1654648307
transform 1 0 56200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1323
timestamp 1654648307
transform 1 0 65200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1322
timestamp 1654648307
transform 1 0 62200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1273
timestamp 1654648307
transform 1 0 65200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1272
timestamp 1654648307
transform 1 0 62200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1325
timestamp 1654648307
transform 1 0 71200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1324
timestamp 1654648307
transform 1 0 68200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1275
timestamp 1654648307
transform 1 0 71200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1274
timestamp 1654648307
transform 1 0 68200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1327
timestamp 1654648307
transform 1 0 77200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1326
timestamp 1654648307
transform 1 0 74200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1277
timestamp 1654648307
transform 1 0 77200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1276
timestamp 1654648307
transform 1 0 74200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1329
timestamp 1654648307
transform 1 0 83200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1328
timestamp 1654648307
transform 1 0 80200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1279
timestamp 1654648307
transform 1 0 83200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1278
timestamp 1654648307
transform 1 0 80200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1331
timestamp 1654648307
transform 1 0 89200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1330
timestamp 1654648307
transform 1 0 86200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1281
timestamp 1654648307
transform 1 0 89200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1280
timestamp 1654648307
transform 1 0 86200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1332
timestamp 1654648307
transform 1 0 92200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1333
timestamp 1654648307
transform 1 0 95200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1282
timestamp 1654648307
transform 1 0 92200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1283
timestamp 1654648307
transform 1 0 95200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1334
timestamp 1654648307
transform 1 0 98200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1335
timestamp 1654648307
transform 1 0 101200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1284
timestamp 1654648307
transform 1 0 98200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1285
timestamp 1654648307
transform 1 0 101200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1336
timestamp 1654648307
transform 1 0 104200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1337
timestamp 1654648307
transform 1 0 107200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1286
timestamp 1654648307
transform 1 0 104200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1287
timestamp 1654648307
transform 1 0 107200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1338
timestamp 1654648307
transform 1 0 110200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1339
timestamp 1654648307
transform 1 0 113200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1288
timestamp 1654648307
transform 1 0 110200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1289
timestamp 1654648307
transform 1 0 113200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1340
timestamp 1654648307
transform 1 0 116200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1341
timestamp 1654648307
transform 1 0 119200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1290
timestamp 1654648307
transform 1 0 116200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1291
timestamp 1654648307
transform 1 0 119200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1342
timestamp 1654648307
transform 1 0 122200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1343
timestamp 1654648307
transform 1 0 125200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1292
timestamp 1654648307
transform 1 0 122200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1293
timestamp 1654648307
transform 1 0 125200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1344
timestamp 1654648307
transform 1 0 128200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1345
timestamp 1654648307
transform 1 0 131200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1294
timestamp 1654648307
transform 1 0 128200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1295
timestamp 1654648307
transform 1 0 131200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1346
timestamp 1654648307
transform 1 0 134200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1347
timestamp 1654648307
transform 1 0 137200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1296
timestamp 1654648307
transform 1 0 134200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1297
timestamp 1654648307
transform 1 0 137200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1348
timestamp 1654648307
transform 1 0 140200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1349
timestamp 1654648307
transform 1 0 143200 0 1 -75300
box 3640 -2860 6960 460
use pixel  pixel_1298
timestamp 1654648307
transform 1 0 140200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1299
timestamp 1654648307
transform 1 0 143200 0 1 -72300
box 3640 -2860 6960 460
use pixel  pixel_1201
timestamp 1654648307
transform 1 0 -800 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1200
timestamp 1654648307
transform 1 0 -3800 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1151
timestamp 1654648307
transform 1 0 -800 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1150
timestamp 1654648307
transform 1 0 -3800 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1203
timestamp 1654648307
transform 1 0 5200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1202
timestamp 1654648307
transform 1 0 2200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1153
timestamp 1654648307
transform 1 0 5200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1152
timestamp 1654648307
transform 1 0 2200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1205
timestamp 1654648307
transform 1 0 11200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1204
timestamp 1654648307
transform 1 0 8200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1155
timestamp 1654648307
transform 1 0 11200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1154
timestamp 1654648307
transform 1 0 8200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1207
timestamp 1654648307
transform 1 0 17200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1206
timestamp 1654648307
transform 1 0 14200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1157
timestamp 1654648307
transform 1 0 17200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1156
timestamp 1654648307
transform 1 0 14200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1209
timestamp 1654648307
transform 1 0 23200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1208
timestamp 1654648307
transform 1 0 20200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1159
timestamp 1654648307
transform 1 0 23200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1158
timestamp 1654648307
transform 1 0 20200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1211
timestamp 1654648307
transform 1 0 29200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1210
timestamp 1654648307
transform 1 0 26200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1161
timestamp 1654648307
transform 1 0 29200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1160
timestamp 1654648307
transform 1 0 26200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1213
timestamp 1654648307
transform 1 0 35200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1212
timestamp 1654648307
transform 1 0 32200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1163
timestamp 1654648307
transform 1 0 35200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1162
timestamp 1654648307
transform 1 0 32200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1214
timestamp 1654648307
transform 1 0 38200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1215
timestamp 1654648307
transform 1 0 41200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1164
timestamp 1654648307
transform 1 0 38200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1165
timestamp 1654648307
transform 1 0 41200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1216
timestamp 1654648307
transform 1 0 44200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1217
timestamp 1654648307
transform 1 0 47200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1166
timestamp 1654648307
transform 1 0 44200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1167
timestamp 1654648307
transform 1 0 47200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1218
timestamp 1654648307
transform 1 0 50200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1219
timestamp 1654648307
transform 1 0 53200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1168
timestamp 1654648307
transform 1 0 50200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1169
timestamp 1654648307
transform 1 0 53200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1220
timestamp 1654648307
transform 1 0 56200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1221
timestamp 1654648307
transform 1 0 59200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1170
timestamp 1654648307
transform 1 0 56200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1171
timestamp 1654648307
transform 1 0 59200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1222
timestamp 1654648307
transform 1 0 62200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1223
timestamp 1654648307
transform 1 0 65200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1172
timestamp 1654648307
transform 1 0 62200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1173
timestamp 1654648307
transform 1 0 65200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1224
timestamp 1654648307
transform 1 0 68200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1225
timestamp 1654648307
transform 1 0 71200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1174
timestamp 1654648307
transform 1 0 68200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1175
timestamp 1654648307
transform 1 0 71200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1226
timestamp 1654648307
transform 1 0 74200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1227
timestamp 1654648307
transform 1 0 77200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1176
timestamp 1654648307
transform 1 0 74200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1177
timestamp 1654648307
transform 1 0 77200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1228
timestamp 1654648307
transform 1 0 80200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1229
timestamp 1654648307
transform 1 0 83200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1178
timestamp 1654648307
transform 1 0 80200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1179
timestamp 1654648307
transform 1 0 83200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1230
timestamp 1654648307
transform 1 0 86200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1231
timestamp 1654648307
transform 1 0 89200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1180
timestamp 1654648307
transform 1 0 86200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1181
timestamp 1654648307
transform 1 0 89200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1232
timestamp 1654648307
transform 1 0 92200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1233
timestamp 1654648307
transform 1 0 95200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1182
timestamp 1654648307
transform 1 0 92200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1183
timestamp 1654648307
transform 1 0 95200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1234
timestamp 1654648307
transform 1 0 98200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1235
timestamp 1654648307
transform 1 0 101200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1184
timestamp 1654648307
transform 1 0 98200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1185
timestamp 1654648307
transform 1 0 101200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1236
timestamp 1654648307
transform 1 0 104200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1237
timestamp 1654648307
transform 1 0 107200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1186
timestamp 1654648307
transform 1 0 104200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1187
timestamp 1654648307
transform 1 0 107200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1238
timestamp 1654648307
transform 1 0 110200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1239
timestamp 1654648307
transform 1 0 113200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1188
timestamp 1654648307
transform 1 0 110200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1189
timestamp 1654648307
transform 1 0 113200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1240
timestamp 1654648307
transform 1 0 116200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1241
timestamp 1654648307
transform 1 0 119200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1190
timestamp 1654648307
transform 1 0 116200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1191
timestamp 1654648307
transform 1 0 119200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1242
timestamp 1654648307
transform 1 0 122200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1243
timestamp 1654648307
transform 1 0 125200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1192
timestamp 1654648307
transform 1 0 122200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1193
timestamp 1654648307
transform 1 0 125200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1244
timestamp 1654648307
transform 1 0 128200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1245
timestamp 1654648307
transform 1 0 131200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1194
timestamp 1654648307
transform 1 0 128200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1195
timestamp 1654648307
transform 1 0 131200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1246
timestamp 1654648307
transform 1 0 134200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1247
timestamp 1654648307
transform 1 0 137200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1196
timestamp 1654648307
transform 1 0 134200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1197
timestamp 1654648307
transform 1 0 137200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1248
timestamp 1654648307
transform 1 0 140200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1249
timestamp 1654648307
transform 1 0 143200 0 1 -69300
box 3640 -2860 6960 460
use pixel  pixel_1198
timestamp 1654648307
transform 1 0 140200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1199
timestamp 1654648307
transform 1 0 143200 0 1 -66300
box 3640 -2860 6960 460
use pixel  pixel_1101
timestamp 1654648307
transform 1 0 -800 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1100
timestamp 1654648307
transform 1 0 -3800 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1051
timestamp 1654648307
transform 1 0 -800 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1050
timestamp 1654648307
transform 1 0 -3800 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1103
timestamp 1654648307
transform 1 0 5200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1102
timestamp 1654648307
transform 1 0 2200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1053
timestamp 1654648307
transform 1 0 5200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1052
timestamp 1654648307
transform 1 0 2200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1105
timestamp 1654648307
transform 1 0 11200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1104
timestamp 1654648307
transform 1 0 8200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1055
timestamp 1654648307
transform 1 0 11200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1054
timestamp 1654648307
transform 1 0 8200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1107
timestamp 1654648307
transform 1 0 17200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1106
timestamp 1654648307
transform 1 0 14200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1057
timestamp 1654648307
transform 1 0 17200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1056
timestamp 1654648307
transform 1 0 14200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1109
timestamp 1654648307
transform 1 0 23200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1108
timestamp 1654648307
transform 1 0 20200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1059
timestamp 1654648307
transform 1 0 23200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1058
timestamp 1654648307
transform 1 0 20200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1111
timestamp 1654648307
transform 1 0 29200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1110
timestamp 1654648307
transform 1 0 26200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1061
timestamp 1654648307
transform 1 0 29200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1060
timestamp 1654648307
transform 1 0 26200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1113
timestamp 1654648307
transform 1 0 35200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1112
timestamp 1654648307
transform 1 0 32200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1063
timestamp 1654648307
transform 1 0 35200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1062
timestamp 1654648307
transform 1 0 32200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1114
timestamp 1654648307
transform 1 0 38200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1115
timestamp 1654648307
transform 1 0 41200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1064
timestamp 1654648307
transform 1 0 38200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1065
timestamp 1654648307
transform 1 0 41200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1116
timestamp 1654648307
transform 1 0 44200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1117
timestamp 1654648307
transform 1 0 47200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1066
timestamp 1654648307
transform 1 0 44200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1067
timestamp 1654648307
transform 1 0 47200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1118
timestamp 1654648307
transform 1 0 50200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1119
timestamp 1654648307
transform 1 0 53200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1068
timestamp 1654648307
transform 1 0 50200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1069
timestamp 1654648307
transform 1 0 53200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1120
timestamp 1654648307
transform 1 0 56200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1121
timestamp 1654648307
transform 1 0 59200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1070
timestamp 1654648307
transform 1 0 56200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1071
timestamp 1654648307
transform 1 0 59200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1122
timestamp 1654648307
transform 1 0 62200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1123
timestamp 1654648307
transform 1 0 65200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1072
timestamp 1654648307
transform 1 0 62200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1073
timestamp 1654648307
transform 1 0 65200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1124
timestamp 1654648307
transform 1 0 68200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1125
timestamp 1654648307
transform 1 0 71200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1074
timestamp 1654648307
transform 1 0 68200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1075
timestamp 1654648307
transform 1 0 71200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1126
timestamp 1654648307
transform 1 0 74200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1127
timestamp 1654648307
transform 1 0 77200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1076
timestamp 1654648307
transform 1 0 74200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1077
timestamp 1654648307
transform 1 0 77200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1128
timestamp 1654648307
transform 1 0 80200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1129
timestamp 1654648307
transform 1 0 83200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1078
timestamp 1654648307
transform 1 0 80200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1079
timestamp 1654648307
transform 1 0 83200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1130
timestamp 1654648307
transform 1 0 86200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1131
timestamp 1654648307
transform 1 0 89200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1080
timestamp 1654648307
transform 1 0 86200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1081
timestamp 1654648307
transform 1 0 89200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1132
timestamp 1654648307
transform 1 0 92200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1133
timestamp 1654648307
transform 1 0 95200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1082
timestamp 1654648307
transform 1 0 92200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1083
timestamp 1654648307
transform 1 0 95200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1134
timestamp 1654648307
transform 1 0 98200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1135
timestamp 1654648307
transform 1 0 101200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1084
timestamp 1654648307
transform 1 0 98200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1085
timestamp 1654648307
transform 1 0 101200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1136
timestamp 1654648307
transform 1 0 104200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1137
timestamp 1654648307
transform 1 0 107200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1086
timestamp 1654648307
transform 1 0 104200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1087
timestamp 1654648307
transform 1 0 107200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1138
timestamp 1654648307
transform 1 0 110200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1139
timestamp 1654648307
transform 1 0 113200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1088
timestamp 1654648307
transform 1 0 110200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1089
timestamp 1654648307
transform 1 0 113200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1140
timestamp 1654648307
transform 1 0 116200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1141
timestamp 1654648307
transform 1 0 119200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1090
timestamp 1654648307
transform 1 0 116200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1091
timestamp 1654648307
transform 1 0 119200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1142
timestamp 1654648307
transform 1 0 122200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1143
timestamp 1654648307
transform 1 0 125200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1092
timestamp 1654648307
transform 1 0 122200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1093
timestamp 1654648307
transform 1 0 125200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1144
timestamp 1654648307
transform 1 0 128200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1145
timestamp 1654648307
transform 1 0 131200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1094
timestamp 1654648307
transform 1 0 128200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1095
timestamp 1654648307
transform 1 0 131200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1146
timestamp 1654648307
transform 1 0 134200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1147
timestamp 1654648307
transform 1 0 137200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1096
timestamp 1654648307
transform 1 0 134200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1097
timestamp 1654648307
transform 1 0 137200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1148
timestamp 1654648307
transform 1 0 140200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1149
timestamp 1654648307
transform 1 0 143200 0 1 -63300
box 3640 -2860 6960 460
use pixel  pixel_1098
timestamp 1654648307
transform 1 0 140200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1099
timestamp 1654648307
transform 1 0 143200 0 1 -60300
box 3640 -2860 6960 460
use pixel  pixel_1001
timestamp 1654648307
transform 1 0 -800 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_1000
timestamp 1654648307
transform 1 0 -3800 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_951
timestamp 1654648307
transform 1 0 -800 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_950
timestamp 1654648307
transform 1 0 -3800 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1003
timestamp 1654648307
transform 1 0 5200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_1002
timestamp 1654648307
transform 1 0 2200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_953
timestamp 1654648307
transform 1 0 5200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_952
timestamp 1654648307
transform 1 0 2200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1005
timestamp 1654648307
transform 1 0 11200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_1004
timestamp 1654648307
transform 1 0 8200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_955
timestamp 1654648307
transform 1 0 11200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_954
timestamp 1654648307
transform 1 0 8200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1007
timestamp 1654648307
transform 1 0 17200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_1006
timestamp 1654648307
transform 1 0 14200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_957
timestamp 1654648307
transform 1 0 17200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_956
timestamp 1654648307
transform 1 0 14200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1009
timestamp 1654648307
transform 1 0 23200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_1008
timestamp 1654648307
transform 1 0 20200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_959
timestamp 1654648307
transform 1 0 23200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_958
timestamp 1654648307
transform 1 0 20200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1011
timestamp 1654648307
transform 1 0 29200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_1010
timestamp 1654648307
transform 1 0 26200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_961
timestamp 1654648307
transform 1 0 29200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_960
timestamp 1654648307
transform 1 0 26200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1013
timestamp 1654648307
transform 1 0 35200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_1012
timestamp 1654648307
transform 1 0 32200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_963
timestamp 1654648307
transform 1 0 35200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_962
timestamp 1654648307
transform 1 0 32200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1014
timestamp 1654648307
transform 1 0 38200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_1015
timestamp 1654648307
transform 1 0 41200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_964
timestamp 1654648307
transform 1 0 38200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_965
timestamp 1654648307
transform 1 0 41200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1016
timestamp 1654648307
transform 1 0 44200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_1017
timestamp 1654648307
transform 1 0 47200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_966
timestamp 1654648307
transform 1 0 44200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_967
timestamp 1654648307
transform 1 0 47200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1018
timestamp 1654648307
transform 1 0 50200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_1019
timestamp 1654648307
transform 1 0 53200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_968
timestamp 1654648307
transform 1 0 50200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_969
timestamp 1654648307
transform 1 0 53200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1020
timestamp 1654648307
transform 1 0 56200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_1021
timestamp 1654648307
transform 1 0 59200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_970
timestamp 1654648307
transform 1 0 56200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_971
timestamp 1654648307
transform 1 0 59200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1022
timestamp 1654648307
transform 1 0 62200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_1023
timestamp 1654648307
transform 1 0 65200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_972
timestamp 1654648307
transform 1 0 62200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_973
timestamp 1654648307
transform 1 0 65200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1024
timestamp 1654648307
transform 1 0 68200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_1025
timestamp 1654648307
transform 1 0 71200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_974
timestamp 1654648307
transform 1 0 68200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_975
timestamp 1654648307
transform 1 0 71200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1026
timestamp 1654648307
transform 1 0 74200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_1027
timestamp 1654648307
transform 1 0 77200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_976
timestamp 1654648307
transform 1 0 74200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_977
timestamp 1654648307
transform 1 0 77200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1028
timestamp 1654648307
transform 1 0 80200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_1029
timestamp 1654648307
transform 1 0 83200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_978
timestamp 1654648307
transform 1 0 80200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_979
timestamp 1654648307
transform 1 0 83200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1030
timestamp 1654648307
transform 1 0 86200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_1031
timestamp 1654648307
transform 1 0 89200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_980
timestamp 1654648307
transform 1 0 86200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_981
timestamp 1654648307
transform 1 0 89200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1032
timestamp 1654648307
transform 1 0 92200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_1033
timestamp 1654648307
transform 1 0 95200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_982
timestamp 1654648307
transform 1 0 92200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_983
timestamp 1654648307
transform 1 0 95200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1034
timestamp 1654648307
transform 1 0 98200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_1035
timestamp 1654648307
transform 1 0 101200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_984
timestamp 1654648307
transform 1 0 98200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_985
timestamp 1654648307
transform 1 0 101200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1036
timestamp 1654648307
transform 1 0 104200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_1037
timestamp 1654648307
transform 1 0 107200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_986
timestamp 1654648307
transform 1 0 104200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_987
timestamp 1654648307
transform 1 0 107200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1038
timestamp 1654648307
transform 1 0 110200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_1039
timestamp 1654648307
transform 1 0 113200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_988
timestamp 1654648307
transform 1 0 110200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_989
timestamp 1654648307
transform 1 0 113200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1040
timestamp 1654648307
transform 1 0 116200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_1041
timestamp 1654648307
transform 1 0 119200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_990
timestamp 1654648307
transform 1 0 116200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_991
timestamp 1654648307
transform 1 0 119200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1042
timestamp 1654648307
transform 1 0 122200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_1043
timestamp 1654648307
transform 1 0 125200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_992
timestamp 1654648307
transform 1 0 122200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_993
timestamp 1654648307
transform 1 0 125200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1044
timestamp 1654648307
transform 1 0 128200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_1045
timestamp 1654648307
transform 1 0 131200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_994
timestamp 1654648307
transform 1 0 128200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_995
timestamp 1654648307
transform 1 0 131200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1046
timestamp 1654648307
transform 1 0 134200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_1047
timestamp 1654648307
transform 1 0 137200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_996
timestamp 1654648307
transform 1 0 134200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_997
timestamp 1654648307
transform 1 0 137200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_1048
timestamp 1654648307
transform 1 0 140200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_1049
timestamp 1654648307
transform 1 0 143200 0 1 -57300
box 3640 -2860 6960 460
use pixel  pixel_998
timestamp 1654648307
transform 1 0 140200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_999
timestamp 1654648307
transform 1 0 143200 0 1 -54300
box 3640 -2860 6960 460
use pixel  pixel_901
timestamp 1654648307
transform 1 0 -800 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_900
timestamp 1654648307
transform 1 0 -3800 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_851
timestamp 1654648307
transform 1 0 -800 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_850
timestamp 1654648307
transform 1 0 -3800 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_903
timestamp 1654648307
transform 1 0 5200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_902
timestamp 1654648307
transform 1 0 2200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_853
timestamp 1654648307
transform 1 0 5200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_852
timestamp 1654648307
transform 1 0 2200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_905
timestamp 1654648307
transform 1 0 11200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_904
timestamp 1654648307
transform 1 0 8200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_855
timestamp 1654648307
transform 1 0 11200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_854
timestamp 1654648307
transform 1 0 8200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_907
timestamp 1654648307
transform 1 0 17200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_906
timestamp 1654648307
transform 1 0 14200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_857
timestamp 1654648307
transform 1 0 17200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_856
timestamp 1654648307
transform 1 0 14200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_909
timestamp 1654648307
transform 1 0 23200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_908
timestamp 1654648307
transform 1 0 20200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_859
timestamp 1654648307
transform 1 0 23200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_858
timestamp 1654648307
transform 1 0 20200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_911
timestamp 1654648307
transform 1 0 29200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_910
timestamp 1654648307
transform 1 0 26200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_861
timestamp 1654648307
transform 1 0 29200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_860
timestamp 1654648307
transform 1 0 26200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_913
timestamp 1654648307
transform 1 0 35200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_912
timestamp 1654648307
transform 1 0 32200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_863
timestamp 1654648307
transform 1 0 35200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_862
timestamp 1654648307
transform 1 0 32200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_914
timestamp 1654648307
transform 1 0 38200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_915
timestamp 1654648307
transform 1 0 41200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_864
timestamp 1654648307
transform 1 0 38200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_865
timestamp 1654648307
transform 1 0 41200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_916
timestamp 1654648307
transform 1 0 44200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_917
timestamp 1654648307
transform 1 0 47200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_866
timestamp 1654648307
transform 1 0 44200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_867
timestamp 1654648307
transform 1 0 47200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_918
timestamp 1654648307
transform 1 0 50200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_919
timestamp 1654648307
transform 1 0 53200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_868
timestamp 1654648307
transform 1 0 50200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_869
timestamp 1654648307
transform 1 0 53200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_920
timestamp 1654648307
transform 1 0 56200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_921
timestamp 1654648307
transform 1 0 59200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_870
timestamp 1654648307
transform 1 0 56200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_871
timestamp 1654648307
transform 1 0 59200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_922
timestamp 1654648307
transform 1 0 62200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_923
timestamp 1654648307
transform 1 0 65200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_872
timestamp 1654648307
transform 1 0 62200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_873
timestamp 1654648307
transform 1 0 65200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_924
timestamp 1654648307
transform 1 0 68200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_925
timestamp 1654648307
transform 1 0 71200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_874
timestamp 1654648307
transform 1 0 68200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_875
timestamp 1654648307
transform 1 0 71200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_926
timestamp 1654648307
transform 1 0 74200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_927
timestamp 1654648307
transform 1 0 77200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_876
timestamp 1654648307
transform 1 0 74200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_877
timestamp 1654648307
transform 1 0 77200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_928
timestamp 1654648307
transform 1 0 80200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_929
timestamp 1654648307
transform 1 0 83200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_878
timestamp 1654648307
transform 1 0 80200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_879
timestamp 1654648307
transform 1 0 83200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_930
timestamp 1654648307
transform 1 0 86200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_931
timestamp 1654648307
transform 1 0 89200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_880
timestamp 1654648307
transform 1 0 86200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_881
timestamp 1654648307
transform 1 0 89200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_932
timestamp 1654648307
transform 1 0 92200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_933
timestamp 1654648307
transform 1 0 95200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_882
timestamp 1654648307
transform 1 0 92200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_883
timestamp 1654648307
transform 1 0 95200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_934
timestamp 1654648307
transform 1 0 98200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_935
timestamp 1654648307
transform 1 0 101200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_884
timestamp 1654648307
transform 1 0 98200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_885
timestamp 1654648307
transform 1 0 101200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_936
timestamp 1654648307
transform 1 0 104200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_937
timestamp 1654648307
transform 1 0 107200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_886
timestamp 1654648307
transform 1 0 104200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_887
timestamp 1654648307
transform 1 0 107200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_938
timestamp 1654648307
transform 1 0 110200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_939
timestamp 1654648307
transform 1 0 113200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_888
timestamp 1654648307
transform 1 0 110200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_889
timestamp 1654648307
transform 1 0 113200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_940
timestamp 1654648307
transform 1 0 116200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_941
timestamp 1654648307
transform 1 0 119200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_890
timestamp 1654648307
transform 1 0 116200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_891
timestamp 1654648307
transform 1 0 119200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_942
timestamp 1654648307
transform 1 0 122200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_943
timestamp 1654648307
transform 1 0 125200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_892
timestamp 1654648307
transform 1 0 122200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_893
timestamp 1654648307
transform 1 0 125200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_944
timestamp 1654648307
transform 1 0 128200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_945
timestamp 1654648307
transform 1 0 131200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_894
timestamp 1654648307
transform 1 0 128200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_895
timestamp 1654648307
transform 1 0 131200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_946
timestamp 1654648307
transform 1 0 134200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_947
timestamp 1654648307
transform 1 0 137200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_896
timestamp 1654648307
transform 1 0 134200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_897
timestamp 1654648307
transform 1 0 137200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_948
timestamp 1654648307
transform 1 0 140200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_949
timestamp 1654648307
transform 1 0 143200 0 1 -51300
box 3640 -2860 6960 460
use pixel  pixel_898
timestamp 1654648307
transform 1 0 140200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_899
timestamp 1654648307
transform 1 0 143200 0 1 -48300
box 3640 -2860 6960 460
use pixel  pixel_801
timestamp 1654648307
transform 1 0 -800 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_800
timestamp 1654648307
transform 1 0 -3800 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_750
timestamp 1654648307
transform 1 0 -3800 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_751
timestamp 1654648307
transform 1 0 -800 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_803
timestamp 1654648307
transform 1 0 5200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_802
timestamp 1654648307
transform 1 0 2200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_752
timestamp 1654648307
transform 1 0 2200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_753
timestamp 1654648307
transform 1 0 5200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_805
timestamp 1654648307
transform 1 0 11200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_804
timestamp 1654648307
transform 1 0 8200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_754
timestamp 1654648307
transform 1 0 8200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_755
timestamp 1654648307
transform 1 0 11200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_807
timestamp 1654648307
transform 1 0 17200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_806
timestamp 1654648307
transform 1 0 14200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_756
timestamp 1654648307
transform 1 0 14200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_757
timestamp 1654648307
transform 1 0 17200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_809
timestamp 1654648307
transform 1 0 23200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_808
timestamp 1654648307
transform 1 0 20200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_758
timestamp 1654648307
transform 1 0 20200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_759
timestamp 1654648307
transform 1 0 23200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_811
timestamp 1654648307
transform 1 0 29200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_810
timestamp 1654648307
transform 1 0 26200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_760
timestamp 1654648307
transform 1 0 26200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_761
timestamp 1654648307
transform 1 0 29200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_813
timestamp 1654648307
transform 1 0 35200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_812
timestamp 1654648307
transform 1 0 32200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_762
timestamp 1654648307
transform 1 0 32200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_763
timestamp 1654648307
transform 1 0 35200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_814
timestamp 1654648307
transform 1 0 38200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_815
timestamp 1654648307
transform 1 0 41200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_764
timestamp 1654648307
transform 1 0 38200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_765
timestamp 1654648307
transform 1 0 41200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_816
timestamp 1654648307
transform 1 0 44200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_817
timestamp 1654648307
transform 1 0 47200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_766
timestamp 1654648307
transform 1 0 44200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_767
timestamp 1654648307
transform 1 0 47200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_818
timestamp 1654648307
transform 1 0 50200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_819
timestamp 1654648307
transform 1 0 53200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_768
timestamp 1654648307
transform 1 0 50200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_769
timestamp 1654648307
transform 1 0 53200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_820
timestamp 1654648307
transform 1 0 56200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_821
timestamp 1654648307
transform 1 0 59200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_770
timestamp 1654648307
transform 1 0 56200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_771
timestamp 1654648307
transform 1 0 59200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_822
timestamp 1654648307
transform 1 0 62200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_823
timestamp 1654648307
transform 1 0 65200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_772
timestamp 1654648307
transform 1 0 62200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_773
timestamp 1654648307
transform 1 0 65200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_824
timestamp 1654648307
transform 1 0 68200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_825
timestamp 1654648307
transform 1 0 71200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_774
timestamp 1654648307
transform 1 0 68200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_775
timestamp 1654648307
transform 1 0 71200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_826
timestamp 1654648307
transform 1 0 74200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_827
timestamp 1654648307
transform 1 0 77200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_776
timestamp 1654648307
transform 1 0 74200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_777
timestamp 1654648307
transform 1 0 77200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_828
timestamp 1654648307
transform 1 0 80200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_829
timestamp 1654648307
transform 1 0 83200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_778
timestamp 1654648307
transform 1 0 80200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_779
timestamp 1654648307
transform 1 0 83200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_830
timestamp 1654648307
transform 1 0 86200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_831
timestamp 1654648307
transform 1 0 89200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_780
timestamp 1654648307
transform 1 0 86200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_781
timestamp 1654648307
transform 1 0 89200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_832
timestamp 1654648307
transform 1 0 92200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_833
timestamp 1654648307
transform 1 0 95200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_782
timestamp 1654648307
transform 1 0 92200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_783
timestamp 1654648307
transform 1 0 95200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_834
timestamp 1654648307
transform 1 0 98200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_835
timestamp 1654648307
transform 1 0 101200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_784
timestamp 1654648307
transform 1 0 98200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_785
timestamp 1654648307
transform 1 0 101200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_836
timestamp 1654648307
transform 1 0 104200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_837
timestamp 1654648307
transform 1 0 107200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_786
timestamp 1654648307
transform 1 0 104200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_787
timestamp 1654648307
transform 1 0 107200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_838
timestamp 1654648307
transform 1 0 110200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_839
timestamp 1654648307
transform 1 0 113200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_788
timestamp 1654648307
transform 1 0 110200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_789
timestamp 1654648307
transform 1 0 113200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_840
timestamp 1654648307
transform 1 0 116200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_841
timestamp 1654648307
transform 1 0 119200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_790
timestamp 1654648307
transform 1 0 116200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_791
timestamp 1654648307
transform 1 0 119200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_842
timestamp 1654648307
transform 1 0 122200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_843
timestamp 1654648307
transform 1 0 125200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_792
timestamp 1654648307
transform 1 0 122200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_793
timestamp 1654648307
transform 1 0 125200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_844
timestamp 1654648307
transform 1 0 128200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_845
timestamp 1654648307
transform 1 0 131200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_794
timestamp 1654648307
transform 1 0 128200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_795
timestamp 1654648307
transform 1 0 131200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_846
timestamp 1654648307
transform 1 0 134200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_847
timestamp 1654648307
transform 1 0 137200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_796
timestamp 1654648307
transform 1 0 134200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_797
timestamp 1654648307
transform 1 0 137200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_848
timestamp 1654648307
transform 1 0 140200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_849
timestamp 1654648307
transform 1 0 143200 0 1 -45300
box 3640 -2860 6960 460
use pixel  pixel_798
timestamp 1654648307
transform 1 0 140200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_799
timestamp 1654648307
transform 1 0 143200 0 1 -42300
box 3640 -2860 6960 460
use pixel  pixel_700
timestamp 1654648307
transform 1 0 -3800 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_701
timestamp 1654648307
transform 1 0 -800 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_650
timestamp 1654648307
transform 1 0 -3800 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_651
timestamp 1654648307
transform 1 0 -800 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_702
timestamp 1654648307
transform 1 0 2200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_703
timestamp 1654648307
transform 1 0 5200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_652
timestamp 1654648307
transform 1 0 2200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_653
timestamp 1654648307
transform 1 0 5200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_704
timestamp 1654648307
transform 1 0 8200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_705
timestamp 1654648307
transform 1 0 11200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_654
timestamp 1654648307
transform 1 0 8200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_655
timestamp 1654648307
transform 1 0 11200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_706
timestamp 1654648307
transform 1 0 14200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_707
timestamp 1654648307
transform 1 0 17200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_656
timestamp 1654648307
transform 1 0 14200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_657
timestamp 1654648307
transform 1 0 17200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_708
timestamp 1654648307
transform 1 0 20200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_709
timestamp 1654648307
transform 1 0 23200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_658
timestamp 1654648307
transform 1 0 20200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_659
timestamp 1654648307
transform 1 0 23200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_710
timestamp 1654648307
transform 1 0 26200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_711
timestamp 1654648307
transform 1 0 29200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_660
timestamp 1654648307
transform 1 0 26200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_661
timestamp 1654648307
transform 1 0 29200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_712
timestamp 1654648307
transform 1 0 32200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_713
timestamp 1654648307
transform 1 0 35200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_662
timestamp 1654648307
transform 1 0 32200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_663
timestamp 1654648307
transform 1 0 35200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_714
timestamp 1654648307
transform 1 0 38200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_715
timestamp 1654648307
transform 1 0 41200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_664
timestamp 1654648307
transform 1 0 38200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_665
timestamp 1654648307
transform 1 0 41200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_716
timestamp 1654648307
transform 1 0 44200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_717
timestamp 1654648307
transform 1 0 47200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_666
timestamp 1654648307
transform 1 0 44200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_667
timestamp 1654648307
transform 1 0 47200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_718
timestamp 1654648307
transform 1 0 50200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_719
timestamp 1654648307
transform 1 0 53200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_668
timestamp 1654648307
transform 1 0 50200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_669
timestamp 1654648307
transform 1 0 53200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_720
timestamp 1654648307
transform 1 0 56200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_721
timestamp 1654648307
transform 1 0 59200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_670
timestamp 1654648307
transform 1 0 56200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_671
timestamp 1654648307
transform 1 0 59200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_722
timestamp 1654648307
transform 1 0 62200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_723
timestamp 1654648307
transform 1 0 65200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_672
timestamp 1654648307
transform 1 0 62200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_673
timestamp 1654648307
transform 1 0 65200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_724
timestamp 1654648307
transform 1 0 68200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_725
timestamp 1654648307
transform 1 0 71200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_674
timestamp 1654648307
transform 1 0 68200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_675
timestamp 1654648307
transform 1 0 71200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_726
timestamp 1654648307
transform 1 0 74200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_727
timestamp 1654648307
transform 1 0 77200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_676
timestamp 1654648307
transform 1 0 74200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_677
timestamp 1654648307
transform 1 0 77200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_728
timestamp 1654648307
transform 1 0 80200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_729
timestamp 1654648307
transform 1 0 83200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_678
timestamp 1654648307
transform 1 0 80200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_679
timestamp 1654648307
transform 1 0 83200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_730
timestamp 1654648307
transform 1 0 86200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_731
timestamp 1654648307
transform 1 0 89200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_680
timestamp 1654648307
transform 1 0 86200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_681
timestamp 1654648307
transform 1 0 89200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_732
timestamp 1654648307
transform 1 0 92200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_733
timestamp 1654648307
transform 1 0 95200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_682
timestamp 1654648307
transform 1 0 92200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_683
timestamp 1654648307
transform 1 0 95200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_734
timestamp 1654648307
transform 1 0 98200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_735
timestamp 1654648307
transform 1 0 101200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_684
timestamp 1654648307
transform 1 0 98200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_685
timestamp 1654648307
transform 1 0 101200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_736
timestamp 1654648307
transform 1 0 104200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_737
timestamp 1654648307
transform 1 0 107200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_686
timestamp 1654648307
transform 1 0 104200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_687
timestamp 1654648307
transform 1 0 107200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_738
timestamp 1654648307
transform 1 0 110200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_739
timestamp 1654648307
transform 1 0 113200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_688
timestamp 1654648307
transform 1 0 110200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_689
timestamp 1654648307
transform 1 0 113200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_740
timestamp 1654648307
transform 1 0 116200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_741
timestamp 1654648307
transform 1 0 119200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_690
timestamp 1654648307
transform 1 0 116200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_691
timestamp 1654648307
transform 1 0 119200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_742
timestamp 1654648307
transform 1 0 122200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_743
timestamp 1654648307
transform 1 0 125200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_692
timestamp 1654648307
transform 1 0 122200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_693
timestamp 1654648307
transform 1 0 125200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_744
timestamp 1654648307
transform 1 0 128200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_745
timestamp 1654648307
transform 1 0 131200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_694
timestamp 1654648307
transform 1 0 128200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_695
timestamp 1654648307
transform 1 0 131200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_746
timestamp 1654648307
transform 1 0 134200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_747
timestamp 1654648307
transform 1 0 137200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_696
timestamp 1654648307
transform 1 0 134200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_697
timestamp 1654648307
transform 1 0 137200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_748
timestamp 1654648307
transform 1 0 140200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_749
timestamp 1654648307
transform 1 0 143200 0 1 -39300
box 3640 -2860 6960 460
use pixel  pixel_698
timestamp 1654648307
transform 1 0 140200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_699
timestamp 1654648307
transform 1 0 143200 0 1 -36300
box 3640 -2860 6960 460
use pixel  pixel_600
timestamp 1654648307
transform 1 0 -3800 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_601
timestamp 1654648307
transform 1 0 -800 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_550
timestamp 1654648307
transform 1 0 -3800 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_551
timestamp 1654648307
transform 1 0 -800 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_602
timestamp 1654648307
transform 1 0 2200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_603
timestamp 1654648307
transform 1 0 5200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_552
timestamp 1654648307
transform 1 0 2200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_553
timestamp 1654648307
transform 1 0 5200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_604
timestamp 1654648307
transform 1 0 8200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_605
timestamp 1654648307
transform 1 0 11200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_554
timestamp 1654648307
transform 1 0 8200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_555
timestamp 1654648307
transform 1 0 11200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_606
timestamp 1654648307
transform 1 0 14200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_607
timestamp 1654648307
transform 1 0 17200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_556
timestamp 1654648307
transform 1 0 14200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_557
timestamp 1654648307
transform 1 0 17200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_608
timestamp 1654648307
transform 1 0 20200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_609
timestamp 1654648307
transform 1 0 23200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_558
timestamp 1654648307
transform 1 0 20200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_559
timestamp 1654648307
transform 1 0 23200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_610
timestamp 1654648307
transform 1 0 26200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_611
timestamp 1654648307
transform 1 0 29200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_560
timestamp 1654648307
transform 1 0 26200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_561
timestamp 1654648307
transform 1 0 29200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_612
timestamp 1654648307
transform 1 0 32200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_613
timestamp 1654648307
transform 1 0 35200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_562
timestamp 1654648307
transform 1 0 32200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_563
timestamp 1654648307
transform 1 0 35200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_614
timestamp 1654648307
transform 1 0 38200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_615
timestamp 1654648307
transform 1 0 41200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_564
timestamp 1654648307
transform 1 0 38200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_565
timestamp 1654648307
transform 1 0 41200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_616
timestamp 1654648307
transform 1 0 44200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_617
timestamp 1654648307
transform 1 0 47200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_566
timestamp 1654648307
transform 1 0 44200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_567
timestamp 1654648307
transform 1 0 47200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_618
timestamp 1654648307
transform 1 0 50200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_619
timestamp 1654648307
transform 1 0 53200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_568
timestamp 1654648307
transform 1 0 50200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_569
timestamp 1654648307
transform 1 0 53200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_620
timestamp 1654648307
transform 1 0 56200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_621
timestamp 1654648307
transform 1 0 59200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_570
timestamp 1654648307
transform 1 0 56200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_571
timestamp 1654648307
transform 1 0 59200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_622
timestamp 1654648307
transform 1 0 62200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_623
timestamp 1654648307
transform 1 0 65200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_572
timestamp 1654648307
transform 1 0 62200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_573
timestamp 1654648307
transform 1 0 65200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_624
timestamp 1654648307
transform 1 0 68200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_625
timestamp 1654648307
transform 1 0 71200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_574
timestamp 1654648307
transform 1 0 68200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_575
timestamp 1654648307
transform 1 0 71200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_626
timestamp 1654648307
transform 1 0 74200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_627
timestamp 1654648307
transform 1 0 77200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_576
timestamp 1654648307
transform 1 0 74200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_577
timestamp 1654648307
transform 1 0 77200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_628
timestamp 1654648307
transform 1 0 80200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_629
timestamp 1654648307
transform 1 0 83200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_578
timestamp 1654648307
transform 1 0 80200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_579
timestamp 1654648307
transform 1 0 83200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_630
timestamp 1654648307
transform 1 0 86200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_631
timestamp 1654648307
transform 1 0 89200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_580
timestamp 1654648307
transform 1 0 86200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_581
timestamp 1654648307
transform 1 0 89200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_632
timestamp 1654648307
transform 1 0 92200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_633
timestamp 1654648307
transform 1 0 95200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_582
timestamp 1654648307
transform 1 0 92200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_583
timestamp 1654648307
transform 1 0 95200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_634
timestamp 1654648307
transform 1 0 98200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_635
timestamp 1654648307
transform 1 0 101200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_584
timestamp 1654648307
transform 1 0 98200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_585
timestamp 1654648307
transform 1 0 101200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_636
timestamp 1654648307
transform 1 0 104200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_637
timestamp 1654648307
transform 1 0 107200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_586
timestamp 1654648307
transform 1 0 104200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_587
timestamp 1654648307
transform 1 0 107200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_638
timestamp 1654648307
transform 1 0 110200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_639
timestamp 1654648307
transform 1 0 113200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_588
timestamp 1654648307
transform 1 0 110200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_589
timestamp 1654648307
transform 1 0 113200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_640
timestamp 1654648307
transform 1 0 116200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_641
timestamp 1654648307
transform 1 0 119200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_590
timestamp 1654648307
transform 1 0 116200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_591
timestamp 1654648307
transform 1 0 119200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_642
timestamp 1654648307
transform 1 0 122200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_643
timestamp 1654648307
transform 1 0 125200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_592
timestamp 1654648307
transform 1 0 122200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_593
timestamp 1654648307
transform 1 0 125200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_644
timestamp 1654648307
transform 1 0 128200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_645
timestamp 1654648307
transform 1 0 131200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_594
timestamp 1654648307
transform 1 0 128200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_595
timestamp 1654648307
transform 1 0 131200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_646
timestamp 1654648307
transform 1 0 134200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_647
timestamp 1654648307
transform 1 0 137200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_596
timestamp 1654648307
transform 1 0 134200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_597
timestamp 1654648307
transform 1 0 137200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_648
timestamp 1654648307
transform 1 0 140200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_649
timestamp 1654648307
transform 1 0 143200 0 1 -33300
box 3640 -2860 6960 460
use pixel  pixel_598
timestamp 1654648307
transform 1 0 140200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_599
timestamp 1654648307
transform 1 0 143200 0 1 -30300
box 3640 -2860 6960 460
use pixel  pixel_500
timestamp 1654648307
transform 1 0 -3800 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_501
timestamp 1654648307
transform 1 0 -800 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_450
timestamp 1654648307
transform 1 0 -3800 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_451
timestamp 1654648307
transform 1 0 -800 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_502
timestamp 1654648307
transform 1 0 2200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_503
timestamp 1654648307
transform 1 0 5200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_452
timestamp 1654648307
transform 1 0 2200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_453
timestamp 1654648307
transform 1 0 5200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_504
timestamp 1654648307
transform 1 0 8200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_505
timestamp 1654648307
transform 1 0 11200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_454
timestamp 1654648307
transform 1 0 8200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_455
timestamp 1654648307
transform 1 0 11200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_506
timestamp 1654648307
transform 1 0 14200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_507
timestamp 1654648307
transform 1 0 17200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_456
timestamp 1654648307
transform 1 0 14200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_457
timestamp 1654648307
transform 1 0 17200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_508
timestamp 1654648307
transform 1 0 20200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_509
timestamp 1654648307
transform 1 0 23200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_458
timestamp 1654648307
transform 1 0 20200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_459
timestamp 1654648307
transform 1 0 23200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_510
timestamp 1654648307
transform 1 0 26200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_511
timestamp 1654648307
transform 1 0 29200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_460
timestamp 1654648307
transform 1 0 26200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_461
timestamp 1654648307
transform 1 0 29200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_512
timestamp 1654648307
transform 1 0 32200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_513
timestamp 1654648307
transform 1 0 35200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_462
timestamp 1654648307
transform 1 0 32200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_463
timestamp 1654648307
transform 1 0 35200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_514
timestamp 1654648307
transform 1 0 38200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_515
timestamp 1654648307
transform 1 0 41200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_464
timestamp 1654648307
transform 1 0 38200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_465
timestamp 1654648307
transform 1 0 41200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_516
timestamp 1654648307
transform 1 0 44200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_517
timestamp 1654648307
transform 1 0 47200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_466
timestamp 1654648307
transform 1 0 44200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_467
timestamp 1654648307
transform 1 0 47200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_518
timestamp 1654648307
transform 1 0 50200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_519
timestamp 1654648307
transform 1 0 53200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_468
timestamp 1654648307
transform 1 0 50200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_469
timestamp 1654648307
transform 1 0 53200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_520
timestamp 1654648307
transform 1 0 56200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_521
timestamp 1654648307
transform 1 0 59200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_470
timestamp 1654648307
transform 1 0 56200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_471
timestamp 1654648307
transform 1 0 59200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_522
timestamp 1654648307
transform 1 0 62200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_523
timestamp 1654648307
transform 1 0 65200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_472
timestamp 1654648307
transform 1 0 62200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_473
timestamp 1654648307
transform 1 0 65200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_524
timestamp 1654648307
transform 1 0 68200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_525
timestamp 1654648307
transform 1 0 71200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_474
timestamp 1654648307
transform 1 0 68200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_475
timestamp 1654648307
transform 1 0 71200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_526
timestamp 1654648307
transform 1 0 74200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_527
timestamp 1654648307
transform 1 0 77200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_476
timestamp 1654648307
transform 1 0 74200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_477
timestamp 1654648307
transform 1 0 77200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_528
timestamp 1654648307
transform 1 0 80200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_529
timestamp 1654648307
transform 1 0 83200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_478
timestamp 1654648307
transform 1 0 80200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_479
timestamp 1654648307
transform 1 0 83200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_530
timestamp 1654648307
transform 1 0 86200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_531
timestamp 1654648307
transform 1 0 89200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_480
timestamp 1654648307
transform 1 0 86200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_481
timestamp 1654648307
transform 1 0 89200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_532
timestamp 1654648307
transform 1 0 92200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_533
timestamp 1654648307
transform 1 0 95200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_482
timestamp 1654648307
transform 1 0 92200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_483
timestamp 1654648307
transform 1 0 95200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_534
timestamp 1654648307
transform 1 0 98200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_535
timestamp 1654648307
transform 1 0 101200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_484
timestamp 1654648307
transform 1 0 98200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_485
timestamp 1654648307
transform 1 0 101200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_536
timestamp 1654648307
transform 1 0 104200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_537
timestamp 1654648307
transform 1 0 107200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_486
timestamp 1654648307
transform 1 0 104200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_487
timestamp 1654648307
transform 1 0 107200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_538
timestamp 1654648307
transform 1 0 110200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_539
timestamp 1654648307
transform 1 0 113200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_488
timestamp 1654648307
transform 1 0 110200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_489
timestamp 1654648307
transform 1 0 113200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_540
timestamp 1654648307
transform 1 0 116200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_541
timestamp 1654648307
transform 1 0 119200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_490
timestamp 1654648307
transform 1 0 116200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_491
timestamp 1654648307
transform 1 0 119200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_542
timestamp 1654648307
transform 1 0 122200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_543
timestamp 1654648307
transform 1 0 125200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_492
timestamp 1654648307
transform 1 0 122200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_493
timestamp 1654648307
transform 1 0 125200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_544
timestamp 1654648307
transform 1 0 128200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_545
timestamp 1654648307
transform 1 0 131200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_494
timestamp 1654648307
transform 1 0 128200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_495
timestamp 1654648307
transform 1 0 131200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_546
timestamp 1654648307
transform 1 0 134200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_547
timestamp 1654648307
transform 1 0 137200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_496
timestamp 1654648307
transform 1 0 134200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_497
timestamp 1654648307
transform 1 0 137200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_548
timestamp 1654648307
transform 1 0 140200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_549
timestamp 1654648307
transform 1 0 143200 0 1 -27300
box 3640 -2860 6960 460
use pixel  pixel_498
timestamp 1654648307
transform 1 0 140200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_499
timestamp 1654648307
transform 1 0 143200 0 1 -24300
box 3640 -2860 6960 460
use pixel  pixel_400
timestamp 1654648307
transform 1 0 -3800 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_401
timestamp 1654648307
transform 1 0 -800 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_350
timestamp 1654648307
transform 1 0 -3800 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_351
timestamp 1654648307
transform 1 0 -800 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_402
timestamp 1654648307
transform 1 0 2200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_403
timestamp 1654648307
transform 1 0 5200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_352
timestamp 1654648307
transform 1 0 2200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_353
timestamp 1654648307
transform 1 0 5200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_404
timestamp 1654648307
transform 1 0 8200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_405
timestamp 1654648307
transform 1 0 11200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_354
timestamp 1654648307
transform 1 0 8200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_355
timestamp 1654648307
transform 1 0 11200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_406
timestamp 1654648307
transform 1 0 14200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_407
timestamp 1654648307
transform 1 0 17200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_356
timestamp 1654648307
transform 1 0 14200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_357
timestamp 1654648307
transform 1 0 17200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_408
timestamp 1654648307
transform 1 0 20200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_409
timestamp 1654648307
transform 1 0 23200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_358
timestamp 1654648307
transform 1 0 20200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_359
timestamp 1654648307
transform 1 0 23200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_410
timestamp 1654648307
transform 1 0 26200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_411
timestamp 1654648307
transform 1 0 29200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_360
timestamp 1654648307
transform 1 0 26200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_361
timestamp 1654648307
transform 1 0 29200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_412
timestamp 1654648307
transform 1 0 32200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_413
timestamp 1654648307
transform 1 0 35200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_362
timestamp 1654648307
transform 1 0 32200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_363
timestamp 1654648307
transform 1 0 35200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_414
timestamp 1654648307
transform 1 0 38200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_415
timestamp 1654648307
transform 1 0 41200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_364
timestamp 1654648307
transform 1 0 38200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_365
timestamp 1654648307
transform 1 0 41200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_416
timestamp 1654648307
transform 1 0 44200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_417
timestamp 1654648307
transform 1 0 47200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_366
timestamp 1654648307
transform 1 0 44200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_367
timestamp 1654648307
transform 1 0 47200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_418
timestamp 1654648307
transform 1 0 50200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_419
timestamp 1654648307
transform 1 0 53200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_368
timestamp 1654648307
transform 1 0 50200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_369
timestamp 1654648307
transform 1 0 53200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_420
timestamp 1654648307
transform 1 0 56200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_421
timestamp 1654648307
transform 1 0 59200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_370
timestamp 1654648307
transform 1 0 56200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_371
timestamp 1654648307
transform 1 0 59200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_422
timestamp 1654648307
transform 1 0 62200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_423
timestamp 1654648307
transform 1 0 65200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_372
timestamp 1654648307
transform 1 0 62200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_373
timestamp 1654648307
transform 1 0 65200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_424
timestamp 1654648307
transform 1 0 68200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_425
timestamp 1654648307
transform 1 0 71200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_374
timestamp 1654648307
transform 1 0 68200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_375
timestamp 1654648307
transform 1 0 71200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_426
timestamp 1654648307
transform 1 0 74200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_427
timestamp 1654648307
transform 1 0 77200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_376
timestamp 1654648307
transform 1 0 74200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_377
timestamp 1654648307
transform 1 0 77200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_428
timestamp 1654648307
transform 1 0 80200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_429
timestamp 1654648307
transform 1 0 83200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_378
timestamp 1654648307
transform 1 0 80200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_379
timestamp 1654648307
transform 1 0 83200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_430
timestamp 1654648307
transform 1 0 86200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_431
timestamp 1654648307
transform 1 0 89200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_380
timestamp 1654648307
transform 1 0 86200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_381
timestamp 1654648307
transform 1 0 89200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_432
timestamp 1654648307
transform 1 0 92200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_433
timestamp 1654648307
transform 1 0 95200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_382
timestamp 1654648307
transform 1 0 92200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_383
timestamp 1654648307
transform 1 0 95200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_434
timestamp 1654648307
transform 1 0 98200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_435
timestamp 1654648307
transform 1 0 101200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_384
timestamp 1654648307
transform 1 0 98200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_385
timestamp 1654648307
transform 1 0 101200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_436
timestamp 1654648307
transform 1 0 104200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_437
timestamp 1654648307
transform 1 0 107200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_386
timestamp 1654648307
transform 1 0 104200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_387
timestamp 1654648307
transform 1 0 107200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_438
timestamp 1654648307
transform 1 0 110200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_439
timestamp 1654648307
transform 1 0 113200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_388
timestamp 1654648307
transform 1 0 110200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_389
timestamp 1654648307
transform 1 0 113200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_440
timestamp 1654648307
transform 1 0 116200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_441
timestamp 1654648307
transform 1 0 119200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_390
timestamp 1654648307
transform 1 0 116200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_391
timestamp 1654648307
transform 1 0 119200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_442
timestamp 1654648307
transform 1 0 122200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_443
timestamp 1654648307
transform 1 0 125200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_392
timestamp 1654648307
transform 1 0 122200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_393
timestamp 1654648307
transform 1 0 125200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_444
timestamp 1654648307
transform 1 0 128200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_445
timestamp 1654648307
transform 1 0 131200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_394
timestamp 1654648307
transform 1 0 128200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_395
timestamp 1654648307
transform 1 0 131200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_446
timestamp 1654648307
transform 1 0 134200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_447
timestamp 1654648307
transform 1 0 137200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_396
timestamp 1654648307
transform 1 0 134200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_397
timestamp 1654648307
transform 1 0 137200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_448
timestamp 1654648307
transform 1 0 140200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_449
timestamp 1654648307
transform 1 0 143200 0 1 -21300
box 3640 -2860 6960 460
use pixel  pixel_398
timestamp 1654648307
transform 1 0 140200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_399
timestamp 1654648307
transform 1 0 143200 0 1 -18300
box 3640 -2860 6960 460
use pixel  pixel_300
timestamp 1654648307
transform 1 0 -3800 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_301
timestamp 1654648307
transform 1 0 -800 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_250
timestamp 1654648307
transform 1 0 -3800 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_251
timestamp 1654648307
transform 1 0 -800 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_302
timestamp 1654648307
transform 1 0 2200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_303
timestamp 1654648307
transform 1 0 5200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_252
timestamp 1654648307
transform 1 0 2200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_253
timestamp 1654648307
transform 1 0 5200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_304
timestamp 1654648307
transform 1 0 8200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_305
timestamp 1654648307
transform 1 0 11200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_254
timestamp 1654648307
transform 1 0 8200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_255
timestamp 1654648307
transform 1 0 11200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_306
timestamp 1654648307
transform 1 0 14200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_307
timestamp 1654648307
transform 1 0 17200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_256
timestamp 1654648307
transform 1 0 14200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_257
timestamp 1654648307
transform 1 0 17200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_308
timestamp 1654648307
transform 1 0 20200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_309
timestamp 1654648307
transform 1 0 23200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_258
timestamp 1654648307
transform 1 0 20200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_259
timestamp 1654648307
transform 1 0 23200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_310
timestamp 1654648307
transform 1 0 26200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_311
timestamp 1654648307
transform 1 0 29200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_260
timestamp 1654648307
transform 1 0 26200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_261
timestamp 1654648307
transform 1 0 29200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_312
timestamp 1654648307
transform 1 0 32200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_313
timestamp 1654648307
transform 1 0 35200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_262
timestamp 1654648307
transform 1 0 32200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_263
timestamp 1654648307
transform 1 0 35200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_314
timestamp 1654648307
transform 1 0 38200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_315
timestamp 1654648307
transform 1 0 41200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_264
timestamp 1654648307
transform 1 0 38200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_265
timestamp 1654648307
transform 1 0 41200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_316
timestamp 1654648307
transform 1 0 44200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_317
timestamp 1654648307
transform 1 0 47200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_266
timestamp 1654648307
transform 1 0 44200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_267
timestamp 1654648307
transform 1 0 47200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_318
timestamp 1654648307
transform 1 0 50200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_319
timestamp 1654648307
transform 1 0 53200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_268
timestamp 1654648307
transform 1 0 50200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_269
timestamp 1654648307
transform 1 0 53200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_320
timestamp 1654648307
transform 1 0 56200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_321
timestamp 1654648307
transform 1 0 59200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_270
timestamp 1654648307
transform 1 0 56200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_271
timestamp 1654648307
transform 1 0 59200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_322
timestamp 1654648307
transform 1 0 62200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_323
timestamp 1654648307
transform 1 0 65200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_272
timestamp 1654648307
transform 1 0 62200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_273
timestamp 1654648307
transform 1 0 65200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_324
timestamp 1654648307
transform 1 0 68200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_325
timestamp 1654648307
transform 1 0 71200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_274
timestamp 1654648307
transform 1 0 68200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_275
timestamp 1654648307
transform 1 0 71200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_326
timestamp 1654648307
transform 1 0 74200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_327
timestamp 1654648307
transform 1 0 77200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_276
timestamp 1654648307
transform 1 0 74200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_277
timestamp 1654648307
transform 1 0 77200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_328
timestamp 1654648307
transform 1 0 80200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_329
timestamp 1654648307
transform 1 0 83200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_278
timestamp 1654648307
transform 1 0 80200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_279
timestamp 1654648307
transform 1 0 83200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_330
timestamp 1654648307
transform 1 0 86200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_331
timestamp 1654648307
transform 1 0 89200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_280
timestamp 1654648307
transform 1 0 86200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_281
timestamp 1654648307
transform 1 0 89200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_332
timestamp 1654648307
transform 1 0 92200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_333
timestamp 1654648307
transform 1 0 95200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_282
timestamp 1654648307
transform 1 0 92200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_283
timestamp 1654648307
transform 1 0 95200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_334
timestamp 1654648307
transform 1 0 98200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_335
timestamp 1654648307
transform 1 0 101200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_284
timestamp 1654648307
transform 1 0 98200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_285
timestamp 1654648307
transform 1 0 101200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_336
timestamp 1654648307
transform 1 0 104200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_337
timestamp 1654648307
transform 1 0 107200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_286
timestamp 1654648307
transform 1 0 104200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_287
timestamp 1654648307
transform 1 0 107200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_338
timestamp 1654648307
transform 1 0 110200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_339
timestamp 1654648307
transform 1 0 113200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_288
timestamp 1654648307
transform 1 0 110200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_289
timestamp 1654648307
transform 1 0 113200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_340
timestamp 1654648307
transform 1 0 116200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_341
timestamp 1654648307
transform 1 0 119200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_290
timestamp 1654648307
transform 1 0 116200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_291
timestamp 1654648307
transform 1 0 119200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_342
timestamp 1654648307
transform 1 0 122200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_343
timestamp 1654648307
transform 1 0 125200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_292
timestamp 1654648307
transform 1 0 122200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_293
timestamp 1654648307
transform 1 0 125200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_344
timestamp 1654648307
transform 1 0 128200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_345
timestamp 1654648307
transform 1 0 131200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_294
timestamp 1654648307
transform 1 0 128200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_295
timestamp 1654648307
transform 1 0 131200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_346
timestamp 1654648307
transform 1 0 134200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_347
timestamp 1654648307
transform 1 0 137200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_296
timestamp 1654648307
transform 1 0 134200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_297
timestamp 1654648307
transform 1 0 137200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_348
timestamp 1654648307
transform 1 0 140200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_349
timestamp 1654648307
transform 1 0 143200 0 1 -15300
box 3640 -2860 6960 460
use pixel  pixel_298
timestamp 1654648307
transform 1 0 140200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_299
timestamp 1654648307
transform 1 0 143200 0 1 -12300
box 3640 -2860 6960 460
use pixel  pixel_200
timestamp 1654648307
transform 1 0 -3800 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_201
timestamp 1654648307
transform 1 0 -800 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_150
timestamp 1654648307
transform 1 0 -3800 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_151
timestamp 1654648307
transform 1 0 -800 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_202
timestamp 1654648307
transform 1 0 2200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_203
timestamp 1654648307
transform 1 0 5200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_152
timestamp 1654648307
transform 1 0 2200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_153
timestamp 1654648307
transform 1 0 5200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_204
timestamp 1654648307
transform 1 0 8200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_205
timestamp 1654648307
transform 1 0 11200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_154
timestamp 1654648307
transform 1 0 8200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_155
timestamp 1654648307
transform 1 0 11200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_206
timestamp 1654648307
transform 1 0 14200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_207
timestamp 1654648307
transform 1 0 17200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_156
timestamp 1654648307
transform 1 0 14200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_157
timestamp 1654648307
transform 1 0 17200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_208
timestamp 1654648307
transform 1 0 20200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_209
timestamp 1654648307
transform 1 0 23200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_158
timestamp 1654648307
transform 1 0 20200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_159
timestamp 1654648307
transform 1 0 23200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_210
timestamp 1654648307
transform 1 0 26200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_211
timestamp 1654648307
transform 1 0 29200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_160
timestamp 1654648307
transform 1 0 26200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_161
timestamp 1654648307
transform 1 0 29200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_212
timestamp 1654648307
transform 1 0 32200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_213
timestamp 1654648307
transform 1 0 35200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_162
timestamp 1654648307
transform 1 0 32200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_163
timestamp 1654648307
transform 1 0 35200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_214
timestamp 1654648307
transform 1 0 38200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_215
timestamp 1654648307
transform 1 0 41200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_164
timestamp 1654648307
transform 1 0 38200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_165
timestamp 1654648307
transform 1 0 41200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_216
timestamp 1654648307
transform 1 0 44200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_217
timestamp 1654648307
transform 1 0 47200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_166
timestamp 1654648307
transform 1 0 44200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_167
timestamp 1654648307
transform 1 0 47200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_218
timestamp 1654648307
transform 1 0 50200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_219
timestamp 1654648307
transform 1 0 53200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_168
timestamp 1654648307
transform 1 0 50200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_169
timestamp 1654648307
transform 1 0 53200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_220
timestamp 1654648307
transform 1 0 56200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_221
timestamp 1654648307
transform 1 0 59200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_170
timestamp 1654648307
transform 1 0 56200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_171
timestamp 1654648307
transform 1 0 59200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_222
timestamp 1654648307
transform 1 0 62200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_223
timestamp 1654648307
transform 1 0 65200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_172
timestamp 1654648307
transform 1 0 62200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_173
timestamp 1654648307
transform 1 0 65200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_224
timestamp 1654648307
transform 1 0 68200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_225
timestamp 1654648307
transform 1 0 71200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_174
timestamp 1654648307
transform 1 0 68200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_175
timestamp 1654648307
transform 1 0 71200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_226
timestamp 1654648307
transform 1 0 74200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_227
timestamp 1654648307
transform 1 0 77200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_176
timestamp 1654648307
transform 1 0 74200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_177
timestamp 1654648307
transform 1 0 77200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_228
timestamp 1654648307
transform 1 0 80200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_229
timestamp 1654648307
transform 1 0 83200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_178
timestamp 1654648307
transform 1 0 80200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_179
timestamp 1654648307
transform 1 0 83200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_230
timestamp 1654648307
transform 1 0 86200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_231
timestamp 1654648307
transform 1 0 89200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_180
timestamp 1654648307
transform 1 0 86200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_181
timestamp 1654648307
transform 1 0 89200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_232
timestamp 1654648307
transform 1 0 92200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_233
timestamp 1654648307
transform 1 0 95200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_182
timestamp 1654648307
transform 1 0 92200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_183
timestamp 1654648307
transform 1 0 95200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_234
timestamp 1654648307
transform 1 0 98200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_235
timestamp 1654648307
transform 1 0 101200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_184
timestamp 1654648307
transform 1 0 98200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_185
timestamp 1654648307
transform 1 0 101200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_236
timestamp 1654648307
transform 1 0 104200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_237
timestamp 1654648307
transform 1 0 107200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_186
timestamp 1654648307
transform 1 0 104200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_187
timestamp 1654648307
transform 1 0 107200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_238
timestamp 1654648307
transform 1 0 110200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_239
timestamp 1654648307
transform 1 0 113200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_188
timestamp 1654648307
transform 1 0 110200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_189
timestamp 1654648307
transform 1 0 113200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_240
timestamp 1654648307
transform 1 0 116200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_241
timestamp 1654648307
transform 1 0 119200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_190
timestamp 1654648307
transform 1 0 116200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_191
timestamp 1654648307
transform 1 0 119200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_242
timestamp 1654648307
transform 1 0 122200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_243
timestamp 1654648307
transform 1 0 125200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_192
timestamp 1654648307
transform 1 0 122200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_193
timestamp 1654648307
transform 1 0 125200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_244
timestamp 1654648307
transform 1 0 128200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_245
timestamp 1654648307
transform 1 0 131200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_194
timestamp 1654648307
transform 1 0 128200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_195
timestamp 1654648307
transform 1 0 131200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_246
timestamp 1654648307
transform 1 0 134200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_247
timestamp 1654648307
transform 1 0 137200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_196
timestamp 1654648307
transform 1 0 134200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_197
timestamp 1654648307
transform 1 0 137200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_248
timestamp 1654648307
transform 1 0 140200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_249
timestamp 1654648307
transform 1 0 143200 0 1 -9300
box 3640 -2860 6960 460
use pixel  pixel_198
timestamp 1654648307
transform 1 0 140200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_199
timestamp 1654648307
transform 1 0 143200 0 1 -6300
box 3640 -2860 6960 460
use pixel  pixel_100
timestamp 1654648307
transform 1 0 -3800 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_101
timestamp 1654648307
transform 1 0 -800 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_50
timestamp 1654648307
transform 1 0 -3800 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_51
timestamp 1654648307
transform 1 0 -800 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_102
timestamp 1654648307
transform 1 0 2200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_103
timestamp 1654648307
transform 1 0 5200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_52
timestamp 1654648307
transform 1 0 2200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_53
timestamp 1654648307
transform 1 0 5200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_104
timestamp 1654648307
transform 1 0 8200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_105
timestamp 1654648307
transform 1 0 11200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_54
timestamp 1654648307
transform 1 0 8200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_55
timestamp 1654648307
transform 1 0 11200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_106
timestamp 1654648307
transform 1 0 14200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_107
timestamp 1654648307
transform 1 0 17200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_56
timestamp 1654648307
transform 1 0 14200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_57
timestamp 1654648307
transform 1 0 17200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_108
timestamp 1654648307
transform 1 0 20200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_109
timestamp 1654648307
transform 1 0 23200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_58
timestamp 1654648307
transform 1 0 20200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_59
timestamp 1654648307
transform 1 0 23200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_110
timestamp 1654648307
transform 1 0 26200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_111
timestamp 1654648307
transform 1 0 29200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_60
timestamp 1654648307
transform 1 0 26200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_61
timestamp 1654648307
transform 1 0 29200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_112
timestamp 1654648307
transform 1 0 32200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_113
timestamp 1654648307
transform 1 0 35200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_62
timestamp 1654648307
transform 1 0 32200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_63
timestamp 1654648307
transform 1 0 35200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_114
timestamp 1654648307
transform 1 0 38200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_115
timestamp 1654648307
transform 1 0 41200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_64
timestamp 1654648307
transform 1 0 38200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_65
timestamp 1654648307
transform 1 0 41200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_116
timestamp 1654648307
transform 1 0 44200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_117
timestamp 1654648307
transform 1 0 47200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_66
timestamp 1654648307
transform 1 0 44200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_67
timestamp 1654648307
transform 1 0 47200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_118
timestamp 1654648307
transform 1 0 50200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_119
timestamp 1654648307
transform 1 0 53200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_68
timestamp 1654648307
transform 1 0 50200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_69
timestamp 1654648307
transform 1 0 53200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_120
timestamp 1654648307
transform 1 0 56200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_121
timestamp 1654648307
transform 1 0 59200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_70
timestamp 1654648307
transform 1 0 56200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_71
timestamp 1654648307
transform 1 0 59200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_122
timestamp 1654648307
transform 1 0 62200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_123
timestamp 1654648307
transform 1 0 65200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_72
timestamp 1654648307
transform 1 0 62200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_73
timestamp 1654648307
transform 1 0 65200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_124
timestamp 1654648307
transform 1 0 68200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_125
timestamp 1654648307
transform 1 0 71200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_74
timestamp 1654648307
transform 1 0 68200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_75
timestamp 1654648307
transform 1 0 71200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_126
timestamp 1654648307
transform 1 0 74200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_127
timestamp 1654648307
transform 1 0 77200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_76
timestamp 1654648307
transform 1 0 74200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_77
timestamp 1654648307
transform 1 0 77200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_128
timestamp 1654648307
transform 1 0 80200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_129
timestamp 1654648307
transform 1 0 83200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_78
timestamp 1654648307
transform 1 0 80200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_79
timestamp 1654648307
transform 1 0 83200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_130
timestamp 1654648307
transform 1 0 86200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_131
timestamp 1654648307
transform 1 0 89200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_80
timestamp 1654648307
transform 1 0 86200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_81
timestamp 1654648307
transform 1 0 89200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_132
timestamp 1654648307
transform 1 0 92200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_133
timestamp 1654648307
transform 1 0 95200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_82
timestamp 1654648307
transform 1 0 92200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_83
timestamp 1654648307
transform 1 0 95200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_134
timestamp 1654648307
transform 1 0 98200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_135
timestamp 1654648307
transform 1 0 101200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_84
timestamp 1654648307
transform 1 0 98200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_85
timestamp 1654648307
transform 1 0 101200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_136
timestamp 1654648307
transform 1 0 104200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_137
timestamp 1654648307
transform 1 0 107200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_86
timestamp 1654648307
transform 1 0 104200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_87
timestamp 1654648307
transform 1 0 107200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_138
timestamp 1654648307
transform 1 0 110200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_139
timestamp 1654648307
transform 1 0 113200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_88
timestamp 1654648307
transform 1 0 110200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_89
timestamp 1654648307
transform 1 0 113200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_140
timestamp 1654648307
transform 1 0 116200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_141
timestamp 1654648307
transform 1 0 119200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_90
timestamp 1654648307
transform 1 0 116200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_91
timestamp 1654648307
transform 1 0 119200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_142
timestamp 1654648307
transform 1 0 122200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_143
timestamp 1654648307
transform 1 0 125200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_92
timestamp 1654648307
transform 1 0 122200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_93
timestamp 1654648307
transform 1 0 125200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_144
timestamp 1654648307
transform 1 0 128200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_145
timestamp 1654648307
transform 1 0 131200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_94
timestamp 1654648307
transform 1 0 128200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_95
timestamp 1654648307
transform 1 0 131200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_146
timestamp 1654648307
transform 1 0 134200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_147
timestamp 1654648307
transform 1 0 137200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_96
timestamp 1654648307
transform 1 0 134200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_97
timestamp 1654648307
transform 1 0 137200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_148
timestamp 1654648307
transform 1 0 140200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_149
timestamp 1654648307
transform 1 0 143200 0 1 -3300
box 3640 -2860 6960 460
use pixel  pixel_98
timestamp 1654648307
transform 1 0 140200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_99
timestamp 1654648307
transform 1 0 143200 0 1 -300
box 3640 -2860 6960 460
use pixel  pixel_0
timestamp 1654648307
transform 1 0 -3800 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_1
timestamp 1654648307
transform 1 0 -800 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_2
timestamp 1654648307
transform 1 0 2200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_3
timestamp 1654648307
transform 1 0 5200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_4
timestamp 1654648307
transform 1 0 8200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_5
timestamp 1654648307
transform 1 0 11200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_6
timestamp 1654648307
transform 1 0 14200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_7
timestamp 1654648307
transform 1 0 17200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_8
timestamp 1654648307
transform 1 0 20200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_9
timestamp 1654648307
transform 1 0 23200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_10
timestamp 1654648307
transform 1 0 26200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_11
timestamp 1654648307
transform 1 0 29200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_12
timestamp 1654648307
transform 1 0 32200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_13
timestamp 1654648307
transform 1 0 35200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_14
timestamp 1654648307
transform 1 0 38200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_15
timestamp 1654648307
transform 1 0 41200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_16
timestamp 1654648307
transform 1 0 44200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_17
timestamp 1654648307
transform 1 0 47200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_18
timestamp 1654648307
transform 1 0 50200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_19
timestamp 1654648307
transform 1 0 53200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_20
timestamp 1654648307
transform 1 0 56200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_21
timestamp 1654648307
transform 1 0 59200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_22
timestamp 1654648307
transform 1 0 62200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_23
timestamp 1654648307
transform 1 0 65200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_24
timestamp 1654648307
transform 1 0 68200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_25
timestamp 1654648307
transform 1 0 71200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_26
timestamp 1654648307
transform 1 0 74200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_27
timestamp 1654648307
transform 1 0 77200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_28
timestamp 1654648307
transform 1 0 80200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_29
timestamp 1654648307
transform 1 0 83200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_30
timestamp 1654648307
transform 1 0 86200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_31
timestamp 1654648307
transform 1 0 89200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_32
timestamp 1654648307
transform 1 0 92200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_33
timestamp 1654648307
transform 1 0 95200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_34
timestamp 1654648307
transform 1 0 98200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_35
timestamp 1654648307
transform 1 0 101200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_36
timestamp 1654648307
transform 1 0 104200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_37
timestamp 1654648307
transform 1 0 107200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_38
timestamp 1654648307
transform 1 0 110200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_39
timestamp 1654648307
transform 1 0 113200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_40
timestamp 1654648307
transform 1 0 116200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_41
timestamp 1654648307
transform 1 0 119200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_42
timestamp 1654648307
transform 1 0 122200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_43
timestamp 1654648307
transform 1 0 125200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_44
timestamp 1654648307
transform 1 0 128200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_45
timestamp 1654648307
transform 1 0 131200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_46
timestamp 1654648307
transform 1 0 134200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_47
timestamp 1654648307
transform 1 0 137200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_48
timestamp 1654648307
transform 1 0 140200 0 1 2700
box 3640 -2860 6960 460
use pixel  pixel_49
timestamp 1654648307
transform 1 0 143200 0 1 2700
box 3640 -2860 6960 460
use opamp_wrapper  opamp_wrapper_0
timestamp 1654646295
transform 1 0 154280 0 1 -146491
box -2280 -1609 26995 13665
use bias  bias_0
timestamp 1654639008
transform 1 0 72210 0 1 7236
box 790 -2236 7180 -220
<< labels >>
rlabel metal5 1040 1040 1240 1240 1 PIX0_IN
port 1 n
rlabel metal4 -3000 3550 -3000 3660 1 VBIAS
port 2 n
rlabel metal2 -3000 3350 -3000 3450 3 VREF
port 3 e
rlabel metal2 0 4040 0 4040 1 NB2
port 4 n
rlabel metal1 -2000 0 -2000 0 1 VDD
port 5 n
rlabel space -1160 5750 -1160 5750 5 SF_IB
port 6 s
rlabel metal2 -740 3560 -740 3560 1 NB1
port 7 n
rlabel metal2 -3000 1480 -3000 1570 3 ROW_SEL0
port 8 e
rlabel metal5 -2000 2840 -2000 2840 1 GRING
port 9 n
rlabel metal5 4040 1040 4240 1240 1 PIX1_IN
port 10 n
rlabel metal5 7040 1040 7240 1240 1 PIX2_IN
port 11 n
rlabel metal5 10040 1040 10240 1240 1 PIX3_IN
port 12 n
rlabel metal5 13040 1040 13240 1240 1 PIX4_IN
port 13 n
rlabel metal5 16040 1040 16240 1240 1 PIX5_IN
port 14 n
rlabel metal5 19040 1040 19240 1240 1 PIX6_IN
port 15 n
rlabel metal5 22040 1040 22240 1240 1 PIX7_IN
port 16 n
rlabel metal5 25040 1040 25240 1240 1 PIX8_IN
port 17 n
rlabel metal5 28040 1040 28240 1240 1 PIX9_IN
port 18 n
rlabel metal5 31040 1040 31240 1240 1 PIX10_IN
port 19 n
rlabel metal5 34040 1040 34240 1240 1 PIX11_IN
port 20 n
rlabel metal5 37040 1040 37240 1240 1 PIX12_IN
port 21 n
rlabel metal5 40040 1040 40240 1240 1 PIX13_IN
port 22 n
rlabel metal5 43040 1040 43240 1240 1 PIX14_IN
port 23 n
rlabel metal5 46040 1040 46240 1240 1 PIX15_IN
port 24 n
rlabel metal5 49040 1040 49240 1240 1 PIX16_IN
port 25 n
rlabel metal5 52040 1040 52240 1240 1 PIX17_IN
port 26 n
rlabel metal5 55040 1040 55240 1240 1 PIX18_IN
port 27 n
rlabel metal5 58040 1040 58240 1240 1 PIX19_IN
port 28 n
rlabel metal5 61040 1040 61240 1240 1 PIX20_IN
port 29 n
rlabel metal5 64040 1040 64240 1240 1 PIX21_IN
port 30 n
rlabel metal5 67040 1040 67240 1240 1 PIX22_IN
port 31 n
rlabel metal5 70040 1040 70240 1240 1 PIX23_IN
port 32 n
rlabel metal5 73040 1040 73240 1240 1 PIX24_IN
port 33 n
rlabel metal5 76040 1040 76240 1240 1 PIX25_IN
port 34 n
rlabel metal5 79040 1040 79240 1240 1 PIX26_IN
port 35 n
rlabel metal5 82040 1040 82240 1240 1 PIX27_IN
port 36 n
rlabel metal5 85040 1040 85240 1240 1 PIX28_IN
port 37 n
rlabel metal5 88040 1040 88240 1240 1 PIX29_IN
port 38 n
rlabel metal5 91040 1040 91240 1240 1 PIX30_IN
port 39 n
rlabel metal5 94040 1040 94240 1240 1 PIX31_IN
port 40 n
rlabel metal5 97040 1040 97240 1240 1 PIX32_IN
port 41 n
rlabel metal5 100040 1040 100240 1240 1 PIX33_IN
port 42 n
rlabel metal5 103040 1040 103240 1240 1 PIX34_IN
port 43 n
rlabel metal5 106040 1040 106240 1240 1 PIX35_IN
port 44 n
rlabel metal5 109040 1040 109240 1240 1 PIX36_IN
port 45 n
rlabel metal5 112040 1040 112240 1240 1 PIX37_IN
port 46 n
rlabel metal5 115040 1040 115240 1240 1 PIX38_IN
port 47 n
rlabel metal5 118040 1040 118240 1240 1 PIX39_IN
port 48 n
rlabel metal5 121040 1040 121240 1240 1 PIX40_IN
port 49 n
rlabel metal5 124040 1040 124240 1240 1 PIX41_IN
port 50 n
rlabel metal5 127040 1040 127240 1240 1 PIX42_IN
port 51 n
rlabel metal5 130040 1040 130240 1240 1 PIX43_IN
port 52 n
rlabel metal5 133040 1040 133240 1240 1 PIX44_IN
port 53 n
rlabel metal5 136040 1040 136240 1240 1 PIX45_IN
port 54 n
rlabel metal5 139040 1040 139240 1240 1 PIX46_IN
port 55 n
rlabel metal5 142040 1040 142240 1240 1 PIX47_IN
port 56 n
rlabel metal5 145040 1040 145240 1240 1 PIX48_IN
port 57 n
rlabel metal5 148040 1040 148240 1240 1 PIX49_IN
port 58 n
rlabel metal1 150400 30 150400 30 1 GND
port 59 n
rlabel metal5 1040 -1960 1240 -1760 1 PIX50_IN
port 60 n
rlabel metal2 -3000 -1520 -3000 -1430 3 ROW_SEL1
port 61 e
rlabel metal5 4040 -1960 4240 -1760 1 PIX51_IN
port 62 n
rlabel metal5 7040 -1960 7240 -1760 1 PIX52_IN
port 63 n
rlabel metal5 10040 -1960 10240 -1760 1 PIX53_IN
port 64 n
rlabel metal5 13040 -1960 13240 -1760 1 PIX54_IN
port 65 n
rlabel metal5 16040 -1960 16240 -1760 1 PIX55_IN
port 66 n
rlabel metal5 19040 -1960 19240 -1760 1 PIX56_IN
port 67 n
rlabel metal5 22040 -1960 22240 -1760 1 PIX57_IN
port 68 n
rlabel metal5 25040 -1960 25240 -1760 1 PIX58_IN
port 69 n
rlabel metal5 28040 -1960 28240 -1760 1 PIX59_IN
port 70 n
rlabel metal5 31040 -1960 31240 -1760 1 PIX60_IN
port 71 n
rlabel metal5 34040 -1960 34240 -1760 1 PIX61_IN
port 72 n
rlabel metal5 37040 -1960 37240 -1760 1 PIX62_IN
port 73 n
rlabel metal5 40040 -1960 40240 -1760 1 PIX63_IN
port 74 n
rlabel metal5 43040 -1960 43240 -1760 1 PIX64_IN
port 75 n
rlabel metal5 46040 -1960 46240 -1760 1 PIX65_IN
port 76 n
rlabel metal5 49040 -1960 49240 -1760 1 PIX66_IN
port 77 n
rlabel metal5 52040 -1960 52240 -1760 1 PIX67_IN
port 78 n
rlabel metal5 55040 -1960 55240 -1760 1 PIX68_IN
port 79 n
rlabel metal5 58040 -1960 58240 -1760 1 PIX69_IN
port 80 n
rlabel metal5 61040 -1960 61240 -1760 1 PIX70_IN
port 81 n
rlabel metal5 64040 -1960 64240 -1760 1 PIX71_IN
port 82 n
rlabel metal5 67040 -1960 67240 -1760 1 PIX72_IN
port 83 n
rlabel metal5 70040 -1960 70240 -1760 1 PIX73_IN
port 84 n
rlabel metal5 73040 -1960 73240 -1760 1 PIX74_IN
port 85 n
rlabel metal5 76040 -1960 76240 -1760 1 PIX75_IN
port 86 n
rlabel metal5 79040 -1960 79240 -1760 1 PIX76_IN
port 87 n
rlabel metal5 82040 -1960 82240 -1760 1 PIX77_IN
port 88 n
rlabel metal5 85040 -1960 85240 -1760 1 PIX78_IN
port 89 n
rlabel metal5 88040 -1960 88240 -1760 1 PIX79_IN
port 90 n
rlabel metal5 91040 -1960 91240 -1760 1 PIX80_IN
port 91 n
rlabel metal5 94040 -1960 94240 -1760 1 PIX81_IN
port 92 n
rlabel metal5 97040 -1960 97240 -1760 1 PIX82_IN
port 93 n
rlabel metal5 100040 -1960 100240 -1760 1 PIX83_IN
port 94 n
rlabel metal5 103040 -1960 103240 -1760 1 PIX84_IN
port 95 n
rlabel metal5 106040 -1960 106240 -1760 1 PIX85_IN
port 96 n
rlabel metal5 109040 -1960 109240 -1760 1 PIX86_IN
port 97 n
rlabel metal5 112040 -1960 112240 -1760 1 PIX87_IN
port 98 n
rlabel metal5 115040 -1960 115240 -1760 1 PIX88_IN
port 99 n
rlabel metal5 118040 -1960 118240 -1760 1 PIX89_IN
port 100 n
rlabel metal5 121040 -1960 121240 -1760 1 PIX90_IN
port 101 n
rlabel metal5 124040 -1960 124240 -1760 1 PIX91_IN
port 102 n
rlabel metal5 127040 -1960 127240 -1760 1 PIX92_IN
port 103 n
rlabel metal5 130040 -1960 130240 -1760 1 PIX93_IN
port 104 n
rlabel metal5 133040 -1960 133240 -1760 1 PIX94_IN
port 105 n
rlabel metal5 136040 -1960 136240 -1760 1 PIX95_IN
port 106 n
rlabel metal5 139040 -1960 139240 -1760 1 PIX96_IN
port 107 n
rlabel metal5 142040 -1960 142240 -1760 1 PIX97_IN
port 108 n
rlabel metal5 145040 -1960 145240 -1760 1 PIX98_IN
port 109 n
rlabel metal5 148040 -1960 148240 -1760 1 PIX99_IN
port 110 n
rlabel metal5 1040 -4960 1240 -4760 1 PIX100_IN
port 111 n
rlabel metal2 -3000 -4520 -3000 -4430 3 ROW_SEL2
port 112 e
rlabel metal5 4040 -4960 4240 -4760 1 PIX101_IN
port 113 n
rlabel metal5 7040 -4960 7240 -4760 1 PIX102_IN
port 114 n
rlabel metal5 10040 -4960 10240 -4760 1 PIX103_IN
port 115 n
rlabel metal5 13040 -4960 13240 -4760 1 PIX104_IN
port 116 n
rlabel metal5 16040 -4960 16240 -4760 1 PIX105_IN
port 117 n
rlabel metal5 19040 -4960 19240 -4760 1 PIX106_IN
port 118 n
rlabel metal5 22040 -4960 22240 -4760 1 PIX107_IN
port 119 n
rlabel metal5 25040 -4960 25240 -4760 1 PIX108_IN
port 120 n
rlabel metal5 28040 -4960 28240 -4760 1 PIX109_IN
port 121 n
rlabel metal5 31040 -4960 31240 -4760 1 PIX110_IN
port 122 n
rlabel metal5 34040 -4960 34240 -4760 1 PIX111_IN
port 123 n
rlabel metal5 37040 -4960 37240 -4760 1 PIX112_IN
port 124 n
rlabel metal5 40040 -4960 40240 -4760 1 PIX113_IN
port 125 n
rlabel metal5 43040 -4960 43240 -4760 1 PIX114_IN
port 126 n
rlabel metal5 46040 -4960 46240 -4760 1 PIX115_IN
port 127 n
rlabel metal5 49040 -4960 49240 -4760 1 PIX116_IN
port 128 n
rlabel metal5 52040 -4960 52240 -4760 1 PIX117_IN
port 129 n
rlabel metal5 55040 -4960 55240 -4760 1 PIX118_IN
port 130 n
rlabel metal5 58040 -4960 58240 -4760 1 PIX119_IN
port 131 n
rlabel metal5 61040 -4960 61240 -4760 1 PIX120_IN
port 132 n
rlabel metal5 64040 -4960 64240 -4760 1 PIX121_IN
port 133 n
rlabel metal5 67040 -4960 67240 -4760 1 PIX122_IN
port 134 n
rlabel metal5 70040 -4960 70240 -4760 1 PIX123_IN
port 135 n
rlabel metal5 73040 -4960 73240 -4760 1 PIX124_IN
port 136 n
rlabel metal5 76040 -4960 76240 -4760 1 PIX125_IN
port 137 n
rlabel metal5 79040 -4960 79240 -4760 1 PIX126_IN
port 138 n
rlabel metal5 82040 -4960 82240 -4760 1 PIX127_IN
port 139 n
rlabel metal5 85040 -4960 85240 -4760 1 PIX128_IN
port 140 n
rlabel metal5 88040 -4960 88240 -4760 1 PIX129_IN
port 141 n
rlabel metal5 91040 -4960 91240 -4760 1 PIX130_IN
port 142 n
rlabel metal5 94040 -4960 94240 -4760 1 PIX131_IN
port 143 n
rlabel metal5 97040 -4960 97240 -4760 1 PIX132_IN
port 144 n
rlabel metal5 100040 -4960 100240 -4760 1 PIX133_IN
port 145 n
rlabel metal5 103040 -4960 103240 -4760 1 PIX134_IN
port 146 n
rlabel metal5 106040 -4960 106240 -4760 1 PIX135_IN
port 147 n
rlabel metal5 109040 -4960 109240 -4760 1 PIX136_IN
port 148 n
rlabel metal5 112040 -4960 112240 -4760 1 PIX137_IN
port 149 n
rlabel metal5 115040 -4960 115240 -4760 1 PIX138_IN
port 150 n
rlabel metal5 118040 -4960 118240 -4760 1 PIX139_IN
port 151 n
rlabel metal5 121040 -4960 121240 -4760 1 PIX140_IN
port 152 n
rlabel metal5 124040 -4960 124240 -4760 1 PIX141_IN
port 153 n
rlabel metal5 127040 -4960 127240 -4760 1 PIX142_IN
port 154 n
rlabel metal5 130040 -4960 130240 -4760 1 PIX143_IN
port 155 n
rlabel metal5 133040 -4960 133240 -4760 1 PIX144_IN
port 156 n
rlabel metal5 136040 -4960 136240 -4760 1 PIX145_IN
port 157 n
rlabel metal5 139040 -4960 139240 -4760 1 PIX146_IN
port 158 n
rlabel metal5 142040 -4960 142240 -4760 1 PIX147_IN
port 159 n
rlabel metal5 145040 -4960 145240 -4760 1 PIX148_IN
port 160 n
rlabel metal5 148040 -4960 148240 -4760 1 PIX149_IN
port 161 n
rlabel metal5 1040 -7960 1240 -7760 1 PIX150_IN
port 162 n
rlabel metal2 -3000 -7520 -3000 -7430 3 ROW_SEL3
port 163 e
rlabel metal5 4040 -7960 4240 -7760 1 PIX151_IN
port 164 n
rlabel metal5 7040 -7960 7240 -7760 1 PIX152_IN
port 165 n
rlabel metal5 10040 -7960 10240 -7760 1 PIX153_IN
port 166 n
rlabel metal5 13040 -7960 13240 -7760 1 PIX154_IN
port 167 n
rlabel metal5 16040 -7960 16240 -7760 1 PIX155_IN
port 168 n
rlabel metal5 19040 -7960 19240 -7760 1 PIX156_IN
port 169 n
rlabel metal5 22040 -7960 22240 -7760 1 PIX157_IN
port 170 n
rlabel metal5 25040 -7960 25240 -7760 1 PIX158_IN
port 171 n
rlabel metal5 28040 -7960 28240 -7760 1 PIX159_IN
port 172 n
rlabel metal5 31040 -7960 31240 -7760 1 PIX160_IN
port 173 n
rlabel metal5 34040 -7960 34240 -7760 1 PIX161_IN
port 174 n
rlabel metal5 37040 -7960 37240 -7760 1 PIX162_IN
port 175 n
rlabel metal5 40040 -7960 40240 -7760 1 PIX163_IN
port 176 n
rlabel metal5 43040 -7960 43240 -7760 1 PIX164_IN
port 177 n
rlabel metal5 46040 -7960 46240 -7760 1 PIX165_IN
port 178 n
rlabel metal5 49040 -7960 49240 -7760 1 PIX166_IN
port 179 n
rlabel metal5 52040 -7960 52240 -7760 1 PIX167_IN
port 180 n
rlabel metal5 55040 -7960 55240 -7760 1 PIX168_IN
port 181 n
rlabel metal5 58040 -7960 58240 -7760 1 PIX169_IN
port 182 n
rlabel metal5 61040 -7960 61240 -7760 1 PIX170_IN
port 183 n
rlabel metal5 64040 -7960 64240 -7760 1 PIX171_IN
port 184 n
rlabel metal5 67040 -7960 67240 -7760 1 PIX172_IN
port 185 n
rlabel metal5 70040 -7960 70240 -7760 1 PIX173_IN
port 186 n
rlabel metal5 73040 -7960 73240 -7760 1 PIX174_IN
port 187 n
rlabel metal5 76040 -7960 76240 -7760 1 PIX175_IN
port 188 n
rlabel metal5 79040 -7960 79240 -7760 1 PIX176_IN
port 189 n
rlabel metal5 82040 -7960 82240 -7760 1 PIX177_IN
port 190 n
rlabel metal5 85040 -7960 85240 -7760 1 PIX178_IN
port 191 n
rlabel metal5 88040 -7960 88240 -7760 1 PIX179_IN
port 192 n
rlabel metal5 91040 -7960 91240 -7760 1 PIX180_IN
port 193 n
rlabel metal5 94040 -7960 94240 -7760 1 PIX181_IN
port 194 n
rlabel metal5 97040 -7960 97240 -7760 1 PIX182_IN
port 195 n
rlabel metal5 100040 -7960 100240 -7760 1 PIX183_IN
port 196 n
rlabel metal5 103040 -7960 103240 -7760 1 PIX184_IN
port 197 n
rlabel metal5 106040 -7960 106240 -7760 1 PIX185_IN
port 198 n
rlabel metal5 109040 -7960 109240 -7760 1 PIX186_IN
port 199 n
rlabel metal5 112040 -7960 112240 -7760 1 PIX187_IN
port 200 n
rlabel metal5 115040 -7960 115240 -7760 1 PIX188_IN
port 201 n
rlabel metal5 118040 -7960 118240 -7760 1 PIX189_IN
port 202 n
rlabel metal5 121040 -7960 121240 -7760 1 PIX190_IN
port 203 n
rlabel metal5 124040 -7960 124240 -7760 1 PIX191_IN
port 204 n
rlabel metal5 127040 -7960 127240 -7760 1 PIX192_IN
port 205 n
rlabel metal5 130040 -7960 130240 -7760 1 PIX193_IN
port 206 n
rlabel metal5 133040 -7960 133240 -7760 1 PIX194_IN
port 207 n
rlabel metal5 136040 -7960 136240 -7760 1 PIX195_IN
port 208 n
rlabel metal5 139040 -7960 139240 -7760 1 PIX196_IN
port 209 n
rlabel metal5 142040 -7960 142240 -7760 1 PIX197_IN
port 210 n
rlabel metal5 145040 -7960 145240 -7760 1 PIX198_IN
port 211 n
rlabel metal5 148040 -7960 148240 -7760 1 PIX199_IN
port 212 n
rlabel metal5 1040 -10960 1240 -10760 1 PIX200_IN
port 213 n
rlabel metal2 -3000 -10520 -3000 -10430 3 ROW_SEL4
port 214 e
rlabel metal5 4040 -10960 4240 -10760 1 PIX201_IN
port 215 n
rlabel metal5 7040 -10960 7240 -10760 1 PIX202_IN
port 216 n
rlabel metal5 10040 -10960 10240 -10760 1 PIX203_IN
port 217 n
rlabel metal5 13040 -10960 13240 -10760 1 PIX204_IN
port 218 n
rlabel metal5 16040 -10960 16240 -10760 1 PIX205_IN
port 219 n
rlabel metal5 19040 -10960 19240 -10760 1 PIX206_IN
port 220 n
rlabel metal5 22040 -10960 22240 -10760 1 PIX207_IN
port 221 n
rlabel metal5 25040 -10960 25240 -10760 1 PIX208_IN
port 222 n
rlabel metal5 28040 -10960 28240 -10760 1 PIX209_IN
port 223 n
rlabel metal5 31040 -10960 31240 -10760 1 PIX210_IN
port 224 n
rlabel metal5 34040 -10960 34240 -10760 1 PIX211_IN
port 225 n
rlabel metal5 37040 -10960 37240 -10760 1 PIX212_IN
port 226 n
rlabel metal5 40040 -10960 40240 -10760 1 PIX213_IN
port 227 n
rlabel metal5 43040 -10960 43240 -10760 1 PIX214_IN
port 228 n
rlabel metal5 46040 -10960 46240 -10760 1 PIX215_IN
port 229 n
rlabel metal5 49040 -10960 49240 -10760 1 PIX216_IN
port 230 n
rlabel metal5 52040 -10960 52240 -10760 1 PIX217_IN
port 231 n
rlabel metal5 55040 -10960 55240 -10760 1 PIX218_IN
port 232 n
rlabel metal5 58040 -10960 58240 -10760 1 PIX219_IN
port 233 n
rlabel metal5 61040 -10960 61240 -10760 1 PIX220_IN
port 234 n
rlabel metal5 64040 -10960 64240 -10760 1 PIX221_IN
port 235 n
rlabel metal5 67040 -10960 67240 -10760 1 PIX222_IN
port 236 n
rlabel metal5 70040 -10960 70240 -10760 1 PIX223_IN
port 237 n
rlabel metal5 73040 -10960 73240 -10760 1 PIX224_IN
port 238 n
rlabel metal5 76040 -10960 76240 -10760 1 PIX225_IN
port 239 n
rlabel metal5 79040 -10960 79240 -10760 1 PIX226_IN
port 240 n
rlabel metal5 82040 -10960 82240 -10760 1 PIX227_IN
port 241 n
rlabel metal5 85040 -10960 85240 -10760 1 PIX228_IN
port 242 n
rlabel metal5 88040 -10960 88240 -10760 1 PIX229_IN
port 243 n
rlabel metal5 91040 -10960 91240 -10760 1 PIX230_IN
port 244 n
rlabel metal5 94040 -10960 94240 -10760 1 PIX231_IN
port 245 n
rlabel metal5 97040 -10960 97240 -10760 1 PIX232_IN
port 246 n
rlabel metal5 100040 -10960 100240 -10760 1 PIX233_IN
port 247 n
rlabel metal5 103040 -10960 103240 -10760 1 PIX234_IN
port 248 n
rlabel metal5 106040 -10960 106240 -10760 1 PIX235_IN
port 249 n
rlabel metal5 109040 -10960 109240 -10760 1 PIX236_IN
port 250 n
rlabel metal5 112040 -10960 112240 -10760 1 PIX237_IN
port 251 n
rlabel metal5 115040 -10960 115240 -10760 1 PIX238_IN
port 252 n
rlabel metal5 118040 -10960 118240 -10760 1 PIX239_IN
port 253 n
rlabel metal5 121040 -10960 121240 -10760 1 PIX240_IN
port 254 n
rlabel metal5 124040 -10960 124240 -10760 1 PIX241_IN
port 255 n
rlabel metal5 127040 -10960 127240 -10760 1 PIX242_IN
port 256 n
rlabel metal5 130040 -10960 130240 -10760 1 PIX243_IN
port 257 n
rlabel metal5 133040 -10960 133240 -10760 1 PIX244_IN
port 258 n
rlabel metal5 136040 -10960 136240 -10760 1 PIX245_IN
port 259 n
rlabel metal5 139040 -10960 139240 -10760 1 PIX246_IN
port 260 n
rlabel metal5 142040 -10960 142240 -10760 1 PIX247_IN
port 261 n
rlabel metal5 145040 -10960 145240 -10760 1 PIX248_IN
port 262 n
rlabel metal5 148040 -10960 148240 -10760 1 PIX249_IN
port 263 n
rlabel metal5 1040 -13960 1240 -13760 1 PIX250_IN
port 264 n
rlabel metal2 -3000 -13520 -3000 -13430 3 ROW_SEL5
port 265 e
rlabel metal5 4040 -13960 4240 -13760 1 PIX251_IN
port 266 n
rlabel metal5 7040 -13960 7240 -13760 1 PIX252_IN
port 267 n
rlabel metal5 10040 -13960 10240 -13760 1 PIX253_IN
port 268 n
rlabel metal5 13040 -13960 13240 -13760 1 PIX254_IN
port 269 n
rlabel metal5 16040 -13960 16240 -13760 1 PIX255_IN
port 270 n
rlabel metal5 19040 -13960 19240 -13760 1 PIX256_IN
port 271 n
rlabel metal5 22040 -13960 22240 -13760 1 PIX257_IN
port 272 n
rlabel metal5 25040 -13960 25240 -13760 1 PIX258_IN
port 273 n
rlabel metal5 28040 -13960 28240 -13760 1 PIX259_IN
port 274 n
rlabel metal5 31040 -13960 31240 -13760 1 PIX260_IN
port 275 n
rlabel metal5 34040 -13960 34240 -13760 1 PIX261_IN
port 276 n
rlabel metal5 37040 -13960 37240 -13760 1 PIX262_IN
port 277 n
rlabel metal5 40040 -13960 40240 -13760 1 PIX263_IN
port 278 n
rlabel metal5 43040 -13960 43240 -13760 1 PIX264_IN
port 279 n
rlabel metal5 46040 -13960 46240 -13760 1 PIX265_IN
port 280 n
rlabel metal5 49040 -13960 49240 -13760 1 PIX266_IN
port 281 n
rlabel metal5 52040 -13960 52240 -13760 1 PIX267_IN
port 282 n
rlabel metal5 55040 -13960 55240 -13760 1 PIX268_IN
port 283 n
rlabel metal5 58040 -13960 58240 -13760 1 PIX269_IN
port 284 n
rlabel metal5 61040 -13960 61240 -13760 1 PIX270_IN
port 285 n
rlabel metal5 64040 -13960 64240 -13760 1 PIX271_IN
port 286 n
rlabel metal5 67040 -13960 67240 -13760 1 PIX272_IN
port 287 n
rlabel metal5 70040 -13960 70240 -13760 1 PIX273_IN
port 288 n
rlabel metal5 73040 -13960 73240 -13760 1 PIX274_IN
port 289 n
rlabel metal5 76040 -13960 76240 -13760 1 PIX275_IN
port 290 n
rlabel metal5 79040 -13960 79240 -13760 1 PIX276_IN
port 291 n
rlabel metal5 82040 -13960 82240 -13760 1 PIX277_IN
port 292 n
rlabel metal5 85040 -13960 85240 -13760 1 PIX278_IN
port 293 n
rlabel metal5 88040 -13960 88240 -13760 1 PIX279_IN
port 294 n
rlabel metal5 91040 -13960 91240 -13760 1 PIX280_IN
port 295 n
rlabel metal5 94040 -13960 94240 -13760 1 PIX281_IN
port 296 n
rlabel metal5 97040 -13960 97240 -13760 1 PIX282_IN
port 297 n
rlabel metal5 100040 -13960 100240 -13760 1 PIX283_IN
port 298 n
rlabel metal5 103040 -13960 103240 -13760 1 PIX284_IN
port 299 n
rlabel metal5 106040 -13960 106240 -13760 1 PIX285_IN
port 300 n
rlabel metal5 109040 -13960 109240 -13760 1 PIX286_IN
port 301 n
rlabel metal5 112040 -13960 112240 -13760 1 PIX287_IN
port 302 n
rlabel metal5 115040 -13960 115240 -13760 1 PIX288_IN
port 303 n
rlabel metal5 118040 -13960 118240 -13760 1 PIX289_IN
port 304 n
rlabel metal5 121040 -13960 121240 -13760 1 PIX290_IN
port 305 n
rlabel metal5 124040 -13960 124240 -13760 1 PIX291_IN
port 306 n
rlabel metal5 127040 -13960 127240 -13760 1 PIX292_IN
port 307 n
rlabel metal5 130040 -13960 130240 -13760 1 PIX293_IN
port 308 n
rlabel metal5 133040 -13960 133240 -13760 1 PIX294_IN
port 309 n
rlabel metal5 136040 -13960 136240 -13760 1 PIX295_IN
port 310 n
rlabel metal5 139040 -13960 139240 -13760 1 PIX296_IN
port 311 n
rlabel metal5 142040 -13960 142240 -13760 1 PIX297_IN
port 312 n
rlabel metal5 145040 -13960 145240 -13760 1 PIX298_IN
port 313 n
rlabel metal5 148040 -13960 148240 -13760 1 PIX299_IN
port 314 n
rlabel metal5 1040 -16960 1240 -16760 1 PIX300_IN
port 315 n
rlabel metal2 -3000 -16520 -3000 -16430 3 ROW_SEL6
port 316 e
rlabel metal5 4040 -16960 4240 -16760 1 PIX301_IN
port 317 n
rlabel metal5 7040 -16960 7240 -16760 1 PIX302_IN
port 318 n
rlabel metal5 10040 -16960 10240 -16760 1 PIX303_IN
port 319 n
rlabel metal5 13040 -16960 13240 -16760 1 PIX304_IN
port 320 n
rlabel metal5 16040 -16960 16240 -16760 1 PIX305_IN
port 321 n
rlabel metal5 19040 -16960 19240 -16760 1 PIX306_IN
port 322 n
rlabel metal5 22040 -16960 22240 -16760 1 PIX307_IN
port 323 n
rlabel metal5 25040 -16960 25240 -16760 1 PIX308_IN
port 324 n
rlabel metal5 28040 -16960 28240 -16760 1 PIX309_IN
port 325 n
rlabel metal5 31040 -16960 31240 -16760 1 PIX310_IN
port 326 n
rlabel metal5 34040 -16960 34240 -16760 1 PIX311_IN
port 327 n
rlabel metal5 37040 -16960 37240 -16760 1 PIX312_IN
port 328 n
rlabel metal5 40040 -16960 40240 -16760 1 PIX313_IN
port 329 n
rlabel metal5 43040 -16960 43240 -16760 1 PIX314_IN
port 330 n
rlabel metal5 46040 -16960 46240 -16760 1 PIX315_IN
port 331 n
rlabel metal5 49040 -16960 49240 -16760 1 PIX316_IN
port 332 n
rlabel metal5 52040 -16960 52240 -16760 1 PIX317_IN
port 333 n
rlabel metal5 55040 -16960 55240 -16760 1 PIX318_IN
port 334 n
rlabel metal5 58040 -16960 58240 -16760 1 PIX319_IN
port 335 n
rlabel metal5 61040 -16960 61240 -16760 1 PIX320_IN
port 336 n
rlabel metal5 64040 -16960 64240 -16760 1 PIX321_IN
port 337 n
rlabel metal5 67040 -16960 67240 -16760 1 PIX322_IN
port 338 n
rlabel metal5 70040 -16960 70240 -16760 1 PIX323_IN
port 339 n
rlabel metal5 73040 -16960 73240 -16760 1 PIX324_IN
port 340 n
rlabel metal5 76040 -16960 76240 -16760 1 PIX325_IN
port 341 n
rlabel metal5 79040 -16960 79240 -16760 1 PIX326_IN
port 342 n
rlabel metal5 82040 -16960 82240 -16760 1 PIX327_IN
port 343 n
rlabel metal5 85040 -16960 85240 -16760 1 PIX328_IN
port 344 n
rlabel metal5 88040 -16960 88240 -16760 1 PIX329_IN
port 345 n
rlabel metal5 91040 -16960 91240 -16760 1 PIX330_IN
port 346 n
rlabel metal5 94040 -16960 94240 -16760 1 PIX331_IN
port 347 n
rlabel metal5 97040 -16960 97240 -16760 1 PIX332_IN
port 348 n
rlabel metal5 100040 -16960 100240 -16760 1 PIX333_IN
port 349 n
rlabel metal5 103040 -16960 103240 -16760 1 PIX334_IN
port 350 n
rlabel metal5 106040 -16960 106240 -16760 1 PIX335_IN
port 351 n
rlabel metal5 109040 -16960 109240 -16760 1 PIX336_IN
port 352 n
rlabel metal5 112040 -16960 112240 -16760 1 PIX337_IN
port 353 n
rlabel metal5 115040 -16960 115240 -16760 1 PIX338_IN
port 354 n
rlabel metal5 118040 -16960 118240 -16760 1 PIX339_IN
port 355 n
rlabel metal5 121040 -16960 121240 -16760 1 PIX340_IN
port 356 n
rlabel metal5 124040 -16960 124240 -16760 1 PIX341_IN
port 357 n
rlabel metal5 127040 -16960 127240 -16760 1 PIX342_IN
port 358 n
rlabel metal5 130040 -16960 130240 -16760 1 PIX343_IN
port 359 n
rlabel metal5 133040 -16960 133240 -16760 1 PIX344_IN
port 360 n
rlabel metal5 136040 -16960 136240 -16760 1 PIX345_IN
port 361 n
rlabel metal5 139040 -16960 139240 -16760 1 PIX346_IN
port 362 n
rlabel metal5 142040 -16960 142240 -16760 1 PIX347_IN
port 363 n
rlabel metal5 145040 -16960 145240 -16760 1 PIX348_IN
port 364 n
rlabel metal5 148040 -16960 148240 -16760 1 PIX349_IN
port 365 n
rlabel metal5 1040 -19960 1240 -19760 1 PIX350_IN
port 366 n
rlabel metal2 -3000 -19520 -3000 -19430 3 ROW_SEL7
port 367 e
rlabel metal5 4040 -19960 4240 -19760 1 PIX351_IN
port 368 n
rlabel metal5 7040 -19960 7240 -19760 1 PIX352_IN
port 369 n
rlabel metal5 10040 -19960 10240 -19760 1 PIX353_IN
port 370 n
rlabel metal5 13040 -19960 13240 -19760 1 PIX354_IN
port 371 n
rlabel metal5 16040 -19960 16240 -19760 1 PIX355_IN
port 372 n
rlabel metal5 19040 -19960 19240 -19760 1 PIX356_IN
port 373 n
rlabel metal5 22040 -19960 22240 -19760 1 PIX357_IN
port 374 n
rlabel metal5 25040 -19960 25240 -19760 1 PIX358_IN
port 375 n
rlabel metal5 28040 -19960 28240 -19760 1 PIX359_IN
port 376 n
rlabel metal5 31040 -19960 31240 -19760 1 PIX360_IN
port 377 n
rlabel metal5 34040 -19960 34240 -19760 1 PIX361_IN
port 378 n
rlabel metal5 37040 -19960 37240 -19760 1 PIX362_IN
port 379 n
rlabel metal5 40040 -19960 40240 -19760 1 PIX363_IN
port 380 n
rlabel metal5 43040 -19960 43240 -19760 1 PIX364_IN
port 381 n
rlabel metal5 46040 -19960 46240 -19760 1 PIX365_IN
port 382 n
rlabel metal5 49040 -19960 49240 -19760 1 PIX366_IN
port 383 n
rlabel metal5 52040 -19960 52240 -19760 1 PIX367_IN
port 384 n
rlabel metal5 55040 -19960 55240 -19760 1 PIX368_IN
port 385 n
rlabel metal5 58040 -19960 58240 -19760 1 PIX369_IN
port 386 n
rlabel metal5 61040 -19960 61240 -19760 1 PIX370_IN
port 387 n
rlabel metal5 64040 -19960 64240 -19760 1 PIX371_IN
port 388 n
rlabel metal5 67040 -19960 67240 -19760 1 PIX372_IN
port 389 n
rlabel metal5 70040 -19960 70240 -19760 1 PIX373_IN
port 390 n
rlabel metal5 73040 -19960 73240 -19760 1 PIX374_IN
port 391 n
rlabel metal5 76040 -19960 76240 -19760 1 PIX375_IN
port 392 n
rlabel metal5 79040 -19960 79240 -19760 1 PIX376_IN
port 393 n
rlabel metal5 82040 -19960 82240 -19760 1 PIX377_IN
port 394 n
rlabel metal5 85040 -19960 85240 -19760 1 PIX378_IN
port 395 n
rlabel metal5 88040 -19960 88240 -19760 1 PIX379_IN
port 396 n
rlabel metal5 91040 -19960 91240 -19760 1 PIX380_IN
port 397 n
rlabel metal5 94040 -19960 94240 -19760 1 PIX381_IN
port 398 n
rlabel metal5 97040 -19960 97240 -19760 1 PIX382_IN
port 399 n
rlabel metal5 100040 -19960 100240 -19760 1 PIX383_IN
port 400 n
rlabel metal5 103040 -19960 103240 -19760 1 PIX384_IN
port 401 n
rlabel metal5 106040 -19960 106240 -19760 1 PIX385_IN
port 402 n
rlabel metal5 109040 -19960 109240 -19760 1 PIX386_IN
port 403 n
rlabel metal5 112040 -19960 112240 -19760 1 PIX387_IN
port 404 n
rlabel metal5 115040 -19960 115240 -19760 1 PIX388_IN
port 405 n
rlabel metal5 118040 -19960 118240 -19760 1 PIX389_IN
port 406 n
rlabel metal5 121040 -19960 121240 -19760 1 PIX390_IN
port 407 n
rlabel metal5 124040 -19960 124240 -19760 1 PIX391_IN
port 408 n
rlabel metal5 127040 -19960 127240 -19760 1 PIX392_IN
port 409 n
rlabel metal5 130040 -19960 130240 -19760 1 PIX393_IN
port 410 n
rlabel metal5 133040 -19960 133240 -19760 1 PIX394_IN
port 411 n
rlabel metal5 136040 -19960 136240 -19760 1 PIX395_IN
port 412 n
rlabel metal5 139040 -19960 139240 -19760 1 PIX396_IN
port 413 n
rlabel metal5 142040 -19960 142240 -19760 1 PIX397_IN
port 414 n
rlabel metal5 145040 -19960 145240 -19760 1 PIX398_IN
port 415 n
rlabel metal5 148040 -19960 148240 -19760 1 PIX399_IN
port 416 n
rlabel metal5 1040 -22960 1240 -22760 1 PIX400_IN
port 417 n
rlabel metal2 -3000 -22520 -3000 -22430 3 ROW_SEL8
port 418 e
rlabel metal5 4040 -22960 4240 -22760 1 PIX401_IN
port 419 n
rlabel metal5 7040 -22960 7240 -22760 1 PIX402_IN
port 420 n
rlabel metal5 10040 -22960 10240 -22760 1 PIX403_IN
port 421 n
rlabel metal5 13040 -22960 13240 -22760 1 PIX404_IN
port 422 n
rlabel metal5 16040 -22960 16240 -22760 1 PIX405_IN
port 423 n
rlabel metal5 19040 -22960 19240 -22760 1 PIX406_IN
port 424 n
rlabel metal5 22040 -22960 22240 -22760 1 PIX407_IN
port 425 n
rlabel metal5 25040 -22960 25240 -22760 1 PIX408_IN
port 426 n
rlabel metal5 28040 -22960 28240 -22760 1 PIX409_IN
port 427 n
rlabel metal5 31040 -22960 31240 -22760 1 PIX410_IN
port 428 n
rlabel metal5 34040 -22960 34240 -22760 1 PIX411_IN
port 429 n
rlabel metal5 37040 -22960 37240 -22760 1 PIX412_IN
port 430 n
rlabel metal5 40040 -22960 40240 -22760 1 PIX413_IN
port 431 n
rlabel metal5 43040 -22960 43240 -22760 1 PIX414_IN
port 432 n
rlabel metal5 46040 -22960 46240 -22760 1 PIX415_IN
port 433 n
rlabel metal5 49040 -22960 49240 -22760 1 PIX416_IN
port 434 n
rlabel metal5 52040 -22960 52240 -22760 1 PIX417_IN
port 435 n
rlabel metal5 55040 -22960 55240 -22760 1 PIX418_IN
port 436 n
rlabel metal5 58040 -22960 58240 -22760 1 PIX419_IN
port 437 n
rlabel metal5 61040 -22960 61240 -22760 1 PIX420_IN
port 438 n
rlabel metal5 64040 -22960 64240 -22760 1 PIX421_IN
port 439 n
rlabel metal5 67040 -22960 67240 -22760 1 PIX422_IN
port 440 n
rlabel metal5 70040 -22960 70240 -22760 1 PIX423_IN
port 441 n
rlabel metal5 73040 -22960 73240 -22760 1 PIX424_IN
port 442 n
rlabel metal5 76040 -22960 76240 -22760 1 PIX425_IN
port 443 n
rlabel metal5 79040 -22960 79240 -22760 1 PIX426_IN
port 444 n
rlabel metal5 82040 -22960 82240 -22760 1 PIX427_IN
port 445 n
rlabel metal5 85040 -22960 85240 -22760 1 PIX428_IN
port 446 n
rlabel metal5 88040 -22960 88240 -22760 1 PIX429_IN
port 447 n
rlabel metal5 91040 -22960 91240 -22760 1 PIX430_IN
port 448 n
rlabel metal5 94040 -22960 94240 -22760 1 PIX431_IN
port 449 n
rlabel metal5 97040 -22960 97240 -22760 1 PIX432_IN
port 450 n
rlabel metal5 100040 -22960 100240 -22760 1 PIX433_IN
port 451 n
rlabel metal5 103040 -22960 103240 -22760 1 PIX434_IN
port 452 n
rlabel metal5 106040 -22960 106240 -22760 1 PIX435_IN
port 453 n
rlabel metal5 109040 -22960 109240 -22760 1 PIX436_IN
port 454 n
rlabel metal5 112040 -22960 112240 -22760 1 PIX437_IN
port 455 n
rlabel metal5 115040 -22960 115240 -22760 1 PIX438_IN
port 456 n
rlabel metal5 118040 -22960 118240 -22760 1 PIX439_IN
port 457 n
rlabel metal5 121040 -22960 121240 -22760 1 PIX440_IN
port 458 n
rlabel metal5 124040 -22960 124240 -22760 1 PIX441_IN
port 459 n
rlabel metal5 127040 -22960 127240 -22760 1 PIX442_IN
port 460 n
rlabel metal5 130040 -22960 130240 -22760 1 PIX443_IN
port 461 n
rlabel metal5 133040 -22960 133240 -22760 1 PIX444_IN
port 462 n
rlabel metal5 136040 -22960 136240 -22760 1 PIX445_IN
port 463 n
rlabel metal5 139040 -22960 139240 -22760 1 PIX446_IN
port 464 n
rlabel metal5 142040 -22960 142240 -22760 1 PIX447_IN
port 465 n
rlabel metal5 145040 -22960 145240 -22760 1 PIX448_IN
port 466 n
rlabel metal5 148040 -22960 148240 -22760 1 PIX449_IN
port 467 n
rlabel metal5 1040 -25960 1240 -25760 1 PIX450_IN
port 468 n
rlabel metal2 -3000 -25520 -3000 -25430 3 ROW_SEL9
port 469 e
rlabel metal5 4040 -25960 4240 -25760 1 PIX451_IN
port 470 n
rlabel metal5 7040 -25960 7240 -25760 1 PIX452_IN
port 471 n
rlabel metal5 10040 -25960 10240 -25760 1 PIX453_IN
port 472 n
rlabel metal5 13040 -25960 13240 -25760 1 PIX454_IN
port 473 n
rlabel metal5 16040 -25960 16240 -25760 1 PIX455_IN
port 474 n
rlabel metal5 19040 -25960 19240 -25760 1 PIX456_IN
port 475 n
rlabel metal5 22040 -25960 22240 -25760 1 PIX457_IN
port 476 n
rlabel metal5 25040 -25960 25240 -25760 1 PIX458_IN
port 477 n
rlabel metal5 28040 -25960 28240 -25760 1 PIX459_IN
port 478 n
rlabel metal5 31040 -25960 31240 -25760 1 PIX460_IN
port 479 n
rlabel metal5 34040 -25960 34240 -25760 1 PIX461_IN
port 480 n
rlabel metal5 37040 -25960 37240 -25760 1 PIX462_IN
port 481 n
rlabel metal5 40040 -25960 40240 -25760 1 PIX463_IN
port 482 n
rlabel metal5 43040 -25960 43240 -25760 1 PIX464_IN
port 483 n
rlabel metal5 46040 -25960 46240 -25760 1 PIX465_IN
port 484 n
rlabel metal5 49040 -25960 49240 -25760 1 PIX466_IN
port 485 n
rlabel metal5 52040 -25960 52240 -25760 1 PIX467_IN
port 486 n
rlabel metal5 55040 -25960 55240 -25760 1 PIX468_IN
port 487 n
rlabel metal5 58040 -25960 58240 -25760 1 PIX469_IN
port 488 n
rlabel metal5 61040 -25960 61240 -25760 1 PIX470_IN
port 489 n
rlabel metal5 64040 -25960 64240 -25760 1 PIX471_IN
port 490 n
rlabel metal5 67040 -25960 67240 -25760 1 PIX472_IN
port 491 n
rlabel metal5 70040 -25960 70240 -25760 1 PIX473_IN
port 492 n
rlabel metal5 73040 -25960 73240 -25760 1 PIX474_IN
port 493 n
rlabel metal5 76040 -25960 76240 -25760 1 PIX475_IN
port 494 n
rlabel metal5 79040 -25960 79240 -25760 1 PIX476_IN
port 495 n
rlabel metal5 82040 -25960 82240 -25760 1 PIX477_IN
port 496 n
rlabel metal5 85040 -25960 85240 -25760 1 PIX478_IN
port 497 n
rlabel metal5 88040 -25960 88240 -25760 1 PIX479_IN
port 498 n
rlabel metal5 91040 -25960 91240 -25760 1 PIX480_IN
port 499 n
rlabel metal5 94040 -25960 94240 -25760 1 PIX481_IN
port 500 n
rlabel metal5 97040 -25960 97240 -25760 1 PIX482_IN
port 501 n
rlabel metal5 100040 -25960 100240 -25760 1 PIX483_IN
port 502 n
rlabel metal5 103040 -25960 103240 -25760 1 PIX484_IN
port 503 n
rlabel metal5 106040 -25960 106240 -25760 1 PIX485_IN
port 504 n
rlabel metal5 109040 -25960 109240 -25760 1 PIX486_IN
port 505 n
rlabel metal5 112040 -25960 112240 -25760 1 PIX487_IN
port 506 n
rlabel metal5 115040 -25960 115240 -25760 1 PIX488_IN
port 507 n
rlabel metal5 118040 -25960 118240 -25760 1 PIX489_IN
port 508 n
rlabel metal5 121040 -25960 121240 -25760 1 PIX490_IN
port 509 n
rlabel metal5 124040 -25960 124240 -25760 1 PIX491_IN
port 510 n
rlabel metal5 127040 -25960 127240 -25760 1 PIX492_IN
port 511 n
rlabel metal5 130040 -25960 130240 -25760 1 PIX493_IN
port 512 n
rlabel metal5 133040 -25960 133240 -25760 1 PIX494_IN
port 513 n
rlabel metal5 136040 -25960 136240 -25760 1 PIX495_IN
port 514 n
rlabel metal5 139040 -25960 139240 -25760 1 PIX496_IN
port 515 n
rlabel metal5 142040 -25960 142240 -25760 1 PIX497_IN
port 516 n
rlabel metal5 145040 -25960 145240 -25760 1 PIX498_IN
port 517 n
rlabel metal5 148040 -25960 148240 -25760 1 PIX499_IN
port 518 n
rlabel metal5 1040 -28960 1240 -28760 1 PIX500_IN
port 519 n
rlabel metal2 -3000 -28520 -3000 -28430 3 ROW_SEL10
port 520 e
rlabel metal5 4040 -28960 4240 -28760 1 PIX501_IN
port 521 n
rlabel metal5 7040 -28960 7240 -28760 1 PIX502_IN
port 522 n
rlabel metal5 10040 -28960 10240 -28760 1 PIX503_IN
port 523 n
rlabel metal5 13040 -28960 13240 -28760 1 PIX504_IN
port 524 n
rlabel metal5 16040 -28960 16240 -28760 1 PIX505_IN
port 525 n
rlabel metal5 19040 -28960 19240 -28760 1 PIX506_IN
port 526 n
rlabel metal5 22040 -28960 22240 -28760 1 PIX507_IN
port 527 n
rlabel metal5 25040 -28960 25240 -28760 1 PIX508_IN
port 528 n
rlabel metal5 28040 -28960 28240 -28760 1 PIX509_IN
port 529 n
rlabel metal5 31040 -28960 31240 -28760 1 PIX510_IN
port 530 n
rlabel metal5 34040 -28960 34240 -28760 1 PIX511_IN
port 531 n
rlabel metal5 37040 -28960 37240 -28760 1 PIX512_IN
port 532 n
rlabel metal5 40040 -28960 40240 -28760 1 PIX513_IN
port 533 n
rlabel metal5 43040 -28960 43240 -28760 1 PIX514_IN
port 534 n
rlabel metal5 46040 -28960 46240 -28760 1 PIX515_IN
port 535 n
rlabel metal5 49040 -28960 49240 -28760 1 PIX516_IN
port 536 n
rlabel metal5 52040 -28960 52240 -28760 1 PIX517_IN
port 537 n
rlabel metal5 55040 -28960 55240 -28760 1 PIX518_IN
port 538 n
rlabel metal5 58040 -28960 58240 -28760 1 PIX519_IN
port 539 n
rlabel metal5 61040 -28960 61240 -28760 1 PIX520_IN
port 540 n
rlabel metal5 64040 -28960 64240 -28760 1 PIX521_IN
port 541 n
rlabel metal5 67040 -28960 67240 -28760 1 PIX522_IN
port 542 n
rlabel metal5 70040 -28960 70240 -28760 1 PIX523_IN
port 543 n
rlabel metal5 73040 -28960 73240 -28760 1 PIX524_IN
port 544 n
rlabel metal5 76040 -28960 76240 -28760 1 PIX525_IN
port 545 n
rlabel metal5 79040 -28960 79240 -28760 1 PIX526_IN
port 546 n
rlabel metal5 82040 -28960 82240 -28760 1 PIX527_IN
port 547 n
rlabel metal5 85040 -28960 85240 -28760 1 PIX528_IN
port 548 n
rlabel metal5 88040 -28960 88240 -28760 1 PIX529_IN
port 549 n
rlabel metal5 91040 -28960 91240 -28760 1 PIX530_IN
port 550 n
rlabel metal5 94040 -28960 94240 -28760 1 PIX531_IN
port 551 n
rlabel metal5 97040 -28960 97240 -28760 1 PIX532_IN
port 552 n
rlabel metal5 100040 -28960 100240 -28760 1 PIX533_IN
port 553 n
rlabel metal5 103040 -28960 103240 -28760 1 PIX534_IN
port 554 n
rlabel metal5 106040 -28960 106240 -28760 1 PIX535_IN
port 555 n
rlabel metal5 109040 -28960 109240 -28760 1 PIX536_IN
port 556 n
rlabel metal5 112040 -28960 112240 -28760 1 PIX537_IN
port 557 n
rlabel metal5 115040 -28960 115240 -28760 1 PIX538_IN
port 558 n
rlabel metal5 118040 -28960 118240 -28760 1 PIX539_IN
port 559 n
rlabel metal5 121040 -28960 121240 -28760 1 PIX540_IN
port 560 n
rlabel metal5 124040 -28960 124240 -28760 1 PIX541_IN
port 561 n
rlabel metal5 127040 -28960 127240 -28760 1 PIX542_IN
port 562 n
rlabel metal5 130040 -28960 130240 -28760 1 PIX543_IN
port 563 n
rlabel metal5 133040 -28960 133240 -28760 1 PIX544_IN
port 564 n
rlabel metal5 136040 -28960 136240 -28760 1 PIX545_IN
port 565 n
rlabel metal5 139040 -28960 139240 -28760 1 PIX546_IN
port 566 n
rlabel metal5 142040 -28960 142240 -28760 1 PIX547_IN
port 567 n
rlabel metal5 145040 -28960 145240 -28760 1 PIX548_IN
port 568 n
rlabel metal5 148040 -28960 148240 -28760 1 PIX549_IN
port 569 n
rlabel metal5 1040 -31960 1240 -31760 1 PIX550_IN
port 570 n
rlabel metal2 -3000 -31520 -3000 -31430 3 ROW_SEL11
port 571 e
rlabel metal5 4040 -31960 4240 -31760 1 PIX551_IN
port 572 n
rlabel metal5 7040 -31960 7240 -31760 1 PIX552_IN
port 573 n
rlabel metal5 10040 -31960 10240 -31760 1 PIX553_IN
port 574 n
rlabel metal5 13040 -31960 13240 -31760 1 PIX554_IN
port 575 n
rlabel metal5 16040 -31960 16240 -31760 1 PIX555_IN
port 576 n
rlabel metal5 19040 -31960 19240 -31760 1 PIX556_IN
port 577 n
rlabel metal5 22040 -31960 22240 -31760 1 PIX557_IN
port 578 n
rlabel metal5 25040 -31960 25240 -31760 1 PIX558_IN
port 579 n
rlabel metal5 28040 -31960 28240 -31760 1 PIX559_IN
port 580 n
rlabel metal5 31040 -31960 31240 -31760 1 PIX560_IN
port 581 n
rlabel metal5 34040 -31960 34240 -31760 1 PIX561_IN
port 582 n
rlabel metal5 37040 -31960 37240 -31760 1 PIX562_IN
port 583 n
rlabel metal5 40040 -31960 40240 -31760 1 PIX563_IN
port 584 n
rlabel metal5 43040 -31960 43240 -31760 1 PIX564_IN
port 585 n
rlabel metal5 46040 -31960 46240 -31760 1 PIX565_IN
port 586 n
rlabel metal5 49040 -31960 49240 -31760 1 PIX566_IN
port 587 n
rlabel metal5 52040 -31960 52240 -31760 1 PIX567_IN
port 588 n
rlabel metal5 55040 -31960 55240 -31760 1 PIX568_IN
port 589 n
rlabel metal5 58040 -31960 58240 -31760 1 PIX569_IN
port 590 n
rlabel metal5 61040 -31960 61240 -31760 1 PIX570_IN
port 591 n
rlabel metal5 64040 -31960 64240 -31760 1 PIX571_IN
port 592 n
rlabel metal5 67040 -31960 67240 -31760 1 PIX572_IN
port 593 n
rlabel metal5 70040 -31960 70240 -31760 1 PIX573_IN
port 594 n
rlabel metal5 73040 -31960 73240 -31760 1 PIX574_IN
port 595 n
rlabel metal5 76040 -31960 76240 -31760 1 PIX575_IN
port 596 n
rlabel metal5 79040 -31960 79240 -31760 1 PIX576_IN
port 597 n
rlabel metal5 82040 -31960 82240 -31760 1 PIX577_IN
port 598 n
rlabel metal5 85040 -31960 85240 -31760 1 PIX578_IN
port 599 n
rlabel metal5 88040 -31960 88240 -31760 1 PIX579_IN
port 600 n
rlabel metal5 91040 -31960 91240 -31760 1 PIX580_IN
port 601 n
rlabel metal5 94040 -31960 94240 -31760 1 PIX581_IN
port 602 n
rlabel metal5 97040 -31960 97240 -31760 1 PIX582_IN
port 603 n
rlabel metal5 100040 -31960 100240 -31760 1 PIX583_IN
port 604 n
rlabel metal5 103040 -31960 103240 -31760 1 PIX584_IN
port 605 n
rlabel metal5 106040 -31960 106240 -31760 1 PIX585_IN
port 606 n
rlabel metal5 109040 -31960 109240 -31760 1 PIX586_IN
port 607 n
rlabel metal5 112040 -31960 112240 -31760 1 PIX587_IN
port 608 n
rlabel metal5 115040 -31960 115240 -31760 1 PIX588_IN
port 609 n
rlabel metal5 118040 -31960 118240 -31760 1 PIX589_IN
port 610 n
rlabel metal5 121040 -31960 121240 -31760 1 PIX590_IN
port 611 n
rlabel metal5 124040 -31960 124240 -31760 1 PIX591_IN
port 612 n
rlabel metal5 127040 -31960 127240 -31760 1 PIX592_IN
port 613 n
rlabel metal5 130040 -31960 130240 -31760 1 PIX593_IN
port 614 n
rlabel metal5 133040 -31960 133240 -31760 1 PIX594_IN
port 615 n
rlabel metal5 136040 -31960 136240 -31760 1 PIX595_IN
port 616 n
rlabel metal5 139040 -31960 139240 -31760 1 PIX596_IN
port 617 n
rlabel metal5 142040 -31960 142240 -31760 1 PIX597_IN
port 618 n
rlabel metal5 145040 -31960 145240 -31760 1 PIX598_IN
port 619 n
rlabel metal5 148040 -31960 148240 -31760 1 PIX599_IN
port 620 n
rlabel metal5 1040 -34960 1240 -34760 1 PIX600_IN
port 621 n
rlabel metal2 -3000 -34520 -3000 -34430 3 ROW_SEL12
port 622 e
rlabel metal5 4040 -34960 4240 -34760 1 PIX601_IN
port 623 n
rlabel metal5 7040 -34960 7240 -34760 1 PIX602_IN
port 624 n
rlabel metal5 10040 -34960 10240 -34760 1 PIX603_IN
port 625 n
rlabel metal5 13040 -34960 13240 -34760 1 PIX604_IN
port 626 n
rlabel metal5 16040 -34960 16240 -34760 1 PIX605_IN
port 627 n
rlabel metal5 19040 -34960 19240 -34760 1 PIX606_IN
port 628 n
rlabel metal5 22040 -34960 22240 -34760 1 PIX607_IN
port 629 n
rlabel metal5 25040 -34960 25240 -34760 1 PIX608_IN
port 630 n
rlabel metal5 28040 -34960 28240 -34760 1 PIX609_IN
port 631 n
rlabel metal5 31040 -34960 31240 -34760 1 PIX610_IN
port 632 n
rlabel metal5 34040 -34960 34240 -34760 1 PIX611_IN
port 633 n
rlabel metal5 37040 -34960 37240 -34760 1 PIX612_IN
port 634 n
rlabel metal5 40040 -34960 40240 -34760 1 PIX613_IN
port 635 n
rlabel metal5 43040 -34960 43240 -34760 1 PIX614_IN
port 636 n
rlabel metal5 46040 -34960 46240 -34760 1 PIX615_IN
port 637 n
rlabel metal5 49040 -34960 49240 -34760 1 PIX616_IN
port 638 n
rlabel metal5 52040 -34960 52240 -34760 1 PIX617_IN
port 639 n
rlabel metal5 55040 -34960 55240 -34760 1 PIX618_IN
port 640 n
rlabel metal5 58040 -34960 58240 -34760 1 PIX619_IN
port 641 n
rlabel metal5 61040 -34960 61240 -34760 1 PIX620_IN
port 642 n
rlabel metal5 64040 -34960 64240 -34760 1 PIX621_IN
port 643 n
rlabel metal5 67040 -34960 67240 -34760 1 PIX622_IN
port 644 n
rlabel metal5 70040 -34960 70240 -34760 1 PIX623_IN
port 645 n
rlabel metal5 73040 -34960 73240 -34760 1 PIX624_IN
port 646 n
rlabel metal5 76040 -34960 76240 -34760 1 PIX625_IN
port 647 n
rlabel metal5 79040 -34960 79240 -34760 1 PIX626_IN
port 648 n
rlabel metal5 82040 -34960 82240 -34760 1 PIX627_IN
port 649 n
rlabel metal5 85040 -34960 85240 -34760 1 PIX628_IN
port 650 n
rlabel metal5 88040 -34960 88240 -34760 1 PIX629_IN
port 651 n
rlabel metal5 91040 -34960 91240 -34760 1 PIX630_IN
port 652 n
rlabel metal5 94040 -34960 94240 -34760 1 PIX631_IN
port 653 n
rlabel metal5 97040 -34960 97240 -34760 1 PIX632_IN
port 654 n
rlabel metal5 100040 -34960 100240 -34760 1 PIX633_IN
port 655 n
rlabel metal5 103040 -34960 103240 -34760 1 PIX634_IN
port 656 n
rlabel metal5 106040 -34960 106240 -34760 1 PIX635_IN
port 657 n
rlabel metal5 109040 -34960 109240 -34760 1 PIX636_IN
port 658 n
rlabel metal5 112040 -34960 112240 -34760 1 PIX637_IN
port 659 n
rlabel metal5 115040 -34960 115240 -34760 1 PIX638_IN
port 660 n
rlabel metal5 118040 -34960 118240 -34760 1 PIX639_IN
port 661 n
rlabel metal5 121040 -34960 121240 -34760 1 PIX640_IN
port 662 n
rlabel metal5 124040 -34960 124240 -34760 1 PIX641_IN
port 663 n
rlabel metal5 127040 -34960 127240 -34760 1 PIX642_IN
port 664 n
rlabel metal5 130040 -34960 130240 -34760 1 PIX643_IN
port 665 n
rlabel metal5 133040 -34960 133240 -34760 1 PIX644_IN
port 666 n
rlabel metal5 136040 -34960 136240 -34760 1 PIX645_IN
port 667 n
rlabel metal5 139040 -34960 139240 -34760 1 PIX646_IN
port 668 n
rlabel metal5 142040 -34960 142240 -34760 1 PIX647_IN
port 669 n
rlabel metal5 145040 -34960 145240 -34760 1 PIX648_IN
port 670 n
rlabel metal5 148040 -34960 148240 -34760 1 PIX649_IN
port 671 n
rlabel metal5 1040 -37960 1240 -37760 1 PIX650_IN
port 672 n
rlabel metal2 -3000 -37520 -3000 -37430 3 ROW_SEL13
port 673 e
rlabel metal5 4040 -37960 4240 -37760 1 PIX651_IN
port 674 n
rlabel metal5 7040 -37960 7240 -37760 1 PIX652_IN
port 675 n
rlabel metal5 10040 -37960 10240 -37760 1 PIX653_IN
port 676 n
rlabel metal5 13040 -37960 13240 -37760 1 PIX654_IN
port 677 n
rlabel metal5 16040 -37960 16240 -37760 1 PIX655_IN
port 678 n
rlabel metal5 19040 -37960 19240 -37760 1 PIX656_IN
port 679 n
rlabel metal5 22040 -37960 22240 -37760 1 PIX657_IN
port 680 n
rlabel metal5 25040 -37960 25240 -37760 1 PIX658_IN
port 681 n
rlabel metal5 28040 -37960 28240 -37760 1 PIX659_IN
port 682 n
rlabel metal5 31040 -37960 31240 -37760 1 PIX660_IN
port 683 n
rlabel metal5 34040 -37960 34240 -37760 1 PIX661_IN
port 684 n
rlabel metal5 37040 -37960 37240 -37760 1 PIX662_IN
port 685 n
rlabel metal5 40040 -37960 40240 -37760 1 PIX663_IN
port 686 n
rlabel metal5 43040 -37960 43240 -37760 1 PIX664_IN
port 687 n
rlabel metal5 46040 -37960 46240 -37760 1 PIX665_IN
port 688 n
rlabel metal5 49040 -37960 49240 -37760 1 PIX666_IN
port 689 n
rlabel metal5 52040 -37960 52240 -37760 1 PIX667_IN
port 690 n
rlabel metal5 55040 -37960 55240 -37760 1 PIX668_IN
port 691 n
rlabel metal5 58040 -37960 58240 -37760 1 PIX669_IN
port 692 n
rlabel metal5 61040 -37960 61240 -37760 1 PIX670_IN
port 693 n
rlabel metal5 64040 -37960 64240 -37760 1 PIX671_IN
port 694 n
rlabel metal5 67040 -37960 67240 -37760 1 PIX672_IN
port 695 n
rlabel metal5 70040 -37960 70240 -37760 1 PIX673_IN
port 696 n
rlabel metal5 73040 -37960 73240 -37760 1 PIX674_IN
port 697 n
rlabel metal5 76040 -37960 76240 -37760 1 PIX675_IN
port 698 n
rlabel metal5 79040 -37960 79240 -37760 1 PIX676_IN
port 699 n
rlabel metal5 82040 -37960 82240 -37760 1 PIX677_IN
port 700 n
rlabel metal5 85040 -37960 85240 -37760 1 PIX678_IN
port 701 n
rlabel metal5 88040 -37960 88240 -37760 1 PIX679_IN
port 702 n
rlabel metal5 91040 -37960 91240 -37760 1 PIX680_IN
port 703 n
rlabel metal5 94040 -37960 94240 -37760 1 PIX681_IN
port 704 n
rlabel metal5 97040 -37960 97240 -37760 1 PIX682_IN
port 705 n
rlabel metal5 100040 -37960 100240 -37760 1 PIX683_IN
port 706 n
rlabel metal5 103040 -37960 103240 -37760 1 PIX684_IN
port 707 n
rlabel metal5 106040 -37960 106240 -37760 1 PIX685_IN
port 708 n
rlabel metal5 109040 -37960 109240 -37760 1 PIX686_IN
port 709 n
rlabel metal5 112040 -37960 112240 -37760 1 PIX687_IN
port 710 n
rlabel metal5 115040 -37960 115240 -37760 1 PIX688_IN
port 711 n
rlabel metal5 118040 -37960 118240 -37760 1 PIX689_IN
port 712 n
rlabel metal5 121040 -37960 121240 -37760 1 PIX690_IN
port 713 n
rlabel metal5 124040 -37960 124240 -37760 1 PIX691_IN
port 714 n
rlabel metal5 127040 -37960 127240 -37760 1 PIX692_IN
port 715 n
rlabel metal5 130040 -37960 130240 -37760 1 PIX693_IN
port 716 n
rlabel metal5 133040 -37960 133240 -37760 1 PIX694_IN
port 717 n
rlabel metal5 136040 -37960 136240 -37760 1 PIX695_IN
port 718 n
rlabel metal5 139040 -37960 139240 -37760 1 PIX696_IN
port 719 n
rlabel metal5 142040 -37960 142240 -37760 1 PIX697_IN
port 720 n
rlabel metal5 145040 -37960 145240 -37760 1 PIX698_IN
port 721 n
rlabel metal5 148040 -37960 148240 -37760 1 PIX699_IN
port 722 n
rlabel metal5 1040 -40960 1240 -40760 1 PIX700_IN
port 723 n
rlabel metal2 -3000 -40520 -3000 -40430 3 ROW_SEL14
port 724 e
rlabel metal5 4040 -40960 4240 -40760 1 PIX701_IN
port 725 n
rlabel metal5 7040 -40960 7240 -40760 1 PIX702_IN
port 726 n
rlabel metal5 10040 -40960 10240 -40760 1 PIX703_IN
port 727 n
rlabel metal5 13040 -40960 13240 -40760 1 PIX704_IN
port 728 n
rlabel metal5 16040 -40960 16240 -40760 1 PIX705_IN
port 729 n
rlabel metal5 19040 -40960 19240 -40760 1 PIX706_IN
port 730 n
rlabel metal5 22040 -40960 22240 -40760 1 PIX707_IN
port 731 n
rlabel metal5 25040 -40960 25240 -40760 1 PIX708_IN
port 732 n
rlabel metal5 28040 -40960 28240 -40760 1 PIX709_IN
port 733 n
rlabel metal5 31040 -40960 31240 -40760 1 PIX710_IN
port 734 n
rlabel metal5 34040 -40960 34240 -40760 1 PIX711_IN
port 735 n
rlabel metal5 37040 -40960 37240 -40760 1 PIX712_IN
port 736 n
rlabel metal5 40040 -40960 40240 -40760 1 PIX713_IN
port 737 n
rlabel metal5 43040 -40960 43240 -40760 1 PIX714_IN
port 738 n
rlabel metal5 46040 -40960 46240 -40760 1 PIX715_IN
port 739 n
rlabel metal5 49040 -40960 49240 -40760 1 PIX716_IN
port 740 n
rlabel metal5 52040 -40960 52240 -40760 1 PIX717_IN
port 741 n
rlabel metal5 55040 -40960 55240 -40760 1 PIX718_IN
port 742 n
rlabel metal5 58040 -40960 58240 -40760 1 PIX719_IN
port 743 n
rlabel metal5 61040 -40960 61240 -40760 1 PIX720_IN
port 744 n
rlabel metal5 64040 -40960 64240 -40760 1 PIX721_IN
port 745 n
rlabel metal5 67040 -40960 67240 -40760 1 PIX722_IN
port 746 n
rlabel metal5 70040 -40960 70240 -40760 1 PIX723_IN
port 747 n
rlabel metal5 73040 -40960 73240 -40760 1 PIX724_IN
port 748 n
rlabel metal5 76040 -40960 76240 -40760 1 PIX725_IN
port 749 n
rlabel metal5 79040 -40960 79240 -40760 1 PIX726_IN
port 750 n
rlabel metal5 82040 -40960 82240 -40760 1 PIX727_IN
port 751 n
rlabel metal5 85040 -40960 85240 -40760 1 PIX728_IN
port 752 n
rlabel metal5 88040 -40960 88240 -40760 1 PIX729_IN
port 753 n
rlabel metal5 91040 -40960 91240 -40760 1 PIX730_IN
port 754 n
rlabel metal5 94040 -40960 94240 -40760 1 PIX731_IN
port 755 n
rlabel metal5 97040 -40960 97240 -40760 1 PIX732_IN
port 756 n
rlabel metal5 100040 -40960 100240 -40760 1 PIX733_IN
port 757 n
rlabel metal5 103040 -40960 103240 -40760 1 PIX734_IN
port 758 n
rlabel metal5 106040 -40960 106240 -40760 1 PIX735_IN
port 759 n
rlabel metal5 109040 -40960 109240 -40760 1 PIX736_IN
port 760 n
rlabel metal5 112040 -40960 112240 -40760 1 PIX737_IN
port 761 n
rlabel metal5 115040 -40960 115240 -40760 1 PIX738_IN
port 762 n
rlabel metal5 118040 -40960 118240 -40760 1 PIX739_IN
port 763 n
rlabel metal5 121040 -40960 121240 -40760 1 PIX740_IN
port 764 n
rlabel metal5 124040 -40960 124240 -40760 1 PIX741_IN
port 765 n
rlabel metal5 127040 -40960 127240 -40760 1 PIX742_IN
port 766 n
rlabel metal5 130040 -40960 130240 -40760 1 PIX743_IN
port 767 n
rlabel metal5 133040 -40960 133240 -40760 1 PIX744_IN
port 768 n
rlabel metal5 136040 -40960 136240 -40760 1 PIX745_IN
port 769 n
rlabel metal5 139040 -40960 139240 -40760 1 PIX746_IN
port 770 n
rlabel metal5 142040 -40960 142240 -40760 1 PIX747_IN
port 771 n
rlabel metal5 145040 -40960 145240 -40760 1 PIX748_IN
port 772 n
rlabel metal5 148040 -40960 148240 -40760 1 PIX749_IN
port 773 n
rlabel metal5 1040 -43960 1240 -43760 1 PIX750_IN
port 774 n
rlabel metal2 -3000 -43520 -3000 -43430 3 ROW_SEL15
port 775 e
rlabel metal5 4040 -43960 4240 -43760 1 PIX751_IN
port 776 n
rlabel metal5 7040 -43960 7240 -43760 1 PIX752_IN
port 777 n
rlabel metal5 10040 -43960 10240 -43760 1 PIX753_IN
port 778 n
rlabel metal5 13040 -43960 13240 -43760 1 PIX754_IN
port 779 n
rlabel metal5 16040 -43960 16240 -43760 1 PIX755_IN
port 780 n
rlabel metal5 19040 -43960 19240 -43760 1 PIX756_IN
port 781 n
rlabel metal5 22040 -43960 22240 -43760 1 PIX757_IN
port 782 n
rlabel metal5 25040 -43960 25240 -43760 1 PIX758_IN
port 783 n
rlabel metal5 28040 -43960 28240 -43760 1 PIX759_IN
port 784 n
rlabel metal5 31040 -43960 31240 -43760 1 PIX760_IN
port 785 n
rlabel metal5 34040 -43960 34240 -43760 1 PIX761_IN
port 786 n
rlabel metal5 37040 -43960 37240 -43760 1 PIX762_IN
port 787 n
rlabel metal5 40040 -43960 40240 -43760 1 PIX763_IN
port 788 n
rlabel metal5 43040 -43960 43240 -43760 1 PIX764_IN
port 789 n
rlabel metal5 46040 -43960 46240 -43760 1 PIX765_IN
port 790 n
rlabel metal5 49040 -43960 49240 -43760 1 PIX766_IN
port 791 n
rlabel metal5 52040 -43960 52240 -43760 1 PIX767_IN
port 792 n
rlabel metal5 55040 -43960 55240 -43760 1 PIX768_IN
port 793 n
rlabel metal5 58040 -43960 58240 -43760 1 PIX769_IN
port 794 n
rlabel metal5 61040 -43960 61240 -43760 1 PIX770_IN
port 795 n
rlabel metal5 64040 -43960 64240 -43760 1 PIX771_IN
port 796 n
rlabel metal5 67040 -43960 67240 -43760 1 PIX772_IN
port 797 n
rlabel metal5 70040 -43960 70240 -43760 1 PIX773_IN
port 798 n
rlabel metal5 73040 -43960 73240 -43760 1 PIX774_IN
port 799 n
rlabel metal5 76040 -43960 76240 -43760 1 PIX775_IN
port 800 n
rlabel metal5 79040 -43960 79240 -43760 1 PIX776_IN
port 801 n
rlabel metal5 82040 -43960 82240 -43760 1 PIX777_IN
port 802 n
rlabel metal5 85040 -43960 85240 -43760 1 PIX778_IN
port 803 n
rlabel metal5 88040 -43960 88240 -43760 1 PIX779_IN
port 804 n
rlabel metal5 91040 -43960 91240 -43760 1 PIX780_IN
port 805 n
rlabel metal5 94040 -43960 94240 -43760 1 PIX781_IN
port 806 n
rlabel metal5 97040 -43960 97240 -43760 1 PIX782_IN
port 807 n
rlabel metal5 100040 -43960 100240 -43760 1 PIX783_IN
port 808 n
rlabel metal5 103040 -43960 103240 -43760 1 PIX784_IN
port 809 n
rlabel metal5 106040 -43960 106240 -43760 1 PIX785_IN
port 810 n
rlabel metal5 109040 -43960 109240 -43760 1 PIX786_IN
port 811 n
rlabel metal5 112040 -43960 112240 -43760 1 PIX787_IN
port 812 n
rlabel metal5 115040 -43960 115240 -43760 1 PIX788_IN
port 813 n
rlabel metal5 118040 -43960 118240 -43760 1 PIX789_IN
port 814 n
rlabel metal5 121040 -43960 121240 -43760 1 PIX790_IN
port 815 n
rlabel metal5 124040 -43960 124240 -43760 1 PIX791_IN
port 816 n
rlabel metal5 127040 -43960 127240 -43760 1 PIX792_IN
port 817 n
rlabel metal5 130040 -43960 130240 -43760 1 PIX793_IN
port 818 n
rlabel metal5 133040 -43960 133240 -43760 1 PIX794_IN
port 819 n
rlabel metal5 136040 -43960 136240 -43760 1 PIX795_IN
port 820 n
rlabel metal5 139040 -43960 139240 -43760 1 PIX796_IN
port 821 n
rlabel metal5 142040 -43960 142240 -43760 1 PIX797_IN
port 822 n
rlabel metal5 145040 -43960 145240 -43760 1 PIX798_IN
port 823 n
rlabel metal5 148040 -43960 148240 -43760 1 PIX799_IN
port 824 n
rlabel metal5 1040 -46960 1240 -46760 1 PIX800_IN
port 825 n
rlabel metal2 -3000 -46520 -3000 -46430 3 ROW_SEL16
port 826 e
rlabel metal5 4040 -46960 4240 -46760 1 PIX801_IN
port 827 n
rlabel metal5 7040 -46960 7240 -46760 1 PIX802_IN
port 828 n
rlabel metal5 10040 -46960 10240 -46760 1 PIX803_IN
port 829 n
rlabel metal5 13040 -46960 13240 -46760 1 PIX804_IN
port 830 n
rlabel metal5 16040 -46960 16240 -46760 1 PIX805_IN
port 831 n
rlabel metal5 19040 -46960 19240 -46760 1 PIX806_IN
port 832 n
rlabel metal5 22040 -46960 22240 -46760 1 PIX807_IN
port 833 n
rlabel metal5 25040 -46960 25240 -46760 1 PIX808_IN
port 834 n
rlabel metal5 28040 -46960 28240 -46760 1 PIX809_IN
port 835 n
rlabel metal5 31040 -46960 31240 -46760 1 PIX810_IN
port 836 n
rlabel metal5 34040 -46960 34240 -46760 1 PIX811_IN
port 837 n
rlabel metal5 37040 -46960 37240 -46760 1 PIX812_IN
port 838 n
rlabel metal5 40040 -46960 40240 -46760 1 PIX813_IN
port 839 n
rlabel metal5 43040 -46960 43240 -46760 1 PIX814_IN
port 840 n
rlabel metal5 46040 -46960 46240 -46760 1 PIX815_IN
port 841 n
rlabel metal5 49040 -46960 49240 -46760 1 PIX816_IN
port 842 n
rlabel metal5 52040 -46960 52240 -46760 1 PIX817_IN
port 843 n
rlabel metal5 55040 -46960 55240 -46760 1 PIX818_IN
port 844 n
rlabel metal5 58040 -46960 58240 -46760 1 PIX819_IN
port 845 n
rlabel metal5 61040 -46960 61240 -46760 1 PIX820_IN
port 846 n
rlabel metal5 64040 -46960 64240 -46760 1 PIX821_IN
port 847 n
rlabel metal5 67040 -46960 67240 -46760 1 PIX822_IN
port 848 n
rlabel metal5 70040 -46960 70240 -46760 1 PIX823_IN
port 849 n
rlabel metal5 73040 -46960 73240 -46760 1 PIX824_IN
port 850 n
rlabel metal5 76040 -46960 76240 -46760 1 PIX825_IN
port 851 n
rlabel metal5 79040 -46960 79240 -46760 1 PIX826_IN
port 852 n
rlabel metal5 82040 -46960 82240 -46760 1 PIX827_IN
port 853 n
rlabel metal5 85040 -46960 85240 -46760 1 PIX828_IN
port 854 n
rlabel metal5 88040 -46960 88240 -46760 1 PIX829_IN
port 855 n
rlabel metal5 91040 -46960 91240 -46760 1 PIX830_IN
port 856 n
rlabel metal5 94040 -46960 94240 -46760 1 PIX831_IN
port 857 n
rlabel metal5 97040 -46960 97240 -46760 1 PIX832_IN
port 858 n
rlabel metal5 100040 -46960 100240 -46760 1 PIX833_IN
port 859 n
rlabel metal5 103040 -46960 103240 -46760 1 PIX834_IN
port 860 n
rlabel metal5 106040 -46960 106240 -46760 1 PIX835_IN
port 861 n
rlabel metal5 109040 -46960 109240 -46760 1 PIX836_IN
port 862 n
rlabel metal5 112040 -46960 112240 -46760 1 PIX837_IN
port 863 n
rlabel metal5 115040 -46960 115240 -46760 1 PIX838_IN
port 864 n
rlabel metal5 118040 -46960 118240 -46760 1 PIX839_IN
port 865 n
rlabel metal5 121040 -46960 121240 -46760 1 PIX840_IN
port 866 n
rlabel metal5 124040 -46960 124240 -46760 1 PIX841_IN
port 867 n
rlabel metal5 127040 -46960 127240 -46760 1 PIX842_IN
port 868 n
rlabel metal5 130040 -46960 130240 -46760 1 PIX843_IN
port 869 n
rlabel metal5 133040 -46960 133240 -46760 1 PIX844_IN
port 870 n
rlabel metal5 136040 -46960 136240 -46760 1 PIX845_IN
port 871 n
rlabel metal5 139040 -46960 139240 -46760 1 PIX846_IN
port 872 n
rlabel metal5 142040 -46960 142240 -46760 1 PIX847_IN
port 873 n
rlabel metal5 145040 -46960 145240 -46760 1 PIX848_IN
port 874 n
rlabel metal5 148040 -46960 148240 -46760 1 PIX849_IN
port 875 n
rlabel metal5 1040 -49960 1240 -49760 1 PIX850_IN
port 876 n
rlabel metal2 -3000 -49520 -3000 -49430 3 ROW_SEL17
port 877 e
rlabel metal5 4040 -49960 4240 -49760 1 PIX851_IN
port 878 n
rlabel metal5 7040 -49960 7240 -49760 1 PIX852_IN
port 879 n
rlabel metal5 10040 -49960 10240 -49760 1 PIX853_IN
port 880 n
rlabel metal5 13040 -49960 13240 -49760 1 PIX854_IN
port 881 n
rlabel metal5 16040 -49960 16240 -49760 1 PIX855_IN
port 882 n
rlabel metal5 19040 -49960 19240 -49760 1 PIX856_IN
port 883 n
rlabel metal5 22040 -49960 22240 -49760 1 PIX857_IN
port 884 n
rlabel metal5 25040 -49960 25240 -49760 1 PIX858_IN
port 885 n
rlabel metal5 28040 -49960 28240 -49760 1 PIX859_IN
port 886 n
rlabel metal5 31040 -49960 31240 -49760 1 PIX860_IN
port 887 n
rlabel metal5 34040 -49960 34240 -49760 1 PIX861_IN
port 888 n
rlabel metal5 37040 -49960 37240 -49760 1 PIX862_IN
port 889 n
rlabel metal5 40040 -49960 40240 -49760 1 PIX863_IN
port 890 n
rlabel metal5 43040 -49960 43240 -49760 1 PIX864_IN
port 891 n
rlabel metal5 46040 -49960 46240 -49760 1 PIX865_IN
port 892 n
rlabel metal5 49040 -49960 49240 -49760 1 PIX866_IN
port 893 n
rlabel metal5 52040 -49960 52240 -49760 1 PIX867_IN
port 894 n
rlabel metal5 55040 -49960 55240 -49760 1 PIX868_IN
port 895 n
rlabel metal5 58040 -49960 58240 -49760 1 PIX869_IN
port 896 n
rlabel metal5 61040 -49960 61240 -49760 1 PIX870_IN
port 897 n
rlabel metal5 64040 -49960 64240 -49760 1 PIX871_IN
port 898 n
rlabel metal5 67040 -49960 67240 -49760 1 PIX872_IN
port 899 n
rlabel metal5 70040 -49960 70240 -49760 1 PIX873_IN
port 900 n
rlabel metal5 73040 -49960 73240 -49760 1 PIX874_IN
port 901 n
rlabel metal5 76040 -49960 76240 -49760 1 PIX875_IN
port 902 n
rlabel metal5 79040 -49960 79240 -49760 1 PIX876_IN
port 903 n
rlabel metal5 82040 -49960 82240 -49760 1 PIX877_IN
port 904 n
rlabel metal5 85040 -49960 85240 -49760 1 PIX878_IN
port 905 n
rlabel metal5 88040 -49960 88240 -49760 1 PIX879_IN
port 906 n
rlabel metal5 91040 -49960 91240 -49760 1 PIX880_IN
port 907 n
rlabel metal5 94040 -49960 94240 -49760 1 PIX881_IN
port 908 n
rlabel metal5 97040 -49960 97240 -49760 1 PIX882_IN
port 909 n
rlabel metal5 100040 -49960 100240 -49760 1 PIX883_IN
port 910 n
rlabel metal5 103040 -49960 103240 -49760 1 PIX884_IN
port 911 n
rlabel metal5 106040 -49960 106240 -49760 1 PIX885_IN
port 912 n
rlabel metal5 109040 -49960 109240 -49760 1 PIX886_IN
port 913 n
rlabel metal5 112040 -49960 112240 -49760 1 PIX887_IN
port 914 n
rlabel metal5 115040 -49960 115240 -49760 1 PIX888_IN
port 915 n
rlabel metal5 118040 -49960 118240 -49760 1 PIX889_IN
port 916 n
rlabel metal5 121040 -49960 121240 -49760 1 PIX890_IN
port 917 n
rlabel metal5 124040 -49960 124240 -49760 1 PIX891_IN
port 918 n
rlabel metal5 127040 -49960 127240 -49760 1 PIX892_IN
port 919 n
rlabel metal5 130040 -49960 130240 -49760 1 PIX893_IN
port 920 n
rlabel metal5 133040 -49960 133240 -49760 1 PIX894_IN
port 921 n
rlabel metal5 136040 -49960 136240 -49760 1 PIX895_IN
port 922 n
rlabel metal5 139040 -49960 139240 -49760 1 PIX896_IN
port 923 n
rlabel metal5 142040 -49960 142240 -49760 1 PIX897_IN
port 924 n
rlabel metal5 145040 -49960 145240 -49760 1 PIX898_IN
port 925 n
rlabel metal5 148040 -49960 148240 -49760 1 PIX899_IN
port 926 n
rlabel metal5 1040 -52960 1240 -52760 1 PIX900_IN
port 927 n
rlabel metal2 -3000 -52520 -3000 -52430 3 ROW_SEL18
port 928 e
rlabel metal5 4040 -52960 4240 -52760 1 PIX901_IN
port 929 n
rlabel metal5 7040 -52960 7240 -52760 1 PIX902_IN
port 930 n
rlabel metal5 10040 -52960 10240 -52760 1 PIX903_IN
port 931 n
rlabel metal5 13040 -52960 13240 -52760 1 PIX904_IN
port 932 n
rlabel metal5 16040 -52960 16240 -52760 1 PIX905_IN
port 933 n
rlabel metal5 19040 -52960 19240 -52760 1 PIX906_IN
port 934 n
rlabel metal5 22040 -52960 22240 -52760 1 PIX907_IN
port 935 n
rlabel metal5 25040 -52960 25240 -52760 1 PIX908_IN
port 936 n
rlabel metal5 28040 -52960 28240 -52760 1 PIX909_IN
port 937 n
rlabel metal5 31040 -52960 31240 -52760 1 PIX910_IN
port 938 n
rlabel metal5 34040 -52960 34240 -52760 1 PIX911_IN
port 939 n
rlabel metal5 37040 -52960 37240 -52760 1 PIX912_IN
port 940 n
rlabel metal5 40040 -52960 40240 -52760 1 PIX913_IN
port 941 n
rlabel metal5 43040 -52960 43240 -52760 1 PIX914_IN
port 942 n
rlabel metal5 46040 -52960 46240 -52760 1 PIX915_IN
port 943 n
rlabel metal5 49040 -52960 49240 -52760 1 PIX916_IN
port 944 n
rlabel metal5 52040 -52960 52240 -52760 1 PIX917_IN
port 945 n
rlabel metal5 55040 -52960 55240 -52760 1 PIX918_IN
port 946 n
rlabel metal5 58040 -52960 58240 -52760 1 PIX919_IN
port 947 n
rlabel metal5 61040 -52960 61240 -52760 1 PIX920_IN
port 948 n
rlabel metal5 64040 -52960 64240 -52760 1 PIX921_IN
port 949 n
rlabel metal5 67040 -52960 67240 -52760 1 PIX922_IN
port 950 n
rlabel metal5 70040 -52960 70240 -52760 1 PIX923_IN
port 951 n
rlabel metal5 73040 -52960 73240 -52760 1 PIX924_IN
port 952 n
rlabel metal5 76040 -52960 76240 -52760 1 PIX925_IN
port 953 n
rlabel metal5 79040 -52960 79240 -52760 1 PIX926_IN
port 954 n
rlabel metal5 82040 -52960 82240 -52760 1 PIX927_IN
port 955 n
rlabel metal5 85040 -52960 85240 -52760 1 PIX928_IN
port 956 n
rlabel metal5 88040 -52960 88240 -52760 1 PIX929_IN
port 957 n
rlabel metal5 91040 -52960 91240 -52760 1 PIX930_IN
port 958 n
rlabel metal5 94040 -52960 94240 -52760 1 PIX931_IN
port 959 n
rlabel metal5 97040 -52960 97240 -52760 1 PIX932_IN
port 960 n
rlabel metal5 100040 -52960 100240 -52760 1 PIX933_IN
port 961 n
rlabel metal5 103040 -52960 103240 -52760 1 PIX934_IN
port 962 n
rlabel metal5 106040 -52960 106240 -52760 1 PIX935_IN
port 963 n
rlabel metal5 109040 -52960 109240 -52760 1 PIX936_IN
port 964 n
rlabel metal5 112040 -52960 112240 -52760 1 PIX937_IN
port 965 n
rlabel metal5 115040 -52960 115240 -52760 1 PIX938_IN
port 966 n
rlabel metal5 118040 -52960 118240 -52760 1 PIX939_IN
port 967 n
rlabel metal5 121040 -52960 121240 -52760 1 PIX940_IN
port 968 n
rlabel metal5 124040 -52960 124240 -52760 1 PIX941_IN
port 969 n
rlabel metal5 127040 -52960 127240 -52760 1 PIX942_IN
port 970 n
rlabel metal5 130040 -52960 130240 -52760 1 PIX943_IN
port 971 n
rlabel metal5 133040 -52960 133240 -52760 1 PIX944_IN
port 972 n
rlabel metal5 136040 -52960 136240 -52760 1 PIX945_IN
port 973 n
rlabel metal5 139040 -52960 139240 -52760 1 PIX946_IN
port 974 n
rlabel metal5 142040 -52960 142240 -52760 1 PIX947_IN
port 975 n
rlabel metal5 145040 -52960 145240 -52760 1 PIX948_IN
port 976 n
rlabel metal5 148040 -52960 148240 -52760 1 PIX949_IN
port 977 n
rlabel metal5 1040 -55960 1240 -55760 1 PIX950_IN
port 978 n
rlabel metal2 -3000 -55520 -3000 -55430 3 ROW_SEL19
port 979 e
rlabel metal5 4040 -55960 4240 -55760 1 PIX951_IN
port 980 n
rlabel metal5 7040 -55960 7240 -55760 1 PIX952_IN
port 981 n
rlabel metal5 10040 -55960 10240 -55760 1 PIX953_IN
port 982 n
rlabel metal5 13040 -55960 13240 -55760 1 PIX954_IN
port 983 n
rlabel metal5 16040 -55960 16240 -55760 1 PIX955_IN
port 984 n
rlabel metal5 19040 -55960 19240 -55760 1 PIX956_IN
port 985 n
rlabel metal5 22040 -55960 22240 -55760 1 PIX957_IN
port 986 n
rlabel metal5 25040 -55960 25240 -55760 1 PIX958_IN
port 987 n
rlabel metal5 28040 -55960 28240 -55760 1 PIX959_IN
port 988 n
rlabel metal5 31040 -55960 31240 -55760 1 PIX960_IN
port 989 n
rlabel metal5 34040 -55960 34240 -55760 1 PIX961_IN
port 990 n
rlabel metal5 37040 -55960 37240 -55760 1 PIX962_IN
port 991 n
rlabel metal5 40040 -55960 40240 -55760 1 PIX963_IN
port 992 n
rlabel metal5 43040 -55960 43240 -55760 1 PIX964_IN
port 993 n
rlabel metal5 46040 -55960 46240 -55760 1 PIX965_IN
port 994 n
rlabel metal5 49040 -55960 49240 -55760 1 PIX966_IN
port 995 n
rlabel metal5 52040 -55960 52240 -55760 1 PIX967_IN
port 996 n
rlabel metal5 55040 -55960 55240 -55760 1 PIX968_IN
port 997 n
rlabel metal5 58040 -55960 58240 -55760 1 PIX969_IN
port 998 n
rlabel metal5 61040 -55960 61240 -55760 1 PIX970_IN
port 999 n
rlabel metal5 64040 -55960 64240 -55760 1 PIX971_IN
port 1000 n
rlabel metal5 67040 -55960 67240 -55760 1 PIX972_IN
port 1001 n
rlabel metal5 70040 -55960 70240 -55760 1 PIX973_IN
port 1002 n
rlabel metal5 73040 -55960 73240 -55760 1 PIX974_IN
port 1003 n
rlabel metal5 76040 -55960 76240 -55760 1 PIX975_IN
port 1004 n
rlabel metal5 79040 -55960 79240 -55760 1 PIX976_IN
port 1005 n
rlabel metal5 82040 -55960 82240 -55760 1 PIX977_IN
port 1006 n
rlabel metal5 85040 -55960 85240 -55760 1 PIX978_IN
port 1007 n
rlabel metal5 88040 -55960 88240 -55760 1 PIX979_IN
port 1008 n
rlabel metal5 91040 -55960 91240 -55760 1 PIX980_IN
port 1009 n
rlabel metal5 94040 -55960 94240 -55760 1 PIX981_IN
port 1010 n
rlabel metal5 97040 -55960 97240 -55760 1 PIX982_IN
port 1011 n
rlabel metal5 100040 -55960 100240 -55760 1 PIX983_IN
port 1012 n
rlabel metal5 103040 -55960 103240 -55760 1 PIX984_IN
port 1013 n
rlabel metal5 106040 -55960 106240 -55760 1 PIX985_IN
port 1014 n
rlabel metal5 109040 -55960 109240 -55760 1 PIX986_IN
port 1015 n
rlabel metal5 112040 -55960 112240 -55760 1 PIX987_IN
port 1016 n
rlabel metal5 115040 -55960 115240 -55760 1 PIX988_IN
port 1017 n
rlabel metal5 118040 -55960 118240 -55760 1 PIX989_IN
port 1018 n
rlabel metal5 121040 -55960 121240 -55760 1 PIX990_IN
port 1019 n
rlabel metal5 124040 -55960 124240 -55760 1 PIX991_IN
port 1020 n
rlabel metal5 127040 -55960 127240 -55760 1 PIX992_IN
port 1021 n
rlabel metal5 130040 -55960 130240 -55760 1 PIX993_IN
port 1022 n
rlabel metal5 133040 -55960 133240 -55760 1 PIX994_IN
port 1023 n
rlabel metal5 136040 -55960 136240 -55760 1 PIX995_IN
port 1024 n
rlabel metal5 139040 -55960 139240 -55760 1 PIX996_IN
port 1025 n
rlabel metal5 142040 -55960 142240 -55760 1 PIX997_IN
port 1026 n
rlabel metal5 145040 -55960 145240 -55760 1 PIX998_IN
port 1027 n
rlabel metal5 148040 -55960 148240 -55760 1 PIX999_IN
port 1028 n
rlabel metal5 1040 -58960 1240 -58760 1 PIX1000_IN
port 1029 n
rlabel metal2 -3000 -58520 -3000 -58430 3 ROW_SEL20
port 1030 e
rlabel metal5 4040 -58960 4240 -58760 1 PIX1001_IN
port 1031 n
rlabel metal5 7040 -58960 7240 -58760 1 PIX1002_IN
port 1032 n
rlabel metal5 10040 -58960 10240 -58760 1 PIX1003_IN
port 1033 n
rlabel metal5 13040 -58960 13240 -58760 1 PIX1004_IN
port 1034 n
rlabel metal5 16040 -58960 16240 -58760 1 PIX1005_IN
port 1035 n
rlabel metal5 19040 -58960 19240 -58760 1 PIX1006_IN
port 1036 n
rlabel metal5 22040 -58960 22240 -58760 1 PIX1007_IN
port 1037 n
rlabel metal5 25040 -58960 25240 -58760 1 PIX1008_IN
port 1038 n
rlabel metal5 28040 -58960 28240 -58760 1 PIX1009_IN
port 1039 n
rlabel metal5 31040 -58960 31240 -58760 1 PIX1010_IN
port 1040 n
rlabel metal5 34040 -58960 34240 -58760 1 PIX1011_IN
port 1041 n
rlabel metal5 37040 -58960 37240 -58760 1 PIX1012_IN
port 1042 n
rlabel metal5 40040 -58960 40240 -58760 1 PIX1013_IN
port 1043 n
rlabel metal5 43040 -58960 43240 -58760 1 PIX1014_IN
port 1044 n
rlabel metal5 46040 -58960 46240 -58760 1 PIX1015_IN
port 1045 n
rlabel metal5 49040 -58960 49240 -58760 1 PIX1016_IN
port 1046 n
rlabel metal5 52040 -58960 52240 -58760 1 PIX1017_IN
port 1047 n
rlabel metal5 55040 -58960 55240 -58760 1 PIX1018_IN
port 1048 n
rlabel metal5 58040 -58960 58240 -58760 1 PIX1019_IN
port 1049 n
rlabel metal5 61040 -58960 61240 -58760 1 PIX1020_IN
port 1050 n
rlabel metal5 64040 -58960 64240 -58760 1 PIX1021_IN
port 1051 n
rlabel metal5 67040 -58960 67240 -58760 1 PIX1022_IN
port 1052 n
rlabel metal5 70040 -58960 70240 -58760 1 PIX1023_IN
port 1053 n
rlabel metal5 73040 -58960 73240 -58760 1 PIX1024_IN
port 1054 n
rlabel metal5 76040 -58960 76240 -58760 1 PIX1025_IN
port 1055 n
rlabel metal5 79040 -58960 79240 -58760 1 PIX1026_IN
port 1056 n
rlabel metal5 82040 -58960 82240 -58760 1 PIX1027_IN
port 1057 n
rlabel metal5 85040 -58960 85240 -58760 1 PIX1028_IN
port 1058 n
rlabel metal5 88040 -58960 88240 -58760 1 PIX1029_IN
port 1059 n
rlabel metal5 91040 -58960 91240 -58760 1 PIX1030_IN
port 1060 n
rlabel metal5 94040 -58960 94240 -58760 1 PIX1031_IN
port 1061 n
rlabel metal5 97040 -58960 97240 -58760 1 PIX1032_IN
port 1062 n
rlabel metal5 100040 -58960 100240 -58760 1 PIX1033_IN
port 1063 n
rlabel metal5 103040 -58960 103240 -58760 1 PIX1034_IN
port 1064 n
rlabel metal5 106040 -58960 106240 -58760 1 PIX1035_IN
port 1065 n
rlabel metal5 109040 -58960 109240 -58760 1 PIX1036_IN
port 1066 n
rlabel metal5 112040 -58960 112240 -58760 1 PIX1037_IN
port 1067 n
rlabel metal5 115040 -58960 115240 -58760 1 PIX1038_IN
port 1068 n
rlabel metal5 118040 -58960 118240 -58760 1 PIX1039_IN
port 1069 n
rlabel metal5 121040 -58960 121240 -58760 1 PIX1040_IN
port 1070 n
rlabel metal5 124040 -58960 124240 -58760 1 PIX1041_IN
port 1071 n
rlabel metal5 127040 -58960 127240 -58760 1 PIX1042_IN
port 1072 n
rlabel metal5 130040 -58960 130240 -58760 1 PIX1043_IN
port 1073 n
rlabel metal5 133040 -58960 133240 -58760 1 PIX1044_IN
port 1074 n
rlabel metal5 136040 -58960 136240 -58760 1 PIX1045_IN
port 1075 n
rlabel metal5 139040 -58960 139240 -58760 1 PIX1046_IN
port 1076 n
rlabel metal5 142040 -58960 142240 -58760 1 PIX1047_IN
port 1077 n
rlabel metal5 145040 -58960 145240 -58760 1 PIX1048_IN
port 1078 n
rlabel metal5 148040 -58960 148240 -58760 1 PIX1049_IN
port 1079 n
rlabel metal5 1040 -61960 1240 -61760 1 PIX1050_IN
port 1080 n
rlabel metal2 -3000 -61520 -3000 -61430 3 ROW_SEL21
port 1081 e
rlabel metal5 4040 -61960 4240 -61760 1 PIX1051_IN
port 1082 n
rlabel metal5 7040 -61960 7240 -61760 1 PIX1052_IN
port 1083 n
rlabel metal5 10040 -61960 10240 -61760 1 PIX1053_IN
port 1084 n
rlabel metal5 13040 -61960 13240 -61760 1 PIX1054_IN
port 1085 n
rlabel metal5 16040 -61960 16240 -61760 1 PIX1055_IN
port 1086 n
rlabel metal5 19040 -61960 19240 -61760 1 PIX1056_IN
port 1087 n
rlabel metal5 22040 -61960 22240 -61760 1 PIX1057_IN
port 1088 n
rlabel metal5 25040 -61960 25240 -61760 1 PIX1058_IN
port 1089 n
rlabel metal5 28040 -61960 28240 -61760 1 PIX1059_IN
port 1090 n
rlabel metal5 31040 -61960 31240 -61760 1 PIX1060_IN
port 1091 n
rlabel metal5 34040 -61960 34240 -61760 1 PIX1061_IN
port 1092 n
rlabel metal5 37040 -61960 37240 -61760 1 PIX1062_IN
port 1093 n
rlabel metal5 40040 -61960 40240 -61760 1 PIX1063_IN
port 1094 n
rlabel metal5 43040 -61960 43240 -61760 1 PIX1064_IN
port 1095 n
rlabel metal5 46040 -61960 46240 -61760 1 PIX1065_IN
port 1096 n
rlabel metal5 49040 -61960 49240 -61760 1 PIX1066_IN
port 1097 n
rlabel metal5 52040 -61960 52240 -61760 1 PIX1067_IN
port 1098 n
rlabel metal5 55040 -61960 55240 -61760 1 PIX1068_IN
port 1099 n
rlabel metal5 58040 -61960 58240 -61760 1 PIX1069_IN
port 1100 n
rlabel metal5 61040 -61960 61240 -61760 1 PIX1070_IN
port 1101 n
rlabel metal5 64040 -61960 64240 -61760 1 PIX1071_IN
port 1102 n
rlabel metal5 67040 -61960 67240 -61760 1 PIX1072_IN
port 1103 n
rlabel metal5 70040 -61960 70240 -61760 1 PIX1073_IN
port 1104 n
rlabel metal5 73040 -61960 73240 -61760 1 PIX1074_IN
port 1105 n
rlabel metal5 76040 -61960 76240 -61760 1 PIX1075_IN
port 1106 n
rlabel metal5 79040 -61960 79240 -61760 1 PIX1076_IN
port 1107 n
rlabel metal5 82040 -61960 82240 -61760 1 PIX1077_IN
port 1108 n
rlabel metal5 85040 -61960 85240 -61760 1 PIX1078_IN
port 1109 n
rlabel metal5 88040 -61960 88240 -61760 1 PIX1079_IN
port 1110 n
rlabel metal5 91040 -61960 91240 -61760 1 PIX1080_IN
port 1111 n
rlabel metal5 94040 -61960 94240 -61760 1 PIX1081_IN
port 1112 n
rlabel metal5 97040 -61960 97240 -61760 1 PIX1082_IN
port 1113 n
rlabel metal5 100040 -61960 100240 -61760 1 PIX1083_IN
port 1114 n
rlabel metal5 103040 -61960 103240 -61760 1 PIX1084_IN
port 1115 n
rlabel metal5 106040 -61960 106240 -61760 1 PIX1085_IN
port 1116 n
rlabel metal5 109040 -61960 109240 -61760 1 PIX1086_IN
port 1117 n
rlabel metal5 112040 -61960 112240 -61760 1 PIX1087_IN
port 1118 n
rlabel metal5 115040 -61960 115240 -61760 1 PIX1088_IN
port 1119 n
rlabel metal5 118040 -61960 118240 -61760 1 PIX1089_IN
port 1120 n
rlabel metal5 121040 -61960 121240 -61760 1 PIX1090_IN
port 1121 n
rlabel metal5 124040 -61960 124240 -61760 1 PIX1091_IN
port 1122 n
rlabel metal5 127040 -61960 127240 -61760 1 PIX1092_IN
port 1123 n
rlabel metal5 130040 -61960 130240 -61760 1 PIX1093_IN
port 1124 n
rlabel metal5 133040 -61960 133240 -61760 1 PIX1094_IN
port 1125 n
rlabel metal5 136040 -61960 136240 -61760 1 PIX1095_IN
port 1126 n
rlabel metal5 139040 -61960 139240 -61760 1 PIX1096_IN
port 1127 n
rlabel metal5 142040 -61960 142240 -61760 1 PIX1097_IN
port 1128 n
rlabel metal5 145040 -61960 145240 -61760 1 PIX1098_IN
port 1129 n
rlabel metal5 148040 -61960 148240 -61760 1 PIX1099_IN
port 1130 n
rlabel metal5 1040 -64960 1240 -64760 1 PIX1100_IN
port 1131 n
rlabel metal2 -3000 -64520 -3000 -64430 3 ROW_SEL22
port 1132 e
rlabel metal5 4040 -64960 4240 -64760 1 PIX1101_IN
port 1133 n
rlabel metal5 7040 -64960 7240 -64760 1 PIX1102_IN
port 1134 n
rlabel metal5 10040 -64960 10240 -64760 1 PIX1103_IN
port 1135 n
rlabel metal5 13040 -64960 13240 -64760 1 PIX1104_IN
port 1136 n
rlabel metal5 16040 -64960 16240 -64760 1 PIX1105_IN
port 1137 n
rlabel metal5 19040 -64960 19240 -64760 1 PIX1106_IN
port 1138 n
rlabel metal5 22040 -64960 22240 -64760 1 PIX1107_IN
port 1139 n
rlabel metal5 25040 -64960 25240 -64760 1 PIX1108_IN
port 1140 n
rlabel metal5 28040 -64960 28240 -64760 1 PIX1109_IN
port 1141 n
rlabel metal5 31040 -64960 31240 -64760 1 PIX1110_IN
port 1142 n
rlabel metal5 34040 -64960 34240 -64760 1 PIX1111_IN
port 1143 n
rlabel metal5 37040 -64960 37240 -64760 1 PIX1112_IN
port 1144 n
rlabel metal5 40040 -64960 40240 -64760 1 PIX1113_IN
port 1145 n
rlabel metal5 43040 -64960 43240 -64760 1 PIX1114_IN
port 1146 n
rlabel metal5 46040 -64960 46240 -64760 1 PIX1115_IN
port 1147 n
rlabel metal5 49040 -64960 49240 -64760 1 PIX1116_IN
port 1148 n
rlabel metal5 52040 -64960 52240 -64760 1 PIX1117_IN
port 1149 n
rlabel metal5 55040 -64960 55240 -64760 1 PIX1118_IN
port 1150 n
rlabel metal5 58040 -64960 58240 -64760 1 PIX1119_IN
port 1151 n
rlabel metal5 61040 -64960 61240 -64760 1 PIX1120_IN
port 1152 n
rlabel metal5 64040 -64960 64240 -64760 1 PIX1121_IN
port 1153 n
rlabel metal5 67040 -64960 67240 -64760 1 PIX1122_IN
port 1154 n
rlabel metal5 70040 -64960 70240 -64760 1 PIX1123_IN
port 1155 n
rlabel metal5 73040 -64960 73240 -64760 1 PIX1124_IN
port 1156 n
rlabel metal5 76040 -64960 76240 -64760 1 PIX1125_IN
port 1157 n
rlabel metal5 79040 -64960 79240 -64760 1 PIX1126_IN
port 1158 n
rlabel metal5 82040 -64960 82240 -64760 1 PIX1127_IN
port 1159 n
rlabel metal5 85040 -64960 85240 -64760 1 PIX1128_IN
port 1160 n
rlabel metal5 88040 -64960 88240 -64760 1 PIX1129_IN
port 1161 n
rlabel metal5 91040 -64960 91240 -64760 1 PIX1130_IN
port 1162 n
rlabel metal5 94040 -64960 94240 -64760 1 PIX1131_IN
port 1163 n
rlabel metal5 97040 -64960 97240 -64760 1 PIX1132_IN
port 1164 n
rlabel metal5 100040 -64960 100240 -64760 1 PIX1133_IN
port 1165 n
rlabel metal5 103040 -64960 103240 -64760 1 PIX1134_IN
port 1166 n
rlabel metal5 106040 -64960 106240 -64760 1 PIX1135_IN
port 1167 n
rlabel metal5 109040 -64960 109240 -64760 1 PIX1136_IN
port 1168 n
rlabel metal5 112040 -64960 112240 -64760 1 PIX1137_IN
port 1169 n
rlabel metal5 115040 -64960 115240 -64760 1 PIX1138_IN
port 1170 n
rlabel metal5 118040 -64960 118240 -64760 1 PIX1139_IN
port 1171 n
rlabel metal5 121040 -64960 121240 -64760 1 PIX1140_IN
port 1172 n
rlabel metal5 124040 -64960 124240 -64760 1 PIX1141_IN
port 1173 n
rlabel metal5 127040 -64960 127240 -64760 1 PIX1142_IN
port 1174 n
rlabel metal5 130040 -64960 130240 -64760 1 PIX1143_IN
port 1175 n
rlabel metal5 133040 -64960 133240 -64760 1 PIX1144_IN
port 1176 n
rlabel metal5 136040 -64960 136240 -64760 1 PIX1145_IN
port 1177 n
rlabel metal5 139040 -64960 139240 -64760 1 PIX1146_IN
port 1178 n
rlabel metal5 142040 -64960 142240 -64760 1 PIX1147_IN
port 1179 n
rlabel metal5 145040 -64960 145240 -64760 1 PIX1148_IN
port 1180 n
rlabel metal5 148040 -64960 148240 -64760 1 PIX1149_IN
port 1181 n
rlabel metal5 1040 -67960 1240 -67760 1 PIX1150_IN
port 1182 n
rlabel metal2 -3000 -67520 -3000 -67430 3 ROW_SEL23
port 1183 e
rlabel metal5 4040 -67960 4240 -67760 1 PIX1151_IN
port 1184 n
rlabel metal5 7040 -67960 7240 -67760 1 PIX1152_IN
port 1185 n
rlabel metal5 10040 -67960 10240 -67760 1 PIX1153_IN
port 1186 n
rlabel metal5 13040 -67960 13240 -67760 1 PIX1154_IN
port 1187 n
rlabel metal5 16040 -67960 16240 -67760 1 PIX1155_IN
port 1188 n
rlabel metal5 19040 -67960 19240 -67760 1 PIX1156_IN
port 1189 n
rlabel metal5 22040 -67960 22240 -67760 1 PIX1157_IN
port 1190 n
rlabel metal5 25040 -67960 25240 -67760 1 PIX1158_IN
port 1191 n
rlabel metal5 28040 -67960 28240 -67760 1 PIX1159_IN
port 1192 n
rlabel metal5 31040 -67960 31240 -67760 1 PIX1160_IN
port 1193 n
rlabel metal5 34040 -67960 34240 -67760 1 PIX1161_IN
port 1194 n
rlabel metal5 37040 -67960 37240 -67760 1 PIX1162_IN
port 1195 n
rlabel metal5 40040 -67960 40240 -67760 1 PIX1163_IN
port 1196 n
rlabel metal5 43040 -67960 43240 -67760 1 PIX1164_IN
port 1197 n
rlabel metal5 46040 -67960 46240 -67760 1 PIX1165_IN
port 1198 n
rlabel metal5 49040 -67960 49240 -67760 1 PIX1166_IN
port 1199 n
rlabel metal5 52040 -67960 52240 -67760 1 PIX1167_IN
port 1200 n
rlabel metal5 55040 -67960 55240 -67760 1 PIX1168_IN
port 1201 n
rlabel metal5 58040 -67960 58240 -67760 1 PIX1169_IN
port 1202 n
rlabel metal5 61040 -67960 61240 -67760 1 PIX1170_IN
port 1203 n
rlabel metal5 64040 -67960 64240 -67760 1 PIX1171_IN
port 1204 n
rlabel metal5 67040 -67960 67240 -67760 1 PIX1172_IN
port 1205 n
rlabel metal5 70040 -67960 70240 -67760 1 PIX1173_IN
port 1206 n
rlabel metal5 73040 -67960 73240 -67760 1 PIX1174_IN
port 1207 n
rlabel metal5 76040 -67960 76240 -67760 1 PIX1175_IN
port 1208 n
rlabel metal5 79040 -67960 79240 -67760 1 PIX1176_IN
port 1209 n
rlabel metal5 82040 -67960 82240 -67760 1 PIX1177_IN
port 1210 n
rlabel metal5 85040 -67960 85240 -67760 1 PIX1178_IN
port 1211 n
rlabel metal5 88040 -67960 88240 -67760 1 PIX1179_IN
port 1212 n
rlabel metal5 91040 -67960 91240 -67760 1 PIX1180_IN
port 1213 n
rlabel metal5 94040 -67960 94240 -67760 1 PIX1181_IN
port 1214 n
rlabel metal5 97040 -67960 97240 -67760 1 PIX1182_IN
port 1215 n
rlabel metal5 100040 -67960 100240 -67760 1 PIX1183_IN
port 1216 n
rlabel metal5 103040 -67960 103240 -67760 1 PIX1184_IN
port 1217 n
rlabel metal5 106040 -67960 106240 -67760 1 PIX1185_IN
port 1218 n
rlabel metal5 109040 -67960 109240 -67760 1 PIX1186_IN
port 1219 n
rlabel metal5 112040 -67960 112240 -67760 1 PIX1187_IN
port 1220 n
rlabel metal5 115040 -67960 115240 -67760 1 PIX1188_IN
port 1221 n
rlabel metal5 118040 -67960 118240 -67760 1 PIX1189_IN
port 1222 n
rlabel metal5 121040 -67960 121240 -67760 1 PIX1190_IN
port 1223 n
rlabel metal5 124040 -67960 124240 -67760 1 PIX1191_IN
port 1224 n
rlabel metal5 127040 -67960 127240 -67760 1 PIX1192_IN
port 1225 n
rlabel metal5 130040 -67960 130240 -67760 1 PIX1193_IN
port 1226 n
rlabel metal5 133040 -67960 133240 -67760 1 PIX1194_IN
port 1227 n
rlabel metal5 136040 -67960 136240 -67760 1 PIX1195_IN
port 1228 n
rlabel metal5 139040 -67960 139240 -67760 1 PIX1196_IN
port 1229 n
rlabel metal5 142040 -67960 142240 -67760 1 PIX1197_IN
port 1230 n
rlabel metal5 145040 -67960 145240 -67760 1 PIX1198_IN
port 1231 n
rlabel metal5 148040 -67960 148240 -67760 1 PIX1199_IN
port 1232 n
rlabel metal5 1040 -70960 1240 -70760 1 PIX1200_IN
port 1233 n
rlabel metal2 -3000 -70520 -3000 -70430 3 ROW_SEL24
port 1234 e
rlabel metal5 4040 -70960 4240 -70760 1 PIX1201_IN
port 1235 n
rlabel metal5 7040 -70960 7240 -70760 1 PIX1202_IN
port 1236 n
rlabel metal5 10040 -70960 10240 -70760 1 PIX1203_IN
port 1237 n
rlabel metal5 13040 -70960 13240 -70760 1 PIX1204_IN
port 1238 n
rlabel metal5 16040 -70960 16240 -70760 1 PIX1205_IN
port 1239 n
rlabel metal5 19040 -70960 19240 -70760 1 PIX1206_IN
port 1240 n
rlabel metal5 22040 -70960 22240 -70760 1 PIX1207_IN
port 1241 n
rlabel metal5 25040 -70960 25240 -70760 1 PIX1208_IN
port 1242 n
rlabel metal5 28040 -70960 28240 -70760 1 PIX1209_IN
port 1243 n
rlabel metal5 31040 -70960 31240 -70760 1 PIX1210_IN
port 1244 n
rlabel metal5 34040 -70960 34240 -70760 1 PIX1211_IN
port 1245 n
rlabel metal5 37040 -70960 37240 -70760 1 PIX1212_IN
port 1246 n
rlabel metal5 40040 -70960 40240 -70760 1 PIX1213_IN
port 1247 n
rlabel metal5 43040 -70960 43240 -70760 1 PIX1214_IN
port 1248 n
rlabel metal5 46040 -70960 46240 -70760 1 PIX1215_IN
port 1249 n
rlabel metal5 49040 -70960 49240 -70760 1 PIX1216_IN
port 1250 n
rlabel metal5 52040 -70960 52240 -70760 1 PIX1217_IN
port 1251 n
rlabel metal5 55040 -70960 55240 -70760 1 PIX1218_IN
port 1252 n
rlabel metal5 58040 -70960 58240 -70760 1 PIX1219_IN
port 1253 n
rlabel metal5 61040 -70960 61240 -70760 1 PIX1220_IN
port 1254 n
rlabel metal5 64040 -70960 64240 -70760 1 PIX1221_IN
port 1255 n
rlabel metal5 67040 -70960 67240 -70760 1 PIX1222_IN
port 1256 n
rlabel metal5 70040 -70960 70240 -70760 1 PIX1223_IN
port 1257 n
rlabel metal5 73040 -70960 73240 -70760 1 PIX1224_IN
port 1258 n
rlabel metal5 76040 -70960 76240 -70760 1 PIX1225_IN
port 1259 n
rlabel metal5 79040 -70960 79240 -70760 1 PIX1226_IN
port 1260 n
rlabel metal5 82040 -70960 82240 -70760 1 PIX1227_IN
port 1261 n
rlabel metal5 85040 -70960 85240 -70760 1 PIX1228_IN
port 1262 n
rlabel metal5 88040 -70960 88240 -70760 1 PIX1229_IN
port 1263 n
rlabel metal5 91040 -70960 91240 -70760 1 PIX1230_IN
port 1264 n
rlabel metal5 94040 -70960 94240 -70760 1 PIX1231_IN
port 1265 n
rlabel metal5 97040 -70960 97240 -70760 1 PIX1232_IN
port 1266 n
rlabel metal5 100040 -70960 100240 -70760 1 PIX1233_IN
port 1267 n
rlabel metal5 103040 -70960 103240 -70760 1 PIX1234_IN
port 1268 n
rlabel metal5 106040 -70960 106240 -70760 1 PIX1235_IN
port 1269 n
rlabel metal5 109040 -70960 109240 -70760 1 PIX1236_IN
port 1270 n
rlabel metal5 112040 -70960 112240 -70760 1 PIX1237_IN
port 1271 n
rlabel metal5 115040 -70960 115240 -70760 1 PIX1238_IN
port 1272 n
rlabel metal5 118040 -70960 118240 -70760 1 PIX1239_IN
port 1273 n
rlabel metal5 121040 -70960 121240 -70760 1 PIX1240_IN
port 1274 n
rlabel metal5 124040 -70960 124240 -70760 1 PIX1241_IN
port 1275 n
rlabel metal5 127040 -70960 127240 -70760 1 PIX1242_IN
port 1276 n
rlabel metal5 130040 -70960 130240 -70760 1 PIX1243_IN
port 1277 n
rlabel metal5 133040 -70960 133240 -70760 1 PIX1244_IN
port 1278 n
rlabel metal5 136040 -70960 136240 -70760 1 PIX1245_IN
port 1279 n
rlabel metal5 139040 -70960 139240 -70760 1 PIX1246_IN
port 1280 n
rlabel metal5 142040 -70960 142240 -70760 1 PIX1247_IN
port 1281 n
rlabel metal5 145040 -70960 145240 -70760 1 PIX1248_IN
port 1282 n
rlabel metal5 148040 -70960 148240 -70760 1 PIX1249_IN
port 1283 n
rlabel metal5 1040 -73960 1240 -73760 1 PIX1250_IN
port 1284 n
rlabel metal2 -3000 -73520 -3000 -73430 3 ROW_SEL25
port 1285 e
rlabel metal5 4040 -73960 4240 -73760 1 PIX1251_IN
port 1286 n
rlabel metal5 7040 -73960 7240 -73760 1 PIX1252_IN
port 1287 n
rlabel metal5 10040 -73960 10240 -73760 1 PIX1253_IN
port 1288 n
rlabel metal5 13040 -73960 13240 -73760 1 PIX1254_IN
port 1289 n
rlabel metal5 16040 -73960 16240 -73760 1 PIX1255_IN
port 1290 n
rlabel metal5 19040 -73960 19240 -73760 1 PIX1256_IN
port 1291 n
rlabel metal5 22040 -73960 22240 -73760 1 PIX1257_IN
port 1292 n
rlabel metal5 25040 -73960 25240 -73760 1 PIX1258_IN
port 1293 n
rlabel metal5 28040 -73960 28240 -73760 1 PIX1259_IN
port 1294 n
rlabel metal5 31040 -73960 31240 -73760 1 PIX1260_IN
port 1295 n
rlabel metal5 34040 -73960 34240 -73760 1 PIX1261_IN
port 1296 n
rlabel metal5 37040 -73960 37240 -73760 1 PIX1262_IN
port 1297 n
rlabel metal5 40040 -73960 40240 -73760 1 PIX1263_IN
port 1298 n
rlabel metal5 43040 -73960 43240 -73760 1 PIX1264_IN
port 1299 n
rlabel metal5 46040 -73960 46240 -73760 1 PIX1265_IN
port 1300 n
rlabel metal5 49040 -73960 49240 -73760 1 PIX1266_IN
port 1301 n
rlabel metal5 52040 -73960 52240 -73760 1 PIX1267_IN
port 1302 n
rlabel metal5 55040 -73960 55240 -73760 1 PIX1268_IN
port 1303 n
rlabel metal5 58040 -73960 58240 -73760 1 PIX1269_IN
port 1304 n
rlabel metal5 61040 -73960 61240 -73760 1 PIX1270_IN
port 1305 n
rlabel metal5 64040 -73960 64240 -73760 1 PIX1271_IN
port 1306 n
rlabel metal5 67040 -73960 67240 -73760 1 PIX1272_IN
port 1307 n
rlabel metal5 70040 -73960 70240 -73760 1 PIX1273_IN
port 1308 n
rlabel metal5 73040 -73960 73240 -73760 1 PIX1274_IN
port 1309 n
rlabel metal5 76040 -73960 76240 -73760 1 PIX1275_IN
port 1310 n
rlabel metal5 79040 -73960 79240 -73760 1 PIX1276_IN
port 1311 n
rlabel metal5 82040 -73960 82240 -73760 1 PIX1277_IN
port 1312 n
rlabel metal5 85040 -73960 85240 -73760 1 PIX1278_IN
port 1313 n
rlabel metal5 88040 -73960 88240 -73760 1 PIX1279_IN
port 1314 n
rlabel metal5 91040 -73960 91240 -73760 1 PIX1280_IN
port 1315 n
rlabel metal5 94040 -73960 94240 -73760 1 PIX1281_IN
port 1316 n
rlabel metal5 97040 -73960 97240 -73760 1 PIX1282_IN
port 1317 n
rlabel metal5 100040 -73960 100240 -73760 1 PIX1283_IN
port 1318 n
rlabel metal5 103040 -73960 103240 -73760 1 PIX1284_IN
port 1319 n
rlabel metal5 106040 -73960 106240 -73760 1 PIX1285_IN
port 1320 n
rlabel metal5 109040 -73960 109240 -73760 1 PIX1286_IN
port 1321 n
rlabel metal5 112040 -73960 112240 -73760 1 PIX1287_IN
port 1322 n
rlabel metal5 115040 -73960 115240 -73760 1 PIX1288_IN
port 1323 n
rlabel metal5 118040 -73960 118240 -73760 1 PIX1289_IN
port 1324 n
rlabel metal5 121040 -73960 121240 -73760 1 PIX1290_IN
port 1325 n
rlabel metal5 124040 -73960 124240 -73760 1 PIX1291_IN
port 1326 n
rlabel metal5 127040 -73960 127240 -73760 1 PIX1292_IN
port 1327 n
rlabel metal5 130040 -73960 130240 -73760 1 PIX1293_IN
port 1328 n
rlabel metal5 133040 -73960 133240 -73760 1 PIX1294_IN
port 1329 n
rlabel metal5 136040 -73960 136240 -73760 1 PIX1295_IN
port 1330 n
rlabel metal5 139040 -73960 139240 -73760 1 PIX1296_IN
port 1331 n
rlabel metal5 142040 -73960 142240 -73760 1 PIX1297_IN
port 1332 n
rlabel metal5 145040 -73960 145240 -73760 1 PIX1298_IN
port 1333 n
rlabel metal5 148040 -73960 148240 -73760 1 PIX1299_IN
port 1334 n
rlabel metal5 1040 -76960 1240 -76760 1 PIX1300_IN
port 1335 n
rlabel metal2 -3000 -76520 -3000 -76430 3 ROW_SEL26
port 1336 e
rlabel metal5 4040 -76960 4240 -76760 1 PIX1301_IN
port 1337 n
rlabel metal5 7040 -76960 7240 -76760 1 PIX1302_IN
port 1338 n
rlabel metal5 10040 -76960 10240 -76760 1 PIX1303_IN
port 1339 n
rlabel metal5 13040 -76960 13240 -76760 1 PIX1304_IN
port 1340 n
rlabel metal5 16040 -76960 16240 -76760 1 PIX1305_IN
port 1341 n
rlabel metal5 19040 -76960 19240 -76760 1 PIX1306_IN
port 1342 n
rlabel metal5 22040 -76960 22240 -76760 1 PIX1307_IN
port 1343 n
rlabel metal5 25040 -76960 25240 -76760 1 PIX1308_IN
port 1344 n
rlabel metal5 28040 -76960 28240 -76760 1 PIX1309_IN
port 1345 n
rlabel metal5 31040 -76960 31240 -76760 1 PIX1310_IN
port 1346 n
rlabel metal5 34040 -76960 34240 -76760 1 PIX1311_IN
port 1347 n
rlabel metal5 37040 -76960 37240 -76760 1 PIX1312_IN
port 1348 n
rlabel metal5 40040 -76960 40240 -76760 1 PIX1313_IN
port 1349 n
rlabel metal5 43040 -76960 43240 -76760 1 PIX1314_IN
port 1350 n
rlabel metal5 46040 -76960 46240 -76760 1 PIX1315_IN
port 1351 n
rlabel metal5 49040 -76960 49240 -76760 1 PIX1316_IN
port 1352 n
rlabel metal5 52040 -76960 52240 -76760 1 PIX1317_IN
port 1353 n
rlabel metal5 55040 -76960 55240 -76760 1 PIX1318_IN
port 1354 n
rlabel metal5 58040 -76960 58240 -76760 1 PIX1319_IN
port 1355 n
rlabel metal5 61040 -76960 61240 -76760 1 PIX1320_IN
port 1356 n
rlabel metal5 64040 -76960 64240 -76760 1 PIX1321_IN
port 1357 n
rlabel metal5 67040 -76960 67240 -76760 1 PIX1322_IN
port 1358 n
rlabel metal5 70040 -76960 70240 -76760 1 PIX1323_IN
port 1359 n
rlabel metal5 73040 -76960 73240 -76760 1 PIX1324_IN
port 1360 n
rlabel metal5 76040 -76960 76240 -76760 1 PIX1325_IN
port 1361 n
rlabel metal5 79040 -76960 79240 -76760 1 PIX1326_IN
port 1362 n
rlabel metal5 82040 -76960 82240 -76760 1 PIX1327_IN
port 1363 n
rlabel metal5 85040 -76960 85240 -76760 1 PIX1328_IN
port 1364 n
rlabel metal5 88040 -76960 88240 -76760 1 PIX1329_IN
port 1365 n
rlabel metal5 91040 -76960 91240 -76760 1 PIX1330_IN
port 1366 n
rlabel metal5 94040 -76960 94240 -76760 1 PIX1331_IN
port 1367 n
rlabel metal5 97040 -76960 97240 -76760 1 PIX1332_IN
port 1368 n
rlabel metal5 100040 -76960 100240 -76760 1 PIX1333_IN
port 1369 n
rlabel metal5 103040 -76960 103240 -76760 1 PIX1334_IN
port 1370 n
rlabel metal5 106040 -76960 106240 -76760 1 PIX1335_IN
port 1371 n
rlabel metal5 109040 -76960 109240 -76760 1 PIX1336_IN
port 1372 n
rlabel metal5 112040 -76960 112240 -76760 1 PIX1337_IN
port 1373 n
rlabel metal5 115040 -76960 115240 -76760 1 PIX1338_IN
port 1374 n
rlabel metal5 118040 -76960 118240 -76760 1 PIX1339_IN
port 1375 n
rlabel metal5 121040 -76960 121240 -76760 1 PIX1340_IN
port 1376 n
rlabel metal5 124040 -76960 124240 -76760 1 PIX1341_IN
port 1377 n
rlabel metal5 127040 -76960 127240 -76760 1 PIX1342_IN
port 1378 n
rlabel metal5 130040 -76960 130240 -76760 1 PIX1343_IN
port 1379 n
rlabel metal5 133040 -76960 133240 -76760 1 PIX1344_IN
port 1380 n
rlabel metal5 136040 -76960 136240 -76760 1 PIX1345_IN
port 1381 n
rlabel metal5 139040 -76960 139240 -76760 1 PIX1346_IN
port 1382 n
rlabel metal5 142040 -76960 142240 -76760 1 PIX1347_IN
port 1383 n
rlabel metal5 145040 -76960 145240 -76760 1 PIX1348_IN
port 1384 n
rlabel metal5 148040 -76960 148240 -76760 1 PIX1349_IN
port 1385 n
rlabel metal5 1040 -79960 1240 -79760 1 PIX1350_IN
port 1386 n
rlabel metal2 -3000 -79520 -3000 -79430 3 ROW_SEL27
port 1387 e
rlabel metal5 4040 -79960 4240 -79760 1 PIX1351_IN
port 1388 n
rlabel metal5 7040 -79960 7240 -79760 1 PIX1352_IN
port 1389 n
rlabel metal5 10040 -79960 10240 -79760 1 PIX1353_IN
port 1390 n
rlabel metal5 13040 -79960 13240 -79760 1 PIX1354_IN
port 1391 n
rlabel metal5 16040 -79960 16240 -79760 1 PIX1355_IN
port 1392 n
rlabel metal5 19040 -79960 19240 -79760 1 PIX1356_IN
port 1393 n
rlabel metal5 22040 -79960 22240 -79760 1 PIX1357_IN
port 1394 n
rlabel metal5 25040 -79960 25240 -79760 1 PIX1358_IN
port 1395 n
rlabel metal5 28040 -79960 28240 -79760 1 PIX1359_IN
port 1396 n
rlabel metal5 31040 -79960 31240 -79760 1 PIX1360_IN
port 1397 n
rlabel metal5 34040 -79960 34240 -79760 1 PIX1361_IN
port 1398 n
rlabel metal5 37040 -79960 37240 -79760 1 PIX1362_IN
port 1399 n
rlabel metal5 40040 -79960 40240 -79760 1 PIX1363_IN
port 1400 n
rlabel metal5 43040 -79960 43240 -79760 1 PIX1364_IN
port 1401 n
rlabel metal5 46040 -79960 46240 -79760 1 PIX1365_IN
port 1402 n
rlabel metal5 49040 -79960 49240 -79760 1 PIX1366_IN
port 1403 n
rlabel metal5 52040 -79960 52240 -79760 1 PIX1367_IN
port 1404 n
rlabel metal5 55040 -79960 55240 -79760 1 PIX1368_IN
port 1405 n
rlabel metal5 58040 -79960 58240 -79760 1 PIX1369_IN
port 1406 n
rlabel metal5 61040 -79960 61240 -79760 1 PIX1370_IN
port 1407 n
rlabel metal5 64040 -79960 64240 -79760 1 PIX1371_IN
port 1408 n
rlabel metal5 67040 -79960 67240 -79760 1 PIX1372_IN
port 1409 n
rlabel metal5 70040 -79960 70240 -79760 1 PIX1373_IN
port 1410 n
rlabel metal5 73040 -79960 73240 -79760 1 PIX1374_IN
port 1411 n
rlabel metal5 76040 -79960 76240 -79760 1 PIX1375_IN
port 1412 n
rlabel metal5 79040 -79960 79240 -79760 1 PIX1376_IN
port 1413 n
rlabel metal5 82040 -79960 82240 -79760 1 PIX1377_IN
port 1414 n
rlabel metal5 85040 -79960 85240 -79760 1 PIX1378_IN
port 1415 n
rlabel metal5 88040 -79960 88240 -79760 1 PIX1379_IN
port 1416 n
rlabel metal5 91040 -79960 91240 -79760 1 PIX1380_IN
port 1417 n
rlabel metal5 94040 -79960 94240 -79760 1 PIX1381_IN
port 1418 n
rlabel metal5 97040 -79960 97240 -79760 1 PIX1382_IN
port 1419 n
rlabel metal5 100040 -79960 100240 -79760 1 PIX1383_IN
port 1420 n
rlabel metal5 103040 -79960 103240 -79760 1 PIX1384_IN
port 1421 n
rlabel metal5 106040 -79960 106240 -79760 1 PIX1385_IN
port 1422 n
rlabel metal5 109040 -79960 109240 -79760 1 PIX1386_IN
port 1423 n
rlabel metal5 112040 -79960 112240 -79760 1 PIX1387_IN
port 1424 n
rlabel metal5 115040 -79960 115240 -79760 1 PIX1388_IN
port 1425 n
rlabel metal5 118040 -79960 118240 -79760 1 PIX1389_IN
port 1426 n
rlabel metal5 121040 -79960 121240 -79760 1 PIX1390_IN
port 1427 n
rlabel metal5 124040 -79960 124240 -79760 1 PIX1391_IN
port 1428 n
rlabel metal5 127040 -79960 127240 -79760 1 PIX1392_IN
port 1429 n
rlabel metal5 130040 -79960 130240 -79760 1 PIX1393_IN
port 1430 n
rlabel metal5 133040 -79960 133240 -79760 1 PIX1394_IN
port 1431 n
rlabel metal5 136040 -79960 136240 -79760 1 PIX1395_IN
port 1432 n
rlabel metal5 139040 -79960 139240 -79760 1 PIX1396_IN
port 1433 n
rlabel metal5 142040 -79960 142240 -79760 1 PIX1397_IN
port 1434 n
rlabel metal5 145040 -79960 145240 -79760 1 PIX1398_IN
port 1435 n
rlabel metal5 148040 -79960 148240 -79760 1 PIX1399_IN
port 1436 n
rlabel metal5 1040 -82960 1240 -82760 1 PIX1400_IN
port 1437 n
rlabel metal2 -3000 -82520 -3000 -82430 3 ROW_SEL28
port 1438 e
rlabel metal5 4040 -82960 4240 -82760 1 PIX1401_IN
port 1439 n
rlabel metal5 7040 -82960 7240 -82760 1 PIX1402_IN
port 1440 n
rlabel metal5 10040 -82960 10240 -82760 1 PIX1403_IN
port 1441 n
rlabel metal5 13040 -82960 13240 -82760 1 PIX1404_IN
port 1442 n
rlabel metal5 16040 -82960 16240 -82760 1 PIX1405_IN
port 1443 n
rlabel metal5 19040 -82960 19240 -82760 1 PIX1406_IN
port 1444 n
rlabel metal5 22040 -82960 22240 -82760 1 PIX1407_IN
port 1445 n
rlabel metal5 25040 -82960 25240 -82760 1 PIX1408_IN
port 1446 n
rlabel metal5 28040 -82960 28240 -82760 1 PIX1409_IN
port 1447 n
rlabel metal5 31040 -82960 31240 -82760 1 PIX1410_IN
port 1448 n
rlabel metal5 34040 -82960 34240 -82760 1 PIX1411_IN
port 1449 n
rlabel metal5 37040 -82960 37240 -82760 1 PIX1412_IN
port 1450 n
rlabel metal5 40040 -82960 40240 -82760 1 PIX1413_IN
port 1451 n
rlabel metal5 43040 -82960 43240 -82760 1 PIX1414_IN
port 1452 n
rlabel metal5 46040 -82960 46240 -82760 1 PIX1415_IN
port 1453 n
rlabel metal5 49040 -82960 49240 -82760 1 PIX1416_IN
port 1454 n
rlabel metal5 52040 -82960 52240 -82760 1 PIX1417_IN
port 1455 n
rlabel metal5 55040 -82960 55240 -82760 1 PIX1418_IN
port 1456 n
rlabel metal5 58040 -82960 58240 -82760 1 PIX1419_IN
port 1457 n
rlabel metal5 61040 -82960 61240 -82760 1 PIX1420_IN
port 1458 n
rlabel metal5 64040 -82960 64240 -82760 1 PIX1421_IN
port 1459 n
rlabel metal5 67040 -82960 67240 -82760 1 PIX1422_IN
port 1460 n
rlabel metal5 70040 -82960 70240 -82760 1 PIX1423_IN
port 1461 n
rlabel metal5 73040 -82960 73240 -82760 1 PIX1424_IN
port 1462 n
rlabel metal5 76040 -82960 76240 -82760 1 PIX1425_IN
port 1463 n
rlabel metal5 79040 -82960 79240 -82760 1 PIX1426_IN
port 1464 n
rlabel metal5 82040 -82960 82240 -82760 1 PIX1427_IN
port 1465 n
rlabel metal5 85040 -82960 85240 -82760 1 PIX1428_IN
port 1466 n
rlabel metal5 88040 -82960 88240 -82760 1 PIX1429_IN
port 1467 n
rlabel metal5 91040 -82960 91240 -82760 1 PIX1430_IN
port 1468 n
rlabel metal5 94040 -82960 94240 -82760 1 PIX1431_IN
port 1469 n
rlabel metal5 97040 -82960 97240 -82760 1 PIX1432_IN
port 1470 n
rlabel metal5 100040 -82960 100240 -82760 1 PIX1433_IN
port 1471 n
rlabel metal5 103040 -82960 103240 -82760 1 PIX1434_IN
port 1472 n
rlabel metal5 106040 -82960 106240 -82760 1 PIX1435_IN
port 1473 n
rlabel metal5 109040 -82960 109240 -82760 1 PIX1436_IN
port 1474 n
rlabel metal5 112040 -82960 112240 -82760 1 PIX1437_IN
port 1475 n
rlabel metal5 115040 -82960 115240 -82760 1 PIX1438_IN
port 1476 n
rlabel metal5 118040 -82960 118240 -82760 1 PIX1439_IN
port 1477 n
rlabel metal5 121040 -82960 121240 -82760 1 PIX1440_IN
port 1478 n
rlabel metal5 124040 -82960 124240 -82760 1 PIX1441_IN
port 1479 n
rlabel metal5 127040 -82960 127240 -82760 1 PIX1442_IN
port 1480 n
rlabel metal5 130040 -82960 130240 -82760 1 PIX1443_IN
port 1481 n
rlabel metal5 133040 -82960 133240 -82760 1 PIX1444_IN
port 1482 n
rlabel metal5 136040 -82960 136240 -82760 1 PIX1445_IN
port 1483 n
rlabel metal5 139040 -82960 139240 -82760 1 PIX1446_IN
port 1484 n
rlabel metal5 142040 -82960 142240 -82760 1 PIX1447_IN
port 1485 n
rlabel metal5 145040 -82960 145240 -82760 1 PIX1448_IN
port 1486 n
rlabel metal5 148040 -82960 148240 -82760 1 PIX1449_IN
port 1487 n
rlabel metal5 1040 -85960 1240 -85760 1 PIX1450_IN
port 1488 n
rlabel metal2 -3000 -85520 -3000 -85430 3 ROW_SEL29
port 1489 e
rlabel metal5 4040 -85960 4240 -85760 1 PIX1451_IN
port 1490 n
rlabel metal5 7040 -85960 7240 -85760 1 PIX1452_IN
port 1491 n
rlabel metal5 10040 -85960 10240 -85760 1 PIX1453_IN
port 1492 n
rlabel metal5 13040 -85960 13240 -85760 1 PIX1454_IN
port 1493 n
rlabel metal5 16040 -85960 16240 -85760 1 PIX1455_IN
port 1494 n
rlabel metal5 19040 -85960 19240 -85760 1 PIX1456_IN
port 1495 n
rlabel metal5 22040 -85960 22240 -85760 1 PIX1457_IN
port 1496 n
rlabel metal5 25040 -85960 25240 -85760 1 PIX1458_IN
port 1497 n
rlabel metal5 28040 -85960 28240 -85760 1 PIX1459_IN
port 1498 n
rlabel metal5 31040 -85960 31240 -85760 1 PIX1460_IN
port 1499 n
rlabel metal5 34040 -85960 34240 -85760 1 PIX1461_IN
port 1500 n
rlabel metal5 37040 -85960 37240 -85760 1 PIX1462_IN
port 1501 n
rlabel metal5 40040 -85960 40240 -85760 1 PIX1463_IN
port 1502 n
rlabel metal5 43040 -85960 43240 -85760 1 PIX1464_IN
port 1503 n
rlabel metal5 46040 -85960 46240 -85760 1 PIX1465_IN
port 1504 n
rlabel metal5 49040 -85960 49240 -85760 1 PIX1466_IN
port 1505 n
rlabel metal5 52040 -85960 52240 -85760 1 PIX1467_IN
port 1506 n
rlabel metal5 55040 -85960 55240 -85760 1 PIX1468_IN
port 1507 n
rlabel metal5 58040 -85960 58240 -85760 1 PIX1469_IN
port 1508 n
rlabel metal5 61040 -85960 61240 -85760 1 PIX1470_IN
port 1509 n
rlabel metal5 64040 -85960 64240 -85760 1 PIX1471_IN
port 1510 n
rlabel metal5 67040 -85960 67240 -85760 1 PIX1472_IN
port 1511 n
rlabel metal5 70040 -85960 70240 -85760 1 PIX1473_IN
port 1512 n
rlabel metal5 73040 -85960 73240 -85760 1 PIX1474_IN
port 1513 n
rlabel metal5 76040 -85960 76240 -85760 1 PIX1475_IN
port 1514 n
rlabel metal5 79040 -85960 79240 -85760 1 PIX1476_IN
port 1515 n
rlabel metal5 82040 -85960 82240 -85760 1 PIX1477_IN
port 1516 n
rlabel metal5 85040 -85960 85240 -85760 1 PIX1478_IN
port 1517 n
rlabel metal5 88040 -85960 88240 -85760 1 PIX1479_IN
port 1518 n
rlabel metal5 91040 -85960 91240 -85760 1 PIX1480_IN
port 1519 n
rlabel metal5 94040 -85960 94240 -85760 1 PIX1481_IN
port 1520 n
rlabel metal5 97040 -85960 97240 -85760 1 PIX1482_IN
port 1521 n
rlabel metal5 100040 -85960 100240 -85760 1 PIX1483_IN
port 1522 n
rlabel metal5 103040 -85960 103240 -85760 1 PIX1484_IN
port 1523 n
rlabel metal5 106040 -85960 106240 -85760 1 PIX1485_IN
port 1524 n
rlabel metal5 109040 -85960 109240 -85760 1 PIX1486_IN
port 1525 n
rlabel metal5 112040 -85960 112240 -85760 1 PIX1487_IN
port 1526 n
rlabel metal5 115040 -85960 115240 -85760 1 PIX1488_IN
port 1527 n
rlabel metal5 118040 -85960 118240 -85760 1 PIX1489_IN
port 1528 n
rlabel metal5 121040 -85960 121240 -85760 1 PIX1490_IN
port 1529 n
rlabel metal5 124040 -85960 124240 -85760 1 PIX1491_IN
port 1530 n
rlabel metal5 127040 -85960 127240 -85760 1 PIX1492_IN
port 1531 n
rlabel metal5 130040 -85960 130240 -85760 1 PIX1493_IN
port 1532 n
rlabel metal5 133040 -85960 133240 -85760 1 PIX1494_IN
port 1533 n
rlabel metal5 136040 -85960 136240 -85760 1 PIX1495_IN
port 1534 n
rlabel metal5 139040 -85960 139240 -85760 1 PIX1496_IN
port 1535 n
rlabel metal5 142040 -85960 142240 -85760 1 PIX1497_IN
port 1536 n
rlabel metal5 145040 -85960 145240 -85760 1 PIX1498_IN
port 1537 n
rlabel metal5 148040 -85960 148240 -85760 1 PIX1499_IN
port 1538 n
rlabel metal5 1040 -88960 1240 -88760 1 PIX1500_IN
port 1539 n
rlabel metal2 -3000 -88520 -3000 -88430 3 ROW_SEL30
port 1540 e
rlabel metal5 4040 -88960 4240 -88760 1 PIX1501_IN
port 1541 n
rlabel metal5 7040 -88960 7240 -88760 1 PIX1502_IN
port 1542 n
rlabel metal5 10040 -88960 10240 -88760 1 PIX1503_IN
port 1543 n
rlabel metal5 13040 -88960 13240 -88760 1 PIX1504_IN
port 1544 n
rlabel metal5 16040 -88960 16240 -88760 1 PIX1505_IN
port 1545 n
rlabel metal5 19040 -88960 19240 -88760 1 PIX1506_IN
port 1546 n
rlabel metal5 22040 -88960 22240 -88760 1 PIX1507_IN
port 1547 n
rlabel metal5 25040 -88960 25240 -88760 1 PIX1508_IN
port 1548 n
rlabel metal5 28040 -88960 28240 -88760 1 PIX1509_IN
port 1549 n
rlabel metal5 31040 -88960 31240 -88760 1 PIX1510_IN
port 1550 n
rlabel metal5 34040 -88960 34240 -88760 1 PIX1511_IN
port 1551 n
rlabel metal5 37040 -88960 37240 -88760 1 PIX1512_IN
port 1552 n
rlabel metal5 40040 -88960 40240 -88760 1 PIX1513_IN
port 1553 n
rlabel metal5 43040 -88960 43240 -88760 1 PIX1514_IN
port 1554 n
rlabel metal5 46040 -88960 46240 -88760 1 PIX1515_IN
port 1555 n
rlabel metal5 49040 -88960 49240 -88760 1 PIX1516_IN
port 1556 n
rlabel metal5 52040 -88960 52240 -88760 1 PIX1517_IN
port 1557 n
rlabel metal5 55040 -88960 55240 -88760 1 PIX1518_IN
port 1558 n
rlabel metal5 58040 -88960 58240 -88760 1 PIX1519_IN
port 1559 n
rlabel metal5 61040 -88960 61240 -88760 1 PIX1520_IN
port 1560 n
rlabel metal5 64040 -88960 64240 -88760 1 PIX1521_IN
port 1561 n
rlabel metal5 67040 -88960 67240 -88760 1 PIX1522_IN
port 1562 n
rlabel metal5 70040 -88960 70240 -88760 1 PIX1523_IN
port 1563 n
rlabel metal5 73040 -88960 73240 -88760 1 PIX1524_IN
port 1564 n
rlabel metal5 76040 -88960 76240 -88760 1 PIX1525_IN
port 1565 n
rlabel metal5 79040 -88960 79240 -88760 1 PIX1526_IN
port 1566 n
rlabel metal5 82040 -88960 82240 -88760 1 PIX1527_IN
port 1567 n
rlabel metal5 85040 -88960 85240 -88760 1 PIX1528_IN
port 1568 n
rlabel metal5 88040 -88960 88240 -88760 1 PIX1529_IN
port 1569 n
rlabel metal5 91040 -88960 91240 -88760 1 PIX1530_IN
port 1570 n
rlabel metal5 94040 -88960 94240 -88760 1 PIX1531_IN
port 1571 n
rlabel metal5 97040 -88960 97240 -88760 1 PIX1532_IN
port 1572 n
rlabel metal5 100040 -88960 100240 -88760 1 PIX1533_IN
port 1573 n
rlabel metal5 103040 -88960 103240 -88760 1 PIX1534_IN
port 1574 n
rlabel metal5 106040 -88960 106240 -88760 1 PIX1535_IN
port 1575 n
rlabel metal5 109040 -88960 109240 -88760 1 PIX1536_IN
port 1576 n
rlabel metal5 112040 -88960 112240 -88760 1 PIX1537_IN
port 1577 n
rlabel metal5 115040 -88960 115240 -88760 1 PIX1538_IN
port 1578 n
rlabel metal5 118040 -88960 118240 -88760 1 PIX1539_IN
port 1579 n
rlabel metal5 121040 -88960 121240 -88760 1 PIX1540_IN
port 1580 n
rlabel metal5 124040 -88960 124240 -88760 1 PIX1541_IN
port 1581 n
rlabel metal5 127040 -88960 127240 -88760 1 PIX1542_IN
port 1582 n
rlabel metal5 130040 -88960 130240 -88760 1 PIX1543_IN
port 1583 n
rlabel metal5 133040 -88960 133240 -88760 1 PIX1544_IN
port 1584 n
rlabel metal5 136040 -88960 136240 -88760 1 PIX1545_IN
port 1585 n
rlabel metal5 139040 -88960 139240 -88760 1 PIX1546_IN
port 1586 n
rlabel metal5 142040 -88960 142240 -88760 1 PIX1547_IN
port 1587 n
rlabel metal5 145040 -88960 145240 -88760 1 PIX1548_IN
port 1588 n
rlabel metal5 148040 -88960 148240 -88760 1 PIX1549_IN
port 1589 n
rlabel metal5 1040 -91960 1240 -91760 1 PIX1550_IN
port 1590 n
rlabel metal2 -3000 -91520 -3000 -91430 3 ROW_SEL31
port 1591 e
rlabel metal5 4040 -91960 4240 -91760 1 PIX1551_IN
port 1592 n
rlabel metal5 7040 -91960 7240 -91760 1 PIX1552_IN
port 1593 n
rlabel metal5 10040 -91960 10240 -91760 1 PIX1553_IN
port 1594 n
rlabel metal5 13040 -91960 13240 -91760 1 PIX1554_IN
port 1595 n
rlabel metal5 16040 -91960 16240 -91760 1 PIX1555_IN
port 1596 n
rlabel metal5 19040 -91960 19240 -91760 1 PIX1556_IN
port 1597 n
rlabel metal5 22040 -91960 22240 -91760 1 PIX1557_IN
port 1598 n
rlabel metal5 25040 -91960 25240 -91760 1 PIX1558_IN
port 1599 n
rlabel metal5 28040 -91960 28240 -91760 1 PIX1559_IN
port 1600 n
rlabel metal5 31040 -91960 31240 -91760 1 PIX1560_IN
port 1601 n
rlabel metal5 34040 -91960 34240 -91760 1 PIX1561_IN
port 1602 n
rlabel metal5 37040 -91960 37240 -91760 1 PIX1562_IN
port 1603 n
rlabel metal5 40040 -91960 40240 -91760 1 PIX1563_IN
port 1604 n
rlabel metal5 43040 -91960 43240 -91760 1 PIX1564_IN
port 1605 n
rlabel metal5 46040 -91960 46240 -91760 1 PIX1565_IN
port 1606 n
rlabel metal5 49040 -91960 49240 -91760 1 PIX1566_IN
port 1607 n
rlabel metal5 52040 -91960 52240 -91760 1 PIX1567_IN
port 1608 n
rlabel metal5 55040 -91960 55240 -91760 1 PIX1568_IN
port 1609 n
rlabel metal5 58040 -91960 58240 -91760 1 PIX1569_IN
port 1610 n
rlabel metal5 61040 -91960 61240 -91760 1 PIX1570_IN
port 1611 n
rlabel metal5 64040 -91960 64240 -91760 1 PIX1571_IN
port 1612 n
rlabel metal5 67040 -91960 67240 -91760 1 PIX1572_IN
port 1613 n
rlabel metal5 70040 -91960 70240 -91760 1 PIX1573_IN
port 1614 n
rlabel metal5 73040 -91960 73240 -91760 1 PIX1574_IN
port 1615 n
rlabel metal5 76040 -91960 76240 -91760 1 PIX1575_IN
port 1616 n
rlabel metal5 79040 -91960 79240 -91760 1 PIX1576_IN
port 1617 n
rlabel metal5 82040 -91960 82240 -91760 1 PIX1577_IN
port 1618 n
rlabel metal5 85040 -91960 85240 -91760 1 PIX1578_IN
port 1619 n
rlabel metal5 88040 -91960 88240 -91760 1 PIX1579_IN
port 1620 n
rlabel metal5 91040 -91960 91240 -91760 1 PIX1580_IN
port 1621 n
rlabel metal5 94040 -91960 94240 -91760 1 PIX1581_IN
port 1622 n
rlabel metal5 97040 -91960 97240 -91760 1 PIX1582_IN
port 1623 n
rlabel metal5 100040 -91960 100240 -91760 1 PIX1583_IN
port 1624 n
rlabel metal5 103040 -91960 103240 -91760 1 PIX1584_IN
port 1625 n
rlabel metal5 106040 -91960 106240 -91760 1 PIX1585_IN
port 1626 n
rlabel metal5 109040 -91960 109240 -91760 1 PIX1586_IN
port 1627 n
rlabel metal5 112040 -91960 112240 -91760 1 PIX1587_IN
port 1628 n
rlabel metal5 115040 -91960 115240 -91760 1 PIX1588_IN
port 1629 n
rlabel metal5 118040 -91960 118240 -91760 1 PIX1589_IN
port 1630 n
rlabel metal5 121040 -91960 121240 -91760 1 PIX1590_IN
port 1631 n
rlabel metal5 124040 -91960 124240 -91760 1 PIX1591_IN
port 1632 n
rlabel metal5 127040 -91960 127240 -91760 1 PIX1592_IN
port 1633 n
rlabel metal5 130040 -91960 130240 -91760 1 PIX1593_IN
port 1634 n
rlabel metal5 133040 -91960 133240 -91760 1 PIX1594_IN
port 1635 n
rlabel metal5 136040 -91960 136240 -91760 1 PIX1595_IN
port 1636 n
rlabel metal5 139040 -91960 139240 -91760 1 PIX1596_IN
port 1637 n
rlabel metal5 142040 -91960 142240 -91760 1 PIX1597_IN
port 1638 n
rlabel metal5 145040 -91960 145240 -91760 1 PIX1598_IN
port 1639 n
rlabel metal5 148040 -91960 148240 -91760 1 PIX1599_IN
port 1640 n
rlabel metal5 1040 -94960 1240 -94760 1 PIX1600_IN
port 1641 n
rlabel metal2 -3000 -94520 -3000 -94430 3 ROW_SEL32
port 1642 e
rlabel metal5 4040 -94960 4240 -94760 1 PIX1601_IN
port 1643 n
rlabel metal5 7040 -94960 7240 -94760 1 PIX1602_IN
port 1644 n
rlabel metal5 10040 -94960 10240 -94760 1 PIX1603_IN
port 1645 n
rlabel metal5 13040 -94960 13240 -94760 1 PIX1604_IN
port 1646 n
rlabel metal5 16040 -94960 16240 -94760 1 PIX1605_IN
port 1647 n
rlabel metal5 19040 -94960 19240 -94760 1 PIX1606_IN
port 1648 n
rlabel metal5 22040 -94960 22240 -94760 1 PIX1607_IN
port 1649 n
rlabel metal5 25040 -94960 25240 -94760 1 PIX1608_IN
port 1650 n
rlabel metal5 28040 -94960 28240 -94760 1 PIX1609_IN
port 1651 n
rlabel metal5 31040 -94960 31240 -94760 1 PIX1610_IN
port 1652 n
rlabel metal5 34040 -94960 34240 -94760 1 PIX1611_IN
port 1653 n
rlabel metal5 37040 -94960 37240 -94760 1 PIX1612_IN
port 1654 n
rlabel metal5 40040 -94960 40240 -94760 1 PIX1613_IN
port 1655 n
rlabel metal5 43040 -94960 43240 -94760 1 PIX1614_IN
port 1656 n
rlabel metal5 46040 -94960 46240 -94760 1 PIX1615_IN
port 1657 n
rlabel metal5 49040 -94960 49240 -94760 1 PIX1616_IN
port 1658 n
rlabel metal5 52040 -94960 52240 -94760 1 PIX1617_IN
port 1659 n
rlabel metal5 55040 -94960 55240 -94760 1 PIX1618_IN
port 1660 n
rlabel metal5 58040 -94960 58240 -94760 1 PIX1619_IN
port 1661 n
rlabel metal5 61040 -94960 61240 -94760 1 PIX1620_IN
port 1662 n
rlabel metal5 64040 -94960 64240 -94760 1 PIX1621_IN
port 1663 n
rlabel metal5 67040 -94960 67240 -94760 1 PIX1622_IN
port 1664 n
rlabel metal5 70040 -94960 70240 -94760 1 PIX1623_IN
port 1665 n
rlabel metal5 73040 -94960 73240 -94760 1 PIX1624_IN
port 1666 n
rlabel metal5 76040 -94960 76240 -94760 1 PIX1625_IN
port 1667 n
rlabel metal5 79040 -94960 79240 -94760 1 PIX1626_IN
port 1668 n
rlabel metal5 82040 -94960 82240 -94760 1 PIX1627_IN
port 1669 n
rlabel metal5 85040 -94960 85240 -94760 1 PIX1628_IN
port 1670 n
rlabel metal5 88040 -94960 88240 -94760 1 PIX1629_IN
port 1671 n
rlabel metal5 91040 -94960 91240 -94760 1 PIX1630_IN
port 1672 n
rlabel metal5 94040 -94960 94240 -94760 1 PIX1631_IN
port 1673 n
rlabel metal5 97040 -94960 97240 -94760 1 PIX1632_IN
port 1674 n
rlabel metal5 100040 -94960 100240 -94760 1 PIX1633_IN
port 1675 n
rlabel metal5 103040 -94960 103240 -94760 1 PIX1634_IN
port 1676 n
rlabel metal5 106040 -94960 106240 -94760 1 PIX1635_IN
port 1677 n
rlabel metal5 109040 -94960 109240 -94760 1 PIX1636_IN
port 1678 n
rlabel metal5 112040 -94960 112240 -94760 1 PIX1637_IN
port 1679 n
rlabel metal5 115040 -94960 115240 -94760 1 PIX1638_IN
port 1680 n
rlabel metal5 118040 -94960 118240 -94760 1 PIX1639_IN
port 1681 n
rlabel metal5 121040 -94960 121240 -94760 1 PIX1640_IN
port 1682 n
rlabel metal5 124040 -94960 124240 -94760 1 PIX1641_IN
port 1683 n
rlabel metal5 127040 -94960 127240 -94760 1 PIX1642_IN
port 1684 n
rlabel metal5 130040 -94960 130240 -94760 1 PIX1643_IN
port 1685 n
rlabel metal5 133040 -94960 133240 -94760 1 PIX1644_IN
port 1686 n
rlabel metal5 136040 -94960 136240 -94760 1 PIX1645_IN
port 1687 n
rlabel metal5 139040 -94960 139240 -94760 1 PIX1646_IN
port 1688 n
rlabel metal5 142040 -94960 142240 -94760 1 PIX1647_IN
port 1689 n
rlabel metal5 145040 -94960 145240 -94760 1 PIX1648_IN
port 1690 n
rlabel metal5 148040 -94960 148240 -94760 1 PIX1649_IN
port 1691 n
rlabel metal5 1040 -97960 1240 -97760 1 PIX1650_IN
port 1692 n
rlabel metal2 -3000 -97520 -3000 -97430 3 ROW_SEL33
port 1693 e
rlabel metal5 4040 -97960 4240 -97760 1 PIX1651_IN
port 1694 n
rlabel metal5 7040 -97960 7240 -97760 1 PIX1652_IN
port 1695 n
rlabel metal5 10040 -97960 10240 -97760 1 PIX1653_IN
port 1696 n
rlabel metal5 13040 -97960 13240 -97760 1 PIX1654_IN
port 1697 n
rlabel metal5 16040 -97960 16240 -97760 1 PIX1655_IN
port 1698 n
rlabel metal5 19040 -97960 19240 -97760 1 PIX1656_IN
port 1699 n
rlabel metal5 22040 -97960 22240 -97760 1 PIX1657_IN
port 1700 n
rlabel metal5 25040 -97960 25240 -97760 1 PIX1658_IN
port 1701 n
rlabel metal5 28040 -97960 28240 -97760 1 PIX1659_IN
port 1702 n
rlabel metal5 31040 -97960 31240 -97760 1 PIX1660_IN
port 1703 n
rlabel metal5 34040 -97960 34240 -97760 1 PIX1661_IN
port 1704 n
rlabel metal5 37040 -97960 37240 -97760 1 PIX1662_IN
port 1705 n
rlabel metal5 40040 -97960 40240 -97760 1 PIX1663_IN
port 1706 n
rlabel metal5 43040 -97960 43240 -97760 1 PIX1664_IN
port 1707 n
rlabel metal5 46040 -97960 46240 -97760 1 PIX1665_IN
port 1708 n
rlabel metal5 49040 -97960 49240 -97760 1 PIX1666_IN
port 1709 n
rlabel metal5 52040 -97960 52240 -97760 1 PIX1667_IN
port 1710 n
rlabel metal5 55040 -97960 55240 -97760 1 PIX1668_IN
port 1711 n
rlabel metal5 58040 -97960 58240 -97760 1 PIX1669_IN
port 1712 n
rlabel metal5 61040 -97960 61240 -97760 1 PIX1670_IN
port 1713 n
rlabel metal5 64040 -97960 64240 -97760 1 PIX1671_IN
port 1714 n
rlabel metal5 67040 -97960 67240 -97760 1 PIX1672_IN
port 1715 n
rlabel metal5 70040 -97960 70240 -97760 1 PIX1673_IN
port 1716 n
rlabel metal5 73040 -97960 73240 -97760 1 PIX1674_IN
port 1717 n
rlabel metal5 76040 -97960 76240 -97760 1 PIX1675_IN
port 1718 n
rlabel metal5 79040 -97960 79240 -97760 1 PIX1676_IN
port 1719 n
rlabel metal5 82040 -97960 82240 -97760 1 PIX1677_IN
port 1720 n
rlabel metal5 85040 -97960 85240 -97760 1 PIX1678_IN
port 1721 n
rlabel metal5 88040 -97960 88240 -97760 1 PIX1679_IN
port 1722 n
rlabel metal5 91040 -97960 91240 -97760 1 PIX1680_IN
port 1723 n
rlabel metal5 94040 -97960 94240 -97760 1 PIX1681_IN
port 1724 n
rlabel metal5 97040 -97960 97240 -97760 1 PIX1682_IN
port 1725 n
rlabel metal5 100040 -97960 100240 -97760 1 PIX1683_IN
port 1726 n
rlabel metal5 103040 -97960 103240 -97760 1 PIX1684_IN
port 1727 n
rlabel metal5 106040 -97960 106240 -97760 1 PIX1685_IN
port 1728 n
rlabel metal5 109040 -97960 109240 -97760 1 PIX1686_IN
port 1729 n
rlabel metal5 112040 -97960 112240 -97760 1 PIX1687_IN
port 1730 n
rlabel metal5 115040 -97960 115240 -97760 1 PIX1688_IN
port 1731 n
rlabel metal5 118040 -97960 118240 -97760 1 PIX1689_IN
port 1732 n
rlabel metal5 121040 -97960 121240 -97760 1 PIX1690_IN
port 1733 n
rlabel metal5 124040 -97960 124240 -97760 1 PIX1691_IN
port 1734 n
rlabel metal5 127040 -97960 127240 -97760 1 PIX1692_IN
port 1735 n
rlabel metal5 130040 -97960 130240 -97760 1 PIX1693_IN
port 1736 n
rlabel metal5 133040 -97960 133240 -97760 1 PIX1694_IN
port 1737 n
rlabel metal5 136040 -97960 136240 -97760 1 PIX1695_IN
port 1738 n
rlabel metal5 139040 -97960 139240 -97760 1 PIX1696_IN
port 1739 n
rlabel metal5 142040 -97960 142240 -97760 1 PIX1697_IN
port 1740 n
rlabel metal5 145040 -97960 145240 -97760 1 PIX1698_IN
port 1741 n
rlabel metal5 148040 -97960 148240 -97760 1 PIX1699_IN
port 1742 n
rlabel metal5 1040 -100960 1240 -100760 1 PIX1700_IN
port 1743 n
rlabel metal2 -3000 -100520 -3000 -100430 3 ROW_SEL34
port 1744 e
rlabel metal5 4040 -100960 4240 -100760 1 PIX1701_IN
port 1745 n
rlabel metal5 7040 -100960 7240 -100760 1 PIX1702_IN
port 1746 n
rlabel metal5 10040 -100960 10240 -100760 1 PIX1703_IN
port 1747 n
rlabel metal5 13040 -100960 13240 -100760 1 PIX1704_IN
port 1748 n
rlabel metal5 16040 -100960 16240 -100760 1 PIX1705_IN
port 1749 n
rlabel metal5 19040 -100960 19240 -100760 1 PIX1706_IN
port 1750 n
rlabel metal5 22040 -100960 22240 -100760 1 PIX1707_IN
port 1751 n
rlabel metal5 25040 -100960 25240 -100760 1 PIX1708_IN
port 1752 n
rlabel metal5 28040 -100960 28240 -100760 1 PIX1709_IN
port 1753 n
rlabel metal5 31040 -100960 31240 -100760 1 PIX1710_IN
port 1754 n
rlabel metal5 34040 -100960 34240 -100760 1 PIX1711_IN
port 1755 n
rlabel metal5 37040 -100960 37240 -100760 1 PIX1712_IN
port 1756 n
rlabel metal5 40040 -100960 40240 -100760 1 PIX1713_IN
port 1757 n
rlabel metal5 43040 -100960 43240 -100760 1 PIX1714_IN
port 1758 n
rlabel metal5 46040 -100960 46240 -100760 1 PIX1715_IN
port 1759 n
rlabel metal5 49040 -100960 49240 -100760 1 PIX1716_IN
port 1760 n
rlabel metal5 52040 -100960 52240 -100760 1 PIX1717_IN
port 1761 n
rlabel metal5 55040 -100960 55240 -100760 1 PIX1718_IN
port 1762 n
rlabel metal5 58040 -100960 58240 -100760 1 PIX1719_IN
port 1763 n
rlabel metal5 61040 -100960 61240 -100760 1 PIX1720_IN
port 1764 n
rlabel metal5 64040 -100960 64240 -100760 1 PIX1721_IN
port 1765 n
rlabel metal5 67040 -100960 67240 -100760 1 PIX1722_IN
port 1766 n
rlabel metal5 70040 -100960 70240 -100760 1 PIX1723_IN
port 1767 n
rlabel metal5 73040 -100960 73240 -100760 1 PIX1724_IN
port 1768 n
rlabel metal5 76040 -100960 76240 -100760 1 PIX1725_IN
port 1769 n
rlabel metal5 79040 -100960 79240 -100760 1 PIX1726_IN
port 1770 n
rlabel metal5 82040 -100960 82240 -100760 1 PIX1727_IN
port 1771 n
rlabel metal5 85040 -100960 85240 -100760 1 PIX1728_IN
port 1772 n
rlabel metal5 88040 -100960 88240 -100760 1 PIX1729_IN
port 1773 n
rlabel metal5 91040 -100960 91240 -100760 1 PIX1730_IN
port 1774 n
rlabel metal5 94040 -100960 94240 -100760 1 PIX1731_IN
port 1775 n
rlabel metal5 97040 -100960 97240 -100760 1 PIX1732_IN
port 1776 n
rlabel metal5 100040 -100960 100240 -100760 1 PIX1733_IN
port 1777 n
rlabel metal5 103040 -100960 103240 -100760 1 PIX1734_IN
port 1778 n
rlabel metal5 106040 -100960 106240 -100760 1 PIX1735_IN
port 1779 n
rlabel metal5 109040 -100960 109240 -100760 1 PIX1736_IN
port 1780 n
rlabel metal5 112040 -100960 112240 -100760 1 PIX1737_IN
port 1781 n
rlabel metal5 115040 -100960 115240 -100760 1 PIX1738_IN
port 1782 n
rlabel metal5 118040 -100960 118240 -100760 1 PIX1739_IN
port 1783 n
rlabel metal5 121040 -100960 121240 -100760 1 PIX1740_IN
port 1784 n
rlabel metal5 124040 -100960 124240 -100760 1 PIX1741_IN
port 1785 n
rlabel metal5 127040 -100960 127240 -100760 1 PIX1742_IN
port 1786 n
rlabel metal5 130040 -100960 130240 -100760 1 PIX1743_IN
port 1787 n
rlabel metal5 133040 -100960 133240 -100760 1 PIX1744_IN
port 1788 n
rlabel metal5 136040 -100960 136240 -100760 1 PIX1745_IN
port 1789 n
rlabel metal5 139040 -100960 139240 -100760 1 PIX1746_IN
port 1790 n
rlabel metal5 142040 -100960 142240 -100760 1 PIX1747_IN
port 1791 n
rlabel metal5 145040 -100960 145240 -100760 1 PIX1748_IN
port 1792 n
rlabel metal5 148040 -100960 148240 -100760 1 PIX1749_IN
port 1793 n
rlabel metal5 1040 -103960 1240 -103760 1 PIX1750_IN
port 1794 n
rlabel metal2 -3000 -103520 -3000 -103430 3 ROW_SEL35
port 1795 e
rlabel metal5 4040 -103960 4240 -103760 1 PIX1751_IN
port 1796 n
rlabel metal5 7040 -103960 7240 -103760 1 PIX1752_IN
port 1797 n
rlabel metal5 10040 -103960 10240 -103760 1 PIX1753_IN
port 1798 n
rlabel metal5 13040 -103960 13240 -103760 1 PIX1754_IN
port 1799 n
rlabel metal5 16040 -103960 16240 -103760 1 PIX1755_IN
port 1800 n
rlabel metal5 19040 -103960 19240 -103760 1 PIX1756_IN
port 1801 n
rlabel metal5 22040 -103960 22240 -103760 1 PIX1757_IN
port 1802 n
rlabel metal5 25040 -103960 25240 -103760 1 PIX1758_IN
port 1803 n
rlabel metal5 28040 -103960 28240 -103760 1 PIX1759_IN
port 1804 n
rlabel metal5 31040 -103960 31240 -103760 1 PIX1760_IN
port 1805 n
rlabel metal5 34040 -103960 34240 -103760 1 PIX1761_IN
port 1806 n
rlabel metal5 37040 -103960 37240 -103760 1 PIX1762_IN
port 1807 n
rlabel metal5 40040 -103960 40240 -103760 1 PIX1763_IN
port 1808 n
rlabel metal5 43040 -103960 43240 -103760 1 PIX1764_IN
port 1809 n
rlabel metal5 46040 -103960 46240 -103760 1 PIX1765_IN
port 1810 n
rlabel metal5 49040 -103960 49240 -103760 1 PIX1766_IN
port 1811 n
rlabel metal5 52040 -103960 52240 -103760 1 PIX1767_IN
port 1812 n
rlabel metal5 55040 -103960 55240 -103760 1 PIX1768_IN
port 1813 n
rlabel metal5 58040 -103960 58240 -103760 1 PIX1769_IN
port 1814 n
rlabel metal5 61040 -103960 61240 -103760 1 PIX1770_IN
port 1815 n
rlabel metal5 64040 -103960 64240 -103760 1 PIX1771_IN
port 1816 n
rlabel metal5 67040 -103960 67240 -103760 1 PIX1772_IN
port 1817 n
rlabel metal5 70040 -103960 70240 -103760 1 PIX1773_IN
port 1818 n
rlabel metal5 73040 -103960 73240 -103760 1 PIX1774_IN
port 1819 n
rlabel metal5 76040 -103960 76240 -103760 1 PIX1775_IN
port 1820 n
rlabel metal5 79040 -103960 79240 -103760 1 PIX1776_IN
port 1821 n
rlabel metal5 82040 -103960 82240 -103760 1 PIX1777_IN
port 1822 n
rlabel metal5 85040 -103960 85240 -103760 1 PIX1778_IN
port 1823 n
rlabel metal5 88040 -103960 88240 -103760 1 PIX1779_IN
port 1824 n
rlabel metal5 91040 -103960 91240 -103760 1 PIX1780_IN
port 1825 n
rlabel metal5 94040 -103960 94240 -103760 1 PIX1781_IN
port 1826 n
rlabel metal5 97040 -103960 97240 -103760 1 PIX1782_IN
port 1827 n
rlabel metal5 100040 -103960 100240 -103760 1 PIX1783_IN
port 1828 n
rlabel metal5 103040 -103960 103240 -103760 1 PIX1784_IN
port 1829 n
rlabel metal5 106040 -103960 106240 -103760 1 PIX1785_IN
port 1830 n
rlabel metal5 109040 -103960 109240 -103760 1 PIX1786_IN
port 1831 n
rlabel metal5 112040 -103960 112240 -103760 1 PIX1787_IN
port 1832 n
rlabel metal5 115040 -103960 115240 -103760 1 PIX1788_IN
port 1833 n
rlabel metal5 118040 -103960 118240 -103760 1 PIX1789_IN
port 1834 n
rlabel metal5 121040 -103960 121240 -103760 1 PIX1790_IN
port 1835 n
rlabel metal5 124040 -103960 124240 -103760 1 PIX1791_IN
port 1836 n
rlabel metal5 127040 -103960 127240 -103760 1 PIX1792_IN
port 1837 n
rlabel metal5 130040 -103960 130240 -103760 1 PIX1793_IN
port 1838 n
rlabel metal5 133040 -103960 133240 -103760 1 PIX1794_IN
port 1839 n
rlabel metal5 136040 -103960 136240 -103760 1 PIX1795_IN
port 1840 n
rlabel metal5 139040 -103960 139240 -103760 1 PIX1796_IN
port 1841 n
rlabel metal5 142040 -103960 142240 -103760 1 PIX1797_IN
port 1842 n
rlabel metal5 145040 -103960 145240 -103760 1 PIX1798_IN
port 1843 n
rlabel metal5 148040 -103960 148240 -103760 1 PIX1799_IN
port 1844 n
rlabel metal5 1040 -106960 1240 -106760 1 PIX1800_IN
port 1845 n
rlabel metal2 -3000 -106520 -3000 -106430 3 ROW_SEL36
port 1846 e
rlabel metal5 4040 -106960 4240 -106760 1 PIX1801_IN
port 1847 n
rlabel metal5 7040 -106960 7240 -106760 1 PIX1802_IN
port 1848 n
rlabel metal5 10040 -106960 10240 -106760 1 PIX1803_IN
port 1849 n
rlabel metal5 13040 -106960 13240 -106760 1 PIX1804_IN
port 1850 n
rlabel metal5 16040 -106960 16240 -106760 1 PIX1805_IN
port 1851 n
rlabel metal5 19040 -106960 19240 -106760 1 PIX1806_IN
port 1852 n
rlabel metal5 22040 -106960 22240 -106760 1 PIX1807_IN
port 1853 n
rlabel metal5 25040 -106960 25240 -106760 1 PIX1808_IN
port 1854 n
rlabel metal5 28040 -106960 28240 -106760 1 PIX1809_IN
port 1855 n
rlabel metal5 31040 -106960 31240 -106760 1 PIX1810_IN
port 1856 n
rlabel metal5 34040 -106960 34240 -106760 1 PIX1811_IN
port 1857 n
rlabel metal5 37040 -106960 37240 -106760 1 PIX1812_IN
port 1858 n
rlabel metal5 40040 -106960 40240 -106760 1 PIX1813_IN
port 1859 n
rlabel metal5 43040 -106960 43240 -106760 1 PIX1814_IN
port 1860 n
rlabel metal5 46040 -106960 46240 -106760 1 PIX1815_IN
port 1861 n
rlabel metal5 49040 -106960 49240 -106760 1 PIX1816_IN
port 1862 n
rlabel metal5 52040 -106960 52240 -106760 1 PIX1817_IN
port 1863 n
rlabel metal5 55040 -106960 55240 -106760 1 PIX1818_IN
port 1864 n
rlabel metal5 58040 -106960 58240 -106760 1 PIX1819_IN
port 1865 n
rlabel metal5 61040 -106960 61240 -106760 1 PIX1820_IN
port 1866 n
rlabel metal5 64040 -106960 64240 -106760 1 PIX1821_IN
port 1867 n
rlabel metal5 67040 -106960 67240 -106760 1 PIX1822_IN
port 1868 n
rlabel metal5 70040 -106960 70240 -106760 1 PIX1823_IN
port 1869 n
rlabel metal5 73040 -106960 73240 -106760 1 PIX1824_IN
port 1870 n
rlabel metal5 76040 -106960 76240 -106760 1 PIX1825_IN
port 1871 n
rlabel metal5 79040 -106960 79240 -106760 1 PIX1826_IN
port 1872 n
rlabel metal5 82040 -106960 82240 -106760 1 PIX1827_IN
port 1873 n
rlabel metal5 85040 -106960 85240 -106760 1 PIX1828_IN
port 1874 n
rlabel metal5 88040 -106960 88240 -106760 1 PIX1829_IN
port 1875 n
rlabel metal5 91040 -106960 91240 -106760 1 PIX1830_IN
port 1876 n
rlabel metal5 94040 -106960 94240 -106760 1 PIX1831_IN
port 1877 n
rlabel metal5 97040 -106960 97240 -106760 1 PIX1832_IN
port 1878 n
rlabel metal5 100040 -106960 100240 -106760 1 PIX1833_IN
port 1879 n
rlabel metal5 103040 -106960 103240 -106760 1 PIX1834_IN
port 1880 n
rlabel metal5 106040 -106960 106240 -106760 1 PIX1835_IN
port 1881 n
rlabel metal5 109040 -106960 109240 -106760 1 PIX1836_IN
port 1882 n
rlabel metal5 112040 -106960 112240 -106760 1 PIX1837_IN
port 1883 n
rlabel metal5 115040 -106960 115240 -106760 1 PIX1838_IN
port 1884 n
rlabel metal5 118040 -106960 118240 -106760 1 PIX1839_IN
port 1885 n
rlabel metal5 121040 -106960 121240 -106760 1 PIX1840_IN
port 1886 n
rlabel metal5 124040 -106960 124240 -106760 1 PIX1841_IN
port 1887 n
rlabel metal5 127040 -106960 127240 -106760 1 PIX1842_IN
port 1888 n
rlabel metal5 130040 -106960 130240 -106760 1 PIX1843_IN
port 1889 n
rlabel metal5 133040 -106960 133240 -106760 1 PIX1844_IN
port 1890 n
rlabel metal5 136040 -106960 136240 -106760 1 PIX1845_IN
port 1891 n
rlabel metal5 139040 -106960 139240 -106760 1 PIX1846_IN
port 1892 n
rlabel metal5 142040 -106960 142240 -106760 1 PIX1847_IN
port 1893 n
rlabel metal5 145040 -106960 145240 -106760 1 PIX1848_IN
port 1894 n
rlabel metal5 148040 -106960 148240 -106760 1 PIX1849_IN
port 1895 n
rlabel metal5 1040 -109960 1240 -109760 1 PIX1850_IN
port 1896 n
rlabel metal2 -3000 -109520 -3000 -109430 3 ROW_SEL37
port 1897 e
rlabel metal5 4040 -109960 4240 -109760 1 PIX1851_IN
port 1898 n
rlabel metal5 7040 -109960 7240 -109760 1 PIX1852_IN
port 1899 n
rlabel metal5 10040 -109960 10240 -109760 1 PIX1853_IN
port 1900 n
rlabel metal5 13040 -109960 13240 -109760 1 PIX1854_IN
port 1901 n
rlabel metal5 16040 -109960 16240 -109760 1 PIX1855_IN
port 1902 n
rlabel metal5 19040 -109960 19240 -109760 1 PIX1856_IN
port 1903 n
rlabel metal5 22040 -109960 22240 -109760 1 PIX1857_IN
port 1904 n
rlabel metal5 25040 -109960 25240 -109760 1 PIX1858_IN
port 1905 n
rlabel metal5 28040 -109960 28240 -109760 1 PIX1859_IN
port 1906 n
rlabel metal5 31040 -109960 31240 -109760 1 PIX1860_IN
port 1907 n
rlabel metal5 34040 -109960 34240 -109760 1 PIX1861_IN
port 1908 n
rlabel metal5 37040 -109960 37240 -109760 1 PIX1862_IN
port 1909 n
rlabel metal5 40040 -109960 40240 -109760 1 PIX1863_IN
port 1910 n
rlabel metal5 43040 -109960 43240 -109760 1 PIX1864_IN
port 1911 n
rlabel metal5 46040 -109960 46240 -109760 1 PIX1865_IN
port 1912 n
rlabel metal5 49040 -109960 49240 -109760 1 PIX1866_IN
port 1913 n
rlabel metal5 52040 -109960 52240 -109760 1 PIX1867_IN
port 1914 n
rlabel metal5 55040 -109960 55240 -109760 1 PIX1868_IN
port 1915 n
rlabel metal5 58040 -109960 58240 -109760 1 PIX1869_IN
port 1916 n
rlabel metal5 61040 -109960 61240 -109760 1 PIX1870_IN
port 1917 n
rlabel metal5 64040 -109960 64240 -109760 1 PIX1871_IN
port 1918 n
rlabel metal5 67040 -109960 67240 -109760 1 PIX1872_IN
port 1919 n
rlabel metal5 70040 -109960 70240 -109760 1 PIX1873_IN
port 1920 n
rlabel metal5 73040 -109960 73240 -109760 1 PIX1874_IN
port 1921 n
rlabel metal5 76040 -109960 76240 -109760 1 PIX1875_IN
port 1922 n
rlabel metal5 79040 -109960 79240 -109760 1 PIX1876_IN
port 1923 n
rlabel metal5 82040 -109960 82240 -109760 1 PIX1877_IN
port 1924 n
rlabel metal5 85040 -109960 85240 -109760 1 PIX1878_IN
port 1925 n
rlabel metal5 88040 -109960 88240 -109760 1 PIX1879_IN
port 1926 n
rlabel metal5 91040 -109960 91240 -109760 1 PIX1880_IN
port 1927 n
rlabel metal5 94040 -109960 94240 -109760 1 PIX1881_IN
port 1928 n
rlabel metal5 97040 -109960 97240 -109760 1 PIX1882_IN
port 1929 n
rlabel metal5 100040 -109960 100240 -109760 1 PIX1883_IN
port 1930 n
rlabel metal5 103040 -109960 103240 -109760 1 PIX1884_IN
port 1931 n
rlabel metal5 106040 -109960 106240 -109760 1 PIX1885_IN
port 1932 n
rlabel metal5 109040 -109960 109240 -109760 1 PIX1886_IN
port 1933 n
rlabel metal5 112040 -109960 112240 -109760 1 PIX1887_IN
port 1934 n
rlabel metal5 115040 -109960 115240 -109760 1 PIX1888_IN
port 1935 n
rlabel metal5 118040 -109960 118240 -109760 1 PIX1889_IN
port 1936 n
rlabel metal5 121040 -109960 121240 -109760 1 PIX1890_IN
port 1937 n
rlabel metal5 124040 -109960 124240 -109760 1 PIX1891_IN
port 1938 n
rlabel metal5 127040 -109960 127240 -109760 1 PIX1892_IN
port 1939 n
rlabel metal5 130040 -109960 130240 -109760 1 PIX1893_IN
port 1940 n
rlabel metal5 133040 -109960 133240 -109760 1 PIX1894_IN
port 1941 n
rlabel metal5 136040 -109960 136240 -109760 1 PIX1895_IN
port 1942 n
rlabel metal5 139040 -109960 139240 -109760 1 PIX1896_IN
port 1943 n
rlabel metal5 142040 -109960 142240 -109760 1 PIX1897_IN
port 1944 n
rlabel metal5 145040 -109960 145240 -109760 1 PIX1898_IN
port 1945 n
rlabel metal5 148040 -109960 148240 -109760 1 PIX1899_IN
port 1946 n
rlabel metal5 1040 -112960 1240 -112760 1 PIX1900_IN
port 1947 n
rlabel metal2 -3000 -112520 -3000 -112430 3 ROW_SEL38
port 1948 e
rlabel metal5 4040 -112960 4240 -112760 1 PIX1901_IN
port 1949 n
rlabel metal5 7040 -112960 7240 -112760 1 PIX1902_IN
port 1950 n
rlabel metal5 10040 -112960 10240 -112760 1 PIX1903_IN
port 1951 n
rlabel metal5 13040 -112960 13240 -112760 1 PIX1904_IN
port 1952 n
rlabel metal5 16040 -112960 16240 -112760 1 PIX1905_IN
port 1953 n
rlabel metal5 19040 -112960 19240 -112760 1 PIX1906_IN
port 1954 n
rlabel metal5 22040 -112960 22240 -112760 1 PIX1907_IN
port 1955 n
rlabel metal5 25040 -112960 25240 -112760 1 PIX1908_IN
port 1956 n
rlabel metal5 28040 -112960 28240 -112760 1 PIX1909_IN
port 1957 n
rlabel metal5 31040 -112960 31240 -112760 1 PIX1910_IN
port 1958 n
rlabel metal5 34040 -112960 34240 -112760 1 PIX1911_IN
port 1959 n
rlabel metal5 37040 -112960 37240 -112760 1 PIX1912_IN
port 1960 n
rlabel metal5 40040 -112960 40240 -112760 1 PIX1913_IN
port 1961 n
rlabel metal5 43040 -112960 43240 -112760 1 PIX1914_IN
port 1962 n
rlabel metal5 46040 -112960 46240 -112760 1 PIX1915_IN
port 1963 n
rlabel metal5 49040 -112960 49240 -112760 1 PIX1916_IN
port 1964 n
rlabel metal5 52040 -112960 52240 -112760 1 PIX1917_IN
port 1965 n
rlabel metal5 55040 -112960 55240 -112760 1 PIX1918_IN
port 1966 n
rlabel metal5 58040 -112960 58240 -112760 1 PIX1919_IN
port 1967 n
rlabel metal5 61040 -112960 61240 -112760 1 PIX1920_IN
port 1968 n
rlabel metal5 64040 -112960 64240 -112760 1 PIX1921_IN
port 1969 n
rlabel metal5 67040 -112960 67240 -112760 1 PIX1922_IN
port 1970 n
rlabel metal5 70040 -112960 70240 -112760 1 PIX1923_IN
port 1971 n
rlabel metal5 73040 -112960 73240 -112760 1 PIX1924_IN
port 1972 n
rlabel metal5 76040 -112960 76240 -112760 1 PIX1925_IN
port 1973 n
rlabel metal5 79040 -112960 79240 -112760 1 PIX1926_IN
port 1974 n
rlabel metal5 82040 -112960 82240 -112760 1 PIX1927_IN
port 1975 n
rlabel metal5 85040 -112960 85240 -112760 1 PIX1928_IN
port 1976 n
rlabel metal5 88040 -112960 88240 -112760 1 PIX1929_IN
port 1977 n
rlabel metal5 91040 -112960 91240 -112760 1 PIX1930_IN
port 1978 n
rlabel metal5 94040 -112960 94240 -112760 1 PIX1931_IN
port 1979 n
rlabel metal5 97040 -112960 97240 -112760 1 PIX1932_IN
port 1980 n
rlabel metal5 100040 -112960 100240 -112760 1 PIX1933_IN
port 1981 n
rlabel metal5 103040 -112960 103240 -112760 1 PIX1934_IN
port 1982 n
rlabel metal5 106040 -112960 106240 -112760 1 PIX1935_IN
port 1983 n
rlabel metal5 109040 -112960 109240 -112760 1 PIX1936_IN
port 1984 n
rlabel metal5 112040 -112960 112240 -112760 1 PIX1937_IN
port 1985 n
rlabel metal5 115040 -112960 115240 -112760 1 PIX1938_IN
port 1986 n
rlabel metal5 118040 -112960 118240 -112760 1 PIX1939_IN
port 1987 n
rlabel metal5 121040 -112960 121240 -112760 1 PIX1940_IN
port 1988 n
rlabel metal5 124040 -112960 124240 -112760 1 PIX1941_IN
port 1989 n
rlabel metal5 127040 -112960 127240 -112760 1 PIX1942_IN
port 1990 n
rlabel metal5 130040 -112960 130240 -112760 1 PIX1943_IN
port 1991 n
rlabel metal5 133040 -112960 133240 -112760 1 PIX1944_IN
port 1992 n
rlabel metal5 136040 -112960 136240 -112760 1 PIX1945_IN
port 1993 n
rlabel metal5 139040 -112960 139240 -112760 1 PIX1946_IN
port 1994 n
rlabel metal5 142040 -112960 142240 -112760 1 PIX1947_IN
port 1995 n
rlabel metal5 145040 -112960 145240 -112760 1 PIX1948_IN
port 1996 n
rlabel metal5 148040 -112960 148240 -112760 1 PIX1949_IN
port 1997 n
rlabel metal5 1040 -115960 1240 -115760 1 PIX1950_IN
port 1998 n
rlabel metal2 -3000 -115520 -3000 -115430 3 ROW_SEL39
port 1999 e
rlabel metal5 4040 -115960 4240 -115760 1 PIX1951_IN
port 2000 n
rlabel metal5 7040 -115960 7240 -115760 1 PIX1952_IN
port 2001 n
rlabel metal5 10040 -115960 10240 -115760 1 PIX1953_IN
port 2002 n
rlabel metal5 13040 -115960 13240 -115760 1 PIX1954_IN
port 2003 n
rlabel metal5 16040 -115960 16240 -115760 1 PIX1955_IN
port 2004 n
rlabel metal5 19040 -115960 19240 -115760 1 PIX1956_IN
port 2005 n
rlabel metal5 22040 -115960 22240 -115760 1 PIX1957_IN
port 2006 n
rlabel metal5 25040 -115960 25240 -115760 1 PIX1958_IN
port 2007 n
rlabel metal5 28040 -115960 28240 -115760 1 PIX1959_IN
port 2008 n
rlabel metal5 31040 -115960 31240 -115760 1 PIX1960_IN
port 2009 n
rlabel metal5 34040 -115960 34240 -115760 1 PIX1961_IN
port 2010 n
rlabel metal5 37040 -115960 37240 -115760 1 PIX1962_IN
port 2011 n
rlabel metal5 40040 -115960 40240 -115760 1 PIX1963_IN
port 2012 n
rlabel metal5 43040 -115960 43240 -115760 1 PIX1964_IN
port 2013 n
rlabel metal5 46040 -115960 46240 -115760 1 PIX1965_IN
port 2014 n
rlabel metal5 49040 -115960 49240 -115760 1 PIX1966_IN
port 2015 n
rlabel metal5 52040 -115960 52240 -115760 1 PIX1967_IN
port 2016 n
rlabel metal5 55040 -115960 55240 -115760 1 PIX1968_IN
port 2017 n
rlabel metal5 58040 -115960 58240 -115760 1 PIX1969_IN
port 2018 n
rlabel metal5 61040 -115960 61240 -115760 1 PIX1970_IN
port 2019 n
rlabel metal5 64040 -115960 64240 -115760 1 PIX1971_IN
port 2020 n
rlabel metal5 67040 -115960 67240 -115760 1 PIX1972_IN
port 2021 n
rlabel metal5 70040 -115960 70240 -115760 1 PIX1973_IN
port 2022 n
rlabel metal5 73040 -115960 73240 -115760 1 PIX1974_IN
port 2023 n
rlabel metal5 76040 -115960 76240 -115760 1 PIX1975_IN
port 2024 n
rlabel metal5 79040 -115960 79240 -115760 1 PIX1976_IN
port 2025 n
rlabel metal5 82040 -115960 82240 -115760 1 PIX1977_IN
port 2026 n
rlabel metal5 85040 -115960 85240 -115760 1 PIX1978_IN
port 2027 n
rlabel metal5 88040 -115960 88240 -115760 1 PIX1979_IN
port 2028 n
rlabel metal5 91040 -115960 91240 -115760 1 PIX1980_IN
port 2029 n
rlabel metal5 94040 -115960 94240 -115760 1 PIX1981_IN
port 2030 n
rlabel metal5 97040 -115960 97240 -115760 1 PIX1982_IN
port 2031 n
rlabel metal5 100040 -115960 100240 -115760 1 PIX1983_IN
port 2032 n
rlabel metal5 103040 -115960 103240 -115760 1 PIX1984_IN
port 2033 n
rlabel metal5 106040 -115960 106240 -115760 1 PIX1985_IN
port 2034 n
rlabel metal5 109040 -115960 109240 -115760 1 PIX1986_IN
port 2035 n
rlabel metal5 112040 -115960 112240 -115760 1 PIX1987_IN
port 2036 n
rlabel metal5 115040 -115960 115240 -115760 1 PIX1988_IN
port 2037 n
rlabel metal5 118040 -115960 118240 -115760 1 PIX1989_IN
port 2038 n
rlabel metal5 121040 -115960 121240 -115760 1 PIX1990_IN
port 2039 n
rlabel metal5 124040 -115960 124240 -115760 1 PIX1991_IN
port 2040 n
rlabel metal5 127040 -115960 127240 -115760 1 PIX1992_IN
port 2041 n
rlabel metal5 130040 -115960 130240 -115760 1 PIX1993_IN
port 2042 n
rlabel metal5 133040 -115960 133240 -115760 1 PIX1994_IN
port 2043 n
rlabel metal5 136040 -115960 136240 -115760 1 PIX1995_IN
port 2044 n
rlabel metal5 139040 -115960 139240 -115760 1 PIX1996_IN
port 2045 n
rlabel metal5 142040 -115960 142240 -115760 1 PIX1997_IN
port 2046 n
rlabel metal5 145040 -115960 145240 -115760 1 PIX1998_IN
port 2047 n
rlabel metal5 148040 -115960 148240 -115760 1 PIX1999_IN
port 2048 n
rlabel metal5 1040 -118960 1240 -118760 1 PIX2000_IN
port 2049 n
rlabel metal2 -3000 -118520 -3000 -118430 3 ROW_SEL40
port 2050 e
rlabel metal5 4040 -118960 4240 -118760 1 PIX2001_IN
port 2051 n
rlabel metal5 7040 -118960 7240 -118760 1 PIX2002_IN
port 2052 n
rlabel metal5 10040 -118960 10240 -118760 1 PIX2003_IN
port 2053 n
rlabel metal5 13040 -118960 13240 -118760 1 PIX2004_IN
port 2054 n
rlabel metal5 16040 -118960 16240 -118760 1 PIX2005_IN
port 2055 n
rlabel metal5 19040 -118960 19240 -118760 1 PIX2006_IN
port 2056 n
rlabel metal5 22040 -118960 22240 -118760 1 PIX2007_IN
port 2057 n
rlabel metal5 25040 -118960 25240 -118760 1 PIX2008_IN
port 2058 n
rlabel metal5 28040 -118960 28240 -118760 1 PIX2009_IN
port 2059 n
rlabel metal5 31040 -118960 31240 -118760 1 PIX2010_IN
port 2060 n
rlabel metal5 34040 -118960 34240 -118760 1 PIX2011_IN
port 2061 n
rlabel metal5 37040 -118960 37240 -118760 1 PIX2012_IN
port 2062 n
rlabel metal5 40040 -118960 40240 -118760 1 PIX2013_IN
port 2063 n
rlabel metal5 43040 -118960 43240 -118760 1 PIX2014_IN
port 2064 n
rlabel metal5 46040 -118960 46240 -118760 1 PIX2015_IN
port 2065 n
rlabel metal5 49040 -118960 49240 -118760 1 PIX2016_IN
port 2066 n
rlabel metal5 52040 -118960 52240 -118760 1 PIX2017_IN
port 2067 n
rlabel metal5 55040 -118960 55240 -118760 1 PIX2018_IN
port 2068 n
rlabel metal5 58040 -118960 58240 -118760 1 PIX2019_IN
port 2069 n
rlabel metal5 61040 -118960 61240 -118760 1 PIX2020_IN
port 2070 n
rlabel metal5 64040 -118960 64240 -118760 1 PIX2021_IN
port 2071 n
rlabel metal5 67040 -118960 67240 -118760 1 PIX2022_IN
port 2072 n
rlabel metal5 70040 -118960 70240 -118760 1 PIX2023_IN
port 2073 n
rlabel metal5 73040 -118960 73240 -118760 1 PIX2024_IN
port 2074 n
rlabel metal5 76040 -118960 76240 -118760 1 PIX2025_IN
port 2075 n
rlabel metal5 79040 -118960 79240 -118760 1 PIX2026_IN
port 2076 n
rlabel metal5 82040 -118960 82240 -118760 1 PIX2027_IN
port 2077 n
rlabel metal5 85040 -118960 85240 -118760 1 PIX2028_IN
port 2078 n
rlabel metal5 88040 -118960 88240 -118760 1 PIX2029_IN
port 2079 n
rlabel metal5 91040 -118960 91240 -118760 1 PIX2030_IN
port 2080 n
rlabel metal5 94040 -118960 94240 -118760 1 PIX2031_IN
port 2081 n
rlabel metal5 97040 -118960 97240 -118760 1 PIX2032_IN
port 2082 n
rlabel metal5 100040 -118960 100240 -118760 1 PIX2033_IN
port 2083 n
rlabel metal5 103040 -118960 103240 -118760 1 PIX2034_IN
port 2084 n
rlabel metal5 106040 -118960 106240 -118760 1 PIX2035_IN
port 2085 n
rlabel metal5 109040 -118960 109240 -118760 1 PIX2036_IN
port 2086 n
rlabel metal5 112040 -118960 112240 -118760 1 PIX2037_IN
port 2087 n
rlabel metal5 115040 -118960 115240 -118760 1 PIX2038_IN
port 2088 n
rlabel metal5 118040 -118960 118240 -118760 1 PIX2039_IN
port 2089 n
rlabel metal5 121040 -118960 121240 -118760 1 PIX2040_IN
port 2090 n
rlabel metal5 124040 -118960 124240 -118760 1 PIX2041_IN
port 2091 n
rlabel metal5 127040 -118960 127240 -118760 1 PIX2042_IN
port 2092 n
rlabel metal5 130040 -118960 130240 -118760 1 PIX2043_IN
port 2093 n
rlabel metal5 133040 -118960 133240 -118760 1 PIX2044_IN
port 2094 n
rlabel metal5 136040 -118960 136240 -118760 1 PIX2045_IN
port 2095 n
rlabel metal5 139040 -118960 139240 -118760 1 PIX2046_IN
port 2096 n
rlabel metal5 142040 -118960 142240 -118760 1 PIX2047_IN
port 2097 n
rlabel metal5 145040 -118960 145240 -118760 1 PIX2048_IN
port 2098 n
rlabel metal5 148040 -118960 148240 -118760 1 PIX2049_IN
port 2099 n
rlabel metal5 1040 -121960 1240 -121760 1 PIX2050_IN
port 2100 n
rlabel metal2 -3000 -121520 -3000 -121430 3 ROW_SEL41
port 2101 e
rlabel metal5 4040 -121960 4240 -121760 1 PIX2051_IN
port 2102 n
rlabel metal5 7040 -121960 7240 -121760 1 PIX2052_IN
port 2103 n
rlabel metal5 10040 -121960 10240 -121760 1 PIX2053_IN
port 2104 n
rlabel metal5 13040 -121960 13240 -121760 1 PIX2054_IN
port 2105 n
rlabel metal5 16040 -121960 16240 -121760 1 PIX2055_IN
port 2106 n
rlabel metal5 19040 -121960 19240 -121760 1 PIX2056_IN
port 2107 n
rlabel metal5 22040 -121960 22240 -121760 1 PIX2057_IN
port 2108 n
rlabel metal5 25040 -121960 25240 -121760 1 PIX2058_IN
port 2109 n
rlabel metal5 28040 -121960 28240 -121760 1 PIX2059_IN
port 2110 n
rlabel metal5 31040 -121960 31240 -121760 1 PIX2060_IN
port 2111 n
rlabel metal5 34040 -121960 34240 -121760 1 PIX2061_IN
port 2112 n
rlabel metal5 37040 -121960 37240 -121760 1 PIX2062_IN
port 2113 n
rlabel metal5 40040 -121960 40240 -121760 1 PIX2063_IN
port 2114 n
rlabel metal5 43040 -121960 43240 -121760 1 PIX2064_IN
port 2115 n
rlabel metal5 46040 -121960 46240 -121760 1 PIX2065_IN
port 2116 n
rlabel metal5 49040 -121960 49240 -121760 1 PIX2066_IN
port 2117 n
rlabel metal5 52040 -121960 52240 -121760 1 PIX2067_IN
port 2118 n
rlabel metal5 55040 -121960 55240 -121760 1 PIX2068_IN
port 2119 n
rlabel metal5 58040 -121960 58240 -121760 1 PIX2069_IN
port 2120 n
rlabel metal5 61040 -121960 61240 -121760 1 PIX2070_IN
port 2121 n
rlabel metal5 64040 -121960 64240 -121760 1 PIX2071_IN
port 2122 n
rlabel metal5 67040 -121960 67240 -121760 1 PIX2072_IN
port 2123 n
rlabel metal5 70040 -121960 70240 -121760 1 PIX2073_IN
port 2124 n
rlabel metal5 73040 -121960 73240 -121760 1 PIX2074_IN
port 2125 n
rlabel metal5 76040 -121960 76240 -121760 1 PIX2075_IN
port 2126 n
rlabel metal5 79040 -121960 79240 -121760 1 PIX2076_IN
port 2127 n
rlabel metal5 82040 -121960 82240 -121760 1 PIX2077_IN
port 2128 n
rlabel metal5 85040 -121960 85240 -121760 1 PIX2078_IN
port 2129 n
rlabel metal5 88040 -121960 88240 -121760 1 PIX2079_IN
port 2130 n
rlabel metal5 91040 -121960 91240 -121760 1 PIX2080_IN
port 2131 n
rlabel metal5 94040 -121960 94240 -121760 1 PIX2081_IN
port 2132 n
rlabel metal5 97040 -121960 97240 -121760 1 PIX2082_IN
port 2133 n
rlabel metal5 100040 -121960 100240 -121760 1 PIX2083_IN
port 2134 n
rlabel metal5 103040 -121960 103240 -121760 1 PIX2084_IN
port 2135 n
rlabel metal5 106040 -121960 106240 -121760 1 PIX2085_IN
port 2136 n
rlabel metal5 109040 -121960 109240 -121760 1 PIX2086_IN
port 2137 n
rlabel metal5 112040 -121960 112240 -121760 1 PIX2087_IN
port 2138 n
rlabel metal5 115040 -121960 115240 -121760 1 PIX2088_IN
port 2139 n
rlabel metal5 118040 -121960 118240 -121760 1 PIX2089_IN
port 2140 n
rlabel metal5 121040 -121960 121240 -121760 1 PIX2090_IN
port 2141 n
rlabel metal5 124040 -121960 124240 -121760 1 PIX2091_IN
port 2142 n
rlabel metal5 127040 -121960 127240 -121760 1 PIX2092_IN
port 2143 n
rlabel metal5 130040 -121960 130240 -121760 1 PIX2093_IN
port 2144 n
rlabel metal5 133040 -121960 133240 -121760 1 PIX2094_IN
port 2145 n
rlabel metal5 136040 -121960 136240 -121760 1 PIX2095_IN
port 2146 n
rlabel metal5 139040 -121960 139240 -121760 1 PIX2096_IN
port 2147 n
rlabel metal5 142040 -121960 142240 -121760 1 PIX2097_IN
port 2148 n
rlabel metal5 145040 -121960 145240 -121760 1 PIX2098_IN
port 2149 n
rlabel metal5 148040 -121960 148240 -121760 1 PIX2099_IN
port 2150 n
rlabel metal5 1040 -124960 1240 -124760 1 PIX2100_IN
port 2151 n
rlabel metal2 -3000 -124520 -3000 -124430 3 ROW_SEL42
port 2152 e
rlabel metal5 4040 -124960 4240 -124760 1 PIX2101_IN
port 2153 n
rlabel metal5 7040 -124960 7240 -124760 1 PIX2102_IN
port 2154 n
rlabel metal5 10040 -124960 10240 -124760 1 PIX2103_IN
port 2155 n
rlabel metal5 13040 -124960 13240 -124760 1 PIX2104_IN
port 2156 n
rlabel metal5 16040 -124960 16240 -124760 1 PIX2105_IN
port 2157 n
rlabel metal5 19040 -124960 19240 -124760 1 PIX2106_IN
port 2158 n
rlabel metal5 22040 -124960 22240 -124760 1 PIX2107_IN
port 2159 n
rlabel metal5 25040 -124960 25240 -124760 1 PIX2108_IN
port 2160 n
rlabel metal5 28040 -124960 28240 -124760 1 PIX2109_IN
port 2161 n
rlabel metal5 31040 -124960 31240 -124760 1 PIX2110_IN
port 2162 n
rlabel metal5 34040 -124960 34240 -124760 1 PIX2111_IN
port 2163 n
rlabel metal5 37040 -124960 37240 -124760 1 PIX2112_IN
port 2164 n
rlabel metal5 40040 -124960 40240 -124760 1 PIX2113_IN
port 2165 n
rlabel metal5 43040 -124960 43240 -124760 1 PIX2114_IN
port 2166 n
rlabel metal5 46040 -124960 46240 -124760 1 PIX2115_IN
port 2167 n
rlabel metal5 49040 -124960 49240 -124760 1 PIX2116_IN
port 2168 n
rlabel metal5 52040 -124960 52240 -124760 1 PIX2117_IN
port 2169 n
rlabel metal5 55040 -124960 55240 -124760 1 PIX2118_IN
port 2170 n
rlabel metal5 58040 -124960 58240 -124760 1 PIX2119_IN
port 2171 n
rlabel metal5 61040 -124960 61240 -124760 1 PIX2120_IN
port 2172 n
rlabel metal5 64040 -124960 64240 -124760 1 PIX2121_IN
port 2173 n
rlabel metal5 67040 -124960 67240 -124760 1 PIX2122_IN
port 2174 n
rlabel metal5 70040 -124960 70240 -124760 1 PIX2123_IN
port 2175 n
rlabel metal5 73040 -124960 73240 -124760 1 PIX2124_IN
port 2176 n
rlabel metal5 76040 -124960 76240 -124760 1 PIX2125_IN
port 2177 n
rlabel metal5 79040 -124960 79240 -124760 1 PIX2126_IN
port 2178 n
rlabel metal5 82040 -124960 82240 -124760 1 PIX2127_IN
port 2179 n
rlabel metal5 85040 -124960 85240 -124760 1 PIX2128_IN
port 2180 n
rlabel metal5 88040 -124960 88240 -124760 1 PIX2129_IN
port 2181 n
rlabel metal5 91040 -124960 91240 -124760 1 PIX2130_IN
port 2182 n
rlabel metal5 94040 -124960 94240 -124760 1 PIX2131_IN
port 2183 n
rlabel metal5 97040 -124960 97240 -124760 1 PIX2132_IN
port 2184 n
rlabel metal5 100040 -124960 100240 -124760 1 PIX2133_IN
port 2185 n
rlabel metal5 103040 -124960 103240 -124760 1 PIX2134_IN
port 2186 n
rlabel metal5 106040 -124960 106240 -124760 1 PIX2135_IN
port 2187 n
rlabel metal5 109040 -124960 109240 -124760 1 PIX2136_IN
port 2188 n
rlabel metal5 112040 -124960 112240 -124760 1 PIX2137_IN
port 2189 n
rlabel metal5 115040 -124960 115240 -124760 1 PIX2138_IN
port 2190 n
rlabel metal5 118040 -124960 118240 -124760 1 PIX2139_IN
port 2191 n
rlabel metal5 121040 -124960 121240 -124760 1 PIX2140_IN
port 2192 n
rlabel metal5 124040 -124960 124240 -124760 1 PIX2141_IN
port 2193 n
rlabel metal5 127040 -124960 127240 -124760 1 PIX2142_IN
port 2194 n
rlabel metal5 130040 -124960 130240 -124760 1 PIX2143_IN
port 2195 n
rlabel metal5 133040 -124960 133240 -124760 1 PIX2144_IN
port 2196 n
rlabel metal5 136040 -124960 136240 -124760 1 PIX2145_IN
port 2197 n
rlabel metal5 139040 -124960 139240 -124760 1 PIX2146_IN
port 2198 n
rlabel metal5 142040 -124960 142240 -124760 1 PIX2147_IN
port 2199 n
rlabel metal5 145040 -124960 145240 -124760 1 PIX2148_IN
port 2200 n
rlabel metal5 148040 -124960 148240 -124760 1 PIX2149_IN
port 2201 n
rlabel metal5 1040 -127960 1240 -127760 1 PIX2150_IN
port 2202 n
rlabel metal2 -3000 -127520 -3000 -127430 3 ROW_SEL43
port 2203 e
rlabel metal5 4040 -127960 4240 -127760 1 PIX2151_IN
port 2204 n
rlabel metal5 7040 -127960 7240 -127760 1 PIX2152_IN
port 2205 n
rlabel metal5 10040 -127960 10240 -127760 1 PIX2153_IN
port 2206 n
rlabel metal5 13040 -127960 13240 -127760 1 PIX2154_IN
port 2207 n
rlabel metal5 16040 -127960 16240 -127760 1 PIX2155_IN
port 2208 n
rlabel metal5 19040 -127960 19240 -127760 1 PIX2156_IN
port 2209 n
rlabel metal5 22040 -127960 22240 -127760 1 PIX2157_IN
port 2210 n
rlabel metal5 25040 -127960 25240 -127760 1 PIX2158_IN
port 2211 n
rlabel metal5 28040 -127960 28240 -127760 1 PIX2159_IN
port 2212 n
rlabel metal5 31040 -127960 31240 -127760 1 PIX2160_IN
port 2213 n
rlabel metal5 34040 -127960 34240 -127760 1 PIX2161_IN
port 2214 n
rlabel metal5 37040 -127960 37240 -127760 1 PIX2162_IN
port 2215 n
rlabel metal5 40040 -127960 40240 -127760 1 PIX2163_IN
port 2216 n
rlabel metal5 43040 -127960 43240 -127760 1 PIX2164_IN
port 2217 n
rlabel metal5 46040 -127960 46240 -127760 1 PIX2165_IN
port 2218 n
rlabel metal5 49040 -127960 49240 -127760 1 PIX2166_IN
port 2219 n
rlabel metal5 52040 -127960 52240 -127760 1 PIX2167_IN
port 2220 n
rlabel metal5 55040 -127960 55240 -127760 1 PIX2168_IN
port 2221 n
rlabel metal5 58040 -127960 58240 -127760 1 PIX2169_IN
port 2222 n
rlabel metal5 61040 -127960 61240 -127760 1 PIX2170_IN
port 2223 n
rlabel metal5 64040 -127960 64240 -127760 1 PIX2171_IN
port 2224 n
rlabel metal5 67040 -127960 67240 -127760 1 PIX2172_IN
port 2225 n
rlabel metal5 70040 -127960 70240 -127760 1 PIX2173_IN
port 2226 n
rlabel metal5 73040 -127960 73240 -127760 1 PIX2174_IN
port 2227 n
rlabel metal5 76040 -127960 76240 -127760 1 PIX2175_IN
port 2228 n
rlabel metal5 79040 -127960 79240 -127760 1 PIX2176_IN
port 2229 n
rlabel metal5 82040 -127960 82240 -127760 1 PIX2177_IN
port 2230 n
rlabel metal5 85040 -127960 85240 -127760 1 PIX2178_IN
port 2231 n
rlabel metal5 88040 -127960 88240 -127760 1 PIX2179_IN
port 2232 n
rlabel metal5 91040 -127960 91240 -127760 1 PIX2180_IN
port 2233 n
rlabel metal5 94040 -127960 94240 -127760 1 PIX2181_IN
port 2234 n
rlabel metal5 97040 -127960 97240 -127760 1 PIX2182_IN
port 2235 n
rlabel metal5 100040 -127960 100240 -127760 1 PIX2183_IN
port 2236 n
rlabel metal5 103040 -127960 103240 -127760 1 PIX2184_IN
port 2237 n
rlabel metal5 106040 -127960 106240 -127760 1 PIX2185_IN
port 2238 n
rlabel metal5 109040 -127960 109240 -127760 1 PIX2186_IN
port 2239 n
rlabel metal5 112040 -127960 112240 -127760 1 PIX2187_IN
port 2240 n
rlabel metal5 115040 -127960 115240 -127760 1 PIX2188_IN
port 2241 n
rlabel metal5 118040 -127960 118240 -127760 1 PIX2189_IN
port 2242 n
rlabel metal5 121040 -127960 121240 -127760 1 PIX2190_IN
port 2243 n
rlabel metal5 124040 -127960 124240 -127760 1 PIX2191_IN
port 2244 n
rlabel metal5 127040 -127960 127240 -127760 1 PIX2192_IN
port 2245 n
rlabel metal5 130040 -127960 130240 -127760 1 PIX2193_IN
port 2246 n
rlabel metal5 133040 -127960 133240 -127760 1 PIX2194_IN
port 2247 n
rlabel metal5 136040 -127960 136240 -127760 1 PIX2195_IN
port 2248 n
rlabel metal5 139040 -127960 139240 -127760 1 PIX2196_IN
port 2249 n
rlabel metal5 142040 -127960 142240 -127760 1 PIX2197_IN
port 2250 n
rlabel metal5 145040 -127960 145240 -127760 1 PIX2198_IN
port 2251 n
rlabel metal5 148040 -127960 148240 -127760 1 PIX2199_IN
port 2252 n
rlabel metal5 1040 -130960 1240 -130760 1 PIX2200_IN
port 2253 n
rlabel metal2 -3000 -130520 -3000 -130430 3 ROW_SEL44
port 2254 e
rlabel metal5 4040 -130960 4240 -130760 1 PIX2201_IN
port 2255 n
rlabel metal5 7040 -130960 7240 -130760 1 PIX2202_IN
port 2256 n
rlabel metal5 10040 -130960 10240 -130760 1 PIX2203_IN
port 2257 n
rlabel metal5 13040 -130960 13240 -130760 1 PIX2204_IN
port 2258 n
rlabel metal5 16040 -130960 16240 -130760 1 PIX2205_IN
port 2259 n
rlabel metal5 19040 -130960 19240 -130760 1 PIX2206_IN
port 2260 n
rlabel metal5 22040 -130960 22240 -130760 1 PIX2207_IN
port 2261 n
rlabel metal5 25040 -130960 25240 -130760 1 PIX2208_IN
port 2262 n
rlabel metal5 28040 -130960 28240 -130760 1 PIX2209_IN
port 2263 n
rlabel metal5 31040 -130960 31240 -130760 1 PIX2210_IN
port 2264 n
rlabel metal5 34040 -130960 34240 -130760 1 PIX2211_IN
port 2265 n
rlabel metal5 37040 -130960 37240 -130760 1 PIX2212_IN
port 2266 n
rlabel metal5 40040 -130960 40240 -130760 1 PIX2213_IN
port 2267 n
rlabel metal5 43040 -130960 43240 -130760 1 PIX2214_IN
port 2268 n
rlabel metal5 46040 -130960 46240 -130760 1 PIX2215_IN
port 2269 n
rlabel metal5 49040 -130960 49240 -130760 1 PIX2216_IN
port 2270 n
rlabel metal5 52040 -130960 52240 -130760 1 PIX2217_IN
port 2271 n
rlabel metal5 55040 -130960 55240 -130760 1 PIX2218_IN
port 2272 n
rlabel metal5 58040 -130960 58240 -130760 1 PIX2219_IN
port 2273 n
rlabel metal5 61040 -130960 61240 -130760 1 PIX2220_IN
port 2274 n
rlabel metal5 64040 -130960 64240 -130760 1 PIX2221_IN
port 2275 n
rlabel metal5 67040 -130960 67240 -130760 1 PIX2222_IN
port 2276 n
rlabel metal5 70040 -130960 70240 -130760 1 PIX2223_IN
port 2277 n
rlabel metal5 73040 -130960 73240 -130760 1 PIX2224_IN
port 2278 n
rlabel metal5 76040 -130960 76240 -130760 1 PIX2225_IN
port 2279 n
rlabel metal5 79040 -130960 79240 -130760 1 PIX2226_IN
port 2280 n
rlabel metal5 82040 -130960 82240 -130760 1 PIX2227_IN
port 2281 n
rlabel metal5 85040 -130960 85240 -130760 1 PIX2228_IN
port 2282 n
rlabel metal5 88040 -130960 88240 -130760 1 PIX2229_IN
port 2283 n
rlabel metal5 91040 -130960 91240 -130760 1 PIX2230_IN
port 2284 n
rlabel metal5 94040 -130960 94240 -130760 1 PIX2231_IN
port 2285 n
rlabel metal5 97040 -130960 97240 -130760 1 PIX2232_IN
port 2286 n
rlabel metal5 100040 -130960 100240 -130760 1 PIX2233_IN
port 2287 n
rlabel metal5 103040 -130960 103240 -130760 1 PIX2234_IN
port 2288 n
rlabel metal5 106040 -130960 106240 -130760 1 PIX2235_IN
port 2289 n
rlabel metal5 109040 -130960 109240 -130760 1 PIX2236_IN
port 2290 n
rlabel metal5 112040 -130960 112240 -130760 1 PIX2237_IN
port 2291 n
rlabel metal5 115040 -130960 115240 -130760 1 PIX2238_IN
port 2292 n
rlabel metal5 118040 -130960 118240 -130760 1 PIX2239_IN
port 2293 n
rlabel metal5 121040 -130960 121240 -130760 1 PIX2240_IN
port 2294 n
rlabel metal5 124040 -130960 124240 -130760 1 PIX2241_IN
port 2295 n
rlabel metal5 127040 -130960 127240 -130760 1 PIX2242_IN
port 2296 n
rlabel metal5 130040 -130960 130240 -130760 1 PIX2243_IN
port 2297 n
rlabel metal5 133040 -130960 133240 -130760 1 PIX2244_IN
port 2298 n
rlabel metal5 136040 -130960 136240 -130760 1 PIX2245_IN
port 2299 n
rlabel metal5 139040 -130960 139240 -130760 1 PIX2246_IN
port 2300 n
rlabel metal5 142040 -130960 142240 -130760 1 PIX2247_IN
port 2301 n
rlabel metal5 145040 -130960 145240 -130760 1 PIX2248_IN
port 2302 n
rlabel metal5 148040 -130960 148240 -130760 1 PIX2249_IN
port 2303 n
rlabel metal5 1040 -133960 1240 -133760 1 PIX2250_IN
port 2304 n
rlabel metal2 -3000 -133520 -3000 -133430 3 ROW_SEL45
port 2305 e
rlabel metal5 4040 -133960 4240 -133760 1 PIX2251_IN
port 2306 n
rlabel metal5 7040 -133960 7240 -133760 1 PIX2252_IN
port 2307 n
rlabel metal5 10040 -133960 10240 -133760 1 PIX2253_IN
port 2308 n
rlabel metal5 13040 -133960 13240 -133760 1 PIX2254_IN
port 2309 n
rlabel metal5 16040 -133960 16240 -133760 1 PIX2255_IN
port 2310 n
rlabel metal5 19040 -133960 19240 -133760 1 PIX2256_IN
port 2311 n
rlabel metal5 22040 -133960 22240 -133760 1 PIX2257_IN
port 2312 n
rlabel metal5 25040 -133960 25240 -133760 1 PIX2258_IN
port 2313 n
rlabel metal5 28040 -133960 28240 -133760 1 PIX2259_IN
port 2314 n
rlabel metal5 31040 -133960 31240 -133760 1 PIX2260_IN
port 2315 n
rlabel metal5 34040 -133960 34240 -133760 1 PIX2261_IN
port 2316 n
rlabel metal5 37040 -133960 37240 -133760 1 PIX2262_IN
port 2317 n
rlabel metal5 40040 -133960 40240 -133760 1 PIX2263_IN
port 2318 n
rlabel metal5 43040 -133960 43240 -133760 1 PIX2264_IN
port 2319 n
rlabel metal5 46040 -133960 46240 -133760 1 PIX2265_IN
port 2320 n
rlabel metal5 49040 -133960 49240 -133760 1 PIX2266_IN
port 2321 n
rlabel metal5 52040 -133960 52240 -133760 1 PIX2267_IN
port 2322 n
rlabel metal5 55040 -133960 55240 -133760 1 PIX2268_IN
port 2323 n
rlabel metal5 58040 -133960 58240 -133760 1 PIX2269_IN
port 2324 n
rlabel metal5 61040 -133960 61240 -133760 1 PIX2270_IN
port 2325 n
rlabel metal5 64040 -133960 64240 -133760 1 PIX2271_IN
port 2326 n
rlabel metal5 67040 -133960 67240 -133760 1 PIX2272_IN
port 2327 n
rlabel metal5 70040 -133960 70240 -133760 1 PIX2273_IN
port 2328 n
rlabel metal5 73040 -133960 73240 -133760 1 PIX2274_IN
port 2329 n
rlabel metal5 76040 -133960 76240 -133760 1 PIX2275_IN
port 2330 n
rlabel metal5 79040 -133960 79240 -133760 1 PIX2276_IN
port 2331 n
rlabel metal5 82040 -133960 82240 -133760 1 PIX2277_IN
port 2332 n
rlabel metal5 85040 -133960 85240 -133760 1 PIX2278_IN
port 2333 n
rlabel metal5 88040 -133960 88240 -133760 1 PIX2279_IN
port 2334 n
rlabel metal5 91040 -133960 91240 -133760 1 PIX2280_IN
port 2335 n
rlabel metal5 94040 -133960 94240 -133760 1 PIX2281_IN
port 2336 n
rlabel metal5 97040 -133960 97240 -133760 1 PIX2282_IN
port 2337 n
rlabel metal5 100040 -133960 100240 -133760 1 PIX2283_IN
port 2338 n
rlabel metal5 103040 -133960 103240 -133760 1 PIX2284_IN
port 2339 n
rlabel metal5 106040 -133960 106240 -133760 1 PIX2285_IN
port 2340 n
rlabel metal5 109040 -133960 109240 -133760 1 PIX2286_IN
port 2341 n
rlabel metal5 112040 -133960 112240 -133760 1 PIX2287_IN
port 2342 n
rlabel metal5 115040 -133960 115240 -133760 1 PIX2288_IN
port 2343 n
rlabel metal5 118040 -133960 118240 -133760 1 PIX2289_IN
port 2344 n
rlabel metal5 121040 -133960 121240 -133760 1 PIX2290_IN
port 2345 n
rlabel metal5 124040 -133960 124240 -133760 1 PIX2291_IN
port 2346 n
rlabel metal5 127040 -133960 127240 -133760 1 PIX2292_IN
port 2347 n
rlabel metal5 130040 -133960 130240 -133760 1 PIX2293_IN
port 2348 n
rlabel metal5 133040 -133960 133240 -133760 1 PIX2294_IN
port 2349 n
rlabel metal5 136040 -133960 136240 -133760 1 PIX2295_IN
port 2350 n
rlabel metal5 139040 -133960 139240 -133760 1 PIX2296_IN
port 2351 n
rlabel metal5 142040 -133960 142240 -133760 1 PIX2297_IN
port 2352 n
rlabel metal5 145040 -133960 145240 -133760 1 PIX2298_IN
port 2353 n
rlabel metal5 148040 -133960 148240 -133760 1 PIX2299_IN
port 2354 n
rlabel metal5 1040 -136960 1240 -136760 1 PIX2300_IN
port 2355 n
rlabel metal2 -3000 -136520 -3000 -136430 3 ROW_SEL46
port 2356 e
rlabel metal5 4040 -136960 4240 -136760 1 PIX2301_IN
port 2357 n
rlabel metal5 7040 -136960 7240 -136760 1 PIX2302_IN
port 2358 n
rlabel metal5 10040 -136960 10240 -136760 1 PIX2303_IN
port 2359 n
rlabel metal5 13040 -136960 13240 -136760 1 PIX2304_IN
port 2360 n
rlabel metal5 16040 -136960 16240 -136760 1 PIX2305_IN
port 2361 n
rlabel metal5 19040 -136960 19240 -136760 1 PIX2306_IN
port 2362 n
rlabel metal5 22040 -136960 22240 -136760 1 PIX2307_IN
port 2363 n
rlabel metal5 25040 -136960 25240 -136760 1 PIX2308_IN
port 2364 n
rlabel metal5 28040 -136960 28240 -136760 1 PIX2309_IN
port 2365 n
rlabel metal5 31040 -136960 31240 -136760 1 PIX2310_IN
port 2366 n
rlabel metal5 34040 -136960 34240 -136760 1 PIX2311_IN
port 2367 n
rlabel metal5 37040 -136960 37240 -136760 1 PIX2312_IN
port 2368 n
rlabel metal5 40040 -136960 40240 -136760 1 PIX2313_IN
port 2369 n
rlabel metal5 43040 -136960 43240 -136760 1 PIX2314_IN
port 2370 n
rlabel metal5 46040 -136960 46240 -136760 1 PIX2315_IN
port 2371 n
rlabel metal5 49040 -136960 49240 -136760 1 PIX2316_IN
port 2372 n
rlabel metal5 52040 -136960 52240 -136760 1 PIX2317_IN
port 2373 n
rlabel metal5 55040 -136960 55240 -136760 1 PIX2318_IN
port 2374 n
rlabel metal5 58040 -136960 58240 -136760 1 PIX2319_IN
port 2375 n
rlabel metal5 61040 -136960 61240 -136760 1 PIX2320_IN
port 2376 n
rlabel metal5 64040 -136960 64240 -136760 1 PIX2321_IN
port 2377 n
rlabel metal5 67040 -136960 67240 -136760 1 PIX2322_IN
port 2378 n
rlabel metal5 70040 -136960 70240 -136760 1 PIX2323_IN
port 2379 n
rlabel metal5 73040 -136960 73240 -136760 1 PIX2324_IN
port 2380 n
rlabel metal5 76040 -136960 76240 -136760 1 PIX2325_IN
port 2381 n
rlabel metal5 79040 -136960 79240 -136760 1 PIX2326_IN
port 2382 n
rlabel metal5 82040 -136960 82240 -136760 1 PIX2327_IN
port 2383 n
rlabel metal5 85040 -136960 85240 -136760 1 PIX2328_IN
port 2384 n
rlabel metal5 88040 -136960 88240 -136760 1 PIX2329_IN
port 2385 n
rlabel metal5 91040 -136960 91240 -136760 1 PIX2330_IN
port 2386 n
rlabel metal5 94040 -136960 94240 -136760 1 PIX2331_IN
port 2387 n
rlabel metal5 97040 -136960 97240 -136760 1 PIX2332_IN
port 2388 n
rlabel metal5 100040 -136960 100240 -136760 1 PIX2333_IN
port 2389 n
rlabel metal5 103040 -136960 103240 -136760 1 PIX2334_IN
port 2390 n
rlabel metal5 106040 -136960 106240 -136760 1 PIX2335_IN
port 2391 n
rlabel metal5 109040 -136960 109240 -136760 1 PIX2336_IN
port 2392 n
rlabel metal5 112040 -136960 112240 -136760 1 PIX2337_IN
port 2393 n
rlabel metal5 115040 -136960 115240 -136760 1 PIX2338_IN
port 2394 n
rlabel metal5 118040 -136960 118240 -136760 1 PIX2339_IN
port 2395 n
rlabel metal5 121040 -136960 121240 -136760 1 PIX2340_IN
port 2396 n
rlabel metal5 124040 -136960 124240 -136760 1 PIX2341_IN
port 2397 n
rlabel metal5 127040 -136960 127240 -136760 1 PIX2342_IN
port 2398 n
rlabel metal5 130040 -136960 130240 -136760 1 PIX2343_IN
port 2399 n
rlabel metal5 133040 -136960 133240 -136760 1 PIX2344_IN
port 2400 n
rlabel metal5 136040 -136960 136240 -136760 1 PIX2345_IN
port 2401 n
rlabel metal5 139040 -136960 139240 -136760 1 PIX2346_IN
port 2402 n
rlabel metal5 142040 -136960 142240 -136760 1 PIX2347_IN
port 2403 n
rlabel metal5 145040 -136960 145240 -136760 1 PIX2348_IN
port 2404 n
rlabel metal5 148040 -136960 148240 -136760 1 PIX2349_IN
port 2405 n
rlabel metal5 1040 -139960 1240 -139760 1 PIX2350_IN
port 2406 n
rlabel metal2 -3000 -139520 -3000 -139430 3 ROW_SEL47
port 2407 e
rlabel metal5 4040 -139960 4240 -139760 1 PIX2351_IN
port 2408 n
rlabel metal5 7040 -139960 7240 -139760 1 PIX2352_IN
port 2409 n
rlabel metal5 10040 -139960 10240 -139760 1 PIX2353_IN
port 2410 n
rlabel metal5 13040 -139960 13240 -139760 1 PIX2354_IN
port 2411 n
rlabel metal5 16040 -139960 16240 -139760 1 PIX2355_IN
port 2412 n
rlabel metal5 19040 -139960 19240 -139760 1 PIX2356_IN
port 2413 n
rlabel metal5 22040 -139960 22240 -139760 1 PIX2357_IN
port 2414 n
rlabel metal5 25040 -139960 25240 -139760 1 PIX2358_IN
port 2415 n
rlabel metal5 28040 -139960 28240 -139760 1 PIX2359_IN
port 2416 n
rlabel metal5 31040 -139960 31240 -139760 1 PIX2360_IN
port 2417 n
rlabel metal5 34040 -139960 34240 -139760 1 PIX2361_IN
port 2418 n
rlabel metal5 37040 -139960 37240 -139760 1 PIX2362_IN
port 2419 n
rlabel metal5 40040 -139960 40240 -139760 1 PIX2363_IN
port 2420 n
rlabel metal5 43040 -139960 43240 -139760 1 PIX2364_IN
port 2421 n
rlabel metal5 46040 -139960 46240 -139760 1 PIX2365_IN
port 2422 n
rlabel metal5 49040 -139960 49240 -139760 1 PIX2366_IN
port 2423 n
rlabel metal5 52040 -139960 52240 -139760 1 PIX2367_IN
port 2424 n
rlabel metal5 55040 -139960 55240 -139760 1 PIX2368_IN
port 2425 n
rlabel metal5 58040 -139960 58240 -139760 1 PIX2369_IN
port 2426 n
rlabel metal5 61040 -139960 61240 -139760 1 PIX2370_IN
port 2427 n
rlabel metal5 64040 -139960 64240 -139760 1 PIX2371_IN
port 2428 n
rlabel metal5 67040 -139960 67240 -139760 1 PIX2372_IN
port 2429 n
rlabel metal5 70040 -139960 70240 -139760 1 PIX2373_IN
port 2430 n
rlabel metal5 73040 -139960 73240 -139760 1 PIX2374_IN
port 2431 n
rlabel metal5 76040 -139960 76240 -139760 1 PIX2375_IN
port 2432 n
rlabel metal5 79040 -139960 79240 -139760 1 PIX2376_IN
port 2433 n
rlabel metal5 82040 -139960 82240 -139760 1 PIX2377_IN
port 2434 n
rlabel metal5 85040 -139960 85240 -139760 1 PIX2378_IN
port 2435 n
rlabel metal5 88040 -139960 88240 -139760 1 PIX2379_IN
port 2436 n
rlabel metal5 91040 -139960 91240 -139760 1 PIX2380_IN
port 2437 n
rlabel metal5 94040 -139960 94240 -139760 1 PIX2381_IN
port 2438 n
rlabel metal5 97040 -139960 97240 -139760 1 PIX2382_IN
port 2439 n
rlabel metal5 100040 -139960 100240 -139760 1 PIX2383_IN
port 2440 n
rlabel metal5 103040 -139960 103240 -139760 1 PIX2384_IN
port 2441 n
rlabel metal5 106040 -139960 106240 -139760 1 PIX2385_IN
port 2442 n
rlabel metal5 109040 -139960 109240 -139760 1 PIX2386_IN
port 2443 n
rlabel metal5 112040 -139960 112240 -139760 1 PIX2387_IN
port 2444 n
rlabel metal5 115040 -139960 115240 -139760 1 PIX2388_IN
port 2445 n
rlabel metal5 118040 -139960 118240 -139760 1 PIX2389_IN
port 2446 n
rlabel metal5 121040 -139960 121240 -139760 1 PIX2390_IN
port 2447 n
rlabel metal5 124040 -139960 124240 -139760 1 PIX2391_IN
port 2448 n
rlabel metal5 127040 -139960 127240 -139760 1 PIX2392_IN
port 2449 n
rlabel metal5 130040 -139960 130240 -139760 1 PIX2393_IN
port 2450 n
rlabel metal5 133040 -139960 133240 -139760 1 PIX2394_IN
port 2451 n
rlabel metal5 136040 -139960 136240 -139760 1 PIX2395_IN
port 2452 n
rlabel metal5 139040 -139960 139240 -139760 1 PIX2396_IN
port 2453 n
rlabel metal5 142040 -139960 142240 -139760 1 PIX2397_IN
port 2454 n
rlabel metal5 145040 -139960 145240 -139760 1 PIX2398_IN
port 2455 n
rlabel metal5 148040 -139960 148240 -139760 1 PIX2399_IN
port 2456 n
rlabel metal5 1040 -142960 1240 -142760 1 PIX2400_IN
port 2457 n
rlabel metal2 -3000 -142520 -3000 -142430 3 ROW_SEL48
port 2458 e
rlabel metal5 4040 -142960 4240 -142760 1 PIX2401_IN
port 2459 n
rlabel metal5 7040 -142960 7240 -142760 1 PIX2402_IN
port 2460 n
rlabel metal5 10040 -142960 10240 -142760 1 PIX2403_IN
port 2461 n
rlabel metal5 13040 -142960 13240 -142760 1 PIX2404_IN
port 2462 n
rlabel metal5 16040 -142960 16240 -142760 1 PIX2405_IN
port 2463 n
rlabel metal5 19040 -142960 19240 -142760 1 PIX2406_IN
port 2464 n
rlabel metal5 22040 -142960 22240 -142760 1 PIX2407_IN
port 2465 n
rlabel metal5 25040 -142960 25240 -142760 1 PIX2408_IN
port 2466 n
rlabel metal5 28040 -142960 28240 -142760 1 PIX2409_IN
port 2467 n
rlabel metal5 31040 -142960 31240 -142760 1 PIX2410_IN
port 2468 n
rlabel metal5 34040 -142960 34240 -142760 1 PIX2411_IN
port 2469 n
rlabel metal5 37040 -142960 37240 -142760 1 PIX2412_IN
port 2470 n
rlabel metal5 40040 -142960 40240 -142760 1 PIX2413_IN
port 2471 n
rlabel metal5 43040 -142960 43240 -142760 1 PIX2414_IN
port 2472 n
rlabel metal5 46040 -142960 46240 -142760 1 PIX2415_IN
port 2473 n
rlabel metal5 49040 -142960 49240 -142760 1 PIX2416_IN
port 2474 n
rlabel metal5 52040 -142960 52240 -142760 1 PIX2417_IN
port 2475 n
rlabel metal5 55040 -142960 55240 -142760 1 PIX2418_IN
port 2476 n
rlabel metal5 58040 -142960 58240 -142760 1 PIX2419_IN
port 2477 n
rlabel metal5 61040 -142960 61240 -142760 1 PIX2420_IN
port 2478 n
rlabel metal5 64040 -142960 64240 -142760 1 PIX2421_IN
port 2479 n
rlabel metal5 67040 -142960 67240 -142760 1 PIX2422_IN
port 2480 n
rlabel metal5 70040 -142960 70240 -142760 1 PIX2423_IN
port 2481 n
rlabel metal5 73040 -142960 73240 -142760 1 PIX2424_IN
port 2482 n
rlabel metal5 76040 -142960 76240 -142760 1 PIX2425_IN
port 2483 n
rlabel metal5 79040 -142960 79240 -142760 1 PIX2426_IN
port 2484 n
rlabel metal5 82040 -142960 82240 -142760 1 PIX2427_IN
port 2485 n
rlabel metal5 85040 -142960 85240 -142760 1 PIX2428_IN
port 2486 n
rlabel metal5 88040 -142960 88240 -142760 1 PIX2429_IN
port 2487 n
rlabel metal5 91040 -142960 91240 -142760 1 PIX2430_IN
port 2488 n
rlabel metal5 94040 -142960 94240 -142760 1 PIX2431_IN
port 2489 n
rlabel metal5 97040 -142960 97240 -142760 1 PIX2432_IN
port 2490 n
rlabel metal5 100040 -142960 100240 -142760 1 PIX2433_IN
port 2491 n
rlabel metal5 103040 -142960 103240 -142760 1 PIX2434_IN
port 2492 n
rlabel metal5 106040 -142960 106240 -142760 1 PIX2435_IN
port 2493 n
rlabel metal5 109040 -142960 109240 -142760 1 PIX2436_IN
port 2494 n
rlabel metal5 112040 -142960 112240 -142760 1 PIX2437_IN
port 2495 n
rlabel metal5 115040 -142960 115240 -142760 1 PIX2438_IN
port 2496 n
rlabel metal5 118040 -142960 118240 -142760 1 PIX2439_IN
port 2497 n
rlabel metal5 121040 -142960 121240 -142760 1 PIX2440_IN
port 2498 n
rlabel metal5 124040 -142960 124240 -142760 1 PIX2441_IN
port 2499 n
rlabel metal5 127040 -142960 127240 -142760 1 PIX2442_IN
port 2500 n
rlabel metal5 130040 -142960 130240 -142760 1 PIX2443_IN
port 2501 n
rlabel metal5 133040 -142960 133240 -142760 1 PIX2444_IN
port 2502 n
rlabel metal5 136040 -142960 136240 -142760 1 PIX2445_IN
port 2503 n
rlabel metal5 139040 -142960 139240 -142760 1 PIX2446_IN
port 2504 n
rlabel metal5 142040 -142960 142240 -142760 1 PIX2447_IN
port 2505 n
rlabel metal5 145040 -142960 145240 -142760 1 PIX2448_IN
port 2506 n
rlabel metal5 148040 -142960 148240 -142760 1 PIX2449_IN
port 2507 n
rlabel metal5 1040 -145960 1240 -145760 1 PIX2450_IN
port 2508 n
rlabel metal4 2630 -147200 2780 -147000 1 PIX_OUT0
port 2509 n
rlabel metal4 220 -148100 440 -147700 1 COL_SEL0
port 2510 n
rlabel metal4 -480 -148600 -480 -148600 1 CSA_VREF
port 2511 n
rlabel metal2 -3000 -145520 -3000 -145430 3 ROW_SEL49
port 2512 e
rlabel metal5 4040 -145960 4240 -145760 1 PIX2451_IN
port 2513 n
rlabel metal4 5630 -147200 5780 -147000 1 PIX_OUT1
port 2514 n
rlabel metal4 3220 -148100 3440 -147700 1 COL_SEL1
port 2515 n
rlabel metal5 7040 -145960 7240 -145760 1 PIX2452_IN
port 2516 n
rlabel metal4 8630 -147200 8780 -147000 1 PIX_OUT2
port 2517 n
rlabel metal4 6220 -148100 6440 -147700 1 COL_SEL2
port 2518 n
rlabel metal5 10040 -145960 10240 -145760 1 PIX2453_IN
port 2519 n
rlabel metal4 11630 -147200 11780 -147000 1 PIX_OUT3
port 2520 n
rlabel metal4 9220 -148100 9440 -147700 1 COL_SEL3
port 2521 n
rlabel metal5 13040 -145960 13240 -145760 1 PIX2454_IN
port 2522 n
rlabel metal4 14630 -147200 14780 -147000 1 PIX_OUT4
port 2523 n
rlabel metal4 12220 -148100 12440 -147700 1 COL_SEL4
port 2524 n
rlabel metal5 16040 -145960 16240 -145760 1 PIX2455_IN
port 2525 n
rlabel metal4 17630 -147200 17780 -147000 1 PIX_OUT5
port 2526 n
rlabel metal4 15220 -148100 15440 -147700 1 COL_SEL5
port 2527 n
rlabel metal5 19040 -145960 19240 -145760 1 PIX2456_IN
port 2528 n
rlabel metal4 20630 -147200 20780 -147000 1 PIX_OUT6
port 2529 n
rlabel metal4 18220 -148100 18440 -147700 1 COL_SEL6
port 2530 n
rlabel metal5 22040 -145960 22240 -145760 1 PIX2457_IN
port 2531 n
rlabel metal4 23630 -147200 23780 -147000 1 PIX_OUT7
port 2532 n
rlabel metal4 21220 -148100 21440 -147700 1 COL_SEL7
port 2533 n
rlabel metal5 25040 -145960 25240 -145760 1 PIX2458_IN
port 2534 n
rlabel metal4 26630 -147200 26780 -147000 1 PIX_OUT8
port 2535 n
rlabel metal4 24220 -148100 24440 -147700 1 COL_SEL8
port 2536 n
rlabel metal5 28040 -145960 28240 -145760 1 PIX2459_IN
port 2537 n
rlabel metal4 29630 -147200 29780 -147000 1 PIX_OUT9
port 2538 n
rlabel metal4 27220 -148100 27440 -147700 1 COL_SEL9
port 2539 n
rlabel metal5 31040 -145960 31240 -145760 1 PIX2460_IN
port 2540 n
rlabel metal4 32630 -147200 32780 -147000 1 PIX_OUT10
port 2541 n
rlabel metal4 30220 -148100 30440 -147700 1 COL_SEL10
port 2542 n
rlabel metal5 34040 -145960 34240 -145760 1 PIX2461_IN
port 2543 n
rlabel metal4 35630 -147200 35780 -147000 1 PIX_OUT11
port 2544 n
rlabel metal4 33220 -148100 33440 -147700 1 COL_SEL11
port 2545 n
rlabel metal5 37040 -145960 37240 -145760 1 PIX2462_IN
port 2546 n
rlabel metal4 38630 -147200 38780 -147000 1 PIX_OUT12
port 2547 n
rlabel metal4 36220 -148100 36440 -147700 1 COL_SEL12
port 2548 n
rlabel metal5 40040 -145960 40240 -145760 1 PIX2463_IN
port 2549 n
rlabel metal4 41630 -147200 41780 -147000 1 PIX_OUT13
port 2550 n
rlabel metal4 39220 -148100 39440 -147700 1 COL_SEL13
port 2551 n
rlabel metal5 43040 -145960 43240 -145760 1 PIX2464_IN
port 2552 n
rlabel metal4 44630 -147200 44780 -147000 1 PIX_OUT14
port 2553 n
rlabel metal4 42220 -148100 42440 -147700 1 COL_SEL14
port 2554 n
rlabel metal5 46040 -145960 46240 -145760 1 PIX2465_IN
port 2555 n
rlabel metal4 47630 -147200 47780 -147000 1 PIX_OUT15
port 2556 n
rlabel metal4 45220 -148100 45440 -147700 1 COL_SEL15
port 2557 n
rlabel metal5 49040 -145960 49240 -145760 1 PIX2466_IN
port 2558 n
rlabel metal4 50630 -147200 50780 -147000 1 PIX_OUT16
port 2559 n
rlabel metal4 48220 -148100 48440 -147700 1 COL_SEL16
port 2560 n
rlabel metal5 52040 -145960 52240 -145760 1 PIX2467_IN
port 2561 n
rlabel metal4 53630 -147200 53780 -147000 1 PIX_OUT17
port 2562 n
rlabel metal4 51220 -148100 51440 -147700 1 COL_SEL17
port 2563 n
rlabel metal5 55040 -145960 55240 -145760 1 PIX2468_IN
port 2564 n
rlabel metal4 56630 -147200 56780 -147000 1 PIX_OUT18
port 2565 n
rlabel metal4 54220 -148100 54440 -147700 1 COL_SEL18
port 2566 n
rlabel metal5 58040 -145960 58240 -145760 1 PIX2469_IN
port 2567 n
rlabel metal4 59630 -147200 59780 -147000 1 PIX_OUT19
port 2568 n
rlabel metal4 57220 -148100 57440 -147700 1 COL_SEL19
port 2569 n
rlabel metal5 61040 -145960 61240 -145760 1 PIX2470_IN
port 2570 n
rlabel metal4 62630 -147200 62780 -147000 1 PIX_OUT20
port 2571 n
rlabel metal4 60220 -148100 60440 -147700 1 COL_SEL20
port 2572 n
rlabel metal5 64040 -145960 64240 -145760 1 PIX2471_IN
port 2573 n
rlabel metal4 65630 -147200 65780 -147000 1 PIX_OUT21
port 2574 n
rlabel metal4 63220 -148100 63440 -147700 1 COL_SEL21
port 2575 n
rlabel metal5 67040 -145960 67240 -145760 1 PIX2472_IN
port 2576 n
rlabel metal4 68630 -147200 68780 -147000 1 PIX_OUT22
port 2577 n
rlabel metal4 66220 -148100 66440 -147700 1 COL_SEL22
port 2578 n
rlabel metal5 70040 -145960 70240 -145760 1 PIX2473_IN
port 2579 n
rlabel metal4 71630 -147200 71780 -147000 1 PIX_OUT23
port 2580 n
rlabel metal4 69220 -148100 69440 -147700 1 COL_SEL23
port 2581 n
rlabel metal5 73040 -145960 73240 -145760 1 PIX2474_IN
port 2582 n
rlabel metal4 74630 -147200 74780 -147000 1 PIX_OUT24
port 2583 n
rlabel metal4 72220 -148100 72440 -147700 1 COL_SEL24
port 2584 n
rlabel metal5 76040 -145960 76240 -145760 1 PIX2475_IN
port 2585 n
rlabel metal4 77630 -147200 77780 -147000 1 PIX_OUT25
port 2586 n
rlabel metal4 75220 -148100 75440 -147700 1 COL_SEL25
port 2587 n
rlabel metal5 79040 -145960 79240 -145760 1 PIX2476_IN
port 2588 n
rlabel metal4 80630 -147200 80780 -147000 1 PIX_OUT26
port 2589 n
rlabel metal4 78220 -148100 78440 -147700 1 COL_SEL26
port 2590 n
rlabel metal5 82040 -145960 82240 -145760 1 PIX2477_IN
port 2591 n
rlabel metal4 83630 -147200 83780 -147000 1 PIX_OUT27
port 2592 n
rlabel metal4 81220 -148100 81440 -147700 1 COL_SEL27
port 2593 n
rlabel metal5 85040 -145960 85240 -145760 1 PIX2478_IN
port 2594 n
rlabel metal4 86630 -147200 86780 -147000 1 PIX_OUT28
port 2595 n
rlabel metal4 84220 -148100 84440 -147700 1 COL_SEL28
port 2596 n
rlabel metal5 88040 -145960 88240 -145760 1 PIX2479_IN
port 2597 n
rlabel metal4 89630 -147200 89780 -147000 1 PIX_OUT29
port 2598 n
rlabel metal4 87220 -148100 87440 -147700 1 COL_SEL29
port 2599 n
rlabel metal5 91040 -145960 91240 -145760 1 PIX2480_IN
port 2600 n
rlabel metal4 92630 -147200 92780 -147000 1 PIX_OUT30
port 2601 n
rlabel metal4 90220 -148100 90440 -147700 1 COL_SEL30
port 2602 n
rlabel metal5 94040 -145960 94240 -145760 1 PIX2481_IN
port 2603 n
rlabel metal4 95630 -147200 95780 -147000 1 PIX_OUT31
port 2604 n
rlabel metal4 93220 -148100 93440 -147700 1 COL_SEL31
port 2605 n
rlabel metal5 97040 -145960 97240 -145760 1 PIX2482_IN
port 2606 n
rlabel metal4 98630 -147200 98780 -147000 1 PIX_OUT32
port 2607 n
rlabel metal4 96220 -148100 96440 -147700 1 COL_SEL32
port 2608 n
rlabel metal5 100040 -145960 100240 -145760 1 PIX2483_IN
port 2609 n
rlabel metal4 101630 -147200 101780 -147000 1 PIX_OUT33
port 2610 n
rlabel metal4 99220 -148100 99440 -147700 1 COL_SEL33
port 2611 n
rlabel metal5 103040 -145960 103240 -145760 1 PIX2484_IN
port 2612 n
rlabel metal4 104630 -147200 104780 -147000 1 PIX_OUT34
port 2613 n
rlabel metal4 102220 -148100 102440 -147700 1 COL_SEL34
port 2614 n
rlabel metal5 106040 -145960 106240 -145760 1 PIX2485_IN
port 2615 n
rlabel metal4 107630 -147200 107780 -147000 1 PIX_OUT35
port 2616 n
rlabel metal4 105220 -148100 105440 -147700 1 COL_SEL35
port 2617 n
rlabel metal5 109040 -145960 109240 -145760 1 PIX2486_IN
port 2618 n
rlabel metal4 110630 -147200 110780 -147000 1 PIX_OUT36
port 2619 n
rlabel metal4 108220 -148100 108440 -147700 1 COL_SEL36
port 2620 n
rlabel metal5 112040 -145960 112240 -145760 1 PIX2487_IN
port 2621 n
rlabel metal4 113630 -147200 113780 -147000 1 PIX_OUT37
port 2622 n
rlabel metal4 111220 -148100 111440 -147700 1 COL_SEL37
port 2623 n
rlabel metal5 115040 -145960 115240 -145760 1 PIX2488_IN
port 2624 n
rlabel metal4 116630 -147200 116780 -147000 1 PIX_OUT38
port 2625 n
rlabel metal4 114220 -148100 114440 -147700 1 COL_SEL38
port 2626 n
rlabel metal5 118040 -145960 118240 -145760 1 PIX2489_IN
port 2627 n
rlabel metal4 119630 -147200 119780 -147000 1 PIX_OUT39
port 2628 n
rlabel metal4 117220 -148100 117440 -147700 1 COL_SEL39
port 2629 n
rlabel metal5 121040 -145960 121240 -145760 1 PIX2490_IN
port 2630 n
rlabel metal4 122630 -147200 122780 -147000 1 PIX_OUT40
port 2631 n
rlabel metal4 120220 -148100 120440 -147700 1 COL_SEL40
port 2632 n
rlabel metal5 124040 -145960 124240 -145760 1 PIX2491_IN
port 2633 n
rlabel metal4 125630 -147200 125780 -147000 1 PIX_OUT41
port 2634 n
rlabel metal4 123220 -148100 123440 -147700 1 COL_SEL41
port 2635 n
rlabel metal5 127040 -145960 127240 -145760 1 PIX2492_IN
port 2636 n
rlabel metal4 128630 -147200 128780 -147000 1 PIX_OUT42
port 2637 n
rlabel metal4 126220 -148100 126440 -147700 1 COL_SEL42
port 2638 n
rlabel metal5 130040 -145960 130240 -145760 1 PIX2493_IN
port 2639 n
rlabel metal4 131630 -147200 131780 -147000 1 PIX_OUT43
port 2640 n
rlabel metal4 129220 -148100 129440 -147700 1 COL_SEL43
port 2641 n
rlabel metal5 133040 -145960 133240 -145760 1 PIX2494_IN
port 2642 n
rlabel metal4 134630 -147200 134780 -147000 1 PIX_OUT44
port 2643 n
rlabel metal4 132220 -148100 132440 -147700 1 COL_SEL44
port 2644 n
rlabel metal5 136040 -145960 136240 -145760 1 PIX2495_IN
port 2645 n
rlabel metal4 137630 -147200 137780 -147000 1 PIX_OUT45
port 2646 n
rlabel metal4 135220 -148100 135440 -147700 1 COL_SEL45
port 2647 n
rlabel metal5 139040 -145960 139240 -145760 1 PIX2496_IN
port 2648 n
rlabel metal4 140630 -147200 140780 -147000 1 PIX_OUT46
port 2649 n
rlabel metal4 138220 -148100 138440 -147700 1 COL_SEL46
port 2650 n
rlabel metal5 142040 -145960 142240 -145760 1 PIX2497_IN
port 2651 n
rlabel metal4 143630 -147200 143780 -147000 1 PIX_OUT47
port 2652 n
rlabel metal4 141220 -148100 141440 -147700 1 COL_SEL47
port 2653 n
rlabel metal5 145040 -145960 145240 -145760 1 PIX2498_IN
port 2654 n
rlabel metal4 146630 -147200 146780 -147000 1 PIX_OUT48
port 2655 n
rlabel metal4 144220 -148100 144440 -147700 1 COL_SEL48
port 2656 n
rlabel metal5 148040 -145960 148240 -145760 1 PIX2499_IN
port 2657 n
rlabel metal4 149630 -147200 149780 -147000 1 PIX_OUT49
port 2658 n
rlabel metal2 149940 -148100 149940 -148100 1 ARRAY_OUT
port 2659 n
rlabel metal4 147220 -148100 147440 -147700 1 COL_SEL49
port 2660 n
<< end >>
