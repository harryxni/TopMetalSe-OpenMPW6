magic
tech sky130A
magscale 1 2
timestamp 1654625306
<< nmoslvt >>
rect -950 9870 650 10270
rect 280 -850 1880 -450
<< ndiff >>
rect -950 10620 650 10670
rect -950 10290 -930 10620
rect 630 10290 650 10620
rect -950 10270 650 10290
rect -950 9840 650 9870
rect -950 9620 -930 9840
rect 630 9620 650 9840
rect -950 9610 650 9620
rect 280 -140 1880 -120
rect 280 -420 300 -140
rect 1860 -420 1880 -140
rect 280 -450 1880 -420
rect 280 -880 1880 -850
rect 280 -1050 300 -880
rect 1860 -1050 1880 -880
rect 280 -1080 1880 -1050
<< ndiffc >>
rect -930 10290 630 10620
rect -930 9620 630 9840
rect 300 -420 1860 -140
rect 300 -1050 1860 -880
<< psubdiff >>
rect -950 9560 650 9610
rect -950 9320 -920 9560
rect 620 9320 650 9560
rect -950 9270 650 9320
rect 280 -1110 1880 -1080
rect 280 -1360 310 -1110
rect 1850 -1360 1880 -1110
rect 280 -1560 1880 -1360
<< psubdiffcont >>
rect -920 9320 620 9560
rect 310 -1360 1850 -1110
<< poly >>
rect -980 10080 -950 10270
rect -1370 10060 -950 10080
rect -1370 9890 -1350 10060
rect -1130 9890 -950 10060
rect -1370 9870 -950 9890
rect 650 9870 680 10270
rect -110 -240 100 -230
rect -110 -410 -90 -240
rect 60 -410 100 -240
rect -110 -450 100 -410
rect -110 -500 280 -450
rect 250 -850 280 -500
rect 1880 -850 1910 -450
<< polycont >>
rect -1350 9890 -1130 10060
rect -90 -410 60 -240
<< locali >>
rect -950 10620 650 10650
rect -950 10290 -930 10620
rect 630 10290 650 10620
rect -950 10270 650 10290
rect -1690 10050 -1350 10060
rect -1130 10050 -1020 10060
rect -1690 9900 -1670 10050
rect -1040 9900 -1020 10050
rect -1690 9890 -1350 9900
rect -1130 9890 -1020 9900
rect -950 9840 650 9850
rect -950 9300 -930 9840
rect 630 9300 650 9840
rect -950 9270 650 9300
rect -400 -250 -90 -240
rect -400 -400 -390 -250
rect -110 -400 -90 -250
rect -400 -410 -90 -400
rect 60 -410 100 -240
rect 280 -420 300 60
rect 1860 -420 1880 60
rect 280 -430 1880 -420
rect 280 -880 1880 -870
rect 280 -1050 300 -880
rect 1860 -1050 1880 -880
rect 280 -1110 1880 -1050
rect 280 -1300 310 -1110
rect 1850 -1300 1880 -1110
rect 280 -1530 300 -1300
rect 1860 -1530 1880 -1300
rect 280 -1550 1880 -1530
<< viali >>
rect -930 10290 630 10620
rect -1670 9900 -1350 10050
rect -1350 9900 -1130 10050
rect -1130 9900 -1040 10050
rect -930 9620 630 9770
rect -930 9560 630 9620
rect -930 9320 -920 9560
rect -920 9320 620 9560
rect 620 9320 630 9560
rect -930 9300 630 9320
rect -390 -400 -110 -250
rect 300 -140 1860 60
rect 300 -420 1860 -140
rect 300 -1360 310 -1300
rect 310 -1360 1850 -1300
rect 1850 -1360 1860 -1300
rect 300 -1530 1860 -1360
<< metal1 >>
rect 23020 11280 26995 11570
rect -950 10620 650 10630
rect -950 10290 -930 10620
rect 630 10290 650 10620
rect -950 10270 650 10290
rect -2280 10050 -1020 10060
rect -2280 9900 -1670 10050
rect -1040 9900 -1020 10050
rect -2280 9890 -1020 9900
rect -960 9770 650 9850
rect -960 9300 -930 9770
rect 630 9300 650 9770
rect -960 9220 650 9300
rect 280 60 1880 180
rect -500 -250 100 -240
rect -500 -400 -490 -250
rect -500 -410 -390 -400
rect -110 -410 100 -250
rect 280 -420 300 60
rect 1860 -420 1880 60
rect 280 -430 1880 -420
rect -950 -1290 2500 -1280
rect -950 -1550 -920 -1290
rect 2280 -1550 2500 -1290
rect -950 -1560 2500 -1550
rect 24530 -1570 26980 -1270
<< via1 >>
rect -930 10290 630 10620
rect -930 9300 630 9770
rect -490 -400 -390 -250
rect -390 -400 -110 -250
rect -390 -410 -110 -400
rect 300 -420 1860 60
rect -920 -1300 2280 -1290
rect -920 -1530 300 -1300
rect 300 -1530 1860 -1300
rect 1860 -1530 2280 -1300
rect -920 -1550 2280 -1530
<< metal2 >>
rect -950 10620 650 10630
rect -950 10290 -930 10620
rect 630 10290 650 10620
rect -950 10270 650 10290
rect -950 10269 529 10270
rect -960 9770 650 9850
rect -960 9300 -930 9770
rect 630 9300 650 9770
rect -960 9220 650 9300
rect 1300 8370 2520 8450
rect 1300 7710 1320 8370
rect 2490 7710 2520 8370
rect 1300 7620 2520 7710
rect 280 3859 1890 3870
rect -1688 3611 2174 3859
rect 280 60 1890 3611
rect -1190 -250 -100 -240
rect -1190 -400 -490 -250
rect -1190 -410 -390 -400
rect -110 -410 -100 -250
rect 280 -420 300 60
rect 1860 -420 1890 60
rect 280 -430 1890 -420
rect -950 -1290 2490 -1280
rect -950 -1550 -920 -1290
rect 2280 -1550 2490 -1290
rect -950 -1560 2490 -1550
<< via2 >>
rect -930 9300 630 9770
rect 1320 7710 2490 8370
rect -920 -1550 2280 -1290
<< metal3 >>
rect -960 9770 650 9850
rect -960 9300 -930 9770
rect 630 9300 650 9770
rect -960 9220 650 9300
rect -950 -1280 -265 9220
rect 1300 8370 2520 8450
rect 1300 7710 1320 8370
rect 2490 7710 2520 8370
rect 1300 7620 2520 7710
rect -950 -1290 2490 -1280
rect -950 -1550 -920 -1290
rect 2280 -1550 2490 -1290
rect -950 -1560 2490 -1550
<< via3 >>
rect 1320 7710 2490 8370
<< metal4 >>
rect -2205 12835 26620 13665
rect -2205 8455 -1375 12835
rect -2205 8370 2515 8455
rect -2205 7710 1320 8370
rect 2490 7710 2515 8370
rect -2205 7625 2515 7710
rect 25795 7690 26620 12835
rect 24850 6830 26620 7690
use opamp_diego  opamp_diego_0 ~/CMOS/TopmetalSe/magic
timestamp 1654624193
transform 1 0 -1719 0 1 8388
box 2069 -10028 26971 3199
<< labels >>
rlabel metal1 26870 -1360 26870 -1360 1 GND
port 6 n
rlabel metal1 26840 11440 26840 11440 1 VDD
port 1 n
rlabel metal4 26418 7258 26418 7258 1 AOUT
port 2 n
rlabel metal1 -2240 9968 -2240 9968 1 AMP_IB
port 4 n
rlabel metal2 -1576 3762 -1576 3762 1 ARRAY_OUT
port 5 n
rlabel metal2 -1078 -314 -1078 -314 1 OUT_IB
port 3 n
<< end >>
