magic
tech sky130A
magscale 1 2
timestamp 1654709766
<< error_p >>
rect 313959 -286004 313993 -285428
rect 319297 -286005 319331 -285429
rect 319415 -286005 319449 -285429
rect 319533 -286005 319567 -285429
rect 319651 -286005 319685 -285429
rect 319769 -286005 319803 -285429
rect 319887 -286005 319921 -285429
rect 320005 -286005 320039 -285429
rect 320123 -286005 320157 -285429
rect 320241 -286005 320275 -285429
rect 320359 -286005 320393 -285429
rect 320477 -286005 320511 -285429
rect 320595 -286005 320629 -285429
rect 320713 -286005 320747 -285429
rect 320831 -286005 320865 -285429
rect 320949 -286005 320983 -285429
rect 321067 -286005 321101 -285429
rect 321185 -286005 321219 -285429
rect 321303 -286005 321337 -285429
rect 321421 -286005 321455 -285429
rect 321539 -286005 321573 -285429
rect 321657 -286005 321691 -285429
rect 321775 -286005 321809 -285429
rect 321893 -286005 321927 -285429
rect 322011 -286005 322045 -285429
rect 323420 -286005 323454 -285429
rect 323538 -286005 323572 -285429
rect 323656 -286005 323690 -285429
rect 323774 -286005 323808 -285429
rect 323892 -286005 323926 -285429
rect 324010 -286005 324044 -285429
rect 324128 -286005 324162 -285429
rect 324246 -286005 324280 -285429
rect 324364 -286005 324398 -285429
rect 324482 -286005 324516 -285429
rect 324600 -286005 324634 -285429
rect 324718 -286005 324752 -285429
rect 324836 -286005 324870 -285429
rect 324954 -286005 324988 -285429
rect 325072 -286005 325106 -285429
rect 325190 -286005 325224 -285429
rect 325308 -286005 325342 -285429
rect 325426 -286005 325460 -285429
rect 325544 -286005 325578 -285429
rect 325662 -286005 325696 -285429
rect 325780 -286005 325814 -285429
rect 325898 -286005 325932 -285429
rect 326016 -286005 326050 -285429
rect 326134 -286005 326168 -285429
rect 327543 -286005 327577 -285429
rect 327661 -286005 327695 -285429
rect 327779 -286005 327813 -285429
rect 327897 -286005 327931 -285429
rect 328015 -286005 328049 -285429
rect 328133 -286005 328167 -285429
rect 328251 -286005 328285 -285429
rect 328369 -286005 328403 -285429
rect 328487 -286005 328521 -285429
rect 328605 -286005 328639 -285429
rect 328723 -286005 328757 -285429
rect 328841 -286005 328875 -285429
rect 328959 -286005 328993 -285429
rect 329077 -286005 329111 -285429
rect 329195 -286005 329229 -285429
rect 329313 -286005 329347 -285429
rect 329431 -286005 329465 -285429
rect 329549 -286005 329583 -285429
rect 329667 -286005 329701 -285429
rect 329785 -286005 329819 -285429
rect 329903 -286005 329937 -285429
rect 330021 -286005 330055 -285429
rect 330139 -286005 330173 -285429
rect 330257 -286005 330291 -285429
rect 311353 -286764 317323 -286730
rect 311257 -288436 311291 -286826
rect 311371 -287501 311405 -286925
rect 311489 -287501 311523 -286925
rect 311607 -287501 311641 -286925
rect 311725 -287501 311759 -286925
rect 311843 -287501 311877 -286925
rect 311961 -287501 311995 -286925
rect 312079 -287501 312113 -286925
rect 312197 -287501 312231 -286925
rect 312315 -287501 312349 -286925
rect 312433 -287501 312467 -286925
rect 312551 -287501 312585 -286925
rect 312669 -287501 312703 -286925
rect 312787 -287501 312821 -286925
rect 312905 -287501 312939 -286925
rect 313023 -287501 313057 -286925
rect 313141 -287501 313175 -286925
rect 313259 -287501 313293 -286925
rect 313377 -287501 313411 -286925
rect 313495 -287501 313529 -286925
rect 313613 -287501 313647 -286925
rect 313731 -287501 313765 -286925
rect 313849 -287501 313883 -286925
rect 313967 -287501 314001 -286925
rect 314085 -287501 314119 -286925
rect 314203 -287501 314237 -286925
rect 314321 -287501 314355 -286925
rect 314439 -287501 314473 -286925
rect 314557 -287501 314591 -286925
rect 314675 -287501 314709 -286925
rect 314793 -287501 314827 -286925
rect 314911 -287501 314945 -286925
rect 315029 -287501 315063 -286925
rect 315147 -287501 315181 -286925
rect 315265 -287501 315299 -286925
rect 315383 -287501 315417 -286925
rect 315501 -287501 315535 -286925
rect 315619 -287501 315653 -286925
rect 315737 -287501 315771 -286925
rect 315855 -287501 315889 -286925
rect 315973 -287501 316007 -286925
rect 316091 -287501 316125 -286925
rect 316209 -287501 316243 -286925
rect 316327 -287501 316361 -286925
rect 316445 -287501 316479 -286925
rect 316563 -287501 316597 -286925
rect 316681 -287501 316715 -286925
rect 316799 -287501 316833 -286925
rect 316917 -287501 316951 -286925
rect 317035 -287501 317069 -286925
rect 317153 -287501 317187 -286925
rect 317271 -287501 317305 -286925
rect 311371 -288337 311405 -287761
rect 311489 -288337 311523 -287761
rect 311607 -288337 311641 -287761
rect 311725 -288337 311759 -287761
rect 311843 -288337 311877 -287761
rect 311961 -288337 311995 -287761
rect 312079 -288337 312113 -287761
rect 312197 -288337 312231 -287761
rect 312315 -288337 312349 -287761
rect 312433 -288337 312467 -287761
rect 312551 -288337 312585 -287761
rect 312669 -288337 312703 -287761
rect 312787 -288337 312821 -287761
rect 312905 -288337 312939 -287761
rect 313023 -288337 313057 -287761
rect 313141 -288337 313175 -287761
rect 313259 -288337 313293 -287761
rect 313377 -288337 313411 -287761
rect 313495 -288337 313529 -287761
rect 313613 -288337 313647 -287761
rect 313731 -288337 313765 -287761
rect 313849 -288337 313883 -287761
rect 313967 -288337 314001 -287761
rect 314085 -288337 314119 -287761
rect 314203 -288337 314237 -287761
rect 314321 -288337 314355 -287761
rect 314439 -288337 314473 -287761
rect 314557 -288337 314591 -287761
rect 314675 -288337 314709 -287761
rect 314793 -288337 314827 -287761
rect 314911 -288337 314945 -287761
rect 315029 -288337 315063 -287761
rect 315147 -288337 315181 -287761
rect 315265 -288337 315299 -287761
rect 315383 -288337 315417 -287761
rect 315501 -288337 315535 -287761
rect 315619 -288337 315653 -287761
rect 315737 -288337 315771 -287761
rect 315855 -288337 315889 -287761
rect 315973 -288337 316007 -287761
rect 316091 -288337 316125 -287761
rect 316209 -288337 316243 -287761
rect 316327 -288337 316361 -287761
rect 316445 -288337 316479 -287761
rect 316563 -288337 316597 -287761
rect 316681 -288337 316715 -287761
rect 316799 -288337 316833 -287761
rect 316917 -288337 316951 -287761
rect 317035 -288337 317069 -287761
rect 317153 -288337 317187 -287761
rect 317271 -288337 317305 -287761
rect 317385 -288436 317419 -286826
rect 319061 -286841 319095 -286265
rect 319179 -286841 319213 -286265
rect 319297 -286841 319331 -286265
rect 319415 -286841 319449 -286265
rect 319533 -286841 319567 -286265
rect 319651 -286841 319685 -286265
rect 319769 -286841 319803 -286265
rect 319887 -286841 319921 -286265
rect 320005 -286841 320039 -286265
rect 320123 -286841 320157 -286265
rect 320241 -286841 320275 -286265
rect 320359 -286841 320393 -286265
rect 320477 -286841 320511 -286265
rect 320595 -286841 320629 -286265
rect 320713 -286841 320747 -286265
rect 320831 -286841 320865 -286265
rect 320949 -286841 320983 -286265
rect 321067 -286841 321101 -286265
rect 321185 -286841 321219 -286265
rect 321303 -286841 321337 -286265
rect 321421 -286841 321455 -286265
rect 321539 -286841 321573 -286265
rect 321657 -286841 321691 -286265
rect 321775 -286841 321809 -286265
rect 321893 -286841 321927 -286265
rect 322011 -286841 322045 -286265
rect 323184 -286841 323218 -286265
rect 323302 -286841 323336 -286265
rect 323420 -286841 323454 -286265
rect 323538 -286841 323572 -286265
rect 323656 -286841 323690 -286265
rect 323774 -286841 323808 -286265
rect 323892 -286841 323926 -286265
rect 324010 -286841 324044 -286265
rect 324128 -286841 324162 -286265
rect 324246 -286841 324280 -286265
rect 324364 -286841 324398 -286265
rect 324482 -286841 324516 -286265
rect 324600 -286841 324634 -286265
rect 324718 -286841 324752 -286265
rect 324836 -286841 324870 -286265
rect 324954 -286841 324988 -286265
rect 325072 -286841 325106 -286265
rect 325190 -286841 325224 -286265
rect 325308 -286841 325342 -286265
rect 325426 -286841 325460 -286265
rect 325544 -286841 325578 -286265
rect 325662 -286841 325696 -286265
rect 325780 -286841 325814 -286265
rect 325898 -286841 325932 -286265
rect 326016 -286841 326050 -286265
rect 326134 -286841 326168 -286265
rect 327307 -286841 327341 -286265
rect 327425 -286841 327459 -286265
rect 327543 -286841 327577 -286265
rect 327661 -286841 327695 -286265
rect 327779 -286841 327813 -286265
rect 327897 -286841 327931 -286265
rect 328015 -286841 328049 -286265
rect 328133 -286841 328167 -286265
rect 328251 -286841 328285 -286265
rect 328369 -286841 328403 -286265
rect 328487 -286841 328521 -286265
rect 328605 -286841 328639 -286265
rect 328723 -286841 328757 -286265
rect 328841 -286841 328875 -286265
rect 328959 -286841 328993 -286265
rect 329077 -286841 329111 -286265
rect 329195 -286841 329229 -286265
rect 329313 -286841 329347 -286265
rect 329431 -286841 329465 -286265
rect 329549 -286841 329583 -286265
rect 329667 -286841 329701 -286265
rect 329785 -286841 329819 -286265
rect 329903 -286841 329937 -286265
rect 330021 -286841 330055 -286265
rect 330139 -286841 330173 -286265
rect 330257 -286841 330291 -286265
rect 311353 -288532 317323 -288498
rect 311353 -288814 317323 -288780
rect 311257 -290486 311291 -288876
rect 311371 -289551 311405 -288975
rect 311489 -289551 311523 -288975
rect 311607 -289551 311641 -288975
rect 311725 -289551 311759 -288975
rect 311843 -289551 311877 -288975
rect 311961 -289551 311995 -288975
rect 312079 -289551 312113 -288975
rect 312197 -289551 312231 -288975
rect 312315 -289551 312349 -288975
rect 312433 -289551 312467 -288975
rect 312551 -289551 312585 -288975
rect 312669 -289551 312703 -288975
rect 312787 -289551 312821 -288975
rect 312905 -289551 312939 -288975
rect 313023 -289551 313057 -288975
rect 313141 -289551 313175 -288975
rect 313259 -289551 313293 -288975
rect 313377 -289551 313411 -288975
rect 313495 -289551 313529 -288975
rect 313613 -289551 313647 -288975
rect 313731 -289551 313765 -288975
rect 313849 -289551 313883 -288975
rect 313967 -289551 314001 -288975
rect 314085 -289551 314119 -288975
rect 314203 -289551 314237 -288975
rect 314321 -289551 314355 -288975
rect 314439 -289551 314473 -288975
rect 314557 -289551 314591 -288975
rect 314675 -289551 314709 -288975
rect 314793 -289551 314827 -288975
rect 314911 -289551 314945 -288975
rect 315029 -289551 315063 -288975
rect 315147 -289551 315181 -288975
rect 315265 -289551 315299 -288975
rect 315383 -289551 315417 -288975
rect 315501 -289551 315535 -288975
rect 315619 -289551 315653 -288975
rect 315737 -289551 315771 -288975
rect 315855 -289551 315889 -288975
rect 315973 -289551 316007 -288975
rect 316091 -289551 316125 -288975
rect 316209 -289551 316243 -288975
rect 316327 -289551 316361 -288975
rect 316445 -289551 316479 -288975
rect 316563 -289551 316597 -288975
rect 316681 -289551 316715 -288975
rect 316799 -289551 316833 -288975
rect 316917 -289551 316951 -288975
rect 317035 -289551 317069 -288975
rect 317153 -289551 317187 -288975
rect 317271 -289551 317305 -288975
rect 311371 -290387 311405 -289811
rect 311489 -290387 311523 -289811
rect 311607 -290387 311641 -289811
rect 311725 -290387 311759 -289811
rect 311843 -290387 311877 -289811
rect 311961 -290387 311995 -289811
rect 312079 -290387 312113 -289811
rect 312197 -290387 312231 -289811
rect 312315 -290387 312349 -289811
rect 312433 -290387 312467 -289811
rect 312551 -290387 312585 -289811
rect 312669 -290387 312703 -289811
rect 312787 -290387 312821 -289811
rect 312905 -290387 312939 -289811
rect 313023 -290387 313057 -289811
rect 313141 -290387 313175 -289811
rect 313259 -290387 313293 -289811
rect 313377 -290387 313411 -289811
rect 313495 -290387 313529 -289811
rect 313613 -290387 313647 -289811
rect 313731 -290387 313765 -289811
rect 313849 -290387 313883 -289811
rect 313967 -290387 314001 -289811
rect 314085 -290387 314119 -289811
rect 314203 -290387 314237 -289811
rect 314321 -290387 314355 -289811
rect 314439 -290387 314473 -289811
rect 314557 -290387 314591 -289811
rect 314675 -290387 314709 -289811
rect 314793 -290387 314827 -289811
rect 314911 -290387 314945 -289811
rect 315029 -290387 315063 -289811
rect 315147 -290387 315181 -289811
rect 315265 -290387 315299 -289811
rect 315383 -290387 315417 -289811
rect 315501 -290387 315535 -289811
rect 315619 -290387 315653 -289811
rect 315737 -290387 315771 -289811
rect 315855 -290387 315889 -289811
rect 315973 -290387 316007 -289811
rect 316091 -290387 316125 -289811
rect 316209 -290387 316243 -289811
rect 316327 -290387 316361 -289811
rect 316445 -290387 316479 -289811
rect 316563 -290387 316597 -289811
rect 316681 -290387 316715 -289811
rect 316799 -290387 316833 -289811
rect 316917 -290387 316951 -289811
rect 317035 -290387 317069 -289811
rect 317153 -290387 317187 -289811
rect 317271 -290387 317305 -289811
rect 317385 -290486 317419 -288876
rect 311353 -290582 317323 -290548
rect 311353 -290864 317323 -290830
rect 311257 -292536 311291 -290926
rect 311371 -291601 311405 -291025
rect 311489 -291601 311523 -291025
rect 311607 -291601 311641 -291025
rect 311725 -291601 311759 -291025
rect 311843 -291601 311877 -291025
rect 311961 -291601 311995 -291025
rect 312079 -291601 312113 -291025
rect 312197 -291601 312231 -291025
rect 312315 -291601 312349 -291025
rect 312433 -291601 312467 -291025
rect 312551 -291601 312585 -291025
rect 312669 -291601 312703 -291025
rect 312787 -291601 312821 -291025
rect 312905 -291601 312939 -291025
rect 313023 -291601 313057 -291025
rect 313141 -291601 313175 -291025
rect 313259 -291601 313293 -291025
rect 313377 -291601 313411 -291025
rect 313495 -291601 313529 -291025
rect 313613 -291601 313647 -291025
rect 313731 -291601 313765 -291025
rect 313849 -291601 313883 -291025
rect 313967 -291601 314001 -291025
rect 314085 -291601 314119 -291025
rect 314203 -291601 314237 -291025
rect 314321 -291601 314355 -291025
rect 314439 -291601 314473 -291025
rect 314557 -291601 314591 -291025
rect 314675 -291601 314709 -291025
rect 314793 -291601 314827 -291025
rect 314911 -291601 314945 -291025
rect 315029 -291601 315063 -291025
rect 315147 -291601 315181 -291025
rect 315265 -291601 315299 -291025
rect 315383 -291601 315417 -291025
rect 315501 -291601 315535 -291025
rect 315619 -291601 315653 -291025
rect 315737 -291601 315771 -291025
rect 315855 -291601 315889 -291025
rect 315973 -291601 316007 -291025
rect 316091 -291601 316125 -291025
rect 316209 -291601 316243 -291025
rect 316327 -291601 316361 -291025
rect 316445 -291601 316479 -291025
rect 316563 -291601 316597 -291025
rect 316681 -291601 316715 -291025
rect 316799 -291601 316833 -291025
rect 316917 -291601 316951 -291025
rect 317035 -291601 317069 -291025
rect 317153 -291601 317187 -291025
rect 317271 -291601 317305 -291025
rect 311371 -292437 311405 -291861
rect 311489 -292437 311523 -291861
rect 311607 -292437 311641 -291861
rect 311725 -292437 311759 -291861
rect 311843 -292437 311877 -291861
rect 311961 -292437 311995 -291861
rect 312079 -292437 312113 -291861
rect 312197 -292437 312231 -291861
rect 312315 -292437 312349 -291861
rect 312433 -292437 312467 -291861
rect 312551 -292437 312585 -291861
rect 312669 -292437 312703 -291861
rect 312787 -292437 312821 -291861
rect 312905 -292437 312939 -291861
rect 313023 -292437 313057 -291861
rect 313141 -292437 313175 -291861
rect 313259 -292437 313293 -291861
rect 313377 -292437 313411 -291861
rect 313495 -292437 313529 -291861
rect 313613 -292437 313647 -291861
rect 313731 -292437 313765 -291861
rect 313849 -292437 313883 -291861
rect 313967 -292437 314001 -291861
rect 314085 -292437 314119 -291861
rect 314203 -292437 314237 -291861
rect 314321 -292437 314355 -291861
rect 314439 -292437 314473 -291861
rect 314557 -292437 314591 -291861
rect 314675 -292437 314709 -291861
rect 314793 -292437 314827 -291861
rect 314911 -292437 314945 -291861
rect 315029 -292437 315063 -291861
rect 315147 -292437 315181 -291861
rect 315265 -292437 315299 -291861
rect 315383 -292437 315417 -291861
rect 315501 -292437 315535 -291861
rect 315619 -292437 315653 -291861
rect 315737 -292437 315771 -291861
rect 315855 -292437 315889 -291861
rect 315973 -292437 316007 -291861
rect 316091 -292437 316125 -291861
rect 316209 -292437 316243 -291861
rect 316327 -292437 316361 -291861
rect 316445 -292437 316479 -291861
rect 316563 -292437 316597 -291861
rect 316681 -292437 316715 -291861
rect 316799 -292437 316833 -291861
rect 316917 -292437 316951 -291861
rect 317035 -292437 317069 -291861
rect 317153 -292437 317187 -291861
rect 317271 -292437 317305 -291861
rect 317385 -292536 317419 -290926
rect 311353 -292632 317323 -292598
rect 311607 -293651 311641 -293075
rect 311725 -293651 311759 -293075
rect 311843 -293651 311877 -293075
rect 311961 -293651 311995 -293075
rect 312079 -293651 312113 -293075
rect 312197 -293651 312231 -293075
rect 312315 -293651 312349 -293075
rect 312433 -293651 312467 -293075
rect 312551 -293651 312585 -293075
rect 312669 -293651 312703 -293075
rect 312787 -293651 312821 -293075
rect 312905 -293651 312939 -293075
rect 313023 -293651 313057 -293075
rect 313141 -293651 313175 -293075
rect 313259 -293651 313293 -293075
rect 313377 -293651 313411 -293075
rect 313495 -293651 313529 -293075
rect 313613 -293651 313647 -293075
rect 313731 -293651 313765 -293075
rect 313849 -293651 313883 -293075
rect 313967 -293651 314001 -293075
rect 314085 -293651 314119 -293075
rect 314203 -293651 314237 -293075
rect 314321 -293651 314355 -293075
rect 314439 -293651 314473 -293075
rect 314557 -293651 314591 -293075
rect 314675 -293651 314709 -293075
rect 314793 -293651 314827 -293075
rect 314911 -293651 314945 -293075
rect 315029 -293651 315063 -293075
rect 315147 -293651 315181 -293075
rect 315265 -293651 315299 -293075
rect 315383 -293651 315417 -293075
rect 315501 -293651 315535 -293075
rect 315619 -293651 315653 -293075
rect 315737 -293651 315771 -293075
rect 315855 -293651 315889 -293075
rect 315973 -293651 316007 -293075
rect 316091 -293651 316125 -293075
rect 316209 -293651 316243 -293075
rect 316327 -293651 316361 -293075
rect 316445 -293651 316479 -293075
rect 316563 -293651 316597 -293075
rect 316681 -293651 316715 -293075
rect 316799 -293651 316833 -293075
rect 316917 -293651 316951 -293075
rect 317035 -293651 317069 -293075
rect 317153 -293651 317187 -293075
rect 317271 -293651 317305 -293075
rect 311371 -294487 311405 -293911
rect 311489 -294487 311523 -293911
rect 311607 -294487 311641 -293911
rect 311725 -294487 311759 -293911
rect 311843 -294487 311877 -293911
rect 311961 -294487 311995 -293911
rect 312079 -294487 312113 -293911
rect 312197 -294487 312231 -293911
rect 312315 -294487 312349 -293911
rect 312433 -294487 312467 -293911
rect 312551 -294487 312585 -293911
rect 312669 -294487 312703 -293911
rect 312787 -294487 312821 -293911
rect 312905 -294487 312939 -293911
rect 313023 -294487 313057 -293911
rect 313141 -294487 313175 -293911
rect 313259 -294487 313293 -293911
rect 313377 -294487 313411 -293911
rect 313495 -294487 313529 -293911
rect 313613 -294487 313647 -293911
rect 313731 -294487 313765 -293911
rect 313849 -294487 313883 -293911
rect 313967 -294487 314001 -293911
rect 314085 -294487 314119 -293911
rect 314203 -294487 314237 -293911
rect 314321 -294487 314355 -293911
rect 314439 -294487 314473 -293911
rect 314557 -294487 314591 -293911
rect 314675 -294487 314709 -293911
rect 314793 -294487 314827 -293911
rect 314911 -294487 314945 -293911
rect 315029 -294487 315063 -293911
rect 315147 -294487 315181 -293911
rect 315265 -294487 315299 -293911
rect 315383 -294487 315417 -293911
rect 315501 -294487 315535 -293911
rect 315619 -294487 315653 -293911
rect 315737 -294487 315771 -293911
rect 315855 -294487 315889 -293911
rect 315973 -294487 316007 -293911
rect 316091 -294487 316125 -293911
rect 316209 -294487 316243 -293911
rect 316327 -294487 316361 -293911
rect 316445 -294487 316479 -293911
rect 316563 -294487 316597 -293911
rect 316681 -294487 316715 -293911
rect 316799 -294487 316833 -293911
rect 316917 -294487 316951 -293911
rect 317035 -294487 317069 -293911
rect 317153 -294487 317187 -293911
rect 317271 -294487 317305 -293911
rect 312673 -295894 312707 -295318
rect 312791 -295894 312825 -295318
rect 312909 -295894 312943 -295318
rect 313027 -295894 313061 -295318
rect 313145 -295894 313179 -295318
rect 313263 -295894 313297 -295318
rect 313381 -295894 313415 -295318
rect 313499 -295894 313533 -295318
rect 313617 -295894 313651 -295318
rect 313735 -295894 313769 -295318
rect 313853 -295894 313887 -295318
rect 313971 -295894 314005 -295318
rect 314089 -295894 314123 -295318
rect 314207 -295894 314241 -295318
rect 314435 -295894 314469 -295318
rect 314553 -295894 314587 -295318
rect 314671 -295894 314705 -295318
rect 314789 -295894 314823 -295318
rect 314907 -295894 314941 -295318
rect 315025 -295894 315059 -295318
rect 315143 -295894 315177 -295318
rect 315261 -295894 315295 -295318
rect 315379 -295894 315413 -295318
rect 315497 -295894 315531 -295318
rect 315615 -295894 315649 -295318
rect 315733 -295894 315767 -295318
rect 315851 -295894 315885 -295318
rect 315969 -295894 316003 -295318
rect 316087 -295894 316121 -295318
rect 316205 -295894 316239 -295318
rect 317298 -295696 317332 -295390
rect 317412 -295606 317446 -295480
rect 317500 -295606 317534 -295480
rect 317614 -295696 317648 -295390
rect 317728 -295606 317762 -295480
rect 317816 -295606 317850 -295480
rect 317930 -295696 317964 -295390
rect 318044 -295606 318078 -295480
rect 318132 -295606 318166 -295480
rect 318246 -295696 318280 -295390
rect 318360 -295606 318394 -295480
rect 318448 -295606 318482 -295480
rect 318562 -295696 318596 -295390
rect 318676 -295606 318710 -295480
rect 318764 -295606 318798 -295480
rect 318878 -295696 318912 -295390
rect 312437 -296712 312471 -296136
rect 312555 -296712 312589 -296136
rect 312673 -296712 312707 -296136
rect 312791 -296712 312825 -296136
rect 312909 -296712 312943 -296136
rect 313027 -296712 313061 -296136
rect 313145 -296712 313179 -296136
rect 313263 -296712 313297 -296136
rect 313381 -296712 313415 -296136
rect 313499 -296712 313533 -296136
rect 313617 -296712 313651 -296136
rect 313735 -296712 313769 -296136
rect 313853 -296712 313887 -296136
rect 313971 -296712 314005 -296136
rect 314089 -296712 314123 -296136
rect 314207 -296712 314241 -296136
rect 314435 -296712 314469 -296136
rect 314553 -296712 314587 -296136
rect 314671 -296712 314705 -296136
rect 314789 -296712 314823 -296136
rect 314907 -296712 314941 -296136
rect 315025 -296712 315059 -296136
rect 315143 -296712 315177 -296136
rect 315261 -296712 315295 -296136
rect 315379 -296712 315413 -296136
rect 315497 -296712 315531 -296136
rect 315615 -296712 315649 -296136
rect 315733 -296712 315767 -296136
rect 315851 -296712 315885 -296136
rect 315969 -296712 316003 -296136
rect 316087 -296712 316121 -296136
rect 316205 -296712 316239 -296136
rect 319095 -296194 319129 -295318
rect 319243 -296194 319277 -295318
rect 319391 -296194 319425 -295318
rect 319539 -296194 319573 -295318
rect 319687 -296194 319721 -295318
rect 319835 -296194 319869 -295318
rect 319983 -296194 320017 -295318
rect 320131 -296194 320165 -295318
rect 320279 -296194 320313 -295318
rect 320427 -296194 320461 -295318
rect 320575 -296194 320609 -295318
rect 320723 -296194 320757 -295318
rect 320871 -296194 320905 -295318
rect 321019 -296194 321053 -295318
rect 321167 -296194 321201 -295318
rect 321315 -296194 321349 -295318
rect 321463 -296194 321497 -295318
rect 321611 -296194 321645 -295318
rect 321759 -296194 321793 -295318
rect 321907 -296194 321941 -295318
rect 322055 -296194 322089 -295318
rect 322203 -296194 322237 -295318
rect 322351 -296194 322385 -295318
rect 322499 -296194 322533 -295318
rect 322647 -296194 322681 -295318
rect 322795 -296194 322829 -295318
rect 322943 -296194 322977 -295318
rect 323091 -296194 323125 -295318
rect 323239 -296194 323273 -295318
rect 323387 -296194 323421 -295318
rect 323535 -296194 323569 -295318
rect 323683 -296194 323717 -295318
rect 323831 -296194 323865 -295318
rect 323979 -296194 324013 -295318
rect 324127 -296194 324161 -295318
rect 324275 -296194 324309 -295318
rect 324423 -296194 324457 -295318
rect 324571 -296194 324605 -295318
rect 324719 -296194 324753 -295318
rect 324867 -296194 324901 -295318
rect 325015 -296194 325049 -295318
rect 325163 -296194 325197 -295318
rect 325311 -296194 325345 -295318
rect 325459 -296194 325493 -295318
rect 325607 -296194 325641 -295318
rect 325755 -296194 325789 -295318
rect 325903 -296194 325937 -295318
rect 326051 -296194 326085 -295318
rect 326199 -296194 326233 -295318
rect 326347 -296194 326381 -295318
rect 326495 -296194 326529 -295318
rect 326643 -296194 326677 -295318
rect 326791 -296194 326825 -295318
rect 326939 -296194 326973 -295318
rect 327087 -296194 327121 -295318
rect 327235 -296194 327269 -295318
rect 327383 -296194 327417 -295318
rect 327531 -296194 327565 -295318
rect 327679 -296194 327713 -295318
rect 327827 -296194 327861 -295318
rect 327975 -296194 328009 -295318
rect 328123 -296194 328157 -295318
rect 328271 -296194 328305 -295318
rect 328419 -296194 328453 -295318
rect 328567 -296194 328601 -295318
rect 328715 -296194 328749 -295318
rect 328863 -296194 328897 -295318
rect 329011 -296194 329045 -295318
rect 329159 -296194 329193 -295318
rect 329307 -296194 329341 -295318
rect 329455 -296194 329489 -295318
rect 329603 -296194 329637 -295318
rect 329751 -296194 329785 -295318
rect 329899 -296194 329933 -295318
rect 330195 -296194 330229 -295318
rect 319305 -296278 319363 -296244
rect 319453 -296278 319511 -296244
rect 319601 -296278 319659 -296244
rect 319749 -296278 319807 -296244
rect 319897 -296278 319955 -296244
rect 320045 -296278 320103 -296244
rect 320193 -296278 320251 -296244
rect 320341 -296278 320399 -296244
rect 320489 -296278 320547 -296244
rect 320637 -296278 320695 -296244
rect 320785 -296278 320843 -296244
rect 320933 -296278 320991 -296244
rect 321081 -296278 321139 -296244
rect 321229 -296278 321287 -296244
rect 321377 -296278 321435 -296244
rect 321525 -296278 321583 -296244
rect 321673 -296278 321731 -296244
rect 321821 -296278 321879 -296244
rect 321969 -296278 322027 -296244
rect 322117 -296278 322175 -296244
rect 322265 -296278 322323 -296244
rect 322413 -296278 322471 -296244
rect 322561 -296278 322619 -296244
rect 322709 -296278 322767 -296244
rect 322857 -296278 322915 -296244
rect 323005 -296278 323063 -296244
rect 323153 -296278 323211 -296244
rect 323301 -296278 323359 -296244
rect 323449 -296278 323507 -296244
rect 323597 -296278 323655 -296244
rect 323745 -296278 323803 -296244
rect 323893 -296278 323951 -296244
rect 324041 -296278 324099 -296244
rect 324189 -296278 324247 -296244
rect 324337 -296278 324395 -296244
rect 324485 -296278 324543 -296244
rect 324633 -296278 324691 -296244
rect 324781 -296278 324839 -296244
rect 324929 -296278 324987 -296244
rect 325077 -296278 325135 -296244
rect 325225 -296278 325283 -296244
rect 325373 -296278 325431 -296244
rect 325521 -296278 325579 -296244
rect 325669 -296278 325727 -296244
rect 325817 -296278 325875 -296244
rect 325965 -296278 326023 -296244
rect 326113 -296278 326171 -296244
rect 326261 -296278 326319 -296244
rect 326409 -296278 326467 -296244
rect 326557 -296278 326615 -296244
rect 326705 -296278 326763 -296244
rect 326853 -296278 326911 -296244
rect 327001 -296278 327059 -296244
rect 327149 -296278 327207 -296244
rect 327297 -296278 327355 -296244
rect 327445 -296278 327503 -296244
rect 327593 -296278 327651 -296244
rect 327741 -296278 327799 -296244
rect 327889 -296278 327947 -296244
rect 328037 -296278 328095 -296244
rect 328185 -296278 328243 -296244
rect 328333 -296278 328391 -296244
rect 328481 -296278 328539 -296244
rect 328629 -296278 328687 -296244
rect 328777 -296278 328835 -296244
rect 328925 -296278 328983 -296244
rect 329073 -296278 329131 -296244
rect 329221 -296278 329279 -296244
rect 329369 -296278 329427 -296244
rect 329517 -296278 329575 -296244
rect 329665 -296278 329723 -296244
rect 329813 -296278 329871 -296244
rect 329961 -296278 330019 -296244
rect 330109 -296278 330167 -296244
rect 319305 -296386 319363 -296352
rect 319453 -296386 319511 -296352
rect 319601 -296386 319659 -296352
rect 319749 -296386 319807 -296352
rect 319897 -296386 319955 -296352
rect 320045 -296386 320103 -296352
rect 320193 -296386 320251 -296352
rect 320341 -296386 320399 -296352
rect 320489 -296386 320547 -296352
rect 320637 -296386 320695 -296352
rect 320785 -296386 320843 -296352
rect 320933 -296386 320991 -296352
rect 321081 -296386 321139 -296352
rect 321229 -296386 321287 -296352
rect 321377 -296386 321435 -296352
rect 321525 -296386 321583 -296352
rect 321673 -296386 321731 -296352
rect 321821 -296386 321879 -296352
rect 321969 -296386 322027 -296352
rect 322117 -296386 322175 -296352
rect 322265 -296386 322323 -296352
rect 322413 -296386 322471 -296352
rect 322561 -296386 322619 -296352
rect 322709 -296386 322767 -296352
rect 322857 -296386 322915 -296352
rect 323005 -296386 323063 -296352
rect 323153 -296386 323211 -296352
rect 323301 -296386 323359 -296352
rect 323449 -296386 323507 -296352
rect 323597 -296386 323655 -296352
rect 323745 -296386 323803 -296352
rect 323893 -296386 323951 -296352
rect 324041 -296386 324099 -296352
rect 324189 -296386 324247 -296352
rect 324337 -296386 324395 -296352
rect 324485 -296386 324543 -296352
rect 324633 -296386 324691 -296352
rect 324781 -296386 324839 -296352
rect 324929 -296386 324987 -296352
rect 325077 -296386 325135 -296352
rect 325225 -296386 325283 -296352
rect 325373 -296386 325431 -296352
rect 325521 -296386 325579 -296352
rect 325669 -296386 325727 -296352
rect 325817 -296386 325875 -296352
rect 325965 -296386 326023 -296352
rect 326113 -296386 326171 -296352
rect 326261 -296386 326319 -296352
rect 326409 -296386 326467 -296352
rect 326557 -296386 326615 -296352
rect 326705 -296386 326763 -296352
rect 326853 -296386 326911 -296352
rect 327001 -296386 327059 -296352
rect 327149 -296386 327207 -296352
rect 327297 -296386 327355 -296352
rect 327445 -296386 327503 -296352
rect 327593 -296386 327651 -296352
rect 327741 -296386 327799 -296352
rect 327889 -296386 327947 -296352
rect 328037 -296386 328095 -296352
rect 328185 -296386 328243 -296352
rect 328333 -296386 328391 -296352
rect 328481 -296386 328539 -296352
rect 328629 -296386 328687 -296352
rect 328777 -296386 328835 -296352
rect 328925 -296386 328983 -296352
rect 329073 -296386 329131 -296352
rect 329221 -296386 329279 -296352
rect 329369 -296386 329427 -296352
rect 329517 -296386 329575 -296352
rect 329665 -296386 329723 -296352
rect 329813 -296386 329871 -296352
rect 329961 -296386 330019 -296352
rect 330109 -296386 330167 -296352
rect 319095 -297312 319129 -296436
rect 319243 -297312 319277 -296436
rect 319391 -297312 319425 -296436
rect 319539 -297312 319573 -296436
rect 319687 -297312 319721 -296436
rect 319835 -297312 319869 -296436
rect 319983 -297312 320017 -296436
rect 320131 -297312 320165 -296436
rect 320279 -297312 320313 -296436
rect 320427 -297312 320461 -296436
rect 320575 -297312 320609 -296436
rect 320723 -297312 320757 -296436
rect 320871 -297312 320905 -296436
rect 321019 -297312 321053 -296436
rect 321167 -297312 321201 -296436
rect 321315 -297312 321349 -296436
rect 321463 -297312 321497 -296436
rect 321611 -297312 321645 -296436
rect 321759 -297312 321793 -296436
rect 321907 -297312 321941 -296436
rect 322055 -297312 322089 -296436
rect 322203 -297312 322237 -296436
rect 322351 -297312 322385 -296436
rect 322499 -297312 322533 -296436
rect 322647 -297312 322681 -296436
rect 322795 -297312 322829 -296436
rect 322943 -297312 322977 -296436
rect 323091 -297312 323125 -296436
rect 323239 -297312 323273 -296436
rect 323387 -297312 323421 -296436
rect 323535 -297312 323569 -296436
rect 323683 -297312 323717 -296436
rect 323831 -297312 323865 -296436
rect 323979 -297312 324013 -296436
rect 324127 -297312 324161 -296436
rect 324275 -297312 324309 -296436
rect 324423 -297312 324457 -296436
rect 324571 -297312 324605 -296436
rect 324719 -297312 324753 -296436
rect 324867 -297312 324901 -296436
rect 325015 -297312 325049 -296436
rect 325163 -297312 325197 -296436
rect 325311 -297312 325345 -296436
rect 325459 -297312 325493 -296436
rect 325607 -297312 325641 -296436
rect 325755 -297312 325789 -296436
rect 325903 -297312 325937 -296436
rect 326051 -297312 326085 -296436
rect 326199 -297312 326233 -296436
rect 326347 -297312 326381 -296436
rect 326495 -297312 326529 -296436
rect 326643 -297312 326677 -296436
rect 326791 -297312 326825 -296436
rect 326939 -297312 326973 -296436
rect 327087 -297312 327121 -296436
rect 327235 -297312 327269 -296436
rect 327383 -297312 327417 -296436
rect 327531 -297312 327565 -296436
rect 327679 -297312 327713 -296436
rect 327827 -297312 327861 -296436
rect 327975 -297312 328009 -296436
rect 328123 -297312 328157 -296436
rect 328271 -297312 328305 -296436
rect 328419 -297312 328453 -296436
rect 328567 -297312 328601 -296436
rect 328715 -297312 328749 -296436
rect 328863 -297312 328897 -296436
rect 329011 -297312 329045 -296436
rect 329159 -297312 329193 -296436
rect 329307 -297312 329341 -296436
rect 329455 -297312 329489 -296436
rect 329603 -297312 329637 -296436
rect 329751 -297312 329785 -296436
rect 329899 -297312 329933 -296436
use opamp_wrapper  opamp_wrapper_0 ~/CMOS/TopMetalSe-OpenMPW6/mag
timestamp 1654646295
transform 1 0 308280 0 1 -296491
box -2280 -1609 26995 13665
use 100pixel_array  100pixel_array_0 ~/CMOS/TopMetalSe-OpenMPW6/mag
timestamp 1654709558
transform 1 0 3000 0 1 -1400
box -3000 -298600 300740 5750
use bias  bias_0 ~/CMOS/TopMetalSe-OpenMPW6/mag
timestamp 1654639008
transform 1 0 147210 0 1 7236
box 790 -2236 7180 -220
<< end >>
