magic
tech sky130A
magscale 1 2
timestamp 1663354353
<< metal1 >>
rect 143673 694385 144063 694391
rect 7012 688094 7332 688100
rect 7332 687774 137381 688094
rect 7012 687768 7332 687774
rect 1919 686010 4379 686016
rect 4379 684464 25503 686010
rect 4379 683550 26802 684464
rect 1919 683544 4379 683550
rect 23043 682004 26802 683550
rect 29262 682004 29268 684464
rect 1919 678115 4379 678121
rect 4379 675655 26510 678115
rect 28970 675655 28976 678115
rect 1919 675649 4379 675655
rect 137061 675252 137381 687774
rect 137061 674899 137381 674932
rect 143673 675660 144063 693995
rect 143673 675270 146631 675660
rect 140626 673664 140632 673734
rect 140702 673664 140708 673734
rect 1919 672893 4379 672899
rect 4379 670433 26343 672893
rect 28803 670433 28809 672893
rect 143673 670736 144063 675270
rect 396231 674830 396401 674836
rect 364539 674660 396231 674830
rect 155835 674103 156205 674109
rect 152191 673733 155835 674103
rect 156205 673733 156980 674103
rect 155835 673727 156205 673733
rect 154966 673475 154972 673585
rect 155082 673475 155088 673585
rect 154972 672526 155082 673475
rect 364863 673430 365033 674660
rect 396231 674654 396401 674660
rect 177593 673260 365033 673430
rect 178695 672526 178865 673260
rect 154972 672416 178922 672526
rect 1919 670427 4379 670433
rect 143673 670340 144063 670346
rect 13647 669652 50982 669972
rect 13647 657326 13967 669652
rect 50662 664728 50982 669652
rect 53663 664728 53983 664734
rect 50662 664408 53663 664728
rect 53663 664402 53983 664408
rect 13647 657000 13967 657006
rect 364863 369194 365033 673260
rect 397829 665127 398129 665133
rect 397829 647181 398129 664827
rect 380293 427751 396171 428041
rect 370560 377472 414098 377762
rect 414388 377472 414394 377762
rect 370560 370704 370850 377472
rect 373560 376785 413990 377075
rect 414280 376785 414286 377075
rect 373560 370704 373850 376785
rect 376560 375918 414243 376208
rect 414533 375918 414539 376208
rect 376560 370704 376850 375918
rect 379560 374363 414026 374653
rect 414316 374363 414322 374653
rect 379560 370704 379850 374363
rect 382560 373764 413994 374054
rect 414284 373764 414290 374054
rect 382560 370704 382850 373764
rect 385560 372904 414352 373194
rect 414642 372904 414648 373194
rect 385560 370704 385850 372904
rect 388560 372187 414245 372477
rect 414535 372187 414541 372477
rect 388560 370704 388850 372187
rect 391560 371542 414352 371832
rect 414642 371542 414648 371832
rect 391560 370704 391850 371542
rect 394587 371295 394877 371329
rect 394587 371005 414776 371295
rect 415066 371005 415072 371295
rect 369997 370414 393348 370704
rect 394587 370414 394877 371005
rect 396070 370414 413772 370704
rect 414062 370414 414068 370704
rect 364863 369024 367371 369194
rect 370011 357564 394617 357864
rect 396287 357564 397617 357864
rect 1919 353279 4379 353285
rect 4379 350819 26650 353279
rect 29110 350819 29116 353279
rect 1919 350813 4379 350819
rect 1919 348750 4379 348756
rect 4379 346290 26576 348750
rect 29036 346290 29042 348750
rect 1919 346284 4379 346290
rect 55307 345756 55627 345762
rect 58307 345756 58627 345762
rect 61307 345756 61627 345762
rect 64307 345756 64627 345762
rect 67307 345756 67627 345762
rect 70307 345756 70627 345762
rect 73307 345756 73627 345762
rect 76307 345756 76627 345762
rect 79307 345756 79627 345762
rect 82307 345756 82627 345762
rect 85307 345756 85627 345762
rect 88307 345756 88627 345762
rect 91307 345756 91627 345762
rect 94307 345756 94627 345762
rect 97307 345756 97627 345762
rect 100307 345756 100627 345762
rect 103307 345756 103627 345762
rect 106307 345756 106627 345762
rect 109307 345756 109627 345762
rect 112307 345756 112627 345762
rect 115307 345756 115627 345762
rect 118307 345756 118627 345762
rect 121307 345756 121627 345762
rect 124307 345756 124627 345762
rect 127307 345756 127627 345762
rect 130307 345756 130627 345762
rect 133307 345756 133627 345762
rect 136307 345756 136627 345762
rect 139307 345756 139627 345762
rect 142307 345756 142627 345762
rect 145307 345756 145627 345762
rect 148307 345756 148627 345762
rect 151307 345756 151627 345762
rect 154307 345756 154627 345762
rect 157307 345756 157627 345762
rect 160307 345756 160627 345762
rect 163307 345756 163627 345762
rect 166307 345756 166627 345762
rect 169307 345756 169627 345762
rect 172307 345756 172627 345762
rect 175307 345756 175627 345762
rect 178307 345756 178627 345762
rect 181307 345756 181627 345762
rect 184307 345756 184627 345762
rect 187307 345756 187627 345762
rect 190307 345756 190627 345762
rect 193307 345756 193627 345762
rect 196307 345756 196627 345762
rect 199307 345756 199627 345762
rect 202307 345756 202627 345762
rect 205307 345756 205627 345762
rect 208307 345756 208627 345762
rect 211307 345756 211627 345762
rect 214307 345756 214627 345762
rect 217307 345756 217627 345762
rect 220307 345756 220627 345762
rect 223307 345756 223627 345762
rect 226307 345756 226627 345762
rect 229307 345756 229627 345762
rect 232307 345756 232627 345762
rect 235307 345756 235627 345762
rect 238307 345756 238627 345762
rect 241307 345756 241627 345762
rect 244307 345756 244627 345762
rect 247307 345756 247627 345762
rect 250307 345756 250627 345762
rect 253307 345756 253627 345762
rect 256307 345756 256627 345762
rect 259307 345756 259627 345762
rect 262307 345756 262627 345762
rect 265307 345756 265627 345762
rect 268307 345756 268627 345762
rect 271307 345756 271627 345762
rect 274307 345756 274627 345762
rect 277307 345756 277627 345762
rect 280307 345756 280627 345762
rect 283307 345756 283627 345762
rect 286307 345756 286627 345762
rect 289307 345756 289627 345762
rect 292307 345756 292627 345762
rect 295307 345756 295627 345762
rect 298307 345756 298627 345762
rect 301307 345756 301627 345762
rect 304307 345756 304627 345762
rect 307307 345756 307627 345762
rect 310307 345756 310627 345762
rect 313307 345756 313627 345762
rect 316307 345756 316627 345762
rect 319307 345756 319627 345762
rect 325307 345756 325627 345762
rect 328307 345756 328627 345762
rect 331307 345756 331627 345762
rect 334307 345756 334627 345762
rect 337307 345756 337627 345762
rect 340307 345756 340627 345762
rect 343307 345756 343627 345762
rect 346307 345756 346627 345762
rect 349307 345756 349627 345762
rect 352307 345756 352627 345762
rect 355307 345756 355627 345762
rect 358307 345756 358627 345762
rect 55301 345436 55307 345756
rect 55627 345436 55633 345756
rect 58301 345436 58307 345756
rect 58627 345436 58633 345756
rect 61301 345436 61307 345756
rect 61627 345436 61633 345756
rect 64301 345436 64307 345756
rect 64627 345436 64633 345756
rect 67301 345436 67307 345756
rect 67627 345436 67633 345756
rect 70301 345436 70307 345756
rect 70627 345436 70633 345756
rect 73301 345436 73307 345756
rect 73627 345436 73633 345756
rect 76301 345436 76307 345756
rect 76627 345436 76633 345756
rect 79301 345436 79307 345756
rect 79627 345436 79633 345756
rect 82301 345436 82307 345756
rect 82627 345436 82633 345756
rect 85301 345436 85307 345756
rect 85627 345436 85633 345756
rect 88301 345436 88307 345756
rect 88627 345436 88633 345756
rect 91301 345436 91307 345756
rect 91627 345436 91633 345756
rect 94301 345436 94307 345756
rect 94627 345436 94633 345756
rect 97301 345436 97307 345756
rect 97627 345436 97633 345756
rect 100301 345436 100307 345756
rect 100627 345436 100633 345756
rect 103301 345436 103307 345756
rect 103627 345436 103633 345756
rect 106301 345436 106307 345756
rect 106627 345436 106633 345756
rect 109301 345436 109307 345756
rect 109627 345436 109633 345756
rect 112301 345436 112307 345756
rect 112627 345436 112633 345756
rect 115301 345436 115307 345756
rect 115627 345436 115633 345756
rect 118301 345436 118307 345756
rect 118627 345436 118633 345756
rect 121301 345436 121307 345756
rect 121627 345436 121633 345756
rect 124301 345436 124307 345756
rect 124627 345436 124633 345756
rect 127301 345436 127307 345756
rect 127627 345436 127633 345756
rect 130301 345436 130307 345756
rect 130627 345436 130633 345756
rect 133301 345436 133307 345756
rect 133627 345436 133633 345756
rect 136301 345436 136307 345756
rect 136627 345436 136633 345756
rect 139301 345436 139307 345756
rect 139627 345436 139633 345756
rect 142301 345436 142307 345756
rect 142627 345436 142633 345756
rect 145301 345436 145307 345756
rect 145627 345436 145633 345756
rect 148301 345436 148307 345756
rect 148627 345436 148633 345756
rect 151301 345436 151307 345756
rect 151627 345436 151633 345756
rect 154301 345436 154307 345756
rect 154627 345436 154633 345756
rect 157301 345436 157307 345756
rect 157627 345436 157633 345756
rect 160301 345436 160307 345756
rect 160627 345436 160633 345756
rect 163301 345436 163307 345756
rect 163627 345436 163633 345756
rect 166301 345436 166307 345756
rect 166627 345436 166633 345756
rect 169301 345436 169307 345756
rect 169627 345436 169633 345756
rect 172301 345436 172307 345756
rect 172627 345436 172633 345756
rect 175301 345436 175307 345756
rect 175627 345436 175633 345756
rect 178301 345436 178307 345756
rect 178627 345436 178633 345756
rect 181301 345436 181307 345756
rect 181627 345436 181633 345756
rect 184301 345436 184307 345756
rect 184627 345436 184633 345756
rect 187301 345436 187307 345756
rect 187627 345436 187633 345756
rect 190301 345436 190307 345756
rect 190627 345436 190633 345756
rect 193301 345436 193307 345756
rect 193627 345436 193633 345756
rect 196301 345436 196307 345756
rect 196627 345436 196633 345756
rect 199301 345436 199307 345756
rect 199627 345436 199633 345756
rect 202301 345436 202307 345756
rect 202627 345436 202633 345756
rect 205301 345436 205307 345756
rect 205627 345436 205633 345756
rect 208301 345436 208307 345756
rect 208627 345436 208633 345756
rect 211301 345436 211307 345756
rect 211627 345436 211633 345756
rect 214301 345436 214307 345756
rect 214627 345436 214633 345756
rect 217301 345436 217307 345756
rect 217627 345436 217633 345756
rect 220301 345436 220307 345756
rect 220627 345436 220633 345756
rect 223301 345436 223307 345756
rect 223627 345436 223633 345756
rect 226301 345436 226307 345756
rect 226627 345436 226633 345756
rect 229301 345436 229307 345756
rect 229627 345436 229633 345756
rect 232301 345436 232307 345756
rect 232627 345436 232633 345756
rect 235301 345436 235307 345756
rect 235627 345436 235633 345756
rect 238301 345436 238307 345756
rect 238627 345436 238633 345756
rect 241301 345436 241307 345756
rect 241627 345436 241633 345756
rect 244301 345436 244307 345756
rect 244627 345436 244633 345756
rect 247301 345436 247307 345756
rect 247627 345436 247633 345756
rect 250301 345436 250307 345756
rect 250627 345436 250633 345756
rect 253301 345436 253307 345756
rect 253627 345436 253633 345756
rect 256301 345436 256307 345756
rect 256627 345436 256633 345756
rect 259301 345436 259307 345756
rect 259627 345436 259633 345756
rect 262301 345436 262307 345756
rect 262627 345436 262633 345756
rect 265301 345436 265307 345756
rect 265627 345436 265633 345756
rect 268301 345436 268307 345756
rect 268627 345436 268633 345756
rect 271301 345436 271307 345756
rect 271627 345436 271633 345756
rect 274301 345436 274307 345756
rect 274627 345436 274633 345756
rect 277301 345436 277307 345756
rect 277627 345436 277633 345756
rect 280301 345436 280307 345756
rect 280627 345436 280633 345756
rect 283301 345436 283307 345756
rect 283627 345436 283633 345756
rect 286301 345436 286307 345756
rect 286627 345436 286633 345756
rect 289301 345436 289307 345756
rect 289627 345436 289633 345756
rect 292301 345436 292307 345756
rect 292627 345436 292633 345756
rect 295301 345436 295307 345756
rect 295627 345436 295633 345756
rect 298301 345436 298307 345756
rect 298627 345436 298633 345756
rect 301301 345436 301307 345756
rect 301627 345436 301633 345756
rect 304301 345436 304307 345756
rect 304627 345436 304633 345756
rect 307301 345436 307307 345756
rect 307627 345436 307633 345756
rect 310301 345436 310307 345756
rect 310627 345436 310633 345756
rect 313301 345436 313307 345756
rect 313627 345436 313633 345756
rect 316301 345436 316307 345756
rect 316627 345436 316633 345756
rect 319301 345436 319307 345756
rect 319627 345436 319633 345756
rect 325301 345436 325307 345756
rect 325627 345436 325633 345756
rect 328301 345436 328307 345756
rect 328627 345436 328633 345756
rect 331301 345436 331307 345756
rect 331627 345436 331633 345756
rect 334301 345436 334307 345756
rect 334627 345436 334633 345756
rect 337301 345436 337307 345756
rect 337627 345436 337633 345756
rect 340301 345436 340307 345756
rect 340627 345436 340633 345756
rect 343301 345436 343307 345756
rect 343627 345436 343633 345756
rect 346301 345436 346307 345756
rect 346627 345436 346633 345756
rect 349301 345436 349307 345756
rect 349627 345436 349633 345756
rect 352301 345436 352307 345756
rect 352627 345436 352633 345756
rect 355301 345436 355307 345756
rect 355627 345436 355633 345756
rect 358301 345436 358307 345756
rect 358627 345436 358633 345756
rect 55307 345430 55627 345436
rect 58307 345430 58627 345436
rect 61307 345430 61627 345436
rect 64307 345430 64627 345436
rect 67307 345430 67627 345436
rect 70307 345430 70627 345436
rect 73307 345430 73627 345436
rect 76307 345430 76627 345436
rect 79307 345430 79627 345436
rect 82307 345430 82627 345436
rect 85307 345430 85627 345436
rect 88307 345430 88627 345436
rect 91307 345430 91627 345436
rect 94307 345430 94627 345436
rect 97307 345430 97627 345436
rect 100307 345430 100627 345436
rect 103307 345430 103627 345436
rect 106307 345430 106627 345436
rect 109307 345430 109627 345436
rect 112307 345430 112627 345436
rect 115307 345430 115627 345436
rect 118307 345430 118627 345436
rect 121307 345430 121627 345436
rect 124307 345430 124627 345436
rect 127307 345430 127627 345436
rect 130307 345430 130627 345436
rect 133307 345430 133627 345436
rect 136307 345430 136627 345436
rect 139307 345430 139627 345436
rect 142307 345430 142627 345436
rect 145307 345430 145627 345436
rect 148307 345430 148627 345436
rect 151307 345430 151627 345436
rect 154307 345430 154627 345436
rect 157307 345430 157627 345436
rect 160307 345430 160627 345436
rect 163307 345430 163627 345436
rect 166307 345430 166627 345436
rect 169307 345430 169627 345436
rect 172307 345430 172627 345436
rect 175307 345430 175627 345436
rect 178307 345430 178627 345436
rect 181307 345430 181627 345436
rect 184307 345430 184627 345436
rect 187307 345430 187627 345436
rect 190307 345430 190627 345436
rect 193307 345430 193627 345436
rect 196307 345430 196627 345436
rect 199307 345430 199627 345436
rect 202307 345430 202627 345436
rect 205307 345430 205627 345436
rect 208307 345430 208627 345436
rect 211307 345430 211627 345436
rect 214307 345430 214627 345436
rect 217307 345430 217627 345436
rect 220307 345430 220627 345436
rect 223307 345430 223627 345436
rect 226307 345430 226627 345436
rect 229307 345430 229627 345436
rect 232307 345430 232627 345436
rect 235307 345430 235627 345436
rect 238307 345430 238627 345436
rect 241307 345430 241627 345436
rect 244307 345430 244627 345436
rect 247307 345430 247627 345436
rect 250307 345430 250627 345436
rect 253307 345430 253627 345436
rect 256307 345430 256627 345436
rect 259307 345430 259627 345436
rect 262307 345430 262627 345436
rect 265307 345430 265627 345436
rect 268307 345430 268627 345436
rect 271307 345430 271627 345436
rect 274307 345430 274627 345436
rect 277307 345430 277627 345436
rect 280307 345430 280627 345436
rect 283307 345430 283627 345436
rect 286307 345430 286627 345436
rect 289307 345430 289627 345436
rect 292307 345430 292627 345436
rect 295307 345430 295627 345436
rect 298307 345430 298627 345436
rect 301307 345430 301627 345436
rect 304307 345430 304627 345436
rect 307307 345430 307627 345436
rect 310307 345430 310627 345436
rect 313307 345430 313627 345436
rect 316307 345430 316627 345436
rect 319307 345430 319627 345436
rect 325307 345430 325627 345436
rect 328307 345430 328627 345436
rect 331307 345430 331627 345436
rect 334307 345430 334627 345436
rect 337307 345430 337627 345436
rect 340307 345430 340627 345436
rect 343307 345430 343627 345436
rect 346307 345430 346627 345436
rect 349307 345430 349627 345436
rect 352307 345430 352627 345436
rect 355307 345430 355627 345436
rect 358307 345430 358627 345436
rect 1919 344240 4379 344246
rect 4379 341780 26576 344240
rect 29036 341780 29042 344240
rect 1919 341774 4379 341780
rect 372481 336904 372781 357564
rect 375481 336904 375781 357564
rect 378481 336904 378781 357564
rect 381481 336904 381781 357564
rect 384481 336904 384781 357564
rect 387481 336904 387781 357564
rect 390481 336904 390781 357564
rect 393481 336904 393781 357564
rect 396481 336904 396781 357564
rect 372475 336604 372481 336904
rect 372781 336604 372787 336904
rect 375475 336604 375481 336904
rect 375781 336604 375787 336904
rect 378475 336604 378481 336904
rect 378781 336604 378787 336904
rect 381475 336604 381481 336904
rect 381781 336604 381787 336904
rect 384475 336604 384481 336904
rect 384781 336604 384787 336904
rect 387475 336604 387481 336904
rect 387781 336604 387787 336904
rect 390475 336604 390481 336904
rect 390781 336604 390787 336904
rect 393475 336604 393481 336904
rect 393781 336604 393787 336904
rect 396475 336604 396481 336904
rect 396781 336604 396787 336904
rect 8362 261315 8493 261350
rect 64639 261315 64709 261321
rect 8362 261245 8387 261315
rect 8457 261245 64639 261315
rect 8362 261225 8493 261245
rect 64639 261239 64709 261245
rect 180921 207290 181211 207296
rect 176363 196612 176533 196618
rect 55930 193224 55936 193314
rect 56026 193224 56032 193314
rect 55936 189794 56026 193224
rect 176363 190937 176533 196442
rect 180921 192157 181211 207000
rect 183921 207290 184211 207296
rect 183921 192157 184211 207000
rect 186921 207290 187211 207296
rect 186921 192157 187211 207000
rect 189921 207290 190211 207296
rect 189921 192157 190211 207000
rect 192921 207290 193211 207296
rect 192921 192157 193211 207000
rect 195921 207290 196211 207296
rect 195921 192157 196211 207000
rect 198921 207290 199211 207296
rect 198921 192157 199211 207000
rect 201921 207290 202211 207296
rect 201921 192157 202211 207000
rect 204921 207290 205211 207296
rect 204921 192157 205211 207000
rect 176363 190767 177243 190937
rect 55936 189698 56026 189704
rect 175758 188178 175764 188348
rect 175934 188178 175940 188348
rect 175764 186637 175934 188178
rect 175764 186461 175934 186467
rect 180877 172819 181177 179607
rect 180877 172513 181177 172519
rect 183877 172819 184177 179607
rect 183877 172513 184177 172519
rect 186877 172819 187177 179607
rect 186877 172513 187177 172519
rect 189877 172819 190177 179607
rect 189877 172513 190177 172519
rect 192877 172819 193177 179607
rect 192877 172513 193177 172519
rect 195877 172819 196177 179607
rect 195877 172513 196177 172519
rect 198877 172819 199177 179607
rect 198877 172513 199177 172519
rect 201877 172819 202177 179607
rect 201877 172513 202177 172519
rect 204877 172819 205177 179607
rect 204877 172513 205177 172519
<< via1 >>
rect 143673 693995 144063 694385
rect 7012 687774 7332 688094
rect 1919 683550 4379 686010
rect 26802 682004 29262 684464
rect 1919 675655 4379 678115
rect 26510 675655 28970 678115
rect 137061 674932 137381 675252
rect 140632 673664 140702 673734
rect 1919 670433 4379 672893
rect 26343 670433 28803 672893
rect 396231 674660 396401 674830
rect 155835 673733 156205 674103
rect 154972 673475 155082 673585
rect 143673 670346 144063 670736
rect 53663 664408 53983 664728
rect 13647 657006 13967 657326
rect 397829 664827 398129 665127
rect 414098 377472 414388 377762
rect 413990 376785 414280 377075
rect 414243 375918 414533 376208
rect 414026 374363 414316 374653
rect 413994 373764 414284 374054
rect 414352 372904 414642 373194
rect 414245 372187 414535 372477
rect 414352 371542 414642 371832
rect 414776 371005 415066 371295
rect 413772 370414 414062 370704
rect 1919 350819 4379 353279
rect 26650 350819 29110 353279
rect 1919 346290 4379 348750
rect 26576 346290 29036 348750
rect 55307 345436 55627 345756
rect 58307 345436 58627 345756
rect 61307 345436 61627 345756
rect 64307 345436 64627 345756
rect 67307 345436 67627 345756
rect 70307 345436 70627 345756
rect 73307 345436 73627 345756
rect 76307 345436 76627 345756
rect 79307 345436 79627 345756
rect 82307 345436 82627 345756
rect 85307 345436 85627 345756
rect 88307 345436 88627 345756
rect 91307 345436 91627 345756
rect 94307 345436 94627 345756
rect 97307 345436 97627 345756
rect 100307 345436 100627 345756
rect 103307 345436 103627 345756
rect 106307 345436 106627 345756
rect 109307 345436 109627 345756
rect 112307 345436 112627 345756
rect 115307 345436 115627 345756
rect 118307 345436 118627 345756
rect 121307 345436 121627 345756
rect 124307 345436 124627 345756
rect 127307 345436 127627 345756
rect 130307 345436 130627 345756
rect 133307 345436 133627 345756
rect 136307 345436 136627 345756
rect 139307 345436 139627 345756
rect 142307 345436 142627 345756
rect 145307 345436 145627 345756
rect 148307 345436 148627 345756
rect 151307 345436 151627 345756
rect 154307 345436 154627 345756
rect 157307 345436 157627 345756
rect 160307 345436 160627 345756
rect 163307 345436 163627 345756
rect 166307 345436 166627 345756
rect 169307 345436 169627 345756
rect 172307 345436 172627 345756
rect 175307 345436 175627 345756
rect 178307 345436 178627 345756
rect 181307 345436 181627 345756
rect 184307 345436 184627 345756
rect 187307 345436 187627 345756
rect 190307 345436 190627 345756
rect 193307 345436 193627 345756
rect 196307 345436 196627 345756
rect 199307 345436 199627 345756
rect 202307 345436 202627 345756
rect 205307 345436 205627 345756
rect 208307 345436 208627 345756
rect 211307 345436 211627 345756
rect 214307 345436 214627 345756
rect 217307 345436 217627 345756
rect 220307 345436 220627 345756
rect 223307 345436 223627 345756
rect 226307 345436 226627 345756
rect 229307 345436 229627 345756
rect 232307 345436 232627 345756
rect 235307 345436 235627 345756
rect 238307 345436 238627 345756
rect 241307 345436 241627 345756
rect 244307 345436 244627 345756
rect 247307 345436 247627 345756
rect 250307 345436 250627 345756
rect 253307 345436 253627 345756
rect 256307 345436 256627 345756
rect 259307 345436 259627 345756
rect 262307 345436 262627 345756
rect 265307 345436 265627 345756
rect 268307 345436 268627 345756
rect 271307 345436 271627 345756
rect 274307 345436 274627 345756
rect 277307 345436 277627 345756
rect 280307 345436 280627 345756
rect 283307 345436 283627 345756
rect 286307 345436 286627 345756
rect 289307 345436 289627 345756
rect 292307 345436 292627 345756
rect 295307 345436 295627 345756
rect 298307 345436 298627 345756
rect 301307 345436 301627 345756
rect 304307 345436 304627 345756
rect 307307 345436 307627 345756
rect 310307 345436 310627 345756
rect 313307 345436 313627 345756
rect 316307 345436 316627 345756
rect 319307 345436 319627 345756
rect 325307 345436 325627 345756
rect 328307 345436 328627 345756
rect 331307 345436 331627 345756
rect 334307 345436 334627 345756
rect 337307 345436 337627 345756
rect 340307 345436 340627 345756
rect 343307 345436 343627 345756
rect 346307 345436 346627 345756
rect 349307 345436 349627 345756
rect 352307 345436 352627 345756
rect 355307 345436 355627 345756
rect 358307 345436 358627 345756
rect 1919 341780 4379 344240
rect 26576 341780 29036 344240
rect 372481 336604 372781 336904
rect 375481 336604 375781 336904
rect 378481 336604 378781 336904
rect 381481 336604 381781 336904
rect 384481 336604 384781 336904
rect 387481 336604 387781 336904
rect 390481 336604 390781 336904
rect 393481 336604 393781 336904
rect 396481 336604 396781 336904
rect 8387 261245 8457 261315
rect 64639 261245 64709 261315
rect 180921 207000 181211 207290
rect 176363 196442 176533 196612
rect 55936 193224 56026 193314
rect 183921 207000 184211 207290
rect 186921 207000 187211 207290
rect 189921 207000 190211 207290
rect 192921 207000 193211 207290
rect 195921 207000 196211 207290
rect 198921 207000 199211 207290
rect 201921 207000 202211 207290
rect 204921 207000 205211 207290
rect 55936 189704 56026 189794
rect 175764 188178 175934 188348
rect 175764 186467 175934 186637
rect 180877 172519 181177 172819
rect 183877 172519 184177 172819
rect 186877 172519 187177 172819
rect 189877 172519 190177 172819
rect 192877 172519 193177 172819
rect 195877 172519 196177 172819
rect 198877 172519 199177 172819
rect 201877 172519 202177 172819
rect 204877 172519 205177 172819
<< metal2 >>
rect 143673 694385 144063 694394
rect 143667 693995 143673 694385
rect 144063 693995 144069 694385
rect 143673 693986 144063 693995
rect 178455 689116 178515 689125
rect 145941 689061 178455 689111
rect 7017 688094 7327 688098
rect 7006 687774 7012 688094
rect 7332 687774 7338 688094
rect 7017 687770 7327 687774
rect 1924 686010 4374 686014
rect 1913 683550 1919 686010
rect 4379 683550 4385 686010
rect 28681 685548 140743 685553
rect 28677 685488 28686 685548
rect 28746 685488 140743 685548
rect 28681 685483 140743 685488
rect 26802 684464 29262 684470
rect 1924 683546 4374 683550
rect 26793 682004 26802 684464
rect 29262 682004 29271 684464
rect 26802 681998 29262 682004
rect 9021 680862 9121 680866
rect 9016 680857 49154 680862
rect 9016 680757 9021 680857
rect 9121 680757 49154 680857
rect 9016 680752 49154 680757
rect 9021 680748 9121 680752
rect 1924 678115 4374 678119
rect 26510 678115 28970 678121
rect 1913 675655 1919 678115
rect 4379 675655 4385 678115
rect 26501 675655 26510 678115
rect 28970 675655 28979 678115
rect 46334 676370 46444 680752
rect 69665 676370 69775 676379
rect 46334 676260 69665 676370
rect 1924 675651 4374 675655
rect 26510 675649 28970 675655
rect 1924 672893 4374 672897
rect 26343 672893 28803 672899
rect 1913 670433 1919 672893
rect 4379 670433 4385 672893
rect 26334 670433 26343 672893
rect 28803 670433 28812 672893
rect 1924 670429 4374 670433
rect 26343 670427 28803 670433
rect 46334 669571 46444 676260
rect 69665 676251 69775 676260
rect 137061 675252 137381 675261
rect 137055 674932 137061 675252
rect 137381 674932 137387 675252
rect 137061 674923 137381 674932
rect 140632 673767 140702 685483
rect 145941 674802 145991 689061
rect 178455 689047 178515 689056
rect 185338 687770 425014 687940
rect 145941 674752 146221 674802
rect 155835 674103 156205 674112
rect 140600 673734 140742 673767
rect 140600 673664 140632 673734
rect 140702 673664 140742 673734
rect 140600 673640 140742 673664
rect 147471 671904 147561 673735
rect 55827 671823 147561 671904
rect 55827 671794 147548 671823
rect 55827 671030 55937 671794
rect 147981 671172 148071 673745
rect 150421 673079 150531 673785
rect 152421 673585 152531 673785
rect 155829 673733 155835 674103
rect 156205 673733 156211 674103
rect 155835 673724 156205 673733
rect 154972 673585 155082 673591
rect 185338 673585 185508 687770
rect 396236 674830 396396 674834
rect 396225 674660 396231 674830
rect 396401 674660 396407 674830
rect 396236 674656 396396 674660
rect 231029 673585 231038 673684
rect 152412 673475 152421 673585
rect 152531 673475 154972 673585
rect 155082 673475 155098 673585
rect 155830 673475 231038 673585
rect 152431 673466 152531 673475
rect 154972 673469 155082 673475
rect 155846 673079 155956 673475
rect 231029 673374 231038 673475
rect 231348 673585 231357 673684
rect 231348 673475 241562 673585
rect 231348 673374 231357 673475
rect 150242 672969 155956 673079
rect 56588 671130 148395 671172
rect 56588 671070 140637 671130
rect 140697 671070 148395 671130
rect 56588 671062 148395 671070
rect 140637 671061 140697 671062
rect 147981 671023 148071 671062
rect 143673 670736 144063 670745
rect 143667 670346 143673 670736
rect 144063 670346 144069 670736
rect 143673 670337 144063 670346
rect 34058 667760 34368 667764
rect 18911 667440 18920 667760
rect 19240 667755 34373 667760
rect 19240 667445 34058 667755
rect 34368 667445 34373 667755
rect 19240 667440 34373 667445
rect 34058 667436 34368 667440
rect 397829 665127 398129 665136
rect 397823 664827 397829 665127
rect 398129 664827 398135 665127
rect 397829 664818 398129 664827
rect 34058 664760 34368 664764
rect 18911 664440 18920 664760
rect 19240 664755 34373 664760
rect 19240 664445 34058 664755
rect 34368 664445 34373 664755
rect 53668 664728 53978 664732
rect 19240 664440 34373 664445
rect 34058 664436 34368 664440
rect 53657 664408 53663 664728
rect 53983 664408 53989 664728
rect 53668 664404 53978 664408
rect 34058 661760 34368 661764
rect 18911 661440 18920 661760
rect 19240 661755 34373 661760
rect 19240 661445 34058 661755
rect 34368 661445 34373 661755
rect 19240 661440 34373 661445
rect 34058 661436 34368 661440
rect 34058 658760 34368 658764
rect 18911 658440 18920 658760
rect 19240 658755 34373 658760
rect 19240 658445 34058 658755
rect 34368 658445 34373 658755
rect 19240 658440 34373 658445
rect 34058 658436 34368 658440
rect 13638 657006 13647 657326
rect 13967 657006 13976 657326
rect 424844 656024 425014 687770
rect 436506 680010 436515 680180
rect 436685 680010 436694 680180
rect 424840 655864 424849 656024
rect 425009 655864 425018 656024
rect 424844 655859 425014 655864
rect 34058 655760 34368 655764
rect 18911 655440 18920 655760
rect 19240 655755 34373 655760
rect 19240 655445 34058 655755
rect 34368 655445 34373 655755
rect 19240 655440 34373 655445
rect 34058 655436 34368 655440
rect 34058 652760 34368 652764
rect 18911 652440 18920 652760
rect 19240 652755 34373 652760
rect 19240 652445 34058 652755
rect 34368 652445 34373 652755
rect 19240 652440 34373 652445
rect 34058 652436 34368 652440
rect 34058 649760 34368 649764
rect 18911 649440 18920 649760
rect 19240 649755 34373 649760
rect 19240 649445 34058 649755
rect 34368 649445 34373 649755
rect 19240 649440 34373 649445
rect 34058 649436 34368 649440
rect 34058 646760 34368 646764
rect 18911 646440 18920 646760
rect 19240 646755 34373 646760
rect 19240 646445 34058 646755
rect 34368 646445 34373 646755
rect 19240 646440 34373 646445
rect 34058 646436 34368 646440
rect 34058 643760 34368 643764
rect 18911 643440 18920 643760
rect 19240 643755 34373 643760
rect 19240 643445 34058 643755
rect 34368 643445 34373 643755
rect 19240 643440 34373 643445
rect 34058 643436 34368 643440
rect 34058 640760 34368 640764
rect 18911 640440 18920 640760
rect 19240 640755 34373 640760
rect 19240 640445 34058 640755
rect 34368 640445 34373 640755
rect 19240 640440 34373 640445
rect 34058 640436 34368 640440
rect 34058 637760 34368 637764
rect 18911 637440 18920 637760
rect 19240 637755 34373 637760
rect 19240 637445 34058 637755
rect 34368 637445 34373 637755
rect 19240 637440 34373 637445
rect 34058 637436 34368 637440
rect 34058 634760 34368 634764
rect 18911 634440 18920 634760
rect 19240 634755 34373 634760
rect 19240 634445 34058 634755
rect 34368 634445 34373 634755
rect 19240 634440 34373 634445
rect 34058 634436 34368 634440
rect 34058 631760 34368 631764
rect 18911 631440 18920 631760
rect 19240 631755 34373 631760
rect 19240 631445 34058 631755
rect 34368 631445 34373 631755
rect 19240 631440 34373 631445
rect 34058 631436 34368 631440
rect 428434 627989 430884 627993
rect 34058 625760 34368 625764
rect 18911 625440 18920 625760
rect 19240 625755 34373 625760
rect 19240 625445 34058 625755
rect 34368 625445 34373 625755
rect 404758 625529 404767 627989
rect 407227 627984 430889 627989
rect 407227 625534 428434 627984
rect 430884 625534 430889 627984
rect 407227 625529 430889 625534
rect 428434 625525 430884 625529
rect 19240 625440 34373 625445
rect 34058 625436 34368 625440
rect 34058 622760 34368 622764
rect 18911 622440 18920 622760
rect 19240 622755 34373 622760
rect 19240 622445 34058 622755
rect 34368 622445 34373 622755
rect 19240 622440 34373 622445
rect 34058 622436 34368 622440
rect 34058 619760 34368 619764
rect 18911 619440 18920 619760
rect 19240 619755 34373 619760
rect 19240 619445 34058 619755
rect 34368 619445 34373 619755
rect 19240 619440 34373 619445
rect 34058 619436 34368 619440
rect 34058 616760 34368 616764
rect 18911 616440 18920 616760
rect 19240 616755 34373 616760
rect 19240 616445 34058 616755
rect 34368 616445 34373 616755
rect 19240 616440 34373 616445
rect 34058 616436 34368 616440
rect 428429 615823 430879 615828
rect 428429 615819 430884 615823
rect 34058 613760 34368 613764
rect 18911 613440 18920 613760
rect 19240 613755 34373 613760
rect 19240 613445 34058 613755
rect 34368 613445 34373 613755
rect 19240 613440 34373 613445
rect 34058 613436 34368 613440
rect 404898 613359 404907 615819
rect 407367 613359 428429 615819
rect 430889 613359 430898 615819
rect 428429 613355 430884 613359
rect 428429 613350 430879 613355
rect 34058 610760 34368 610764
rect 18911 610440 18920 610760
rect 19240 610755 34373 610760
rect 19240 610445 34058 610755
rect 34368 610445 34373 610755
rect 19240 610440 34373 610445
rect 34058 610436 34368 610440
rect 34058 607760 34368 607764
rect 18911 607440 18920 607760
rect 19240 607755 34373 607760
rect 19240 607445 34058 607755
rect 34368 607445 34373 607755
rect 19240 607440 34373 607445
rect 34058 607436 34368 607440
rect 34058 604760 34368 604764
rect 18911 604440 18920 604760
rect 19240 604755 34373 604760
rect 19240 604445 34058 604755
rect 34368 604445 34373 604755
rect 19240 604440 34373 604445
rect 34058 604436 34368 604440
rect 428434 602180 430884 602184
rect 34058 601760 34368 601764
rect 18911 601440 18920 601760
rect 19240 601755 34373 601760
rect 19240 601445 34058 601755
rect 34368 601445 34373 601755
rect 19240 601440 34373 601445
rect 34058 601436 34368 601440
rect 404409 599720 404418 602180
rect 406878 602175 430889 602180
rect 406878 599725 428434 602175
rect 430884 599725 430889 602175
rect 406878 599720 430889 599725
rect 428434 599716 430884 599720
rect 34058 598760 34368 598764
rect 18911 598440 18920 598760
rect 19240 598755 34373 598760
rect 19240 598445 34058 598755
rect 34368 598445 34373 598755
rect 19240 598440 34373 598445
rect 34058 598436 34368 598440
rect 34058 595760 34368 595764
rect 18911 595440 18920 595760
rect 19240 595755 34373 595760
rect 19240 595445 34058 595755
rect 34368 595445 34373 595755
rect 19240 595440 34373 595445
rect 34058 595436 34368 595440
rect 34058 592760 34368 592764
rect 18911 592440 18920 592760
rect 19240 592755 34373 592760
rect 19240 592445 34058 592755
rect 34368 592445 34373 592755
rect 19240 592440 34373 592445
rect 34058 592436 34368 592440
rect 34058 589760 34368 589764
rect 18911 589440 18920 589760
rect 19240 589755 34373 589760
rect 19240 589445 34058 589755
rect 34368 589445 34373 589755
rect 19240 589440 34373 589445
rect 34058 589436 34368 589440
rect 428434 587353 430884 587357
rect 34058 586760 34368 586764
rect 18911 586440 18920 586760
rect 19240 586755 34373 586760
rect 19240 586445 34058 586755
rect 34368 586445 34373 586755
rect 19240 586440 34373 586445
rect 34058 586436 34368 586440
rect 403709 584893 403718 587353
rect 406178 587348 430889 587353
rect 406178 584898 428434 587348
rect 430884 584898 430889 587348
rect 406178 584893 430889 584898
rect 428434 584889 430884 584893
rect 34058 583760 34368 583764
rect 18911 583440 18920 583760
rect 19240 583755 34373 583760
rect 19240 583445 34058 583755
rect 34368 583445 34373 583755
rect 19240 583440 34373 583445
rect 34058 583436 34368 583440
rect 34058 580760 34368 580764
rect 18911 580440 18920 580760
rect 19240 580755 34373 580760
rect 19240 580445 34058 580755
rect 34368 580445 34373 580755
rect 19240 580440 34373 580445
rect 34058 580436 34368 580440
rect 34058 577760 34368 577764
rect 18911 577440 18920 577760
rect 19240 577755 34373 577760
rect 19240 577445 34058 577755
rect 34368 577445 34373 577755
rect 19240 577440 34373 577445
rect 34058 577436 34368 577440
rect 34058 574760 34368 574764
rect 18911 574440 18920 574760
rect 19240 574755 34373 574760
rect 19240 574445 34058 574755
rect 34368 574445 34373 574755
rect 19240 574440 34373 574445
rect 34058 574436 34368 574440
rect 34058 571760 34368 571764
rect 18911 571440 18920 571760
rect 19240 571755 34373 571760
rect 19240 571445 34058 571755
rect 34368 571445 34373 571755
rect 19240 571440 34373 571445
rect 34058 571436 34368 571440
rect 34058 568760 34368 568764
rect 18911 568440 18920 568760
rect 19240 568755 34373 568760
rect 19240 568445 34058 568755
rect 34368 568445 34373 568755
rect 19240 568440 34373 568445
rect 34058 568436 34368 568440
rect 428434 566278 430884 566282
rect 34058 565760 34368 565764
rect 18911 565440 18920 565760
rect 19240 565755 34373 565760
rect 19240 565445 34058 565755
rect 34368 565445 34373 565755
rect 19240 565440 34373 565445
rect 34058 565436 34368 565440
rect 404344 563818 404353 566278
rect 406813 566273 430889 566278
rect 406813 563823 428434 566273
rect 430884 563823 430889 566273
rect 406813 563818 430889 563823
rect 428434 563814 430884 563818
rect 34058 562760 34368 562764
rect 18911 562440 18920 562760
rect 19240 562755 34373 562760
rect 19240 562445 34058 562755
rect 34368 562445 34373 562755
rect 19240 562440 34373 562445
rect 34058 562436 34368 562440
rect 34058 559760 34368 559764
rect 18911 559440 18920 559760
rect 19240 559755 34373 559760
rect 19240 559445 34058 559755
rect 34368 559445 34373 559755
rect 19240 559440 34373 559445
rect 34058 559436 34368 559440
rect 34058 556760 34368 556764
rect 18911 556440 18920 556760
rect 19240 556755 34373 556760
rect 19240 556445 34058 556755
rect 34368 556445 34373 556755
rect 19240 556440 34373 556445
rect 34058 556436 34368 556440
rect 34058 553760 34368 553764
rect 18911 553440 18920 553760
rect 19240 553755 34373 553760
rect 19240 553445 34058 553755
rect 34368 553445 34373 553755
rect 19240 553440 34373 553445
rect 34058 553436 34368 553440
rect 428434 552465 430884 552469
rect 34058 550760 34368 550764
rect 18911 550440 18920 550760
rect 19240 550755 34373 550760
rect 19240 550445 34058 550755
rect 34368 550445 34373 550755
rect 19240 550440 34373 550445
rect 34058 550436 34368 550440
rect 404418 550005 404427 552465
rect 406887 552460 430889 552465
rect 406887 550010 428434 552460
rect 430884 550010 430889 552460
rect 406887 550005 430889 550010
rect 428434 550001 430884 550005
rect 34058 547760 34368 547764
rect 18911 547440 18920 547760
rect 19240 547755 34373 547760
rect 19240 547445 34058 547755
rect 34368 547445 34373 547755
rect 19240 547440 34373 547445
rect 34058 547436 34368 547440
rect 34058 544760 34368 544764
rect 18911 544440 18920 544760
rect 19240 544755 34373 544760
rect 19240 544445 34058 544755
rect 34368 544445 34373 544755
rect 19240 544440 34373 544445
rect 34058 544436 34368 544440
rect 428434 542841 430884 542845
rect 34058 541760 34368 541764
rect 18911 541440 18920 541760
rect 19240 541755 34373 541760
rect 19240 541445 34058 541755
rect 34368 541445 34373 541755
rect 19240 541440 34373 541445
rect 34058 541436 34368 541440
rect 404124 540381 404133 542841
rect 406593 542836 430889 542841
rect 406593 540386 428434 542836
rect 430884 540386 430889 542836
rect 406593 540381 430889 540386
rect 428434 540377 430884 540381
rect 34058 538760 34368 538764
rect 18911 538440 18920 538760
rect 19240 538755 34373 538760
rect 19240 538445 34058 538755
rect 34368 538445 34373 538755
rect 19240 538440 34373 538445
rect 34058 538436 34368 538440
rect 34058 535760 34368 535764
rect 18911 535440 18920 535760
rect 19240 535755 34373 535760
rect 19240 535445 34058 535755
rect 34368 535445 34373 535755
rect 19240 535440 34373 535445
rect 34058 535436 34368 535440
rect 34058 532760 34368 532764
rect 18911 532440 18920 532760
rect 19240 532755 34373 532760
rect 19240 532445 34058 532755
rect 34368 532445 34373 532755
rect 19240 532440 34373 532445
rect 34058 532436 34368 532440
rect 428434 531893 430884 531897
rect 34058 529760 34368 529764
rect 18911 529440 18920 529760
rect 19240 529755 34373 529760
rect 19240 529445 34058 529755
rect 34368 529445 34373 529755
rect 19240 529440 34373 529445
rect 34058 529436 34368 529440
rect 404124 529433 404133 531893
rect 406593 531888 430889 531893
rect 406593 529438 428434 531888
rect 430884 529438 430889 531888
rect 406593 529433 430889 529438
rect 428434 529429 430884 529433
rect 34058 526760 34368 526764
rect 18911 526440 18920 526760
rect 19240 526755 34373 526760
rect 19240 526445 34058 526755
rect 34368 526445 34373 526755
rect 19240 526440 34373 526445
rect 34058 526436 34368 526440
rect 34058 523760 34368 523764
rect 18911 523440 18920 523760
rect 19240 523755 34373 523760
rect 19240 523445 34058 523755
rect 34368 523445 34373 523755
rect 19240 523440 34373 523445
rect 34058 523436 34368 523440
rect 34058 520760 34368 520764
rect 18911 520440 18920 520760
rect 19240 520755 34373 520760
rect 19240 520445 34058 520755
rect 34368 520445 34373 520755
rect 19240 520440 34373 520445
rect 34058 520436 34368 520440
rect 34058 517760 34368 517764
rect 18911 517440 18920 517760
rect 19240 517755 34373 517760
rect 19240 517445 34058 517755
rect 34368 517445 34373 517755
rect 19240 517440 34373 517445
rect 34058 517436 34368 517440
rect 428434 512943 430884 512947
rect 34058 511760 34368 511764
rect 18911 511440 18920 511760
rect 19240 511755 34373 511760
rect 19240 511445 34058 511755
rect 34368 511445 34373 511755
rect 19240 511440 34373 511445
rect 34058 511436 34368 511440
rect 404170 510483 404179 512943
rect 406639 512938 430889 512943
rect 406639 510488 428434 512938
rect 430884 510488 430889 512938
rect 406639 510483 430889 510488
rect 428434 510479 430884 510483
rect 34058 508760 34368 508764
rect 18911 508440 18920 508760
rect 19240 508755 34373 508760
rect 19240 508445 34058 508755
rect 34368 508445 34373 508755
rect 19240 508440 34373 508445
rect 34058 508436 34368 508440
rect 34058 505760 34368 505764
rect 18911 505440 18920 505760
rect 19240 505755 34373 505760
rect 19240 505445 34058 505755
rect 34368 505445 34373 505755
rect 19240 505440 34373 505445
rect 34058 505436 34368 505440
rect 34058 502760 34368 502764
rect 18911 502440 18920 502760
rect 19240 502755 34373 502760
rect 19240 502445 34058 502755
rect 34368 502445 34373 502755
rect 19240 502440 34373 502445
rect 34058 502436 34368 502440
rect 34058 499760 34368 499764
rect 18911 499440 18920 499760
rect 19240 499755 34373 499760
rect 19240 499445 34058 499755
rect 34368 499445 34373 499755
rect 19240 499440 34373 499445
rect 34058 499436 34368 499440
rect 34058 496760 34368 496764
rect 18911 496440 18920 496760
rect 19240 496755 34373 496760
rect 19240 496445 34058 496755
rect 34368 496445 34373 496755
rect 19240 496440 34373 496445
rect 34058 496436 34368 496440
rect 34058 493760 34368 493764
rect 18911 493440 18920 493760
rect 19240 493755 34373 493760
rect 19240 493445 34058 493755
rect 34368 493445 34373 493755
rect 19240 493440 34373 493445
rect 34058 493436 34368 493440
rect 34058 490760 34368 490764
rect 18911 490440 18920 490760
rect 19240 490755 34373 490760
rect 19240 490445 34058 490755
rect 34368 490445 34373 490755
rect 19240 490440 34373 490445
rect 34058 490436 34368 490440
rect 34058 487760 34368 487764
rect 18911 487440 18920 487760
rect 19240 487755 34373 487760
rect 19240 487445 34058 487755
rect 34368 487445 34373 487755
rect 19240 487440 34373 487445
rect 34058 487436 34368 487440
rect 428434 486407 430884 486411
rect 34058 484760 34368 484764
rect 18911 484440 18920 484760
rect 19240 484755 34373 484760
rect 19240 484445 34058 484755
rect 34368 484445 34373 484755
rect 19240 484440 34373 484445
rect 34058 484436 34368 484440
rect 404451 483947 404460 486407
rect 406920 486402 430889 486407
rect 406920 483952 428434 486402
rect 430884 483952 430889 486402
rect 406920 483947 430889 483952
rect 428434 483943 430884 483947
rect 34058 481760 34368 481764
rect 18911 481440 18920 481760
rect 19240 481755 34373 481760
rect 19240 481445 34058 481755
rect 34368 481445 34373 481755
rect 19240 481440 34373 481445
rect 34058 481436 34368 481440
rect 34058 478760 34368 478764
rect 18911 478440 18920 478760
rect 19240 478755 34373 478760
rect 19240 478445 34058 478755
rect 34368 478445 34373 478755
rect 19240 478440 34373 478445
rect 34058 478436 34368 478440
rect 34058 475760 34368 475764
rect 18911 475440 18920 475760
rect 19240 475755 34373 475760
rect 19240 475445 34058 475755
rect 34368 475445 34373 475755
rect 19240 475440 34373 475445
rect 34058 475436 34368 475440
rect 34058 472760 34368 472764
rect 18911 472440 18920 472760
rect 19240 472755 34373 472760
rect 19240 472445 34058 472755
rect 34368 472445 34373 472755
rect 19240 472440 34373 472445
rect 34058 472436 34368 472440
rect 34058 469760 34368 469764
rect 18911 469440 18920 469760
rect 19240 469755 34373 469760
rect 19240 469445 34058 469755
rect 34368 469445 34373 469755
rect 19240 469440 34373 469445
rect 34058 469436 34368 469440
rect 34058 466760 34368 466764
rect 18911 466440 18920 466760
rect 19240 466755 34373 466760
rect 19240 466445 34058 466755
rect 34368 466445 34373 466755
rect 19240 466440 34373 466445
rect 34058 466436 34368 466440
rect 34058 463760 34368 463764
rect 18911 463440 18920 463760
rect 19240 463755 34373 463760
rect 19240 463445 34058 463755
rect 34368 463445 34373 463755
rect 19240 463440 34373 463445
rect 34058 463436 34368 463440
rect 34058 460760 34368 460764
rect 18911 460440 18920 460760
rect 19240 460755 34373 460760
rect 19240 460445 34058 460755
rect 34368 460445 34373 460755
rect 19240 460440 34373 460445
rect 34058 460436 34368 460440
rect 34058 457760 34368 457764
rect 18911 457440 18920 457760
rect 19240 457755 34373 457760
rect 19240 457445 34058 457755
rect 34368 457445 34373 457755
rect 19240 457440 34373 457445
rect 34058 457436 34368 457440
rect 34058 454760 34368 454764
rect 18911 454440 18920 454760
rect 19240 454755 34373 454760
rect 19240 454445 34058 454755
rect 34368 454445 34373 454755
rect 19240 454440 34373 454445
rect 34058 454436 34368 454440
rect 34058 451760 34368 451764
rect 18911 451440 18920 451760
rect 19240 451755 34373 451760
rect 19240 451445 34058 451755
rect 34368 451445 34373 451755
rect 19240 451440 34373 451445
rect 34058 451436 34368 451440
rect 428434 449962 430884 449966
rect 34058 448760 34368 448764
rect 18911 448440 18920 448760
rect 19240 448755 34373 448760
rect 19240 448445 34058 448755
rect 34368 448445 34373 448755
rect 19240 448440 34373 448445
rect 34058 448436 34368 448440
rect 404472 447502 404481 449962
rect 406941 449957 430889 449962
rect 406941 447507 428434 449957
rect 430884 447507 430889 449957
rect 406941 447502 430889 447507
rect 428434 447498 430884 447502
rect 34058 445760 34368 445764
rect 18911 445440 18920 445760
rect 19240 445755 34373 445760
rect 19240 445445 34058 445755
rect 34368 445445 34373 445755
rect 19240 445440 34373 445445
rect 34058 445436 34368 445440
rect 34058 442760 34368 442764
rect 18911 442440 18920 442760
rect 19240 442755 34373 442760
rect 19240 442445 34058 442755
rect 34368 442445 34373 442755
rect 19240 442440 34373 442445
rect 34058 442436 34368 442440
rect 34058 439760 34368 439764
rect 18911 439440 18920 439760
rect 19240 439755 34373 439760
rect 19240 439445 34058 439755
rect 34368 439445 34373 439755
rect 19240 439440 34373 439445
rect 34058 439436 34368 439440
rect 34058 436760 34368 436764
rect 18911 436440 18920 436760
rect 19240 436755 34373 436760
rect 19240 436445 34058 436755
rect 34368 436445 34373 436755
rect 19240 436440 34373 436445
rect 34058 436436 34368 436440
rect 34058 433760 34368 433764
rect 18911 433440 18920 433760
rect 19240 433755 34373 433760
rect 19240 433445 34058 433755
rect 34368 433445 34373 433755
rect 19240 433440 34373 433445
rect 34058 433436 34368 433440
rect 34058 430760 34368 430764
rect 18911 430440 18920 430760
rect 19240 430755 34373 430760
rect 19240 430445 34058 430755
rect 34368 430445 34373 430755
rect 19240 430440 34373 430445
rect 34058 430436 34368 430440
rect 34058 427760 34368 427764
rect 18911 427440 18920 427760
rect 19240 427755 34373 427760
rect 19240 427445 34058 427755
rect 34368 427445 34373 427755
rect 19240 427440 34373 427445
rect 34058 427436 34368 427440
rect 34058 424760 34368 424764
rect 18911 424440 18920 424760
rect 19240 424755 34373 424760
rect 19240 424445 34058 424755
rect 34368 424445 34373 424755
rect 19240 424440 34373 424445
rect 34058 424436 34368 424440
rect 1553 420470 1655 420474
rect 14170 420470 14290 423400
rect 34058 421760 34368 421764
rect 18911 421440 18920 421760
rect 19240 421755 34373 421760
rect 19240 421445 34058 421755
rect 34368 421445 34373 421755
rect 428434 421579 430884 421583
rect 19240 421440 34373 421445
rect 34058 421436 34368 421440
rect 1548 420465 14806 420470
rect 1548 420363 1553 420465
rect 1655 420363 14806 420465
rect 1548 420358 14806 420363
rect 1553 420354 1655 420358
rect 4929 377248 5031 377252
rect 13084 377248 13196 377476
rect 4924 377243 13406 377248
rect 4924 377141 4929 377243
rect 5031 377141 13406 377243
rect 4924 377136 13406 377141
rect 4929 377132 5031 377136
rect 13084 358966 13196 377136
rect 14170 359517 14290 420358
rect 404804 419119 404813 421579
rect 407273 421574 430889 421579
rect 407273 419124 428434 421574
rect 430884 419124 430889 421574
rect 407273 419119 430889 419124
rect 428434 419115 430884 419119
rect 34058 418760 34368 418764
rect 18911 418440 18920 418760
rect 19240 418755 34373 418760
rect 19240 418445 34058 418755
rect 34368 418445 34373 418755
rect 19240 418440 34373 418445
rect 34058 418436 34368 418440
rect 34058 415760 34368 415764
rect 18911 415440 18920 415760
rect 19240 415755 34373 415760
rect 19240 415445 34058 415755
rect 34368 415445 34373 415755
rect 19240 415440 34373 415445
rect 34058 415436 34368 415440
rect 34058 412760 34368 412764
rect 18911 412440 18920 412760
rect 19240 412755 34373 412760
rect 19240 412445 34058 412755
rect 34368 412445 34373 412755
rect 19240 412440 34373 412445
rect 34058 412436 34368 412440
rect 34058 409760 34368 409764
rect 18911 409440 18920 409760
rect 19240 409755 34373 409760
rect 19240 409445 34058 409755
rect 34368 409445 34373 409755
rect 428434 409691 430884 409695
rect 19240 409440 34373 409445
rect 34058 409436 34368 409440
rect 404570 407231 404579 409691
rect 407039 409686 430889 409691
rect 407039 407236 428434 409686
rect 430884 407236 430889 409686
rect 407039 407231 430889 407236
rect 428434 407227 430884 407231
rect 34058 406760 34368 406764
rect 18911 406440 18920 406760
rect 19240 406755 34373 406760
rect 19240 406445 34058 406755
rect 34368 406445 34373 406755
rect 19240 406440 34373 406445
rect 34058 406436 34368 406440
rect 34058 403760 34368 403764
rect 18911 403440 18920 403760
rect 19240 403755 34373 403760
rect 19240 403445 34058 403755
rect 34368 403445 34373 403755
rect 19240 403440 34373 403445
rect 34058 403436 34368 403440
rect 34058 397760 34368 397764
rect 18911 397440 18920 397760
rect 19240 397755 34373 397760
rect 19240 397445 34058 397755
rect 34368 397445 34373 397755
rect 19240 397440 34373 397445
rect 34058 397436 34368 397440
rect 34058 394760 34368 394764
rect 18911 394440 18920 394760
rect 19240 394755 34373 394760
rect 19240 394445 34058 394755
rect 34368 394445 34373 394755
rect 19240 394440 34373 394445
rect 34058 394436 34368 394440
rect 34058 391760 34368 391764
rect 18911 391440 18920 391760
rect 19240 391755 34373 391760
rect 19240 391445 34058 391755
rect 34368 391445 34373 391755
rect 19240 391440 34373 391445
rect 34058 391436 34368 391440
rect 34058 388760 34368 388764
rect 18911 388440 18920 388760
rect 19240 388755 34373 388760
rect 19240 388445 34058 388755
rect 34368 388445 34373 388755
rect 19240 388440 34373 388445
rect 34058 388436 34368 388440
rect 34058 385760 34368 385764
rect 18911 385440 18920 385760
rect 19240 385755 34373 385760
rect 19240 385445 34058 385755
rect 34368 385445 34373 385755
rect 19240 385440 34373 385445
rect 34058 385436 34368 385440
rect 34058 382760 34368 382764
rect 18911 382440 18920 382760
rect 19240 382755 34373 382760
rect 19240 382445 34058 382755
rect 34368 382445 34373 382755
rect 19240 382440 34373 382445
rect 34058 382436 34368 382440
rect 34058 379760 34368 379764
rect 18911 379440 18920 379760
rect 19240 379755 34373 379760
rect 19240 379445 34058 379755
rect 34368 379445 34373 379755
rect 19240 379440 34373 379445
rect 34058 379436 34368 379440
rect 414098 377762 414388 377768
rect 414089 377472 414098 377762
rect 414388 377472 414397 377762
rect 414098 377466 414388 377472
rect 413990 377075 414280 377081
rect 413981 376785 413990 377075
rect 414280 376785 414289 377075
rect 413990 376779 414280 376785
rect 34058 376760 34368 376764
rect 18911 376440 18920 376760
rect 19240 376755 34373 376760
rect 19240 376445 34058 376755
rect 34368 376445 34373 376755
rect 19240 376440 34373 376445
rect 34058 376436 34368 376440
rect 414243 376208 414533 376214
rect 414234 375918 414243 376208
rect 414533 375918 414542 376208
rect 414243 375912 414533 375918
rect 414026 374653 414316 374659
rect 414017 374363 414026 374653
rect 414316 374363 414325 374653
rect 414026 374357 414316 374363
rect 413994 374054 414284 374060
rect 413985 373764 413994 374054
rect 414284 373764 414293 374054
rect 34058 373760 34368 373764
rect 18911 373440 18920 373760
rect 19240 373755 34373 373760
rect 413994 373758 414284 373764
rect 19240 373445 34058 373755
rect 34368 373445 34373 373755
rect 19240 373440 34373 373445
rect 34058 373436 34368 373440
rect 414352 373194 414642 373200
rect 414343 372904 414352 373194
rect 414642 372904 414651 373194
rect 414352 372898 414642 372904
rect 414245 372477 414535 372483
rect 414236 372187 414245 372477
rect 414535 372187 414544 372477
rect 414245 372181 414535 372187
rect 414352 371832 414642 371838
rect 414343 371542 414352 371832
rect 414642 371542 414651 371832
rect 414352 371536 414642 371542
rect 414776 371295 415066 371301
rect 414767 371005 414776 371295
rect 415066 371005 415075 371295
rect 414776 370999 415066 371005
rect 34058 370760 34368 370764
rect 18911 370440 18920 370760
rect 19240 370755 34373 370760
rect 19240 370445 34058 370755
rect 34368 370445 34373 370755
rect 413772 370704 414062 370710
rect 19240 370440 34373 370445
rect 34058 370436 34368 370440
rect 413763 370414 413772 370704
rect 414062 370414 414071 370704
rect 413772 370408 414062 370414
rect 34058 367760 34368 367764
rect 18911 367440 18920 367760
rect 19240 367755 34373 367760
rect 19240 367445 34058 367755
rect 34368 367445 34373 367755
rect 19240 367440 34373 367445
rect 34058 367436 34368 367440
rect 34058 364760 34368 364764
rect 18911 364440 18920 364760
rect 19240 364755 34373 364760
rect 19240 364445 34058 364755
rect 34368 364445 34373 364755
rect 19240 364440 34373 364445
rect 34058 364436 34368 364440
rect 55827 363630 55937 365011
rect 52296 363520 55937 363630
rect 21725 359517 21835 359521
rect 14170 359512 21840 359517
rect 14170 359402 21725 359512
rect 21835 359402 21840 359512
rect 14170 359397 21840 359402
rect 21725 359393 21835 359397
rect 22916 358966 23018 358970
rect 13084 358961 23023 358966
rect 13084 358859 22916 358961
rect 23018 358859 23023 358961
rect 13084 358854 23023 358859
rect 22916 358850 23018 358854
rect 1924 353279 4374 353283
rect 26650 353279 29110 353285
rect 1913 350819 1919 353279
rect 4379 350819 4385 353279
rect 26641 350819 26650 353279
rect 29110 350819 29119 353279
rect 1924 350815 4374 350819
rect 26650 350813 29110 350819
rect 1924 348750 4374 348754
rect 26576 348750 29036 348756
rect 1913 346290 1919 348750
rect 4379 346290 4385 348750
rect 26567 346290 26576 348750
rect 29036 346290 29045 348750
rect 1924 346286 4374 346290
rect 26576 346284 29036 346290
rect 1924 344240 4374 344244
rect 26576 344240 29036 344246
rect 1913 341780 1919 344240
rect 4379 341780 4385 344240
rect 26567 341780 26576 344240
rect 29036 341780 29045 344240
rect 1924 341776 4374 341780
rect 26576 341774 29036 341780
rect 5660 336789 5772 336794
rect 5656 336687 5665 336789
rect 5767 336687 5776 336789
rect 5660 327595 5772 336687
rect 5660 327474 5772 327483
rect 1924 315915 4374 315919
rect 1919 315910 39936 315915
rect 1919 313460 1924 315910
rect 4374 313460 39936 315910
rect 1919 313455 39936 313460
rect 42396 313455 42405 315915
rect 1924 313451 4374 313455
rect 8362 261315 8493 261350
rect 8362 261245 8387 261315
rect 8457 261245 8493 261315
rect 8362 261225 8493 261245
rect 52296 257496 52406 363520
rect 361653 363482 362756 363662
rect 362576 362993 362756 363482
rect 362389 362745 368047 362993
rect 428434 362175 430884 362179
rect 404516 359715 404525 362175
rect 406985 362170 430889 362175
rect 406985 359720 428434 362170
rect 430884 359720 430889 362170
rect 406985 359715 430889 359720
rect 428434 359711 430884 359715
rect 365000 358894 365170 358903
rect 365170 358724 368461 358894
rect 365000 358715 365170 358724
rect 55307 345756 55627 345762
rect 58307 345756 58627 345762
rect 61307 345756 61627 345762
rect 64307 345756 64627 345762
rect 67307 345756 67627 345762
rect 70307 345756 70627 345762
rect 73307 345756 73627 345762
rect 76307 345756 76627 345762
rect 79307 345756 79627 345762
rect 82307 345756 82627 345762
rect 85307 345756 85627 345762
rect 88307 345756 88627 345762
rect 91307 345756 91627 345762
rect 94307 345756 94627 345762
rect 97307 345756 97627 345762
rect 100307 345756 100627 345762
rect 103307 345756 103627 345762
rect 106307 345756 106627 345762
rect 109307 345756 109627 345762
rect 112307 345756 112627 345762
rect 115307 345756 115627 345762
rect 118307 345756 118627 345762
rect 121307 345756 121627 345762
rect 124307 345756 124627 345762
rect 127307 345756 127627 345762
rect 130307 345756 130627 345762
rect 133307 345756 133627 345762
rect 136307 345756 136627 345762
rect 139307 345756 139627 345762
rect 142307 345756 142627 345762
rect 145307 345756 145627 345762
rect 148307 345756 148627 345762
rect 151307 345756 151627 345762
rect 154307 345756 154627 345762
rect 157307 345756 157627 345762
rect 160307 345756 160627 345762
rect 163307 345756 163627 345762
rect 166307 345756 166627 345762
rect 169307 345756 169627 345762
rect 172307 345756 172627 345762
rect 175307 345756 175627 345762
rect 178307 345756 178627 345762
rect 181307 345756 181627 345762
rect 184307 345756 184627 345762
rect 187307 345756 187627 345762
rect 190307 345756 190627 345762
rect 193307 345756 193627 345762
rect 196307 345756 196627 345762
rect 199307 345756 199627 345762
rect 202307 345756 202627 345762
rect 205307 345756 205627 345762
rect 208307 345756 208627 345762
rect 211307 345756 211627 345762
rect 214307 345756 214627 345762
rect 217307 345756 217627 345762
rect 220307 345756 220627 345762
rect 223307 345756 223627 345762
rect 226307 345756 226627 345762
rect 229307 345756 229627 345762
rect 232307 345756 232627 345762
rect 235307 345756 235627 345762
rect 238307 345756 238627 345762
rect 241307 345756 241627 345762
rect 244307 345756 244627 345762
rect 247307 345756 247627 345762
rect 250307 345756 250627 345762
rect 253307 345756 253627 345762
rect 256307 345756 256627 345762
rect 259307 345756 259627 345762
rect 262307 345756 262627 345762
rect 265307 345756 265627 345762
rect 268307 345756 268627 345762
rect 271307 345756 271627 345762
rect 274307 345756 274627 345762
rect 277307 345756 277627 345762
rect 280307 345756 280627 345762
rect 283307 345756 283627 345762
rect 286307 345756 286627 345762
rect 289307 345756 289627 345762
rect 292307 345756 292627 345762
rect 295307 345756 295627 345762
rect 298307 345756 298627 345762
rect 301307 345756 301627 345762
rect 304307 345756 304627 345762
rect 307307 345756 307627 345762
rect 310307 345756 310627 345762
rect 313307 345756 313627 345762
rect 316307 345756 316627 345762
rect 319307 345756 319627 345762
rect 325307 345756 325627 345762
rect 328307 345756 328627 345762
rect 331307 345756 331627 345762
rect 334307 345756 334627 345762
rect 337307 345756 337627 345762
rect 340307 345756 340627 345762
rect 343307 345756 343627 345762
rect 346307 345756 346627 345762
rect 349307 345756 349627 345762
rect 352307 345756 352627 345762
rect 355307 345756 355627 345762
rect 358307 345756 358627 345762
rect 55301 345436 55307 345756
rect 55627 345436 55633 345756
rect 58301 345436 58307 345756
rect 58627 345436 58633 345756
rect 61301 345436 61307 345756
rect 61627 345436 61633 345756
rect 64301 345436 64307 345756
rect 64627 345436 64633 345756
rect 67301 345436 67307 345756
rect 67627 345436 67633 345756
rect 70301 345436 70307 345756
rect 70627 345436 70633 345756
rect 73301 345436 73307 345756
rect 73627 345436 73633 345756
rect 76301 345436 76307 345756
rect 76627 345436 76633 345756
rect 79301 345436 79307 345756
rect 79627 345436 79633 345756
rect 82301 345436 82307 345756
rect 82627 345436 82633 345756
rect 85301 345436 85307 345756
rect 85627 345436 85633 345756
rect 88301 345436 88307 345756
rect 88627 345436 88633 345756
rect 91301 345436 91307 345756
rect 91627 345436 91633 345756
rect 94301 345436 94307 345756
rect 94627 345436 94633 345756
rect 97301 345436 97307 345756
rect 97627 345436 97633 345756
rect 100301 345436 100307 345756
rect 100627 345436 100633 345756
rect 103301 345436 103307 345756
rect 103627 345436 103633 345756
rect 106301 345436 106307 345756
rect 106627 345436 106633 345756
rect 109301 345436 109307 345756
rect 109627 345436 109633 345756
rect 112301 345436 112307 345756
rect 112627 345436 112633 345756
rect 115301 345436 115307 345756
rect 115627 345436 115633 345756
rect 118301 345436 118307 345756
rect 118627 345436 118633 345756
rect 121301 345436 121307 345756
rect 121627 345436 121633 345756
rect 124301 345436 124307 345756
rect 124627 345436 124633 345756
rect 127301 345436 127307 345756
rect 127627 345436 127633 345756
rect 130301 345436 130307 345756
rect 130627 345436 130633 345756
rect 133301 345436 133307 345756
rect 133627 345436 133633 345756
rect 136301 345436 136307 345756
rect 136627 345436 136633 345756
rect 139301 345436 139307 345756
rect 139627 345436 139633 345756
rect 142301 345436 142307 345756
rect 142627 345436 142633 345756
rect 145301 345436 145307 345756
rect 145627 345436 145633 345756
rect 148301 345436 148307 345756
rect 148627 345436 148633 345756
rect 151301 345436 151307 345756
rect 151627 345436 151633 345756
rect 154301 345436 154307 345756
rect 154627 345436 154633 345756
rect 157301 345436 157307 345756
rect 157627 345436 157633 345756
rect 160301 345436 160307 345756
rect 160627 345436 160633 345756
rect 163301 345436 163307 345756
rect 163627 345436 163633 345756
rect 166301 345436 166307 345756
rect 166627 345436 166633 345756
rect 169301 345436 169307 345756
rect 169627 345436 169633 345756
rect 172301 345436 172307 345756
rect 172627 345436 172633 345756
rect 175301 345436 175307 345756
rect 175627 345436 175633 345756
rect 178301 345436 178307 345756
rect 178627 345436 178633 345756
rect 181301 345436 181307 345756
rect 181627 345436 181633 345756
rect 184301 345436 184307 345756
rect 184627 345436 184633 345756
rect 187301 345436 187307 345756
rect 187627 345436 187633 345756
rect 190301 345436 190307 345756
rect 190627 345436 190633 345756
rect 193301 345436 193307 345756
rect 193627 345436 193633 345756
rect 196301 345436 196307 345756
rect 196627 345436 196633 345756
rect 199301 345436 199307 345756
rect 199627 345436 199633 345756
rect 202301 345436 202307 345756
rect 202627 345436 202633 345756
rect 205301 345436 205307 345756
rect 205627 345436 205633 345756
rect 208301 345436 208307 345756
rect 208627 345436 208633 345756
rect 211301 345436 211307 345756
rect 211627 345436 211633 345756
rect 214301 345436 214307 345756
rect 214627 345436 214633 345756
rect 217301 345436 217307 345756
rect 217627 345436 217633 345756
rect 220301 345436 220307 345756
rect 220627 345436 220633 345756
rect 223301 345436 223307 345756
rect 223627 345436 223633 345756
rect 226301 345436 226307 345756
rect 226627 345436 226633 345756
rect 229301 345436 229307 345756
rect 229627 345436 229633 345756
rect 232301 345436 232307 345756
rect 232627 345436 232633 345756
rect 235301 345436 235307 345756
rect 235627 345436 235633 345756
rect 238301 345436 238307 345756
rect 238627 345436 238633 345756
rect 241301 345436 241307 345756
rect 241627 345436 241633 345756
rect 244301 345436 244307 345756
rect 244627 345436 244633 345756
rect 247301 345436 247307 345756
rect 247627 345436 247633 345756
rect 250301 345436 250307 345756
rect 250627 345436 250633 345756
rect 253301 345436 253307 345756
rect 253627 345436 253633 345756
rect 256301 345436 256307 345756
rect 256627 345436 256633 345756
rect 259301 345436 259307 345756
rect 259627 345436 259633 345756
rect 262301 345436 262307 345756
rect 262627 345436 262633 345756
rect 265301 345436 265307 345756
rect 265627 345436 265633 345756
rect 268301 345436 268307 345756
rect 268627 345436 268633 345756
rect 271301 345436 271307 345756
rect 271627 345436 271633 345756
rect 274301 345436 274307 345756
rect 274627 345436 274633 345756
rect 277301 345436 277307 345756
rect 277627 345436 277633 345756
rect 280301 345436 280307 345756
rect 280627 345436 280633 345756
rect 283301 345436 283307 345756
rect 283627 345436 283633 345756
rect 286301 345436 286307 345756
rect 286627 345436 286633 345756
rect 289301 345436 289307 345756
rect 289627 345436 289633 345756
rect 292301 345436 292307 345756
rect 292627 345436 292633 345756
rect 295301 345436 295307 345756
rect 295627 345436 295633 345756
rect 298301 345436 298307 345756
rect 298627 345436 298633 345756
rect 301301 345436 301307 345756
rect 301627 345436 301633 345756
rect 304301 345436 304307 345756
rect 304627 345436 304633 345756
rect 307301 345436 307307 345756
rect 307627 345436 307633 345756
rect 310301 345436 310307 345756
rect 310627 345436 310633 345756
rect 313301 345436 313307 345756
rect 313627 345436 313633 345756
rect 316301 345436 316307 345756
rect 316627 345436 316633 345756
rect 319301 345436 319307 345756
rect 319627 345436 319633 345756
rect 325301 345436 325307 345756
rect 325627 345436 325633 345756
rect 328301 345436 328307 345756
rect 328627 345436 328633 345756
rect 331301 345436 331307 345756
rect 331627 345436 331633 345756
rect 334301 345436 334307 345756
rect 334627 345436 334633 345756
rect 337301 345436 337307 345756
rect 337627 345436 337633 345756
rect 340301 345436 340307 345756
rect 340627 345436 340633 345756
rect 343301 345436 343307 345756
rect 343627 345436 343633 345756
rect 346301 345436 346307 345756
rect 346627 345436 346633 345756
rect 349301 345436 349307 345756
rect 349627 345436 349633 345756
rect 352301 345436 352307 345756
rect 352627 345436 352633 345756
rect 355301 345436 355307 345756
rect 355627 345436 355633 345756
rect 358301 345436 358307 345756
rect 358627 345436 358633 345756
rect 55307 323427 55627 345436
rect 55307 323098 55627 323107
rect 58307 323427 58627 345436
rect 58307 323098 58627 323107
rect 61307 323427 61627 345436
rect 61307 323098 61627 323107
rect 64307 323427 64627 345436
rect 64307 323098 64627 323107
rect 67307 323427 67627 345436
rect 67307 323098 67627 323107
rect 70307 323427 70627 345436
rect 70307 323098 70627 323107
rect 73307 323427 73627 345436
rect 73307 323098 73627 323107
rect 76307 323427 76627 345436
rect 76307 323098 76627 323107
rect 79307 323427 79627 345436
rect 79307 323098 79627 323107
rect 82307 323427 82627 345436
rect 82307 323098 82627 323107
rect 85307 323427 85627 345436
rect 85307 323098 85627 323107
rect 88307 323427 88627 345436
rect 88307 323098 88627 323107
rect 91307 323427 91627 345436
rect 91307 323098 91627 323107
rect 94307 323427 94627 345436
rect 94307 323098 94627 323107
rect 97307 323427 97627 345436
rect 97307 323098 97627 323107
rect 100307 323427 100627 345436
rect 100307 323098 100627 323107
rect 103307 323427 103627 345436
rect 103307 323098 103627 323107
rect 106307 323427 106627 345436
rect 106307 323098 106627 323107
rect 109307 323427 109627 345436
rect 109307 323098 109627 323107
rect 112307 323427 112627 345436
rect 112307 323098 112627 323107
rect 115307 323427 115627 345436
rect 115307 323098 115627 323107
rect 118307 323427 118627 345436
rect 118307 323098 118627 323107
rect 121307 323427 121627 345436
rect 121307 323098 121627 323107
rect 124307 323427 124627 345436
rect 124307 323098 124627 323107
rect 127307 323427 127627 345436
rect 127307 323098 127627 323107
rect 130307 323427 130627 345436
rect 130307 323098 130627 323107
rect 133307 323427 133627 345436
rect 133307 323098 133627 323107
rect 136307 323427 136627 345436
rect 136307 323098 136627 323107
rect 139307 323427 139627 345436
rect 139307 323098 139627 323107
rect 142307 323427 142627 345436
rect 142307 323098 142627 323107
rect 145307 323427 145627 345436
rect 145307 323098 145627 323107
rect 148307 323427 148627 345436
rect 148307 323098 148627 323107
rect 151307 323427 151627 345436
rect 151307 323098 151627 323107
rect 154307 323427 154627 345436
rect 154307 323098 154627 323107
rect 157307 323427 157627 345436
rect 157307 323098 157627 323107
rect 160307 323427 160627 345436
rect 160307 323098 160627 323107
rect 163307 323427 163627 345436
rect 163307 323098 163627 323107
rect 166307 323427 166627 345436
rect 166307 323098 166627 323107
rect 169307 323427 169627 345436
rect 169307 323098 169627 323107
rect 172307 323427 172627 345436
rect 172307 323098 172627 323107
rect 175307 323427 175627 345436
rect 175307 323098 175627 323107
rect 178307 323427 178627 345436
rect 178307 323098 178627 323107
rect 181307 323427 181627 345436
rect 181307 323098 181627 323107
rect 184307 323427 184627 345436
rect 184307 323098 184627 323107
rect 187307 323427 187627 345436
rect 187307 323098 187627 323107
rect 190307 323427 190627 345436
rect 190307 323098 190627 323107
rect 193307 323427 193627 345436
rect 193307 323098 193627 323107
rect 196307 323427 196627 345436
rect 196307 323098 196627 323107
rect 199307 323427 199627 345436
rect 199307 323098 199627 323107
rect 202307 323427 202627 345436
rect 202307 323098 202627 323107
rect 205307 323427 205627 345436
rect 205307 323098 205627 323107
rect 208307 323427 208627 345436
rect 208307 323098 208627 323107
rect 211307 323427 211627 345436
rect 211307 323098 211627 323107
rect 214307 323427 214627 345436
rect 214307 323098 214627 323107
rect 217307 323427 217627 345436
rect 217307 323098 217627 323107
rect 220307 323427 220627 345436
rect 220307 323098 220627 323107
rect 223307 323427 223627 345436
rect 223307 323098 223627 323107
rect 226307 323427 226627 345436
rect 226307 323098 226627 323107
rect 229307 323427 229627 345436
rect 229307 323098 229627 323107
rect 232307 323427 232627 345436
rect 232307 323098 232627 323107
rect 235307 323427 235627 345436
rect 235307 323098 235627 323107
rect 238307 323427 238627 345436
rect 238307 323098 238627 323107
rect 241307 323427 241627 345436
rect 241307 323098 241627 323107
rect 244307 323427 244627 345436
rect 244307 323098 244627 323107
rect 247307 323427 247627 345436
rect 247307 323098 247627 323107
rect 250307 323427 250627 345436
rect 250307 323098 250627 323107
rect 253307 323427 253627 345436
rect 253307 323098 253627 323107
rect 256307 323427 256627 345436
rect 256307 323098 256627 323107
rect 259307 323427 259627 345436
rect 259307 323098 259627 323107
rect 262307 323427 262627 345436
rect 262307 323098 262627 323107
rect 265307 323427 265627 345436
rect 265307 323098 265627 323107
rect 268307 323427 268627 345436
rect 268307 323098 268627 323107
rect 271307 323427 271627 345436
rect 271307 323098 271627 323107
rect 274307 323427 274627 345436
rect 274307 323098 274627 323107
rect 277307 323427 277627 345436
rect 277307 323098 277627 323107
rect 280307 323427 280627 345436
rect 280307 323098 280627 323107
rect 283307 323427 283627 345436
rect 283307 323098 283627 323107
rect 286307 323427 286627 345436
rect 286307 323098 286627 323107
rect 289307 323427 289627 345436
rect 289307 323098 289627 323107
rect 292307 323427 292627 345436
rect 292307 323098 292627 323107
rect 295307 323427 295627 345436
rect 295307 323098 295627 323107
rect 298307 323427 298627 345436
rect 298307 323098 298627 323107
rect 301307 323427 301627 345436
rect 301307 323098 301627 323107
rect 304307 323427 304627 345436
rect 304307 323098 304627 323107
rect 307307 323427 307627 345436
rect 307307 323098 307627 323107
rect 310307 323427 310627 345436
rect 310307 323098 310627 323107
rect 313307 323427 313627 345436
rect 313307 323098 313627 323107
rect 316307 323427 316627 345436
rect 316307 323098 316627 323107
rect 319307 323427 319627 345436
rect 319307 323098 319627 323107
rect 325307 323427 325627 345436
rect 325307 323098 325627 323107
rect 328307 323427 328627 345436
rect 328307 323098 328627 323107
rect 331307 323427 331627 345436
rect 331307 323098 331627 323107
rect 334307 323427 334627 345436
rect 334307 323098 334627 323107
rect 337307 323427 337627 345436
rect 337307 323098 337627 323107
rect 340307 323427 340627 345436
rect 340307 323098 340627 323107
rect 343307 323427 343627 345436
rect 343307 323098 343627 323107
rect 346307 323427 346627 345436
rect 346307 323098 346627 323107
rect 349307 323427 349627 345436
rect 349307 323098 349627 323107
rect 352307 323427 352627 345436
rect 352307 323098 352627 323107
rect 355307 323427 355627 345436
rect 355307 323098 355627 323107
rect 358307 323427 358627 345436
rect 372481 336904 372781 336910
rect 375481 336904 375781 336910
rect 378481 336904 378781 336910
rect 381481 336904 381781 336910
rect 384481 336904 384781 336910
rect 387481 336904 387781 336910
rect 390481 336904 390781 336910
rect 393481 336904 393781 336910
rect 396481 336904 396781 336910
rect 372472 336604 372481 336904
rect 372781 336604 372790 336904
rect 375472 336604 375481 336904
rect 375781 336604 375790 336904
rect 378472 336604 378481 336904
rect 378781 336604 378790 336904
rect 381472 336604 381481 336904
rect 381781 336604 381790 336904
rect 384472 336604 384481 336904
rect 384781 336604 384790 336904
rect 387472 336604 387481 336904
rect 387781 336604 387790 336904
rect 390472 336604 390481 336904
rect 390781 336604 390790 336904
rect 393472 336604 393481 336904
rect 393781 336604 393790 336904
rect 396472 336604 396481 336904
rect 396781 336604 396790 336904
rect 372481 336598 372781 336604
rect 375481 336598 375781 336604
rect 378481 336598 378781 336604
rect 381481 336598 381781 336604
rect 384481 336598 384781 336604
rect 387481 336598 387781 336604
rect 390481 336598 390781 336604
rect 393481 336598 393781 336604
rect 396481 336598 396781 336604
rect 358307 323098 358627 323107
rect 436515 308724 436685 680010
rect 176363 308554 436685 308724
rect 64633 261245 64639 261315
rect 64709 261245 86272 261315
rect 52296 257386 77307 257496
rect 55936 248968 56026 249069
rect 55921 248959 56026 248968
rect 56023 248857 56026 248959
rect 55921 248848 56026 248857
rect 55936 193314 56026 248848
rect 77197 201383 77307 257386
rect 86202 203651 86272 261245
rect 86202 203581 166751 203651
rect 164911 201383 165021 201410
rect 77197 201273 165276 201383
rect 55936 192961 56026 193224
rect 164911 191749 165021 201273
rect 166681 191771 166751 203581
rect 176363 196612 176533 308554
rect 287964 230745 290424 230750
rect 287960 228295 287969 230745
rect 290419 228295 290428 230745
rect 180921 207290 181211 207299
rect 183921 207290 184211 207299
rect 186921 207290 187211 207299
rect 189921 207290 190211 207299
rect 192921 207290 193211 207299
rect 195921 207290 196211 207299
rect 198921 207290 199211 207299
rect 201921 207290 202211 207299
rect 204921 207290 205211 207299
rect 180915 207000 180921 207290
rect 181211 207000 181217 207290
rect 183915 207000 183921 207290
rect 184211 207000 184217 207290
rect 186915 207000 186921 207290
rect 187211 207000 187217 207290
rect 189915 207000 189921 207290
rect 190211 207000 190217 207290
rect 192915 207000 192921 207290
rect 193211 207000 193217 207290
rect 195915 207000 195921 207290
rect 196211 207000 196217 207290
rect 198915 207000 198921 207290
rect 199211 207000 199217 207290
rect 201915 207000 201921 207290
rect 202211 207000 202217 207290
rect 204915 207000 204921 207290
rect 205211 207000 205217 207290
rect 180921 206991 181211 207000
rect 183921 206991 184211 207000
rect 186921 206991 187211 207000
rect 189921 206991 190211 207000
rect 192921 206991 193211 207000
rect 195921 206991 196211 207000
rect 198921 206991 199211 207000
rect 201921 206991 202211 207000
rect 204921 206991 205211 207000
rect 176357 196442 176363 196612
rect 176533 196442 176539 196612
rect 9016 191337 9126 191346
rect 9126 191227 162771 191337
rect 9016 191218 9126 191227
rect 55936 189794 56026 190122
rect 55930 189704 55936 189794
rect 56026 189704 56032 189794
rect 55936 189447 56026 189704
rect 55936 189357 162751 189447
rect 175764 188348 175934 188354
rect 175760 188183 175764 188343
rect 175934 188183 175938 188343
rect 175764 188172 175934 188178
rect 175764 186637 175934 186646
rect 175758 186467 175764 186637
rect 175934 186467 175940 186637
rect 175764 186458 175934 186467
rect 21843 186357 163538 186447
rect 21865 121346 21955 186357
rect 176755 184488 177913 184736
rect 21843 121337 21955 121346
rect 21945 121235 21955 121337
rect 21843 121226 21955 121235
rect 21865 121124 21955 121226
rect 33627 183357 163447 183447
rect 33627 78124 33717 183357
rect 176755 180985 177003 184488
rect 175393 180870 177003 180985
rect 175393 180766 176999 180870
rect 177597 180467 177606 180637
rect 177776 180467 178333 180637
rect 180877 172819 181177 172828
rect 183877 172819 184177 172828
rect 186877 172819 187177 172828
rect 189877 172819 190177 172828
rect 192877 172819 193177 172828
rect 195877 172819 196177 172828
rect 198877 172819 199177 172828
rect 201877 172819 202177 172828
rect 204877 172819 205177 172828
rect 180871 172519 180877 172819
rect 181177 172519 181183 172819
rect 183871 172519 183877 172819
rect 184177 172519 184183 172819
rect 186871 172519 186877 172819
rect 187177 172519 187183 172819
rect 189871 172519 189877 172819
rect 190177 172519 190183 172819
rect 192871 172519 192877 172819
rect 193177 172519 193183 172819
rect 195871 172519 195877 172819
rect 196177 172519 196183 172819
rect 198871 172519 198877 172819
rect 199177 172519 199183 172819
rect 201871 172519 201877 172819
rect 202177 172519 202183 172819
rect 204871 172519 204877 172819
rect 205177 172519 205183 172819
rect 180877 172510 181177 172519
rect 183877 172510 184177 172519
rect 186877 172510 187177 172519
rect 189877 172510 190177 172519
rect 192877 172510 193177 172519
rect 195877 172510 196177 172519
rect 198877 172510 199177 172519
rect 201877 172510 202177 172519
rect 204877 172510 205177 172519
rect 287964 118958 290424 228295
rect 287964 116489 290424 116498
rect 33618 78034 33627 78124
rect 33717 78034 33726 78124
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 143673 693995 144063 694385
rect 7017 687779 7327 688089
rect 1924 683555 4374 686005
rect 28686 685488 28746 685548
rect 26802 682004 29262 684464
rect 9021 680757 9121 680857
rect 1924 675660 4374 678110
rect 26510 675655 28970 678115
rect 69665 676260 69775 676370
rect 1924 670438 4374 672888
rect 26343 670433 28803 672893
rect 137061 674932 137381 675252
rect 178455 689056 178515 689116
rect 140632 673664 140702 673734
rect 155835 673733 156205 674103
rect 396236 674665 396396 674825
rect 152421 673475 152531 673585
rect 231038 673374 231348 673684
rect 140637 671070 140697 671130
rect 143673 670346 144063 670736
rect 18920 667440 19240 667760
rect 34058 667445 34368 667755
rect 397829 664827 398129 665127
rect 18920 664440 19240 664760
rect 34058 664445 34368 664755
rect 53668 664413 53978 664723
rect 18920 661440 19240 661760
rect 34058 661445 34368 661755
rect 18920 658440 19240 658760
rect 34058 658445 34368 658755
rect 13647 657006 13967 657326
rect 436515 680010 436685 680180
rect 424849 655864 425009 656024
rect 18920 655440 19240 655760
rect 34058 655445 34368 655755
rect 18920 652440 19240 652760
rect 34058 652445 34368 652755
rect 18920 649440 19240 649760
rect 34058 649445 34368 649755
rect 18920 646440 19240 646760
rect 34058 646445 34368 646755
rect 18920 643440 19240 643760
rect 34058 643445 34368 643755
rect 18920 640440 19240 640760
rect 34058 640445 34368 640755
rect 18920 637440 19240 637760
rect 34058 637445 34368 637755
rect 18920 634440 19240 634760
rect 34058 634445 34368 634755
rect 18920 631440 19240 631760
rect 34058 631445 34368 631755
rect 18920 625440 19240 625760
rect 34058 625445 34368 625755
rect 404767 625529 407227 627989
rect 428434 625534 430884 627984
rect 18920 622440 19240 622760
rect 34058 622445 34368 622755
rect 18920 619440 19240 619760
rect 34058 619445 34368 619755
rect 18920 616440 19240 616760
rect 34058 616445 34368 616755
rect 18920 613440 19240 613760
rect 34058 613445 34368 613755
rect 404907 613359 407367 615819
rect 428429 613359 430889 615819
rect 18920 610440 19240 610760
rect 34058 610445 34368 610755
rect 18920 607440 19240 607760
rect 34058 607445 34368 607755
rect 18920 604440 19240 604760
rect 34058 604445 34368 604755
rect 18920 601440 19240 601760
rect 34058 601445 34368 601755
rect 404418 599720 406878 602180
rect 428434 599725 430884 602175
rect 18920 598440 19240 598760
rect 34058 598445 34368 598755
rect 18920 595440 19240 595760
rect 34058 595445 34368 595755
rect 18920 592440 19240 592760
rect 34058 592445 34368 592755
rect 18920 589440 19240 589760
rect 34058 589445 34368 589755
rect 18920 586440 19240 586760
rect 34058 586445 34368 586755
rect 403718 584893 406178 587353
rect 428434 584898 430884 587348
rect 18920 583440 19240 583760
rect 34058 583445 34368 583755
rect 18920 580440 19240 580760
rect 34058 580445 34368 580755
rect 18920 577440 19240 577760
rect 34058 577445 34368 577755
rect 18920 574440 19240 574760
rect 34058 574445 34368 574755
rect 18920 571440 19240 571760
rect 34058 571445 34368 571755
rect 18920 568440 19240 568760
rect 34058 568445 34368 568755
rect 18920 565440 19240 565760
rect 34058 565445 34368 565755
rect 404353 563818 406813 566278
rect 428434 563823 430884 566273
rect 18920 562440 19240 562760
rect 34058 562445 34368 562755
rect 18920 559440 19240 559760
rect 34058 559445 34368 559755
rect 18920 556440 19240 556760
rect 34058 556445 34368 556755
rect 18920 553440 19240 553760
rect 34058 553445 34368 553755
rect 18920 550440 19240 550760
rect 34058 550445 34368 550755
rect 404427 550005 406887 552465
rect 428434 550010 430884 552460
rect 18920 547440 19240 547760
rect 34058 547445 34368 547755
rect 18920 544440 19240 544760
rect 34058 544445 34368 544755
rect 18920 541440 19240 541760
rect 34058 541445 34368 541755
rect 404133 540381 406593 542841
rect 428434 540386 430884 542836
rect 18920 538440 19240 538760
rect 34058 538445 34368 538755
rect 18920 535440 19240 535760
rect 34058 535445 34368 535755
rect 18920 532440 19240 532760
rect 34058 532445 34368 532755
rect 18920 529440 19240 529760
rect 34058 529445 34368 529755
rect 404133 529433 406593 531893
rect 428434 529438 430884 531888
rect 18920 526440 19240 526760
rect 34058 526445 34368 526755
rect 18920 523440 19240 523760
rect 34058 523445 34368 523755
rect 18920 520440 19240 520760
rect 34058 520445 34368 520755
rect 18920 517440 19240 517760
rect 34058 517445 34368 517755
rect 18920 511440 19240 511760
rect 34058 511445 34368 511755
rect 404179 510483 406639 512943
rect 428434 510488 430884 512938
rect 18920 508440 19240 508760
rect 34058 508445 34368 508755
rect 18920 505440 19240 505760
rect 34058 505445 34368 505755
rect 18920 502440 19240 502760
rect 34058 502445 34368 502755
rect 18920 499440 19240 499760
rect 34058 499445 34368 499755
rect 18920 496440 19240 496760
rect 34058 496445 34368 496755
rect 18920 493440 19240 493760
rect 34058 493445 34368 493755
rect 18920 490440 19240 490760
rect 34058 490445 34368 490755
rect 18920 487440 19240 487760
rect 34058 487445 34368 487755
rect 18920 484440 19240 484760
rect 34058 484445 34368 484755
rect 404460 483947 406920 486407
rect 428434 483952 430884 486402
rect 18920 481440 19240 481760
rect 34058 481445 34368 481755
rect 18920 478440 19240 478760
rect 34058 478445 34368 478755
rect 18920 475440 19240 475760
rect 34058 475445 34368 475755
rect 18920 472440 19240 472760
rect 34058 472445 34368 472755
rect 18920 469440 19240 469760
rect 34058 469445 34368 469755
rect 18920 466440 19240 466760
rect 34058 466445 34368 466755
rect 18920 463440 19240 463760
rect 34058 463445 34368 463755
rect 18920 460440 19240 460760
rect 34058 460445 34368 460755
rect 18920 457440 19240 457760
rect 34058 457445 34368 457755
rect 18920 454440 19240 454760
rect 34058 454445 34368 454755
rect 18920 451440 19240 451760
rect 34058 451445 34368 451755
rect 18920 448440 19240 448760
rect 34058 448445 34368 448755
rect 404481 447502 406941 449962
rect 428434 447507 430884 449957
rect 18920 445440 19240 445760
rect 34058 445445 34368 445755
rect 18920 442440 19240 442760
rect 34058 442445 34368 442755
rect 18920 439440 19240 439760
rect 34058 439445 34368 439755
rect 18920 436440 19240 436760
rect 34058 436445 34368 436755
rect 18920 433440 19240 433760
rect 34058 433445 34368 433755
rect 18920 430440 19240 430760
rect 34058 430445 34368 430755
rect 18920 427440 19240 427760
rect 34058 427445 34368 427755
rect 18920 424440 19240 424760
rect 34058 424445 34368 424755
rect 18920 421440 19240 421760
rect 34058 421445 34368 421755
rect 1553 420363 1655 420465
rect 4929 377141 5031 377243
rect 404813 419119 407273 421579
rect 428434 419124 430884 421574
rect 18920 418440 19240 418760
rect 34058 418445 34368 418755
rect 18920 415440 19240 415760
rect 34058 415445 34368 415755
rect 18920 412440 19240 412760
rect 34058 412445 34368 412755
rect 18920 409440 19240 409760
rect 34058 409445 34368 409755
rect 404579 407231 407039 409691
rect 428434 407236 430884 409686
rect 18920 406440 19240 406760
rect 34058 406445 34368 406755
rect 18920 403440 19240 403760
rect 34058 403445 34368 403755
rect 18920 397440 19240 397760
rect 34058 397445 34368 397755
rect 18920 394440 19240 394760
rect 34058 394445 34368 394755
rect 18920 391440 19240 391760
rect 34058 391445 34368 391755
rect 18920 388440 19240 388760
rect 34058 388445 34368 388755
rect 18920 385440 19240 385760
rect 34058 385445 34368 385755
rect 18920 382440 19240 382760
rect 34058 382445 34368 382755
rect 18920 379440 19240 379760
rect 34058 379445 34368 379755
rect 414098 377472 414388 377762
rect 413990 376785 414280 377075
rect 18920 376440 19240 376760
rect 34058 376445 34368 376755
rect 414243 375918 414533 376208
rect 414026 374363 414316 374653
rect 413994 373764 414284 374054
rect 18920 373440 19240 373760
rect 34058 373445 34368 373755
rect 414352 372904 414642 373194
rect 414245 372187 414535 372477
rect 414352 371542 414642 371832
rect 414776 371005 415066 371295
rect 18920 370440 19240 370760
rect 34058 370445 34368 370755
rect 413772 370414 414062 370704
rect 18920 367440 19240 367760
rect 34058 367445 34368 367755
rect 18920 364440 19240 364760
rect 34058 364445 34368 364755
rect 21725 359402 21835 359512
rect 22916 358859 23018 358961
rect 1924 350824 4374 353274
rect 26650 350819 29110 353279
rect 1924 346295 4374 348745
rect 26576 346290 29036 348750
rect 1924 341785 4374 344235
rect 26576 341780 29036 344240
rect 5665 336687 5767 336789
rect 5660 327483 5772 327595
rect 1924 313460 4374 315910
rect 39936 313455 42396 315915
rect 8387 261245 8457 261315
rect 404525 359715 406985 362175
rect 428434 359720 430884 362170
rect 365000 358724 365170 358894
rect 55312 345441 55622 345751
rect 58312 345441 58622 345751
rect 61312 345441 61622 345751
rect 64312 345441 64622 345751
rect 67312 345441 67622 345751
rect 70312 345441 70622 345751
rect 73312 345441 73622 345751
rect 76312 345441 76622 345751
rect 79312 345441 79622 345751
rect 82312 345441 82622 345751
rect 85312 345441 85622 345751
rect 88312 345441 88622 345751
rect 91312 345441 91622 345751
rect 94312 345441 94622 345751
rect 97312 345441 97622 345751
rect 100312 345441 100622 345751
rect 103312 345441 103622 345751
rect 106312 345441 106622 345751
rect 109312 345441 109622 345751
rect 112312 345441 112622 345751
rect 115312 345441 115622 345751
rect 118312 345441 118622 345751
rect 121312 345441 121622 345751
rect 124312 345441 124622 345751
rect 127312 345441 127622 345751
rect 130312 345441 130622 345751
rect 133312 345441 133622 345751
rect 136312 345441 136622 345751
rect 139312 345441 139622 345751
rect 142312 345441 142622 345751
rect 145312 345441 145622 345751
rect 148312 345441 148622 345751
rect 151312 345441 151622 345751
rect 154312 345441 154622 345751
rect 157312 345441 157622 345751
rect 160312 345441 160622 345751
rect 163312 345441 163622 345751
rect 166312 345441 166622 345751
rect 169312 345441 169622 345751
rect 172312 345441 172622 345751
rect 175312 345441 175622 345751
rect 178312 345441 178622 345751
rect 181312 345441 181622 345751
rect 184312 345441 184622 345751
rect 187312 345441 187622 345751
rect 190312 345441 190622 345751
rect 193312 345441 193622 345751
rect 196312 345441 196622 345751
rect 199312 345441 199622 345751
rect 202312 345441 202622 345751
rect 205312 345441 205622 345751
rect 208312 345441 208622 345751
rect 211312 345441 211622 345751
rect 214312 345441 214622 345751
rect 217312 345441 217622 345751
rect 220312 345441 220622 345751
rect 223312 345441 223622 345751
rect 226312 345441 226622 345751
rect 229312 345441 229622 345751
rect 232312 345441 232622 345751
rect 235312 345441 235622 345751
rect 238312 345441 238622 345751
rect 241312 345441 241622 345751
rect 244312 345441 244622 345751
rect 247312 345441 247622 345751
rect 250312 345441 250622 345751
rect 253312 345441 253622 345751
rect 256312 345441 256622 345751
rect 259312 345441 259622 345751
rect 262312 345441 262622 345751
rect 265312 345441 265622 345751
rect 268312 345441 268622 345751
rect 271312 345441 271622 345751
rect 274312 345441 274622 345751
rect 277312 345441 277622 345751
rect 280312 345441 280622 345751
rect 283312 345441 283622 345751
rect 286312 345441 286622 345751
rect 289312 345441 289622 345751
rect 292312 345441 292622 345751
rect 295312 345441 295622 345751
rect 298312 345441 298622 345751
rect 301312 345441 301622 345751
rect 304312 345441 304622 345751
rect 307312 345441 307622 345751
rect 310312 345441 310622 345751
rect 313312 345441 313622 345751
rect 316312 345441 316622 345751
rect 319312 345441 319622 345751
rect 325312 345441 325622 345751
rect 328312 345441 328622 345751
rect 331312 345441 331622 345751
rect 334312 345441 334622 345751
rect 337312 345441 337622 345751
rect 340312 345441 340622 345751
rect 343312 345441 343622 345751
rect 346312 345441 346622 345751
rect 349312 345441 349622 345751
rect 352312 345441 352622 345751
rect 355312 345441 355622 345751
rect 358312 345441 358622 345751
rect 55307 323107 55627 323427
rect 58307 323107 58627 323427
rect 61307 323107 61627 323427
rect 64307 323107 64627 323427
rect 67307 323107 67627 323427
rect 70307 323107 70627 323427
rect 73307 323107 73627 323427
rect 76307 323107 76627 323427
rect 79307 323107 79627 323427
rect 82307 323107 82627 323427
rect 85307 323107 85627 323427
rect 88307 323107 88627 323427
rect 91307 323107 91627 323427
rect 94307 323107 94627 323427
rect 97307 323107 97627 323427
rect 100307 323107 100627 323427
rect 103307 323107 103627 323427
rect 106307 323107 106627 323427
rect 109307 323107 109627 323427
rect 112307 323107 112627 323427
rect 115307 323107 115627 323427
rect 118307 323107 118627 323427
rect 121307 323107 121627 323427
rect 124307 323107 124627 323427
rect 127307 323107 127627 323427
rect 130307 323107 130627 323427
rect 133307 323107 133627 323427
rect 136307 323107 136627 323427
rect 139307 323107 139627 323427
rect 142307 323107 142627 323427
rect 145307 323107 145627 323427
rect 148307 323107 148627 323427
rect 151307 323107 151627 323427
rect 154307 323107 154627 323427
rect 157307 323107 157627 323427
rect 160307 323107 160627 323427
rect 163307 323107 163627 323427
rect 166307 323107 166627 323427
rect 169307 323107 169627 323427
rect 172307 323107 172627 323427
rect 175307 323107 175627 323427
rect 178307 323107 178627 323427
rect 181307 323107 181627 323427
rect 184307 323107 184627 323427
rect 187307 323107 187627 323427
rect 190307 323107 190627 323427
rect 193307 323107 193627 323427
rect 196307 323107 196627 323427
rect 199307 323107 199627 323427
rect 202307 323107 202627 323427
rect 205307 323107 205627 323427
rect 208307 323107 208627 323427
rect 211307 323107 211627 323427
rect 214307 323107 214627 323427
rect 217307 323107 217627 323427
rect 220307 323107 220627 323427
rect 223307 323107 223627 323427
rect 226307 323107 226627 323427
rect 229307 323107 229627 323427
rect 232307 323107 232627 323427
rect 235307 323107 235627 323427
rect 238307 323107 238627 323427
rect 241307 323107 241627 323427
rect 244307 323107 244627 323427
rect 247307 323107 247627 323427
rect 250307 323107 250627 323427
rect 253307 323107 253627 323427
rect 256307 323107 256627 323427
rect 259307 323107 259627 323427
rect 262307 323107 262627 323427
rect 265307 323107 265627 323427
rect 268307 323107 268627 323427
rect 271307 323107 271627 323427
rect 274307 323107 274627 323427
rect 277307 323107 277627 323427
rect 280307 323107 280627 323427
rect 283307 323107 283627 323427
rect 286307 323107 286627 323427
rect 289307 323107 289627 323427
rect 292307 323107 292627 323427
rect 295307 323107 295627 323427
rect 298307 323107 298627 323427
rect 301307 323107 301627 323427
rect 304307 323107 304627 323427
rect 307307 323107 307627 323427
rect 310307 323107 310627 323427
rect 313307 323107 313627 323427
rect 316307 323107 316627 323427
rect 319307 323107 319627 323427
rect 325307 323107 325627 323427
rect 328307 323107 328627 323427
rect 331307 323107 331627 323427
rect 334307 323107 334627 323427
rect 337307 323107 337627 323427
rect 340307 323107 340627 323427
rect 343307 323107 343627 323427
rect 346307 323107 346627 323427
rect 349307 323107 349627 323427
rect 352307 323107 352627 323427
rect 355307 323107 355627 323427
rect 372481 336604 372781 336904
rect 375481 336604 375781 336904
rect 378481 336604 378781 336904
rect 381481 336604 381781 336904
rect 384481 336604 384781 336904
rect 387481 336604 387781 336904
rect 390481 336604 390781 336904
rect 393481 336604 393781 336904
rect 396481 336604 396781 336904
rect 358307 323107 358627 323427
rect 55921 248857 56023 248959
rect 287969 228295 290419 230745
rect 180921 207000 181211 207290
rect 183921 207000 184211 207290
rect 186921 207000 187211 207290
rect 189921 207000 190211 207290
rect 192921 207000 193211 207290
rect 195921 207000 196211 207290
rect 198921 207000 199211 207290
rect 201921 207000 202211 207290
rect 204921 207000 205211 207290
rect 9016 191227 9126 191337
rect 175769 188183 175929 188343
rect 175764 186467 175934 186637
rect 21843 121235 21945 121337
rect 177606 180467 177776 180637
rect 180877 172519 181177 172819
rect 183877 172519 184177 172819
rect 186877 172519 187177 172819
rect 189877 172519 190177 172819
rect 192877 172519 193177 172819
rect 195877 172519 196177 172819
rect 198877 172519 199177 172819
rect 201877 172519 202177 172819
rect 204877 172519 205177 172819
rect 287964 116498 290424 118958
rect 33627 78034 33717 78124
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 703390 418394 704800
rect 413394 703190 427730 703390
rect 413394 702300 418394 703190
rect 18694 692120 21194 702300
rect 68940 693513 71440 702300
rect 122330 696788 124830 702300
rect 122330 696678 126146 696788
rect 122330 693513 124830 696678
rect 18694 692119 22220 692120
rect 18694 692011 22111 692119
rect 22219 692011 22225 692119
rect 18694 692010 22220 692011
rect 7013 688094 7331 688099
rect 7012 688093 7332 688094
rect 7012 687775 7013 688093
rect 7331 687775 7332 688093
rect 18694 687950 21194 692010
rect 7012 687774 7332 687775
rect 7013 687769 7331 687774
rect 1920 686010 4378 686015
rect 1919 686009 4379 686010
rect -800 682742 1700 685242
rect 1919 683551 1920 686009
rect 4378 683551 4379 686009
rect 28656 685552 28760 685577
rect 28656 685484 28682 685552
rect 28750 685484 28760 685552
rect 28656 685460 28760 685484
rect 1919 683550 4379 683551
rect 26797 684464 26807 684469
rect 1920 683545 4378 683550
rect -800 680242 8830 682742
rect 26797 682004 26802 684464
rect 26797 681999 26807 682004
rect 29267 681999 29273 684469
rect 9017 680862 9125 680867
rect 9016 680861 9126 680862
rect 9016 680753 9017 680861
rect 9125 680753 9126 680861
rect 9016 680752 9126 680753
rect 9017 680747 9125 680752
rect 1920 678115 4378 678120
rect 1919 678114 4379 678115
rect 1919 675656 1920 678114
rect 4378 675656 4379 678114
rect 1919 675655 4379 675656
rect 1920 675650 4378 675655
rect 1920 672893 4378 672898
rect 1919 672892 4379 672893
rect 1919 670434 1920 672892
rect 4378 670434 4379 672892
rect 1919 670433 4379 670434
rect 1920 670428 4378 670433
rect 6330 658270 8830 680242
rect 26505 678115 26515 678120
rect 26505 675655 26510 678115
rect 26505 675650 26515 675655
rect 28975 675650 28981 678120
rect 69665 676375 69775 693513
rect 69660 676370 69780 676375
rect 69660 676260 69665 676370
rect 69775 676260 69780 676370
rect 69660 676255 69780 676260
rect 10675 675140 10783 675145
rect 10674 675139 50936 675140
rect 10674 675031 10675 675139
rect 10783 675031 50936 675139
rect 10674 675030 50936 675031
rect 10675 675025 10783 675030
rect 50826 674598 50936 675030
rect 126036 674594 126146 696678
rect 143668 694390 144068 694396
rect 143668 693995 143673 694000
rect 144063 693995 144068 694000
rect 143668 693990 144068 693995
rect 177230 693513 179730 702300
rect 228438 698529 229478 698530
rect 228433 697491 228439 698529
rect 229477 697491 229483 698529
rect 331191 698285 332129 698286
rect 178455 689121 178515 693513
rect 178450 689116 178520 689121
rect 178450 689056 178455 689116
rect 178515 689056 178520 689116
rect 178450 689051 178520 689056
rect 228438 686295 229478 697491
rect 331186 697349 331192 698285
rect 332128 697349 332134 698285
rect 147741 686095 233572 686295
rect 137056 675252 137386 675257
rect 137056 674932 137061 675252
rect 137381 674932 137386 675252
rect 147741 675242 147941 686095
rect 228438 685734 229478 686095
rect 331191 685196 332129 697349
rect 148251 684996 334616 685196
rect 148251 675274 148451 684996
rect 331191 684805 332129 684996
rect 427530 683959 427730 703190
rect 465394 702300 470394 704800
rect 150041 683839 433994 683959
rect 150041 675080 150161 683839
rect 427530 683735 427730 683839
rect 152091 683277 152211 683401
rect 466776 683277 469276 702300
rect 510594 698160 515394 704800
rect 520594 698160 525394 704800
rect 566594 702300 571594 704800
rect 566594 690142 571476 702300
rect 553288 689282 571476 690142
rect 152091 683157 471789 683277
rect 152091 675080 152211 683157
rect 466776 681546 469276 683157
rect 436510 680180 436690 680185
rect 396231 680010 436515 680180
rect 436685 680010 436690 680180
rect 137056 674927 137386 674932
rect 50826 674482 50936 674488
rect 126031 674486 126037 674594
rect 126145 674486 126151 674594
rect 126036 674485 126146 674486
rect 137061 672916 137381 674927
rect 396231 674825 396401 680010
rect 436510 680005 436690 680010
rect 396231 674665 396236 674825
rect 396396 674665 396401 674825
rect 396231 674660 396401 674665
rect 155830 674108 156210 674114
rect 140600 673734 140742 673767
rect 231033 673996 231353 673997
rect 140600 673729 140632 673734
rect 140702 673729 140742 673734
rect 140600 673659 140627 673729
rect 140707 673659 140742 673729
rect 140600 673640 140742 673659
rect 147221 672916 147311 673734
rect 155830 673733 155835 673738
rect 156205 673733 156210 673738
rect 155830 673728 156210 673733
rect 231028 673678 231034 673996
rect 231352 673678 231358 673996
rect 152416 673585 152536 673590
rect 152416 673475 152421 673585
rect 152531 673475 152536 673585
rect 152416 673470 152536 673475
rect 231033 673374 231038 673678
rect 231348 673374 231353 673678
rect 231033 673369 231353 673374
rect 26338 672893 26348 672898
rect 26338 670433 26343 672893
rect 26338 670428 26348 670433
rect 28808 670428 28814 672898
rect 55254 672826 147311 672916
rect 55377 671464 55467 672826
rect 137061 672795 137381 672826
rect 403004 672740 403010 675200
rect 405470 672740 508212 675200
rect 140564 671134 140731 671159
rect 140564 671066 140633 671134
rect 140701 671066 140731 671134
rect 140564 671035 140731 671066
rect 402810 670886 405270 670892
rect 492825 670886 495285 671161
rect 501550 670886 504010 670892
rect 143668 670736 144068 670741
rect 143668 670731 143673 670736
rect 144063 670731 144068 670736
rect 143668 670335 144068 670341
rect 386054 668426 395680 670886
rect 401993 668426 402810 670886
rect 405270 668426 501550 670886
rect 504010 668426 508212 670886
rect 18909 667435 18915 667765
rect 19235 667760 19245 667765
rect 34054 667760 34372 667765
rect 19240 667440 19245 667760
rect 34053 667759 34373 667760
rect 34053 667441 34054 667759
rect 34372 667441 34373 667759
rect 34053 667440 34373 667441
rect 19235 667435 19245 667440
rect 34054 667435 34372 667440
rect 18909 664435 18915 664765
rect 19235 664760 19245 664765
rect 34054 664760 34372 664765
rect 19240 664440 19245 664760
rect 34053 664759 34373 664760
rect 34053 664441 34054 664759
rect 34372 664441 34373 664759
rect 53664 664728 53982 664733
rect 34053 664440 34373 664441
rect 53663 664727 53983 664728
rect 19235 664435 19245 664440
rect 34054 664435 34372 664440
rect 53663 664409 53664 664727
rect 53982 664409 53983 664727
rect 53663 664408 53983 664409
rect 53664 664403 53982 664408
rect 32571 662310 32889 662315
rect 18814 661990 18820 662310
rect 19140 662309 32890 662310
rect 19140 661991 32571 662309
rect 32889 661991 32890 662309
rect 19140 661990 32890 661991
rect 32571 661985 32889 661990
rect 18909 661435 18915 661765
rect 19235 661760 19245 661765
rect 34054 661760 34372 661765
rect 19240 661440 19245 661760
rect 34053 661759 34373 661760
rect 34053 661441 34054 661759
rect 34372 661441 34373 661759
rect 34053 661440 34373 661441
rect 19235 661435 19245 661440
rect 34054 661435 34372 661440
rect 32571 659310 32889 659315
rect 18814 658990 18820 659310
rect 19140 659309 32890 659310
rect 19140 658991 32571 659309
rect 32889 658991 32890 659309
rect 19140 658990 32890 658991
rect 32571 658985 32889 658990
rect 18909 658435 18915 658765
rect 19235 658760 19245 658765
rect 34054 658760 34372 658765
rect 19240 658440 19245 658760
rect 34053 658759 34373 658760
rect 34053 658441 34054 658759
rect 34372 658441 34373 658759
rect 34053 658440 34373 658441
rect 19235 658435 19245 658440
rect 34054 658435 34372 658440
rect 6330 657331 14285 658270
rect 6330 657326 13652 657331
rect 6330 657006 13647 657326
rect 6330 657001 13652 657006
rect 13972 657001 14285 657331
rect 6330 655770 14285 657001
rect 32571 656310 32889 656315
rect 18814 655990 18820 656310
rect 19140 656309 32890 656310
rect 19140 655991 32571 656309
rect 32889 655991 32890 656309
rect 19140 655990 32890 655991
rect 32571 655985 32889 655990
rect 18909 655435 18915 655765
rect 19235 655760 19245 655765
rect 34054 655760 34372 655765
rect 19240 655440 19245 655760
rect 34053 655759 34373 655760
rect 34053 655441 34054 655759
rect 34372 655441 34373 655759
rect 34053 655440 34373 655441
rect 19235 655435 19245 655440
rect 34054 655435 34372 655440
rect 32571 653310 32889 653315
rect 18814 652990 18820 653310
rect 19140 653309 32890 653310
rect 19140 652991 32571 653309
rect 32889 652991 32890 653309
rect 19140 652990 32890 652991
rect 32571 652985 32889 652990
rect 18909 652435 18915 652765
rect 19235 652760 19245 652765
rect 34054 652760 34372 652765
rect 19240 652440 19245 652760
rect 34053 652759 34373 652760
rect 34053 652441 34054 652759
rect 34372 652441 34373 652759
rect 34053 652440 34373 652441
rect 19235 652435 19245 652440
rect 34054 652435 34372 652440
rect 11078 649252 14835 651712
rect 17295 649252 17301 651712
rect 32571 650310 32889 650315
rect 18814 649990 18820 650310
rect 19140 650309 32890 650310
rect 19140 649991 32571 650309
rect 32889 649991 32890 650309
rect 19140 649990 32890 649991
rect 32571 649985 32889 649990
rect 18909 649435 18915 649765
rect 19235 649760 19245 649765
rect 34054 649760 34372 649765
rect 19240 649440 19245 649760
rect 34053 649759 34373 649760
rect 34053 649441 34054 649759
rect 34372 649441 34373 649759
rect 34053 649440 34373 649441
rect 19235 649435 19245 649440
rect 34054 649435 34372 649440
rect 11078 648642 13538 649252
rect -800 646302 13538 648642
rect 32571 647310 32889 647315
rect 18814 646990 18820 647310
rect 19140 647309 32890 647310
rect 19140 646991 32571 647309
rect 32889 646991 32890 647309
rect 386054 647181 388514 668426
rect 402810 668420 405270 668426
rect 397829 665132 398129 665265
rect 397824 665127 398134 665132
rect 397824 664827 397829 665127
rect 398129 664827 398134 665127
rect 397824 664822 398134 664827
rect 424844 656028 425014 656029
rect 424839 655860 424845 656028
rect 425013 655860 425019 656028
rect 424844 655859 425014 655860
rect 428429 652869 430889 668426
rect 492825 652599 495285 668426
rect 501550 668420 504010 668426
rect 428429 650403 430889 650409
rect 492820 650141 492826 652599
rect 495284 650141 495290 652599
rect 492825 650140 495285 650141
rect 553288 648399 554148 689282
rect 568976 689047 571476 689282
rect 574600 682984 582176 683000
rect 574600 682800 584800 682984
rect 574440 682402 584800 682800
rect 574440 678818 575238 682402
rect 582000 678818 584800 682402
rect 574440 678370 584800 678818
rect 582300 677984 584800 678370
rect 553283 647541 553289 648399
rect 554147 647541 554153 648399
rect 553288 647540 554148 647541
rect 19140 646990 32890 646991
rect 32571 646985 32889 646990
rect 18909 646435 18915 646765
rect 19235 646760 19245 646765
rect 34054 646760 34372 646765
rect 19240 646440 19245 646760
rect 34053 646759 34373 646760
rect 34053 646441 34054 646759
rect 34372 646441 34373 646759
rect 34053 646440 34373 646441
rect 19235 646435 19245 646440
rect 34054 646435 34372 646440
rect -800 643842 14754 646302
rect 17214 645406 17220 646302
rect 17214 645086 21778 645406
rect 17214 643842 17220 645086
rect 21458 644310 21778 645086
rect 32571 644310 32889 644315
rect 18814 643990 18820 644310
rect 19140 644309 32890 644310
rect 19140 643991 32571 644309
rect 32889 643991 32890 644309
rect 19140 643990 32890 643991
rect 11078 642190 13538 643842
rect 18909 643435 18915 643765
rect 19235 643760 19245 643765
rect 19240 643440 19245 643760
rect 19235 643435 19245 643440
rect 22197 642190 22517 643990
rect 32571 643985 32889 643990
rect 34054 643760 34372 643765
rect 34053 643759 34373 643760
rect 34053 643441 34054 643759
rect 34372 643441 34373 643759
rect 34053 643440 34373 643441
rect 34054 643435 34372 643440
rect 11078 641870 22517 642190
rect 412596 642124 412602 644584
rect 11078 639529 13538 641870
rect 32571 641310 32889 641315
rect 18814 640990 18820 641310
rect 19140 641309 32890 641310
rect 19140 640991 32571 641309
rect 32889 640991 32890 641309
rect 19140 640990 32890 640991
rect 18909 640435 18915 640765
rect 19235 640760 19245 640765
rect 19240 640440 19245 640760
rect 19235 640435 19245 640440
rect 21901 639529 22221 640990
rect 32571 640985 32889 640990
rect 34054 640760 34372 640765
rect 34053 640759 34373 640760
rect 34053 640441 34054 640759
rect 34372 640441 34373 640759
rect 34053 640440 34373 640441
rect 34054 640435 34372 640440
rect 412509 639784 412602 642124
rect 417402 639784 584800 644584
rect 11078 639209 22221 639529
rect 11078 638642 13538 639209
rect -800 636609 13854 638642
rect 32571 638310 32889 638315
rect 18814 637990 18820 638310
rect 19140 638309 32890 638310
rect 19140 637991 32571 638309
rect 32889 637991 32890 638309
rect 19140 637990 32890 637991
rect 18909 637435 18915 637765
rect 19235 637760 19245 637765
rect 19240 637440 19245 637760
rect 19235 637435 19245 637440
rect 22234 636609 22554 637990
rect 32571 637985 32889 637990
rect 34054 637760 34372 637765
rect 34053 637759 34373 637760
rect 34053 637441 34054 637759
rect 34372 637441 34373 637759
rect 34053 637440 34373 637441
rect 34054 637435 34372 637440
rect -800 636289 22554 636609
rect -800 636182 13854 636289
rect -800 633842 13833 636182
rect 32571 635310 32889 635315
rect 18814 634990 18820 635310
rect 19140 635309 32890 635310
rect 19140 634991 32571 635309
rect 32889 634991 32890 635309
rect 19140 634990 32890 634991
rect 18909 634435 18915 634765
rect 19235 634760 19245 634765
rect 19240 634440 19245 634760
rect 19235 634435 19245 634440
rect 11078 633779 13833 633842
rect 22715 633779 23035 634990
rect 32571 634985 32889 634990
rect 34054 634760 34372 634765
rect 34053 634759 34373 634760
rect 34053 634441 34054 634759
rect 34372 634441 34373 634759
rect 451369 634584 456169 634590
rect 460694 634584 465494 634590
rect 480022 634584 484822 639784
rect 34053 634440 34373 634441
rect 34054 634435 34372 634440
rect 11078 633459 23035 633779
rect 11078 631370 13833 633459
rect 32571 632310 32889 632315
rect 18814 631990 18820 632310
rect 19140 632309 32890 632310
rect 19140 631991 32571 632309
rect 32889 631991 32890 632309
rect 412463 632244 412469 634584
rect 19140 631990 32890 631991
rect 32571 631985 32889 631990
rect 18909 631435 18915 631765
rect 19235 631760 19245 631765
rect 34054 631760 34372 631765
rect 19240 631440 19245 631760
rect 34053 631759 34373 631760
rect 34053 631441 34054 631759
rect 34372 631441 34373 631759
rect 34053 631440 34373 631441
rect 19235 631435 19245 631440
rect 34054 631435 34372 631440
rect 11035 630293 13881 631370
rect 11035 627835 11334 630293
rect 13792 627835 13881 630293
rect 412462 629784 412468 632244
rect 417269 629784 451369 634584
rect 456169 629784 460694 634584
rect 465494 629784 584800 634584
rect 451369 629778 456169 629784
rect 460694 629778 465494 629784
rect 11035 627711 13881 627835
rect 11078 624842 13833 627711
rect 18909 625435 18915 625765
rect 19235 625760 19245 625765
rect 34054 625760 34372 625765
rect 19240 625440 19245 625760
rect 34053 625759 34373 625760
rect 34053 625441 34054 625759
rect 34372 625441 34373 625759
rect 404756 625524 404762 627994
rect 407222 627989 407232 627994
rect 428430 627989 430888 627994
rect 407227 625529 407232 627989
rect 428429 627988 430889 627989
rect 428429 625530 428430 627988
rect 430888 625530 430889 627988
rect 428429 625529 430889 625530
rect 407222 625524 407232 625529
rect 428430 625524 430888 625529
rect 34053 625440 34373 625441
rect 19235 625435 19245 625440
rect 34054 625435 34372 625440
rect 11072 622087 11078 624842
rect 13833 622087 13839 624842
rect 32571 623310 32889 623315
rect 18814 622990 18820 623310
rect 19140 623309 32890 623310
rect 19140 622991 32571 623309
rect 32889 622991 32890 623309
rect 19140 622990 32890 622991
rect 32571 622985 32889 622990
rect 18909 622435 18915 622765
rect 19235 622760 19245 622765
rect 34054 622760 34372 622765
rect 19240 622440 19245 622760
rect 34053 622759 34373 622760
rect 34053 622441 34054 622759
rect 34372 622441 34373 622759
rect 34053 622440 34373 622441
rect 19235 622435 19245 622440
rect 34054 622435 34372 622440
rect 11078 617468 13833 622087
rect 32571 620310 32889 620315
rect 18814 619990 18820 620310
rect 19140 620309 32890 620310
rect 19140 619991 32571 620309
rect 32889 619991 32890 620309
rect 19140 619990 32890 619991
rect 32571 619985 32889 619990
rect 18909 619435 18915 619765
rect 19235 619760 19245 619765
rect 34054 619760 34372 619765
rect 19240 619440 19245 619760
rect 34053 619759 34373 619760
rect 34053 619441 34054 619759
rect 34372 619441 34373 619759
rect 34053 619440 34373 619441
rect 19235 619435 19245 619440
rect 34054 619435 34372 619440
rect 11078 614713 15232 617468
rect 17987 614713 17993 617468
rect 32571 617310 32889 617315
rect 18814 616990 18820 617310
rect 19140 617309 32890 617310
rect 19140 616991 32571 617309
rect 32889 616991 32890 617309
rect 19140 616990 32890 616991
rect 32571 616985 32889 616990
rect 18909 616435 18915 616765
rect 19235 616760 19245 616765
rect 34054 616760 34372 616765
rect 19240 616440 19245 616760
rect 34053 616759 34373 616760
rect 34053 616441 34054 616759
rect 34372 616441 34373 616759
rect 34053 616440 34373 616441
rect 19235 616435 19245 616440
rect 34054 616435 34372 616440
rect 11078 610130 13833 614713
rect 32571 614310 32889 614315
rect 18814 613990 18820 614310
rect 19140 614309 32890 614310
rect 19140 613991 32571 614309
rect 32889 613991 32890 614309
rect 19140 613990 32890 613991
rect 32571 613985 32889 613990
rect 18909 613435 18915 613765
rect 19235 613760 19245 613765
rect 34054 613760 34372 613765
rect 19240 613440 19245 613760
rect 34053 613759 34373 613760
rect 34053 613441 34054 613759
rect 34372 613441 34373 613759
rect 34053 613440 34373 613441
rect 19235 613435 19245 613440
rect 34054 613435 34372 613440
rect 404896 613354 404902 615824
rect 407362 615819 407372 615824
rect 407367 613359 407372 615819
rect 407362 613354 407372 613359
rect 428424 615819 430894 615824
rect 428424 613359 428429 615819
rect 430889 613359 430894 615819
rect 428424 613354 430894 613359
rect 32571 611310 32889 611315
rect 18814 610990 18820 611310
rect 19140 611309 32890 611310
rect 19140 610991 32571 611309
rect 32889 610991 32890 611309
rect 19140 610990 32890 610991
rect 32571 610985 32889 610990
rect 18909 610435 18915 610765
rect 19235 610760 19245 610765
rect 34054 610760 34372 610765
rect 19240 610440 19245 610760
rect 34053 610759 34373 610760
rect 34053 610441 34054 610759
rect 34372 610441 34373 610759
rect 34053 610440 34373 610441
rect 19235 610435 19245 610440
rect 34054 610435 34372 610440
rect 11078 607375 13717 610130
rect 16472 607375 16478 610130
rect 32571 608310 32889 608315
rect 18814 607990 18820 608310
rect 19140 608309 32890 608310
rect 19140 607991 32571 608309
rect 32889 607991 32890 608309
rect 19140 607990 32890 607991
rect 32571 607985 32889 607990
rect 18909 607435 18915 607765
rect 19235 607760 19245 607765
rect 34054 607760 34372 607765
rect 19240 607440 19245 607760
rect 34053 607759 34373 607760
rect 34053 607441 34054 607759
rect 34372 607441 34373 607759
rect 34053 607440 34373 607441
rect 19235 607435 19245 607440
rect 34054 607435 34372 607440
rect 11078 605645 13833 607375
rect 11072 602850 11078 605645
rect 13833 602850 13839 605645
rect 32571 605310 32889 605315
rect 18814 604990 18820 605310
rect 19140 605309 32890 605310
rect 19140 604991 32571 605309
rect 32889 604991 32890 605309
rect 19140 604990 32890 604991
rect 32571 604985 32889 604990
rect 18909 604435 18915 604765
rect 19235 604760 19245 604765
rect 34054 604760 34372 604765
rect 19240 604440 19245 604760
rect 34053 604759 34373 604760
rect 34053 604441 34054 604759
rect 34372 604441 34373 604759
rect 34053 604440 34373 604441
rect 19235 604435 19245 604440
rect 34054 604435 34372 604440
rect 11078 597310 13833 602850
rect 32571 602310 32889 602315
rect 18814 601990 18820 602310
rect 19140 602309 32890 602310
rect 19140 601991 32571 602309
rect 32889 601991 32890 602309
rect 19140 601990 32890 601991
rect 32571 601985 32889 601990
rect 18909 601435 18915 601765
rect 19235 601760 19245 601765
rect 34054 601760 34372 601765
rect 19240 601440 19245 601760
rect 34053 601759 34373 601760
rect 34053 601441 34054 601759
rect 34372 601441 34373 601759
rect 34053 601440 34373 601441
rect 19235 601435 19245 601440
rect 34054 601435 34372 601440
rect 404407 599715 404413 602185
rect 406873 602180 406883 602185
rect 428430 602180 430888 602185
rect 406878 599720 406883 602180
rect 428429 602179 430889 602180
rect 428429 599721 428430 602179
rect 430888 599721 430889 602179
rect 428429 599720 430889 599721
rect 406873 599715 406883 599720
rect 428430 599715 430888 599720
rect 32571 599310 32889 599315
rect 18814 598990 18820 599310
rect 19140 599309 32890 599310
rect 19140 598991 32571 599309
rect 32889 598991 32890 599309
rect 19140 598990 32890 598991
rect 32571 598985 32889 598990
rect 18909 598435 18915 598765
rect 19235 598760 19245 598765
rect 34054 598760 34372 598765
rect 19240 598440 19245 598760
rect 34053 598759 34373 598760
rect 34053 598441 34054 598759
rect 34372 598441 34373 598759
rect 34053 598440 34373 598441
rect 19235 598435 19245 598440
rect 34054 598435 34372 598440
rect 11078 594555 14987 597310
rect 17742 594555 17748 597310
rect 413053 596863 415511 596868
rect 480022 596863 484822 629784
rect 413052 596862 484822 596863
rect 32571 596310 32889 596315
rect 18814 595990 18820 596310
rect 19140 596309 32890 596310
rect 19140 595991 32571 596309
rect 32889 595991 32890 596309
rect 19140 595990 32890 595991
rect 32571 595985 32889 595990
rect 18909 595435 18915 595765
rect 19235 595760 19245 595765
rect 34054 595760 34372 595765
rect 19240 595440 19245 595760
rect 34053 595759 34373 595760
rect 34053 595441 34054 595759
rect 34372 595441 34373 595759
rect 34053 595440 34373 595441
rect 19235 595435 19245 595440
rect 34054 595435 34372 595440
rect 11078 589487 13833 594555
rect 413052 594404 413053 596862
rect 415511 594404 484822 596862
rect 413052 594403 484822 594404
rect 413053 594398 415511 594403
rect 32571 593310 32889 593315
rect 18814 592990 18820 593310
rect 19140 593309 32890 593310
rect 19140 592991 32571 593309
rect 32889 592991 32890 593309
rect 19140 592990 32890 592991
rect 32571 592985 32889 592990
rect 18909 592435 18915 592765
rect 19235 592760 19245 592765
rect 34054 592760 34372 592765
rect 19240 592440 19245 592760
rect 34053 592759 34373 592760
rect 34053 592441 34054 592759
rect 34372 592441 34373 592759
rect 34053 592440 34373 592441
rect 19235 592435 19245 592440
rect 34054 592435 34372 592440
rect 32571 590310 32889 590315
rect 18814 589990 18820 590310
rect 19140 590309 32890 590310
rect 19140 589991 32571 590309
rect 32889 589991 32890 590309
rect 19140 589990 32890 589991
rect 32571 589985 32889 589990
rect 11078 586732 14577 589487
rect 17332 586732 17338 589487
rect 18909 589435 18915 589765
rect 19235 589760 19245 589765
rect 34054 589760 34372 589765
rect 19240 589440 19245 589760
rect 34053 589759 34373 589760
rect 34053 589441 34054 589759
rect 34372 589441 34373 589759
rect 34053 589440 34373 589441
rect 19235 589435 19245 589440
rect 34054 589435 34372 589440
rect 32571 587310 32889 587315
rect 18814 586990 18820 587310
rect 19140 587309 32890 587310
rect 19140 586991 32571 587309
rect 32889 586991 32890 587309
rect 19140 586990 32890 586991
rect 32571 586985 32889 586990
rect 11078 584039 13833 586732
rect 18909 586435 18915 586765
rect 19235 586760 19245 586765
rect 34054 586760 34372 586765
rect 19240 586440 19245 586760
rect 34053 586759 34373 586760
rect 34053 586441 34054 586759
rect 34372 586441 34373 586759
rect 34053 586440 34373 586441
rect 19235 586435 19245 586440
rect 34054 586435 34372 586440
rect 403707 584888 403713 587358
rect 406173 587353 406183 587358
rect 428430 587353 430888 587358
rect 406178 584893 406183 587353
rect 428429 587352 430889 587353
rect 428429 584894 428430 587352
rect 430888 584894 430889 587352
rect 428429 584893 430889 584894
rect 406173 584888 406183 584893
rect 428430 584888 430888 584893
rect 32571 584310 32889 584315
rect 11078 581284 14536 584039
rect 17291 581284 17297 584039
rect 18814 583990 18820 584310
rect 19140 584309 32890 584310
rect 19140 583991 32571 584309
rect 32889 583991 32890 584309
rect 19140 583990 32890 583991
rect 32571 583985 32889 583990
rect 18909 583435 18915 583765
rect 19235 583760 19245 583765
rect 34054 583760 34372 583765
rect 19240 583440 19245 583760
rect 34053 583759 34373 583760
rect 34053 583441 34054 583759
rect 34372 583441 34373 583759
rect 34053 583440 34373 583441
rect 19235 583435 19245 583440
rect 34054 583435 34372 583440
rect 32571 581310 32889 581315
rect 11078 578591 13833 581284
rect 18814 580990 18820 581310
rect 19140 581309 32890 581310
rect 19140 580991 32571 581309
rect 32889 580991 32890 581309
rect 19140 580990 32890 580991
rect 32571 580985 32889 580990
rect 18909 580435 18915 580765
rect 19235 580760 19245 580765
rect 34054 580760 34372 580765
rect 19240 580440 19245 580760
rect 34053 580759 34373 580760
rect 34053 580441 34054 580759
rect 34372 580441 34373 580759
rect 34053 580440 34373 580441
rect 19235 580435 19245 580440
rect 34054 580435 34372 580440
rect 11078 575836 14577 578591
rect 17332 575836 17338 578591
rect 32571 578310 32889 578315
rect 18814 577990 18820 578310
rect 19140 578309 32890 578310
rect 19140 577991 32571 578309
rect 32889 577991 32890 578309
rect 19140 577990 32890 577991
rect 32571 577985 32889 577990
rect 18909 577435 18915 577765
rect 19235 577760 19245 577765
rect 34054 577760 34372 577765
rect 19240 577440 19245 577760
rect 34053 577759 34373 577760
rect 34053 577441 34054 577759
rect 34372 577441 34373 577759
rect 34053 577440 34373 577441
rect 19235 577435 19245 577440
rect 34054 577435 34372 577440
rect 11078 571587 13833 575836
rect 32571 575310 32889 575315
rect 18814 574990 18820 575310
rect 19140 575309 32890 575310
rect 19140 574991 32571 575309
rect 32889 574991 32890 575309
rect 19140 574990 32890 574991
rect 32571 574985 32889 574990
rect 18909 574435 18915 574765
rect 19235 574760 19245 574765
rect 34054 574760 34372 574765
rect 19240 574440 19245 574760
rect 34053 574759 34373 574760
rect 34053 574441 34054 574759
rect 34372 574441 34373 574759
rect 34053 574440 34373 574441
rect 19235 574435 19245 574440
rect 34054 574435 34372 574440
rect 480022 573840 484822 594403
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 581085 583562 584800 583674
rect 32571 572310 32889 572315
rect 18814 571990 18820 572310
rect 19140 572309 32890 572310
rect 19140 571991 32571 572309
rect 32889 571991 32890 572309
rect 19140 571990 32890 571991
rect 32571 571985 32889 571990
rect 11078 568832 14946 571587
rect 17701 568832 17707 571587
rect 18909 571435 18915 571765
rect 19235 571760 19245 571765
rect 34054 571760 34372 571765
rect 19240 571440 19245 571760
rect 34053 571759 34373 571760
rect 34053 571441 34054 571759
rect 34372 571441 34373 571759
rect 34053 571440 34373 571441
rect 19235 571435 19245 571440
rect 34054 571435 34372 571440
rect 32571 569310 32889 569315
rect 18814 568990 18820 569310
rect 19140 569309 32890 569310
rect 19140 568991 32571 569309
rect 32889 568991 32890 569309
rect 413169 569040 413175 573840
rect 417975 569040 484822 573840
rect 19140 568990 32890 568991
rect 32571 568985 32889 568990
rect 11078 564870 13833 568832
rect 18909 568435 18915 568765
rect 19235 568760 19245 568765
rect 34054 568760 34372 568765
rect 19240 568440 19245 568760
rect 34053 568759 34373 568760
rect 34053 568441 34054 568759
rect 34372 568441 34373 568759
rect 34053 568440 34373 568441
rect 19235 568435 19245 568440
rect 34054 568435 34372 568440
rect 32571 566310 32889 566315
rect 18814 565990 18820 566310
rect 19140 566309 32890 566310
rect 19140 565991 32571 566309
rect 32889 565991 32890 566309
rect 19140 565990 32890 565991
rect 32571 565985 32889 565990
rect 18909 565435 18915 565765
rect 19235 565760 19245 565765
rect 34054 565760 34372 565765
rect 19240 565440 19245 565760
rect 34053 565759 34373 565760
rect 34053 565441 34054 565759
rect 34372 565441 34373 565759
rect 34053 565440 34373 565441
rect 19235 565435 19245 565440
rect 34054 565435 34372 565440
rect -800 561902 1660 564242
rect 11078 562115 15150 564870
rect 17905 562115 17911 564870
rect 404342 563813 404348 566283
rect 406808 566278 406818 566283
rect 428430 566278 430888 566283
rect 406813 563818 406818 566278
rect 428429 566277 430889 566278
rect 428429 563819 428430 566277
rect 430888 563819 430889 566277
rect 428429 563818 430889 563819
rect 406808 563813 406818 563818
rect 428430 563813 430888 563818
rect 32571 563310 32889 563315
rect 18814 562990 18820 563310
rect 19140 563309 32890 563310
rect 19140 562991 32571 563309
rect 32889 562991 32890 563309
rect 19140 562990 32890 562991
rect 32571 562985 32889 562990
rect 18909 562435 18915 562765
rect 19235 562760 19245 562765
rect 34054 562760 34372 562765
rect 19240 562440 19245 562760
rect 34053 562759 34373 562760
rect 34053 562441 34054 562759
rect 34372 562441 34373 562759
rect 34053 562440 34373 562441
rect 19235 562435 19245 562440
rect 34054 562435 34372 562440
rect 480022 562185 484822 569040
rect -800 559442 1754 561902
rect 11078 560733 13833 562115
rect 11078 557978 15355 560733
rect 18110 557978 18116 560733
rect 32571 560310 32889 560315
rect 18814 559990 18820 560310
rect 19140 560309 32890 560310
rect 19140 559991 32571 560309
rect 32889 559991 32890 560309
rect 19140 559990 32890 559991
rect 32571 559985 32889 559990
rect 18909 559435 18915 559765
rect 19235 559760 19245 559765
rect 34054 559760 34372 559765
rect 19240 559440 19245 559760
rect 34053 559759 34373 559760
rect 34053 559441 34054 559759
rect 34372 559441 34373 559759
rect 34053 559440 34373 559441
rect 19235 559435 19245 559440
rect 34054 559435 34372 559440
rect 11078 554834 13833 557978
rect 413349 557385 413355 562185
rect 418155 557385 484822 562185
rect 32571 557310 32889 557315
rect 18814 556990 18820 557310
rect 19140 557309 32890 557310
rect 19140 556991 32571 557309
rect 32889 556991 32890 557309
rect 19140 556990 32890 556991
rect 32571 556985 32889 556990
rect 18909 556435 18915 556765
rect 19235 556760 19245 556765
rect 34054 556760 34372 556765
rect 19240 556440 19245 556760
rect 34053 556759 34373 556760
rect 34053 556441 34054 556759
rect 34372 556441 34373 556759
rect 34053 556440 34373 556441
rect 19235 556435 19245 556440
rect 34054 556435 34372 556440
rect -800 551902 1660 554242
rect 11078 552079 14659 554834
rect 17414 552079 17420 554834
rect 32571 554310 32889 554315
rect 18814 553990 18820 554310
rect 19140 554309 32890 554310
rect 19140 553991 32571 554309
rect 32889 553991 32890 554309
rect 19140 553990 32890 553991
rect 32571 553985 32889 553990
rect 18909 553435 18915 553765
rect 19235 553760 19245 553765
rect 34054 553760 34372 553765
rect 19240 553440 19245 553760
rect 34053 553759 34373 553760
rect 34053 553441 34054 553759
rect 34372 553441 34373 553759
rect 34053 553440 34373 553441
rect 19235 553435 19245 553440
rect 34054 553435 34372 553440
rect -800 549442 1754 551902
rect 11078 547421 13833 552079
rect 32571 551310 32889 551315
rect 18814 550990 18820 551310
rect 19140 551309 32890 551310
rect 19140 550991 32571 551309
rect 32889 550991 32890 551309
rect 19140 550990 32890 550991
rect 32571 550985 32889 550990
rect 18909 550435 18915 550765
rect 19235 550760 19245 550765
rect 34054 550760 34372 550765
rect 19240 550440 19245 550760
rect 34053 550759 34373 550760
rect 34053 550441 34054 550759
rect 34372 550441 34373 550759
rect 34053 550440 34373 550441
rect 19235 550435 19245 550440
rect 34054 550435 34372 550440
rect 404416 550000 404422 552470
rect 406882 552465 406892 552470
rect 428430 552465 430888 552470
rect 406887 550005 406892 552465
rect 428429 552464 430889 552465
rect 428429 550006 428430 552464
rect 430888 550006 430889 552464
rect 428429 550005 430889 550006
rect 406882 550000 406892 550005
rect 428430 550000 430888 550005
rect 32571 548310 32889 548315
rect 18814 547990 18820 548310
rect 19140 548309 32890 548310
rect 19140 547991 32571 548309
rect 32889 547991 32890 548309
rect 19140 547990 32890 547991
rect 32571 547985 32889 547990
rect 18909 547435 18915 547765
rect 19235 547760 19245 547765
rect 34054 547760 34372 547765
rect 19240 547440 19245 547760
rect 34053 547759 34373 547760
rect 34053 547441 34054 547759
rect 34372 547441 34373 547759
rect 34053 547440 34373 547441
rect 19235 547435 19245 547440
rect 34054 547435 34372 547440
rect 11078 544666 14946 547421
rect 17701 544666 17707 547421
rect 32571 545310 32889 545315
rect 18814 544990 18820 545310
rect 19140 545309 32890 545310
rect 19140 544991 32571 545309
rect 32889 544991 32890 545309
rect 19140 544990 32890 544991
rect 32571 544985 32889 544990
rect 11078 540744 13833 544666
rect 18909 544435 18915 544765
rect 19235 544760 19245 544765
rect 34054 544760 34372 544765
rect 19240 544440 19245 544760
rect 34053 544759 34373 544760
rect 34053 544441 34054 544759
rect 34372 544441 34373 544759
rect 34053 544440 34373 544441
rect 19235 544435 19245 544440
rect 34054 544435 34372 544440
rect 32571 542310 32889 542315
rect 18814 541990 18820 542310
rect 19140 542309 32890 542310
rect 19140 541991 32571 542309
rect 32889 541991 32890 542309
rect 19140 541990 32890 541991
rect 32571 541985 32889 541990
rect 18909 541435 18915 541765
rect 19235 541760 19245 541765
rect 34054 541760 34372 541765
rect 19240 541440 19245 541760
rect 34053 541759 34373 541760
rect 34053 541441 34054 541759
rect 34372 541441 34373 541759
rect 34053 541440 34373 541441
rect 19235 541435 19245 541440
rect 34054 541435 34372 541440
rect 11078 537989 15724 540744
rect 18479 537989 18485 540744
rect 404122 540376 404128 542846
rect 406588 542841 406598 542846
rect 428430 542841 430888 542846
rect 406593 540381 406598 542841
rect 428429 542840 430889 542841
rect 428429 540382 428430 542840
rect 430888 540382 430889 542840
rect 428429 540381 430889 540382
rect 406588 540376 406598 540381
rect 428430 540376 430888 540381
rect 32571 539310 32889 539315
rect 18814 538990 18820 539310
rect 19140 539309 32890 539310
rect 19140 538991 32571 539309
rect 32889 538991 32890 539309
rect 19140 538990 32890 538991
rect 32571 538985 32889 538990
rect 18909 538435 18915 538765
rect 19235 538760 19245 538765
rect 34054 538760 34372 538765
rect 19240 538440 19245 538760
rect 34053 538759 34373 538760
rect 34053 538441 34054 538759
rect 34372 538441 34373 538759
rect 34053 538440 34373 538441
rect 19235 538435 19245 538440
rect 34054 538435 34372 538440
rect 11078 532634 13833 537989
rect 32571 536310 32889 536315
rect 18814 535990 18820 536310
rect 19140 536309 32890 536310
rect 19140 535991 32571 536309
rect 32889 535991 32890 536309
rect 19140 535990 32890 535991
rect 32571 535985 32889 535990
rect 18909 535435 18915 535765
rect 19235 535760 19245 535765
rect 34054 535760 34372 535765
rect 19240 535440 19245 535760
rect 34053 535759 34373 535760
rect 34053 535441 34054 535759
rect 34372 535441 34373 535759
rect 34053 535440 34373 535441
rect 19235 535435 19245 535440
rect 34054 535435 34372 535440
rect 32571 533310 32889 533315
rect 18814 532990 18820 533310
rect 19140 533309 32890 533310
rect 19140 532991 32571 533309
rect 32889 532991 32890 533309
rect 19140 532990 32890 532991
rect 32571 532985 32889 532990
rect 11078 529879 15314 532634
rect 18069 529879 18075 532634
rect 18909 532435 18915 532765
rect 19235 532760 19245 532765
rect 34054 532760 34372 532765
rect 19240 532440 19245 532760
rect 34053 532759 34373 532760
rect 34053 532441 34054 532759
rect 34372 532441 34373 532759
rect 34053 532440 34373 532441
rect 19235 532435 19245 532440
rect 34054 532435 34372 532440
rect 32571 530310 32889 530315
rect 18814 529990 18820 530310
rect 19140 530309 32890 530310
rect 19140 529991 32571 530309
rect 32889 529991 32890 530309
rect 19140 529990 32890 529991
rect 32571 529985 32889 529990
rect 11078 524196 13833 529879
rect 18909 529435 18915 529765
rect 19235 529760 19245 529765
rect 34054 529760 34372 529765
rect 19240 529440 19245 529760
rect 34053 529759 34373 529760
rect 34053 529441 34054 529759
rect 34372 529441 34373 529759
rect 34053 529440 34373 529441
rect 19235 529435 19245 529440
rect 34054 529435 34372 529440
rect 404122 529428 404128 531898
rect 406588 531893 406598 531898
rect 428430 531893 430888 531898
rect 406593 529433 406598 531893
rect 428429 531892 430889 531893
rect 428429 529434 428430 531892
rect 430888 529434 430889 531892
rect 428429 529433 430889 529434
rect 406588 529428 406598 529433
rect 428430 529428 430888 529433
rect 32571 527310 32889 527315
rect 18814 526990 18820 527310
rect 19140 527309 32890 527310
rect 19140 526991 32571 527309
rect 32889 526991 32890 527309
rect 19140 526990 32890 526991
rect 32571 526985 32889 526990
rect 18909 526435 18915 526765
rect 19235 526760 19245 526765
rect 34054 526760 34372 526765
rect 19240 526440 19245 526760
rect 34053 526759 34373 526760
rect 34053 526441 34054 526759
rect 34372 526441 34373 526759
rect 34053 526440 34373 526441
rect 19235 526435 19245 526440
rect 34054 526435 34372 526440
rect 32571 524310 32889 524315
rect 11078 521441 15437 524196
rect 18192 521441 18198 524196
rect 18814 523990 18820 524310
rect 19140 524309 32890 524310
rect 19140 523991 32571 524309
rect 32889 523991 32890 524309
rect 19140 523990 32890 523991
rect 32571 523985 32889 523990
rect 18909 523435 18915 523765
rect 19235 523760 19245 523765
rect 34054 523760 34372 523765
rect 19240 523440 19245 523760
rect 34053 523759 34373 523760
rect 34053 523441 34054 523759
rect 34372 523441 34373 523759
rect 34053 523440 34373 523441
rect 19235 523435 19245 523440
rect 34054 523435 34372 523440
rect 413053 523279 415511 523284
rect 480022 523279 484822 557385
rect 582340 555352 584800 555362
rect 581085 554285 584800 555352
rect 578987 550570 584800 554285
rect 582340 550562 584800 550570
rect 581085 544277 584800 545362
rect 578987 540562 584800 544277
rect 413052 523278 484822 523279
rect 11078 516865 13833 521441
rect 32571 521310 32889 521315
rect 18814 520990 18820 521310
rect 19140 521309 32890 521310
rect 19140 520991 32571 521309
rect 32889 520991 32890 521309
rect 19140 520990 32890 520991
rect 32571 520985 32889 520990
rect 413052 520820 413053 523278
rect 415511 520820 484822 523278
rect 413052 520819 484822 520820
rect 413053 520814 415511 520819
rect 18909 520435 18915 520765
rect 19235 520760 19245 520765
rect 34054 520760 34372 520765
rect 19240 520440 19245 520760
rect 34053 520759 34373 520760
rect 34053 520441 34054 520759
rect 34372 520441 34373 520759
rect 34053 520440 34373 520441
rect 19235 520435 19245 520440
rect 34054 520435 34372 520440
rect 32571 518310 32889 518315
rect 18814 517990 18820 518310
rect 19140 518309 32890 518310
rect 19140 517991 32571 518309
rect 32889 517991 32890 518309
rect 19140 517990 32890 517991
rect 32571 517985 32889 517990
rect 18909 517435 18915 517765
rect 19235 517760 19245 517765
rect 34054 517760 34372 517765
rect 19240 517440 19245 517760
rect 34053 517759 34373 517760
rect 34053 517441 34054 517759
rect 34372 517441 34373 517759
rect 34053 517440 34373 517441
rect 19235 517435 19245 517440
rect 34054 517435 34372 517440
rect 11078 514110 15355 516865
rect 18110 514110 18116 516865
rect 32571 515310 32889 515315
rect 18814 514990 18820 515310
rect 19140 515309 32890 515310
rect 19140 514991 32571 515309
rect 32889 514991 32890 515309
rect 19140 514990 32890 514991
rect 32571 514985 32889 514990
rect 11078 511990 13833 514110
rect 32571 512310 32889 512315
rect 18814 511990 18820 512310
rect 19140 512309 32890 512310
rect 19140 511991 32571 512309
rect 32889 511991 32890 512309
rect 19140 511990 32890 511991
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect 11078 509235 15232 511990
rect 17987 509235 17993 511990
rect 32571 511985 32889 511990
rect 18909 511435 18915 511765
rect 19235 511760 19245 511765
rect 34054 511760 34372 511765
rect 19240 511440 19245 511760
rect 34053 511759 34373 511760
rect 34053 511441 34054 511759
rect 34372 511441 34373 511759
rect 34053 511440 34373 511441
rect 19235 511435 19245 511440
rect 34054 511435 34372 511440
rect 404168 510478 404174 512948
rect 406634 512943 406644 512948
rect 428430 512943 430888 512948
rect 406639 510483 406644 512943
rect 428429 512942 430889 512943
rect 428429 510484 428430 512942
rect 430888 510484 430889 512942
rect 428429 510483 430889 510484
rect 406634 510478 406644 510483
rect 428430 510478 430888 510483
rect 32571 509310 32889 509315
rect 11078 508304 13833 509235
rect 18814 508990 18820 509310
rect 19140 509309 32890 509310
rect 19140 508991 32571 509309
rect 32889 508991 32890 509309
rect 19140 508990 32890 508991
rect 32571 508985 32889 508990
rect 18909 508435 18915 508765
rect 19235 508760 19245 508765
rect 34054 508760 34372 508765
rect 19240 508440 19245 508760
rect 34053 508759 34373 508760
rect 34053 508441 34054 508759
rect 34372 508441 34373 508759
rect 34053 508440 34373 508441
rect 19235 508435 19245 508440
rect 34054 508435 34372 508440
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 11078 505549 15642 508304
rect 18397 505549 18403 508304
rect 32571 506310 32889 506315
rect 18814 505990 18820 506310
rect 19140 506309 32890 506310
rect 19140 505991 32571 506309
rect 32889 505991 32890 506309
rect 19140 505990 32890 505991
rect 32571 505985 32889 505990
rect 11078 499927 13833 505549
rect 18909 505435 18915 505765
rect 19235 505760 19245 505765
rect 34054 505760 34372 505765
rect 19240 505440 19245 505760
rect 34053 505759 34373 505760
rect 34053 505441 34054 505759
rect 34372 505441 34373 505759
rect 34053 505440 34373 505441
rect 19235 505435 19245 505440
rect 34054 505435 34372 505440
rect 32571 503310 32889 503315
rect 18814 502990 18820 503310
rect 19140 503309 32890 503310
rect 19140 502991 32571 503309
rect 32889 502991 32890 503309
rect 19140 502990 32890 502991
rect 32571 502985 32889 502990
rect 18909 502435 18915 502765
rect 19235 502760 19245 502765
rect 34054 502760 34372 502765
rect 19240 502440 19245 502760
rect 34053 502759 34373 502760
rect 34053 502441 34054 502759
rect 34372 502441 34373 502759
rect 34053 502440 34373 502441
rect 19235 502435 19245 502440
rect 34054 502435 34372 502440
rect 32571 500310 32889 500315
rect 18814 499990 18820 500310
rect 19140 500309 32890 500310
rect 19140 499991 32571 500309
rect 32889 499991 32890 500309
rect 19140 499990 32890 499991
rect 32571 499985 32889 499990
rect 11072 497132 11078 499927
rect 13833 497132 13839 499927
rect 18909 499435 18915 499765
rect 19235 499760 19245 499765
rect 34054 499760 34372 499765
rect 19240 499440 19245 499760
rect 34053 499759 34373 499760
rect 34053 499441 34054 499759
rect 34372 499441 34373 499759
rect 34053 499440 34373 499441
rect 19235 499435 19245 499440
rect 34054 499435 34372 499440
rect 32571 497310 32889 497315
rect 11078 492903 13833 497132
rect 18814 496990 18820 497310
rect 19140 497309 32890 497310
rect 19140 496991 32571 497309
rect 32889 496991 32890 497309
rect 413053 497295 415511 497300
rect 480022 497295 484822 520819
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 19140 496990 32890 496991
rect 413052 497294 484822 497295
rect 32571 496985 32889 496990
rect 18909 496435 18915 496765
rect 19235 496760 19245 496765
rect 34054 496760 34372 496765
rect 19240 496440 19245 496760
rect 34053 496759 34373 496760
rect 34053 496441 34054 496759
rect 34372 496441 34373 496759
rect 34053 496440 34373 496441
rect 19235 496435 19245 496440
rect 34054 496435 34372 496440
rect 413052 494836 413053 497294
rect 415511 494836 484822 497294
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 413052 494835 484822 494836
rect 413053 494830 415511 494835
rect 32571 494310 32889 494315
rect 18814 493990 18820 494310
rect 19140 494309 32890 494310
rect 19140 493991 32571 494309
rect 32889 493991 32890 494309
rect 19140 493990 32890 493991
rect 32571 493985 32889 493990
rect 18909 493435 18915 493765
rect 19235 493760 19245 493765
rect 34054 493760 34372 493765
rect 19240 493440 19245 493760
rect 34053 493759 34373 493760
rect 34053 493441 34054 493759
rect 34372 493441 34373 493759
rect 34053 493440 34373 493441
rect 19235 493435 19245 493440
rect 34054 493435 34372 493440
rect 11078 490148 15273 492903
rect 18028 490148 18034 492903
rect 32571 491310 32889 491315
rect 18814 490990 18820 491310
rect 19140 491309 32890 491310
rect 19140 490991 32571 491309
rect 32889 490991 32890 491309
rect 19140 490990 32890 490991
rect 32571 490985 32889 490990
rect 18909 490435 18915 490765
rect 19235 490760 19245 490765
rect 34054 490760 34372 490765
rect 19240 490440 19245 490760
rect 34053 490759 34373 490760
rect 34053 490441 34054 490759
rect 34372 490441 34373 490759
rect 34053 490440 34373 490441
rect 19235 490435 19245 490440
rect 34054 490435 34372 490440
rect 11078 486185 13833 490148
rect 32571 488310 32889 488315
rect 18814 487990 18820 488310
rect 19140 488309 32890 488310
rect 19140 487991 32571 488309
rect 32889 487991 32890 488309
rect 19140 487990 32890 487991
rect 32571 487985 32889 487990
rect 18909 487435 18915 487765
rect 19235 487760 19245 487765
rect 34054 487760 34372 487765
rect 19240 487440 19245 487760
rect 34053 487759 34373 487760
rect 34053 487441 34054 487759
rect 34372 487441 34373 487759
rect 34053 487440 34373 487441
rect 19235 487435 19245 487440
rect 34054 487435 34372 487440
rect 11078 483430 14495 486185
rect 17250 483430 17256 486185
rect 32571 485310 32889 485315
rect 18814 484990 18820 485310
rect 19140 485309 32890 485310
rect 19140 484991 32571 485309
rect 32889 484991 32890 485309
rect 19140 484990 32890 484991
rect 32571 484985 32889 484990
rect 18909 484435 18915 484765
rect 19235 484760 19245 484765
rect 34054 484760 34372 484765
rect 19240 484440 19245 484760
rect 34053 484759 34373 484760
rect 34053 484441 34054 484759
rect 34372 484441 34373 484759
rect 34053 484440 34373 484441
rect 19235 484435 19245 484440
rect 34054 484435 34372 484440
rect 404449 483942 404455 486412
rect 406915 486407 406925 486412
rect 428430 486407 430888 486412
rect 406920 483947 406925 486407
rect 428429 486406 430889 486407
rect 428429 483948 428430 486406
rect 430888 483948 430889 486406
rect 428429 483947 430889 483948
rect 406915 483942 406925 483947
rect 428430 483942 430888 483947
rect -800 468308 891 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect 1366 464931 1478 465323
rect 1366 464874 5772 464931
rect -800 464819 5772 464874
rect -800 464762 1478 464819
rect -800 463580 480 463692
rect -800 462398 480 462510
rect -800 425086 803 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect 1356 421652 1468 421838
rect -800 421540 1468 421652
rect 1356 420470 1468 421540
rect -800 420358 591 420470
rect 1343 420465 1660 420470
rect 1343 420363 1553 420465
rect 1655 420363 1660 420465
rect 1343 420358 1660 420363
rect -800 419176 480 419288
rect -800 381864 979 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect 1356 378430 1468 378793
rect -800 378318 1468 378430
rect 1356 377248 1468 378318
rect -800 377136 824 377248
rect 1285 377243 5036 377248
rect 1285 377141 4929 377243
rect 5031 377141 5036 377243
rect 1285 377136 5036 377141
rect -800 375954 480 376066
rect 1920 353279 4378 353284
rect 1919 353278 4379 353279
rect 1919 350820 1920 353278
rect 4378 350820 4379 353278
rect 1919 350819 4379 350820
rect 1920 350814 4378 350819
rect 1920 348750 4378 348755
rect 1919 348749 4379 348750
rect 1919 346291 1920 348749
rect 4378 346291 4379 348749
rect 1919 346290 4379 346291
rect 1920 346285 4378 346290
rect 1920 344240 4378 344245
rect 1919 344239 4379 344240
rect 1919 341781 1920 344239
rect 4378 341781 4379 344239
rect 1919 341780 4379 341781
rect 1920 341775 4378 341780
rect -800 338642 480 338754
rect -800 337460 480 337572
rect 5660 336789 5772 464819
rect 11078 461424 13833 483430
rect 32571 482310 32889 482315
rect 18814 481990 18820 482310
rect 19140 482309 32890 482310
rect 19140 481991 32571 482309
rect 32889 481991 32890 482309
rect 19140 481990 32890 481991
rect 32571 481985 32889 481990
rect 18909 481435 18915 481765
rect 19235 481760 19245 481765
rect 34054 481760 34372 481765
rect 19240 481440 19245 481760
rect 34053 481759 34373 481760
rect 34053 481441 34054 481759
rect 34372 481441 34373 481759
rect 34053 481440 34373 481441
rect 19235 481435 19245 481440
rect 34054 481435 34372 481440
rect 32571 479310 32889 479315
rect 18814 478990 18820 479310
rect 19140 479309 32890 479310
rect 19140 478991 32571 479309
rect 32889 478991 32890 479309
rect 19140 478990 32890 478991
rect 32571 478985 32889 478990
rect 18909 478435 18915 478765
rect 19235 478760 19245 478765
rect 34054 478760 34372 478765
rect 19240 478440 19245 478760
rect 34053 478759 34373 478760
rect 34053 478441 34054 478759
rect 34372 478441 34373 478759
rect 34053 478440 34373 478441
rect 19235 478435 19245 478440
rect 34054 478435 34372 478440
rect 32571 476310 32889 476315
rect 18814 475990 18820 476310
rect 19140 476309 32890 476310
rect 19140 475991 32571 476309
rect 32889 475991 32890 476309
rect 19140 475990 32890 475991
rect 32571 475985 32889 475990
rect 18909 475435 18915 475765
rect 19235 475760 19245 475765
rect 34054 475760 34372 475765
rect 19240 475440 19245 475760
rect 34053 475759 34373 475760
rect 34053 475441 34054 475759
rect 34372 475441 34373 475759
rect 34053 475440 34373 475441
rect 19235 475435 19245 475440
rect 34054 475435 34372 475440
rect 32571 473310 32889 473315
rect 18814 472990 18820 473310
rect 19140 473309 32890 473310
rect 19140 472991 32571 473309
rect 32889 472991 32890 473309
rect 19140 472990 32890 472991
rect 32571 472985 32889 472990
rect 18909 472435 18915 472765
rect 19235 472760 19245 472765
rect 34054 472760 34372 472765
rect 19240 472440 19245 472760
rect 34053 472759 34373 472760
rect 34053 472441 34054 472759
rect 34372 472441 34373 472759
rect 34053 472440 34373 472441
rect 19235 472435 19245 472440
rect 34054 472435 34372 472440
rect 32571 470310 32889 470315
rect 18814 469990 18820 470310
rect 19140 470309 32890 470310
rect 19140 469991 32571 470309
rect 32889 469991 32890 470309
rect 19140 469990 32890 469991
rect 32571 469985 32889 469990
rect 18909 469435 18915 469765
rect 19235 469760 19245 469765
rect 34054 469760 34372 469765
rect 19240 469440 19245 469760
rect 34053 469759 34373 469760
rect 34053 469441 34054 469759
rect 34372 469441 34373 469759
rect 34053 469440 34373 469441
rect 19235 469435 19245 469440
rect 34054 469435 34372 469440
rect 32571 467310 32889 467315
rect 18814 466990 18820 467310
rect 19140 467309 32890 467310
rect 19140 466991 32571 467309
rect 32889 466991 32890 467309
rect 19140 466990 32890 466991
rect 32571 466985 32889 466990
rect 18909 466435 18915 466765
rect 19235 466760 19245 466765
rect 34054 466760 34372 466765
rect 19240 466440 19245 466760
rect 34053 466759 34373 466760
rect 34053 466441 34054 466759
rect 34372 466441 34373 466759
rect 34053 466440 34373 466441
rect 19235 466435 19245 466440
rect 34054 466435 34372 466440
rect 413053 465331 415511 465336
rect 480022 465331 484822 494835
rect 504833 494140 584800 494252
rect 413052 465330 484822 465331
rect 32571 464310 32889 464315
rect 18814 463990 18820 464310
rect 19140 464309 32890 464310
rect 19140 463991 32571 464309
rect 32889 463991 32890 464309
rect 19140 463990 32890 463991
rect 32571 463985 32889 463990
rect 18909 463435 18915 463765
rect 19235 463760 19245 463765
rect 34054 463760 34372 463765
rect 19240 463440 19245 463760
rect 34053 463759 34373 463760
rect 34053 463441 34054 463759
rect 34372 463441 34373 463759
rect 34053 463440 34373 463441
rect 19235 463435 19245 463440
rect 34054 463435 34372 463440
rect 413052 462872 413053 465330
rect 415511 462872 484822 465330
rect 413052 462871 484822 462872
rect 413053 462866 415511 462871
rect 11072 458587 11078 461424
rect 13833 458587 13839 461424
rect 32571 461310 32889 461315
rect 18814 460990 18820 461310
rect 19140 461309 32890 461310
rect 19140 460991 32571 461309
rect 32889 460991 32890 461309
rect 19140 460990 32890 460991
rect 32571 460985 32889 460990
rect 18909 460435 18915 460765
rect 19235 460760 19245 460765
rect 34054 460760 34372 460765
rect 19240 460440 19245 460760
rect 34053 460759 34373 460760
rect 34053 460441 34054 460759
rect 34372 460441 34373 460759
rect 34053 460440 34373 460441
rect 19235 460435 19245 460440
rect 34054 460435 34372 460440
rect 11078 429929 13833 458587
rect 32571 458310 32889 458315
rect 18814 457990 18820 458310
rect 19140 458309 32890 458310
rect 19140 457991 32571 458309
rect 32889 457991 32890 458309
rect 19140 457990 32890 457991
rect 32571 457985 32889 457990
rect 18909 457435 18915 457765
rect 19235 457760 19245 457765
rect 34054 457760 34372 457765
rect 19240 457440 19245 457760
rect 34053 457759 34373 457760
rect 34053 457441 34054 457759
rect 34372 457441 34373 457759
rect 34053 457440 34373 457441
rect 19235 457435 19245 457440
rect 34054 457435 34372 457440
rect 32571 455310 32889 455315
rect 18814 454990 18820 455310
rect 19140 455309 32890 455310
rect 19140 454991 32571 455309
rect 32889 454991 32890 455309
rect 19140 454990 32890 454991
rect 32571 454985 32889 454990
rect 18909 454435 18915 454765
rect 19235 454760 19245 454765
rect 34054 454760 34372 454765
rect 19240 454440 19245 454760
rect 34053 454759 34373 454760
rect 34053 454441 34054 454759
rect 34372 454441 34373 454759
rect 34053 454440 34373 454441
rect 19235 454435 19245 454440
rect 34054 454435 34372 454440
rect 32571 452310 32889 452315
rect 18814 451990 18820 452310
rect 19140 452309 32890 452310
rect 19140 451991 32571 452309
rect 32889 451991 32890 452309
rect 19140 451990 32890 451991
rect 32571 451985 32889 451990
rect 18909 451435 18915 451765
rect 19235 451760 19245 451765
rect 34054 451760 34372 451765
rect 19240 451440 19245 451760
rect 34053 451759 34373 451760
rect 34053 451441 34054 451759
rect 34372 451441 34373 451759
rect 34053 451440 34373 451441
rect 19235 451435 19245 451440
rect 34054 451435 34372 451440
rect 32571 449310 32889 449315
rect 18814 448990 18820 449310
rect 19140 449309 32890 449310
rect 19140 448991 32571 449309
rect 32889 448991 32890 449309
rect 19140 448990 32890 448991
rect 32571 448985 32889 448990
rect 18909 448435 18915 448765
rect 19235 448760 19245 448765
rect 34054 448760 34372 448765
rect 19240 448440 19245 448760
rect 34053 448759 34373 448760
rect 34053 448441 34054 448759
rect 34372 448441 34373 448759
rect 34053 448440 34373 448441
rect 19235 448435 19245 448440
rect 34054 448435 34372 448440
rect 404470 447497 404476 449967
rect 406936 449962 406946 449967
rect 428430 449962 430888 449967
rect 406941 447502 406946 449962
rect 428429 449961 430889 449962
rect 428429 447503 428430 449961
rect 430888 447503 430889 449961
rect 428429 447502 430889 447503
rect 406936 447497 406946 447502
rect 428430 447497 430888 447502
rect 32571 446310 32889 446315
rect 18814 445990 18820 446310
rect 19140 446309 32890 446310
rect 19140 445991 32571 446309
rect 32889 445991 32890 446309
rect 19140 445990 32890 445991
rect 32571 445985 32889 445990
rect 18909 445435 18915 445765
rect 19235 445760 19245 445765
rect 34054 445760 34372 445765
rect 19240 445440 19245 445760
rect 34053 445759 34373 445760
rect 34053 445441 34054 445759
rect 34372 445441 34373 445759
rect 34053 445440 34373 445441
rect 19235 445435 19245 445440
rect 34054 445435 34372 445440
rect 32571 443310 32889 443315
rect 18814 442990 18820 443310
rect 19140 443309 32890 443310
rect 19140 442991 32571 443309
rect 32889 442991 32890 443309
rect 19140 442990 32890 442991
rect 32571 442985 32889 442990
rect 18909 442435 18915 442765
rect 19235 442760 19245 442765
rect 34054 442760 34372 442765
rect 19240 442440 19245 442760
rect 34053 442759 34373 442760
rect 34053 442441 34054 442759
rect 34372 442441 34373 442759
rect 34053 442440 34373 442441
rect 19235 442435 19245 442440
rect 34054 442435 34372 442440
rect 32571 440310 32889 440315
rect 18814 439990 18820 440310
rect 19140 440309 32890 440310
rect 19140 439991 32571 440309
rect 32889 439991 32890 440309
rect 19140 439990 32890 439991
rect 32571 439985 32889 439990
rect 18909 439435 18915 439765
rect 19235 439760 19245 439765
rect 34054 439760 34372 439765
rect 19240 439440 19245 439760
rect 34053 439759 34373 439760
rect 34053 439441 34054 439759
rect 34372 439441 34373 439759
rect 34053 439440 34373 439441
rect 19235 439435 19245 439440
rect 34054 439435 34372 439440
rect 32571 437310 32889 437315
rect 18814 436990 18820 437310
rect 19140 437309 32890 437310
rect 19140 436991 32571 437309
rect 32889 436991 32890 437309
rect 19140 436990 32890 436991
rect 32571 436985 32889 436990
rect 18909 436435 18915 436765
rect 19235 436760 19245 436765
rect 34054 436760 34372 436765
rect 19240 436440 19245 436760
rect 34053 436759 34373 436760
rect 34053 436441 34054 436759
rect 34372 436441 34373 436759
rect 34053 436440 34373 436441
rect 19235 436435 19245 436440
rect 34054 436435 34372 436440
rect 413053 435898 415511 435903
rect 480022 435898 484822 462871
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 504833 449718 584800 449830
rect 413052 435897 484822 435898
rect 32571 434310 32889 434315
rect 18814 433990 18820 434310
rect 19140 434309 32890 434310
rect 19140 433991 32571 434309
rect 32889 433991 32890 434309
rect 19140 433990 32890 433991
rect 32571 433985 32889 433990
rect 18909 433435 18915 433765
rect 19235 433760 19245 433765
rect 34054 433760 34372 433765
rect 19240 433440 19245 433760
rect 34053 433759 34373 433760
rect 34053 433441 34054 433759
rect 34372 433441 34373 433759
rect 34053 433440 34373 433441
rect 19235 433435 19245 433440
rect 34054 433435 34372 433440
rect 413052 433439 413053 435897
rect 415511 433439 484822 435897
rect 413052 433438 484822 433439
rect 413053 433433 415511 433438
rect 32571 431310 32889 431315
rect 18814 430990 18820 431310
rect 19140 431309 32890 431310
rect 19140 430991 32571 431309
rect 32889 430991 32890 431309
rect 19140 430990 32890 430991
rect 32571 430985 32889 430990
rect 18909 430435 18915 430765
rect 19235 430760 19245 430765
rect 34054 430760 34372 430765
rect 19240 430440 19245 430760
rect 34053 430759 34373 430760
rect 34053 430441 34054 430759
rect 34372 430441 34373 430759
rect 34053 430440 34373 430441
rect 19235 430435 19245 430440
rect 34054 430435 34372 430440
rect 11078 427174 14457 429929
rect 17212 427174 17218 429929
rect 32571 428310 32889 428315
rect 18814 427990 18820 428310
rect 19140 428309 32890 428310
rect 19140 427991 32571 428309
rect 32889 427991 32890 428309
rect 19140 427990 32890 427991
rect 32571 427985 32889 427990
rect 18909 427435 18915 427765
rect 19235 427760 19245 427765
rect 34054 427760 34372 427765
rect 19240 427440 19245 427760
rect 34053 427759 34373 427760
rect 34053 427441 34054 427759
rect 34372 427441 34373 427759
rect 34053 427440 34373 427441
rect 19235 427435 19245 427440
rect 34054 427435 34372 427440
rect 11078 340671 13833 427174
rect 24171 425310 24291 426309
rect 32571 425310 32889 425315
rect 18814 424990 18820 425310
rect 19140 425309 32890 425310
rect 19140 424991 32571 425309
rect 32889 424991 32890 425309
rect 19140 424990 32890 424991
rect 18909 424435 18915 424765
rect 19235 424760 19245 424765
rect 19240 424440 19245 424760
rect 19235 424435 19245 424440
rect 24171 422310 24291 424990
rect 32571 424985 32889 424990
rect 34054 424760 34372 424765
rect 34053 424759 34373 424760
rect 34053 424441 34054 424759
rect 34372 424441 34373 424759
rect 34053 424440 34373 424441
rect 34054 424435 34372 424440
rect 32571 422310 32889 422315
rect 18814 421990 18820 422310
rect 19140 422309 32890 422310
rect 19140 421991 32571 422309
rect 32889 421991 32890 422309
rect 19140 421990 32890 421991
rect 18909 421435 18915 421765
rect 19235 421760 19245 421765
rect 19240 421440 19245 421760
rect 19235 421435 19245 421440
rect 24171 420470 24291 421990
rect 32571 421985 32889 421990
rect 34054 421760 34372 421765
rect 34053 421759 34373 421760
rect 34053 421441 34054 421759
rect 34372 421441 34373 421759
rect 34053 421440 34373 421441
rect 34054 421435 34372 421440
rect 24171 419310 24291 420358
rect 32571 419310 32889 419315
rect 18814 418990 18820 419310
rect 19140 419309 32890 419310
rect 19140 418991 32571 419309
rect 32889 418991 32890 419309
rect 404802 419114 404808 421584
rect 407268 421579 407278 421584
rect 428430 421579 430888 421584
rect 407273 419119 407278 421579
rect 428429 421578 430889 421579
rect 428429 419120 428430 421578
rect 430888 419120 430889 421578
rect 428429 419119 430889 419120
rect 407268 419114 407278 419119
rect 428430 419114 430888 419119
rect 19140 418990 32890 418991
rect 18909 418435 18915 418765
rect 19235 418760 19245 418765
rect 19240 418440 19245 418760
rect 19235 418435 19245 418440
rect 24171 416310 24291 418990
rect 32571 418985 32889 418990
rect 34054 418760 34372 418765
rect 34053 418759 34373 418760
rect 34053 418441 34054 418759
rect 34372 418441 34373 418759
rect 34053 418440 34373 418441
rect 34054 418435 34372 418440
rect 32571 416310 32889 416315
rect 18814 415990 18820 416310
rect 19140 416309 32890 416310
rect 19140 415991 32571 416309
rect 32889 415991 32890 416309
rect 19140 415990 32890 415991
rect 18909 415435 18915 415765
rect 19235 415760 19245 415765
rect 19240 415440 19245 415760
rect 19235 415435 19245 415440
rect 24171 413310 24291 415990
rect 32571 415985 32889 415990
rect 34054 415760 34372 415765
rect 34053 415759 34373 415760
rect 34053 415441 34054 415759
rect 34372 415441 34373 415759
rect 34053 415440 34373 415441
rect 34054 415435 34372 415440
rect 32571 413310 32889 413315
rect 18814 412990 18820 413310
rect 19140 413309 32890 413310
rect 19140 412991 32571 413309
rect 32889 412991 32890 413309
rect 19140 412990 32890 412991
rect 18909 412435 18915 412765
rect 19235 412760 19245 412765
rect 19240 412440 19245 412760
rect 19235 412435 19245 412440
rect 24171 410310 24291 412990
rect 32571 412985 32889 412990
rect 34054 412760 34372 412765
rect 34053 412759 34373 412760
rect 34053 412441 34054 412759
rect 34372 412441 34373 412759
rect 34053 412440 34373 412441
rect 34054 412435 34372 412440
rect 32571 410310 32889 410315
rect 18814 409990 18820 410310
rect 19140 410309 32890 410310
rect 19140 409991 32571 410309
rect 32889 409991 32890 410309
rect 19140 409990 32890 409991
rect 18909 409435 18915 409765
rect 19235 409760 19245 409765
rect 19240 409440 19245 409760
rect 19235 409435 19245 409440
rect 24171 407310 24291 409990
rect 32571 409985 32889 409990
rect 34054 409760 34372 409765
rect 34053 409759 34373 409760
rect 34053 409441 34054 409759
rect 34372 409441 34373 409759
rect 34053 409440 34373 409441
rect 34054 409435 34372 409440
rect 32571 407310 32889 407315
rect 18814 406990 18820 407310
rect 19140 407309 32890 407310
rect 19140 406991 32571 407309
rect 32889 406991 32890 407309
rect 404568 407226 404574 409696
rect 407034 409691 407044 409696
rect 428430 409691 430888 409696
rect 407039 407231 407044 409691
rect 428429 409690 430889 409691
rect 428429 407232 428430 409690
rect 430888 407232 430889 409690
rect 428429 407231 430889 407232
rect 407034 407226 407044 407231
rect 428430 407226 430888 407231
rect 19140 406990 32890 406991
rect 18909 406435 18915 406765
rect 19235 406760 19245 406765
rect 19240 406440 19245 406760
rect 19235 406435 19245 406440
rect 24171 404310 24291 406990
rect 32571 406985 32889 406990
rect 34054 406760 34372 406765
rect 34053 406759 34373 406760
rect 34053 406441 34054 406759
rect 34372 406441 34373 406759
rect 34053 406440 34373 406441
rect 34054 406435 34372 406440
rect 32571 404310 32889 404315
rect 18814 403990 18820 404310
rect 19140 404309 32890 404310
rect 19140 403991 32571 404309
rect 32889 403991 32890 404309
rect 19140 403990 32890 403991
rect 18909 403435 18915 403765
rect 19235 403760 19245 403765
rect 19240 403440 19245 403760
rect 19235 403435 19245 403440
rect 24171 401310 24291 403990
rect 32571 403985 32889 403990
rect 34054 403760 34372 403765
rect 34053 403759 34373 403760
rect 34053 403441 34054 403759
rect 34372 403441 34373 403759
rect 34053 403440 34373 403441
rect 34054 403435 34372 403440
rect 32571 401310 32889 401315
rect 18814 400990 18820 401310
rect 19140 401309 32890 401310
rect 19140 400991 32571 401309
rect 32889 400991 32890 401309
rect 19140 400990 32890 400991
rect 24171 398310 24291 400990
rect 32571 400985 32889 400990
rect 413053 399795 415511 399800
rect 480022 399795 484822 433438
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect 413052 399794 484822 399795
rect 32571 398310 32889 398315
rect 18814 397990 18820 398310
rect 19140 398309 32890 398310
rect 19140 397991 32571 398309
rect 32889 397991 32890 398309
rect 19140 397990 32890 397991
rect 18909 397435 18915 397765
rect 19235 397760 19245 397765
rect 19240 397440 19245 397760
rect 19235 397435 19245 397440
rect 24171 395310 24291 397990
rect 32571 397985 32889 397990
rect 34054 397760 34372 397765
rect 34053 397759 34373 397760
rect 34053 397441 34054 397759
rect 34372 397441 34373 397759
rect 34053 397440 34373 397441
rect 34054 397435 34372 397440
rect 413052 397336 413053 399794
rect 415511 397336 484822 399794
rect 413052 397335 484822 397336
rect 413053 397330 415511 397335
rect 32571 395310 32889 395315
rect 18814 394990 18820 395310
rect 19140 395309 32890 395310
rect 19140 394991 32571 395309
rect 32889 394991 32890 395309
rect 19140 394990 32890 394991
rect 18909 394435 18915 394765
rect 19235 394760 19245 394765
rect 19240 394440 19245 394760
rect 19235 394435 19245 394440
rect 24171 392310 24291 394990
rect 32571 394985 32889 394990
rect 34054 394760 34372 394765
rect 34053 394759 34373 394760
rect 34053 394441 34054 394759
rect 34372 394441 34373 394759
rect 34053 394440 34373 394441
rect 34054 394435 34372 394440
rect 32571 392310 32889 392315
rect 18814 391990 18820 392310
rect 19140 392309 32890 392310
rect 19140 391991 32571 392309
rect 32889 391991 32890 392309
rect 19140 391990 32890 391991
rect 18909 391435 18915 391765
rect 19235 391760 19245 391765
rect 19240 391440 19245 391760
rect 19235 391435 19245 391440
rect 24171 389310 24291 391990
rect 32571 391985 32889 391990
rect 34054 391760 34372 391765
rect 34053 391759 34373 391760
rect 34053 391441 34054 391759
rect 34372 391441 34373 391759
rect 34053 391440 34373 391441
rect 34054 391435 34372 391440
rect 32571 389310 32889 389315
rect 18814 388990 18820 389310
rect 19140 389309 32890 389310
rect 19140 388991 32571 389309
rect 32889 388991 32890 389309
rect 19140 388990 32890 388991
rect 18909 388435 18915 388765
rect 19235 388760 19245 388765
rect 19240 388440 19245 388760
rect 19235 388435 19245 388440
rect 24171 386310 24291 388990
rect 32571 388985 32889 388990
rect 34054 388760 34372 388765
rect 34053 388759 34373 388760
rect 34053 388441 34054 388759
rect 34372 388441 34373 388759
rect 34053 388440 34373 388441
rect 34054 388435 34372 388440
rect 32571 386310 32889 386315
rect 18814 385990 18820 386310
rect 19140 386309 32890 386310
rect 19140 385991 32571 386309
rect 32889 385991 32890 386309
rect 19140 385990 32890 385991
rect 18909 385435 18915 385765
rect 19235 385760 19245 385765
rect 19240 385440 19245 385760
rect 19235 385435 19245 385440
rect 24171 383310 24291 385990
rect 32571 385985 32889 385990
rect 413053 385768 415511 385773
rect 480022 385768 484822 397335
rect 413052 385767 484822 385768
rect 34054 385760 34372 385765
rect 34053 385759 34373 385760
rect 34053 385441 34054 385759
rect 34372 385441 34373 385759
rect 34053 385440 34373 385441
rect 34054 385435 34372 385440
rect 32571 383310 32889 383315
rect 18814 382990 18820 383310
rect 19140 383309 32890 383310
rect 19140 382991 32571 383309
rect 32889 382991 32890 383309
rect 413052 383309 413053 385767
rect 415511 383309 484822 385767
rect 413052 383308 484822 383309
rect 413053 383303 415511 383308
rect 19140 382990 32890 382991
rect 18909 382435 18915 382765
rect 19235 382760 19245 382765
rect 19240 382440 19245 382760
rect 19235 382435 19245 382440
rect 24171 380310 24291 382990
rect 32571 382985 32889 382990
rect 34054 382760 34372 382765
rect 34053 382759 34373 382760
rect 34053 382441 34054 382759
rect 34372 382441 34373 382759
rect 34053 382440 34373 382441
rect 34054 382435 34372 382440
rect 32571 380310 32889 380315
rect 18814 379990 18820 380310
rect 19140 380309 32890 380310
rect 19140 379991 32571 380309
rect 32889 379991 32890 380309
rect 19140 379990 32890 379991
rect 18909 379435 18915 379765
rect 19235 379760 19245 379765
rect 19240 379440 19245 379760
rect 19235 379435 19245 379440
rect 24171 377310 24291 379990
rect 32571 379985 32889 379990
rect 34054 379760 34372 379765
rect 34053 379759 34373 379760
rect 34053 379441 34054 379759
rect 34372 379441 34373 379759
rect 34053 379440 34373 379441
rect 34054 379435 34372 379440
rect 414093 377762 414103 377767
rect 414093 377472 414098 377762
rect 414093 377467 414103 377472
rect 414393 377467 414399 377767
rect 32571 377310 32889 377315
rect 18814 377248 18820 377310
rect 17740 377136 18820 377248
rect 18814 376990 18820 377136
rect 19140 377309 32890 377310
rect 19140 376991 32571 377309
rect 32889 376991 32890 377309
rect 19140 376990 32890 376991
rect 413985 377075 413995 377080
rect 18909 376435 18915 376765
rect 19235 376760 19245 376765
rect 19240 376440 19245 376760
rect 19235 376435 19245 376440
rect 22911 374310 23023 376990
rect 24171 374310 24291 376990
rect 32571 376985 32889 376990
rect 413985 376785 413990 377075
rect 413985 376780 413995 376785
rect 414285 376780 414291 377080
rect 34054 376760 34372 376765
rect 34053 376759 34373 376760
rect 34053 376441 34054 376759
rect 34372 376441 34373 376759
rect 34053 376440 34373 376441
rect 34054 376435 34372 376440
rect 414238 376208 414248 376213
rect 414238 375918 414243 376208
rect 414238 375913 414248 375918
rect 414538 375913 414544 376213
rect 414021 374653 414031 374658
rect 414021 374363 414026 374653
rect 414021 374358 414031 374363
rect 414321 374358 414327 374658
rect 32571 374310 32889 374315
rect 18814 373990 18820 374310
rect 19140 374309 32890 374310
rect 19140 373991 32571 374309
rect 32889 373991 32890 374309
rect 19140 373990 32890 373991
rect 413989 374054 413999 374059
rect 18909 373435 18915 373765
rect 19235 373760 19245 373765
rect 19240 373440 19245 373760
rect 19235 373435 19245 373440
rect 22911 371310 23023 373990
rect 24171 371310 24291 373990
rect 32571 373985 32889 373990
rect 34054 373760 34372 373765
rect 413989 373764 413994 374054
rect 34053 373759 34373 373760
rect 413989 373759 413999 373764
rect 414289 373759 414295 374059
rect 34053 373441 34054 373759
rect 34372 373441 34373 373759
rect 34053 373440 34373 373441
rect 34054 373435 34372 373440
rect 414347 373194 414357 373199
rect 414347 372904 414352 373194
rect 414347 372899 414357 372904
rect 414647 372899 414653 373199
rect 414240 372477 414250 372482
rect 414240 372187 414245 372477
rect 414240 372182 414250 372187
rect 414540 372182 414546 372482
rect 480022 372310 484822 383308
rect 414347 371832 414357 371837
rect 414347 371542 414352 371832
rect 414347 371537 414357 371542
rect 414647 371537 414653 371837
rect 32571 371310 32889 371315
rect 18814 370990 18820 371310
rect 19140 371309 32890 371310
rect 19140 370991 32571 371309
rect 32889 370991 32890 371309
rect 414771 371295 414781 371300
rect 414771 371005 414776 371295
rect 414771 371000 414781 371005
rect 415071 371000 415077 371300
rect 19140 370990 32890 370991
rect 18909 370435 18915 370765
rect 19235 370760 19245 370765
rect 19240 370440 19245 370760
rect 19235 370435 19245 370440
rect 22911 368310 23023 370990
rect 24171 368310 24291 370990
rect 32571 370985 32889 370990
rect 34054 370760 34372 370765
rect 34053 370759 34373 370760
rect 34053 370441 34054 370759
rect 34372 370441 34373 370759
rect 34053 370440 34373 370441
rect 413767 370704 413777 370709
rect 34054 370435 34372 370440
rect 413767 370414 413772 370704
rect 413767 370409 413777 370414
rect 414067 370409 414073 370709
rect 32571 368310 32889 368315
rect 18814 367990 18820 368310
rect 19140 368309 32890 368310
rect 19140 367991 32571 368309
rect 32889 367991 32890 368309
rect 19140 367990 32890 367991
rect 18909 367435 18915 367765
rect 19235 367760 19245 367765
rect 19240 367440 19245 367760
rect 19235 367435 19245 367440
rect 22911 365310 23023 367990
rect 24171 365310 24291 367990
rect 32571 367985 32889 367990
rect 34054 367760 34372 367765
rect 34053 367759 34373 367760
rect 34053 367441 34054 367759
rect 34372 367441 34373 367759
rect 34053 367440 34373 367441
rect 34054 367435 34372 367440
rect 32571 365310 32889 365315
rect 18814 364990 18820 365310
rect 19140 365309 32890 365310
rect 19140 364991 32571 365309
rect 32889 364991 32890 365309
rect 19140 364990 32890 364991
rect 18909 364435 18915 364765
rect 19235 364760 19245 364765
rect 19240 364440 19245 364760
rect 19235 364435 19245 364440
rect 22911 362310 23023 364990
rect 24171 362310 24291 364990
rect 32571 364985 32889 364990
rect 583520 364784 584800 364896
rect 34054 364760 34372 364765
rect 34053 364759 34373 364760
rect 34053 364441 34054 364759
rect 34372 364441 34373 364759
rect 53818 364727 54138 364728
rect 34053 364440 34373 364441
rect 34054 364435 34372 364440
rect 53813 364409 53819 364727
rect 54137 364409 54143 364727
rect 32571 362310 32889 362315
rect 18814 361990 18820 362310
rect 19140 362309 32890 362310
rect 19140 361991 32571 362309
rect 32889 361991 32890 362309
rect 19140 361990 32890 361991
rect 22911 360420 23023 361990
rect 24171 360420 24291 361990
rect 32571 361985 32889 361990
rect 35309 359517 35429 361429
rect 21720 359512 35429 359517
rect 21720 359402 21725 359512
rect 21835 359402 35429 359512
rect 21720 359397 35429 359402
rect 22911 358961 23023 359010
rect 22911 358859 22916 358961
rect 23018 358859 23023 358961
rect 22911 357975 23023 358859
rect 39253 357975 39373 361409
rect 22911 357863 40458 357975
rect 43333 357427 43453 361455
rect 14726 357307 43453 357427
rect 11078 337916 14606 340671
rect 14726 337916 14741 340671
rect 17496 337916 17502 340671
rect 11078 337476 13833 337916
rect 5660 336687 5665 336789
rect 5767 336687 5772 336789
rect 5660 336682 5772 336687
rect -800 336278 480 336390
rect 22555 335208 22675 357307
rect 26645 353279 26655 353284
rect 26645 350819 26650 353279
rect 26645 350814 26655 350819
rect 29115 350814 29121 353284
rect 26571 348750 26581 348755
rect 26571 346290 26576 348750
rect 26571 346285 26581 346290
rect 29041 346285 29047 348755
rect 26571 344240 26581 344245
rect 26571 341780 26576 344240
rect 26571 341775 26581 341780
rect 29041 341775 29047 344245
rect -800 335096 22675 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 22555 330961 22675 335096
rect 5655 327595 5777 327600
rect 5655 327483 5660 327595
rect 5772 327483 5777 327595
rect 5655 327478 5777 327483
rect 1920 315915 4378 315920
rect 1919 315914 4379 315915
rect 1919 313456 1920 315914
rect 4378 313456 4379 315914
rect 1919 313455 4379 313456
rect 1920 313450 4378 313455
rect -800 295420 680 295532
rect -800 294238 480 294350
rect 5660 293381 5772 327478
rect 39931 315915 39941 315920
rect 39931 313455 39936 315915
rect 39931 313450 39941 313455
rect 42401 313450 42407 315920
rect 5660 293263 5772 293269
rect -800 293056 480 293168
rect 3192 291986 3304 292104
rect -800 291874 3840 291986
rect 3694 290804 3806 291874
rect -800 290692 1908 290804
rect 3672 290692 9839 290804
rect -800 289510 480 289622
rect 9727 289082 9839 290692
rect 47277 289082 47397 361377
rect 53818 361159 54138 364409
rect 583520 363602 584800 363714
rect 492062 362420 584800 362532
rect 9482 288962 47397 289082
rect 52612 360839 54138 361159
rect 365000 362221 365170 362227
rect 9727 288921 9839 288962
rect 8362 261320 8493 261350
rect 8362 261250 8382 261320
rect 8462 261250 8493 261320
rect 8362 261245 8387 261250
rect 8457 261245 8493 261250
rect 8362 261225 8493 261245
rect 52612 254006 52932 360839
rect 365000 358899 365170 362051
rect 404514 359710 404520 362180
rect 406980 362175 406990 362180
rect 428430 362175 430888 362180
rect 406985 359715 406990 362175
rect 428429 362174 430889 362175
rect 428429 359716 428430 362174
rect 430888 359716 430889 362174
rect 428429 359715 430889 359716
rect 406980 359710 406990 359715
rect 428430 359710 430888 359715
rect 364995 358894 365175 358899
rect 361284 358660 363551 358780
rect 364995 358724 365000 358894
rect 365170 358724 365175 358894
rect 364995 358719 365175 358724
rect 363431 355489 363551 358660
rect 492062 355489 492174 362420
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583093 358874 584800 358986
rect 363431 355369 493623 355489
rect 361279 354716 444537 354836
rect 361369 350636 441316 350756
rect 361381 346692 435926 346812
rect 55307 345755 55627 345756
rect 58307 345755 58627 345756
rect 61307 345755 61627 345756
rect 64307 345755 64627 345756
rect 67307 345755 67627 345756
rect 70307 345755 70627 345756
rect 73307 345755 73627 345756
rect 76307 345755 76627 345756
rect 79307 345755 79627 345756
rect 82307 345755 82627 345756
rect 85307 345755 85627 345756
rect 88307 345755 88627 345756
rect 91307 345755 91627 345756
rect 94307 345755 94627 345756
rect 97307 345755 97627 345756
rect 100307 345755 100627 345756
rect 103307 345755 103627 345756
rect 106307 345755 106627 345756
rect 109307 345755 109627 345756
rect 112307 345755 112627 345756
rect 115307 345755 115627 345756
rect 118307 345755 118627 345756
rect 121307 345755 121627 345756
rect 124307 345755 124627 345756
rect 127307 345755 127627 345756
rect 130307 345755 130627 345756
rect 133307 345755 133627 345756
rect 136307 345755 136627 345756
rect 139307 345755 139627 345756
rect 142307 345755 142627 345756
rect 145307 345755 145627 345756
rect 148307 345755 148627 345756
rect 151307 345755 151627 345756
rect 154307 345755 154627 345756
rect 157307 345755 157627 345756
rect 160307 345755 160627 345756
rect 163307 345755 163627 345756
rect 166307 345755 166627 345756
rect 169307 345755 169627 345756
rect 172307 345755 172627 345756
rect 175307 345755 175627 345756
rect 178307 345755 178627 345756
rect 181307 345755 181627 345756
rect 184307 345755 184627 345756
rect 187307 345755 187627 345756
rect 190307 345755 190627 345756
rect 193307 345755 193627 345756
rect 196307 345755 196627 345756
rect 199307 345755 199627 345756
rect 202307 345755 202627 345756
rect 205307 345755 205627 345756
rect 208307 345755 208627 345756
rect 211307 345755 211627 345756
rect 214307 345755 214627 345756
rect 217307 345755 217627 345756
rect 220307 345755 220627 345756
rect 223307 345755 223627 345756
rect 226307 345755 226627 345756
rect 229307 345755 229627 345756
rect 232307 345755 232627 345756
rect 235307 345755 235627 345756
rect 238307 345755 238627 345756
rect 241307 345755 241627 345756
rect 244307 345755 244627 345756
rect 247307 345755 247627 345756
rect 250307 345755 250627 345756
rect 253307 345755 253627 345756
rect 256307 345755 256627 345756
rect 259307 345755 259627 345756
rect 262307 345755 262627 345756
rect 265307 345755 265627 345756
rect 268307 345755 268627 345756
rect 271307 345755 271627 345756
rect 274307 345755 274627 345756
rect 277307 345755 277627 345756
rect 280307 345755 280627 345756
rect 283307 345755 283627 345756
rect 286307 345755 286627 345756
rect 289307 345755 289627 345756
rect 292307 345755 292627 345756
rect 295307 345755 295627 345756
rect 298307 345755 298627 345756
rect 301307 345755 301627 345756
rect 304307 345755 304627 345756
rect 307307 345755 307627 345756
rect 310307 345755 310627 345756
rect 313307 345755 313627 345756
rect 316307 345755 316627 345756
rect 319307 345755 319627 345756
rect 325307 345755 325627 345756
rect 328307 345755 328627 345756
rect 331307 345755 331627 345756
rect 334307 345755 334627 345756
rect 337307 345755 337627 345756
rect 340307 345755 340627 345756
rect 343307 345755 343627 345756
rect 346307 345755 346627 345756
rect 349307 345755 349627 345756
rect 352307 345755 352627 345756
rect 355307 345755 355627 345756
rect 358307 345755 358627 345756
rect 55302 345437 55308 345755
rect 55626 345437 55632 345755
rect 58302 345437 58308 345755
rect 58626 345437 58632 345755
rect 61302 345437 61308 345755
rect 61626 345437 61632 345755
rect 64302 345437 64308 345755
rect 64626 345437 64632 345755
rect 67302 345437 67308 345755
rect 67626 345437 67632 345755
rect 70302 345437 70308 345755
rect 70626 345437 70632 345755
rect 73302 345437 73308 345755
rect 73626 345437 73632 345755
rect 76302 345437 76308 345755
rect 76626 345437 76632 345755
rect 79302 345437 79308 345755
rect 79626 345437 79632 345755
rect 82302 345437 82308 345755
rect 82626 345437 82632 345755
rect 85302 345437 85308 345755
rect 85626 345437 85632 345755
rect 88302 345437 88308 345755
rect 88626 345437 88632 345755
rect 91302 345437 91308 345755
rect 91626 345437 91632 345755
rect 94302 345437 94308 345755
rect 94626 345437 94632 345755
rect 97302 345437 97308 345755
rect 97626 345437 97632 345755
rect 100302 345437 100308 345755
rect 100626 345437 100632 345755
rect 103302 345437 103308 345755
rect 103626 345437 103632 345755
rect 106302 345437 106308 345755
rect 106626 345437 106632 345755
rect 109302 345437 109308 345755
rect 109626 345437 109632 345755
rect 112302 345437 112308 345755
rect 112626 345437 112632 345755
rect 115302 345437 115308 345755
rect 115626 345437 115632 345755
rect 118302 345437 118308 345755
rect 118626 345437 118632 345755
rect 121302 345437 121308 345755
rect 121626 345437 121632 345755
rect 124302 345437 124308 345755
rect 124626 345437 124632 345755
rect 127302 345437 127308 345755
rect 127626 345437 127632 345755
rect 130302 345437 130308 345755
rect 130626 345437 130632 345755
rect 133302 345437 133308 345755
rect 133626 345437 133632 345755
rect 136302 345437 136308 345755
rect 136626 345437 136632 345755
rect 139302 345437 139308 345755
rect 139626 345437 139632 345755
rect 142302 345437 142308 345755
rect 142626 345437 142632 345755
rect 145302 345437 145308 345755
rect 145626 345437 145632 345755
rect 148302 345437 148308 345755
rect 148626 345437 148632 345755
rect 151302 345437 151308 345755
rect 151626 345437 151632 345755
rect 154302 345437 154308 345755
rect 154626 345437 154632 345755
rect 157302 345437 157308 345755
rect 157626 345437 157632 345755
rect 160302 345437 160308 345755
rect 160626 345437 160632 345755
rect 163302 345437 163308 345755
rect 163626 345437 163632 345755
rect 166302 345437 166308 345755
rect 166626 345437 166632 345755
rect 169302 345437 169308 345755
rect 169626 345437 169632 345755
rect 172302 345437 172308 345755
rect 172626 345437 172632 345755
rect 175302 345437 175308 345755
rect 175626 345437 175632 345755
rect 178302 345437 178308 345755
rect 178626 345437 178632 345755
rect 181302 345437 181308 345755
rect 181626 345437 181632 345755
rect 184302 345437 184308 345755
rect 184626 345437 184632 345755
rect 187302 345437 187308 345755
rect 187626 345437 187632 345755
rect 190302 345437 190308 345755
rect 190626 345437 190632 345755
rect 193302 345437 193308 345755
rect 193626 345437 193632 345755
rect 196302 345437 196308 345755
rect 196626 345437 196632 345755
rect 199302 345437 199308 345755
rect 199626 345437 199632 345755
rect 202302 345437 202308 345755
rect 202626 345437 202632 345755
rect 205302 345437 205308 345755
rect 205626 345437 205632 345755
rect 208302 345437 208308 345755
rect 208626 345437 208632 345755
rect 211302 345437 211308 345755
rect 211626 345437 211632 345755
rect 214302 345437 214308 345755
rect 214626 345437 214632 345755
rect 217302 345437 217308 345755
rect 217626 345437 217632 345755
rect 220302 345437 220308 345755
rect 220626 345437 220632 345755
rect 223302 345437 223308 345755
rect 223626 345437 223632 345755
rect 226302 345437 226308 345755
rect 226626 345437 226632 345755
rect 229302 345437 229308 345755
rect 229626 345437 229632 345755
rect 232302 345437 232308 345755
rect 232626 345437 232632 345755
rect 235302 345437 235308 345755
rect 235626 345437 235632 345755
rect 238302 345437 238308 345755
rect 238626 345437 238632 345755
rect 241302 345437 241308 345755
rect 241626 345437 241632 345755
rect 244302 345437 244308 345755
rect 244626 345437 244632 345755
rect 247302 345437 247308 345755
rect 247626 345437 247632 345755
rect 250302 345437 250308 345755
rect 250626 345437 250632 345755
rect 253302 345437 253308 345755
rect 253626 345437 253632 345755
rect 256302 345437 256308 345755
rect 256626 345437 256632 345755
rect 259302 345437 259308 345755
rect 259626 345437 259632 345755
rect 262302 345437 262308 345755
rect 262626 345437 262632 345755
rect 265302 345437 265308 345755
rect 265626 345437 265632 345755
rect 268302 345437 268308 345755
rect 268626 345437 268632 345755
rect 271302 345437 271308 345755
rect 271626 345437 271632 345755
rect 274302 345437 274308 345755
rect 274626 345437 274632 345755
rect 277302 345437 277308 345755
rect 277626 345437 277632 345755
rect 280302 345437 280308 345755
rect 280626 345437 280632 345755
rect 283302 345437 283308 345755
rect 283626 345437 283632 345755
rect 286302 345437 286308 345755
rect 286626 345437 286632 345755
rect 289302 345437 289308 345755
rect 289626 345437 289632 345755
rect 292302 345437 292308 345755
rect 292626 345437 292632 345755
rect 295302 345437 295308 345755
rect 295626 345437 295632 345755
rect 298302 345437 298308 345755
rect 298626 345437 298632 345755
rect 301302 345437 301308 345755
rect 301626 345437 301632 345755
rect 304302 345437 304308 345755
rect 304626 345437 304632 345755
rect 307302 345437 307308 345755
rect 307626 345437 307632 345755
rect 310302 345437 310308 345755
rect 310626 345437 310632 345755
rect 313302 345437 313308 345755
rect 313626 345437 313632 345755
rect 316302 345437 316308 345755
rect 316626 345437 316632 345755
rect 319302 345437 319308 345755
rect 319626 345437 319632 345755
rect 325302 345437 325308 345755
rect 325626 345437 325632 345755
rect 328302 345437 328308 345755
rect 328626 345437 328632 345755
rect 331302 345437 331308 345755
rect 331626 345437 331632 345755
rect 334302 345437 334308 345755
rect 334626 345437 334632 345755
rect 337302 345437 337308 345755
rect 337626 345437 337632 345755
rect 340302 345437 340308 345755
rect 340626 345437 340632 345755
rect 343302 345437 343308 345755
rect 343626 345437 343632 345755
rect 346302 345437 346308 345755
rect 346626 345437 346632 345755
rect 349302 345437 349308 345755
rect 349626 345437 349632 345755
rect 352302 345437 352308 345755
rect 352626 345437 352632 345755
rect 355302 345437 355308 345755
rect 355626 345437 355632 345755
rect 358302 345437 358308 345755
rect 358626 345437 358632 345755
rect 55307 345436 55627 345437
rect 58307 345436 58627 345437
rect 61307 345436 61627 345437
rect 64307 345436 64627 345437
rect 67307 345436 67627 345437
rect 70307 345436 70627 345437
rect 73307 345436 73627 345437
rect 76307 345436 76627 345437
rect 79307 345436 79627 345437
rect 82307 345436 82627 345437
rect 85307 345436 85627 345437
rect 88307 345436 88627 345437
rect 91307 345436 91627 345437
rect 94307 345436 94627 345437
rect 97307 345436 97627 345437
rect 100307 345436 100627 345437
rect 103307 345436 103627 345437
rect 106307 345436 106627 345437
rect 109307 345436 109627 345437
rect 112307 345436 112627 345437
rect 115307 345436 115627 345437
rect 118307 345436 118627 345437
rect 121307 345436 121627 345437
rect 124307 345436 124627 345437
rect 127307 345436 127627 345437
rect 130307 345436 130627 345437
rect 133307 345436 133627 345437
rect 136307 345436 136627 345437
rect 139307 345436 139627 345437
rect 142307 345436 142627 345437
rect 145307 345436 145627 345437
rect 148307 345436 148627 345437
rect 151307 345436 151627 345437
rect 154307 345436 154627 345437
rect 157307 345436 157627 345437
rect 160307 345436 160627 345437
rect 163307 345436 163627 345437
rect 166307 345436 166627 345437
rect 169307 345436 169627 345437
rect 172307 345436 172627 345437
rect 175307 345436 175627 345437
rect 178307 345436 178627 345437
rect 181307 345436 181627 345437
rect 184307 345436 184627 345437
rect 187307 345436 187627 345437
rect 190307 345436 190627 345437
rect 193307 345436 193627 345437
rect 196307 345436 196627 345437
rect 199307 345436 199627 345437
rect 202307 345436 202627 345437
rect 205307 345436 205627 345437
rect 208307 345436 208627 345437
rect 211307 345436 211627 345437
rect 214307 345436 214627 345437
rect 217307 345436 217627 345437
rect 220307 345436 220627 345437
rect 223307 345436 223627 345437
rect 226307 345436 226627 345437
rect 229307 345436 229627 345437
rect 232307 345436 232627 345437
rect 235307 345436 235627 345437
rect 238307 345436 238627 345437
rect 241307 345436 241627 345437
rect 244307 345436 244627 345437
rect 247307 345436 247627 345437
rect 250307 345436 250627 345437
rect 253307 345436 253627 345437
rect 256307 345436 256627 345437
rect 259307 345436 259627 345437
rect 262307 345436 262627 345437
rect 265307 345436 265627 345437
rect 268307 345436 268627 345437
rect 271307 345436 271627 345437
rect 274307 345436 274627 345437
rect 277307 345436 277627 345437
rect 280307 345436 280627 345437
rect 283307 345436 283627 345437
rect 286307 345436 286627 345437
rect 289307 345436 289627 345437
rect 292307 345436 292627 345437
rect 295307 345436 295627 345437
rect 298307 345436 298627 345437
rect 301307 345436 301627 345437
rect 304307 345436 304627 345437
rect 307307 345436 307627 345437
rect 310307 345436 310627 345437
rect 313307 345436 313627 345437
rect 316307 345436 316627 345437
rect 319307 345436 319627 345437
rect 325307 345436 325627 345437
rect 328307 345436 328627 345437
rect 331307 345436 331627 345437
rect 334307 345436 334627 345437
rect 337307 345436 337627 345437
rect 340307 345436 340627 345437
rect 343307 345436 343627 345437
rect 346307 345436 346627 345437
rect 349307 345436 349627 345437
rect 352307 345436 352627 345437
rect 355307 345436 355627 345437
rect 358307 345436 358627 345437
rect 372476 336904 372486 336909
rect 372476 336604 372481 336904
rect 372476 336599 372486 336604
rect 372786 336599 372792 336909
rect 375476 336904 375486 336909
rect 375476 336604 375481 336904
rect 375476 336599 375486 336604
rect 375786 336599 375792 336909
rect 378476 336904 378486 336909
rect 378476 336604 378481 336904
rect 378476 336599 378486 336604
rect 378786 336599 378792 336909
rect 381476 336904 381486 336909
rect 381476 336604 381481 336904
rect 381476 336599 381486 336604
rect 381786 336599 381792 336909
rect 384476 336904 384486 336909
rect 384476 336604 384481 336904
rect 384476 336599 384486 336604
rect 384786 336599 384792 336909
rect 387476 336904 387486 336909
rect 387476 336604 387481 336904
rect 387476 336599 387486 336604
rect 387786 336599 387792 336909
rect 390476 336904 390486 336909
rect 390476 336604 390481 336904
rect 390476 336599 390486 336604
rect 390786 336599 390792 336909
rect 393476 336904 393486 336909
rect 393476 336604 393481 336904
rect 393476 336599 393486 336604
rect 393786 336599 393792 336909
rect 396476 336904 396486 336909
rect 396476 336604 396481 336904
rect 396476 336599 396486 336604
rect 396786 336599 396792 336909
rect 55302 323427 55632 323432
rect 55302 323422 55307 323427
rect 55627 323422 55632 323427
rect 55302 323096 55632 323102
rect 58302 323427 58632 323432
rect 58302 323422 58307 323427
rect 58627 323422 58632 323427
rect 58302 323096 58632 323102
rect 61302 323427 61632 323432
rect 61302 323422 61307 323427
rect 61627 323422 61632 323427
rect 61302 323096 61632 323102
rect 64302 323427 64632 323432
rect 64302 323422 64307 323427
rect 64627 323422 64632 323427
rect 64302 323096 64632 323102
rect 67302 323427 67632 323432
rect 67302 323422 67307 323427
rect 67627 323422 67632 323427
rect 67302 323096 67632 323102
rect 70302 323427 70632 323432
rect 70302 323422 70307 323427
rect 70627 323422 70632 323427
rect 70302 323096 70632 323102
rect 73302 323427 73632 323432
rect 73302 323422 73307 323427
rect 73627 323422 73632 323427
rect 73302 323096 73632 323102
rect 76302 323427 76632 323432
rect 76302 323422 76307 323427
rect 76627 323422 76632 323427
rect 76302 323096 76632 323102
rect 79302 323427 79632 323432
rect 79302 323422 79307 323427
rect 79627 323422 79632 323427
rect 79302 323096 79632 323102
rect 82302 323427 82632 323432
rect 82302 323422 82307 323427
rect 82627 323422 82632 323427
rect 82302 323096 82632 323102
rect 85302 323427 85632 323432
rect 85302 323422 85307 323427
rect 85627 323422 85632 323427
rect 85302 323096 85632 323102
rect 88302 323427 88632 323432
rect 88302 323422 88307 323427
rect 88627 323422 88632 323427
rect 88302 323096 88632 323102
rect 91302 323427 91632 323432
rect 91302 323422 91307 323427
rect 91627 323422 91632 323427
rect 91302 323096 91632 323102
rect 94302 323427 94632 323432
rect 94302 323422 94307 323427
rect 94627 323422 94632 323427
rect 94302 323096 94632 323102
rect 97302 323427 97632 323432
rect 97302 323422 97307 323427
rect 97627 323422 97632 323427
rect 97302 323096 97632 323102
rect 100302 323427 100632 323432
rect 100302 323422 100307 323427
rect 100627 323422 100632 323427
rect 100302 323096 100632 323102
rect 103302 323427 103632 323432
rect 103302 323422 103307 323427
rect 103627 323422 103632 323427
rect 103302 323096 103632 323102
rect 106302 323427 106632 323432
rect 106302 323422 106307 323427
rect 106627 323422 106632 323427
rect 106302 323096 106632 323102
rect 109302 323427 109632 323432
rect 109302 323422 109307 323427
rect 109627 323422 109632 323427
rect 109302 323096 109632 323102
rect 112302 323427 112632 323432
rect 112302 323422 112307 323427
rect 112627 323422 112632 323427
rect 112302 323096 112632 323102
rect 115302 323427 115632 323432
rect 115302 323422 115307 323427
rect 115627 323422 115632 323427
rect 115302 323096 115632 323102
rect 118302 323427 118632 323432
rect 118302 323422 118307 323427
rect 118627 323422 118632 323427
rect 118302 323096 118632 323102
rect 121302 323427 121632 323432
rect 121302 323422 121307 323427
rect 121627 323422 121632 323427
rect 121302 323096 121632 323102
rect 124302 323427 124632 323432
rect 124302 323422 124307 323427
rect 124627 323422 124632 323427
rect 124302 323096 124632 323102
rect 127302 323427 127632 323432
rect 127302 323422 127307 323427
rect 127627 323422 127632 323427
rect 127302 323096 127632 323102
rect 130302 323427 130632 323432
rect 130302 323422 130307 323427
rect 130627 323422 130632 323427
rect 130302 323096 130632 323102
rect 133302 323427 133632 323432
rect 133302 323422 133307 323427
rect 133627 323422 133632 323427
rect 133302 323096 133632 323102
rect 136302 323427 136632 323432
rect 136302 323422 136307 323427
rect 136627 323422 136632 323427
rect 136302 323096 136632 323102
rect 139302 323427 139632 323432
rect 139302 323422 139307 323427
rect 139627 323422 139632 323427
rect 139302 323096 139632 323102
rect 142302 323427 142632 323432
rect 142302 323422 142307 323427
rect 142627 323422 142632 323427
rect 142302 323096 142632 323102
rect 145302 323427 145632 323432
rect 145302 323422 145307 323427
rect 145627 323422 145632 323427
rect 145302 323096 145632 323102
rect 148302 323427 148632 323432
rect 148302 323422 148307 323427
rect 148627 323422 148632 323427
rect 148302 323096 148632 323102
rect 151302 323427 151632 323432
rect 151302 323422 151307 323427
rect 151627 323422 151632 323427
rect 151302 323096 151632 323102
rect 154302 323427 154632 323432
rect 154302 323422 154307 323427
rect 154627 323422 154632 323427
rect 154302 323096 154632 323102
rect 157302 323427 157632 323432
rect 157302 323422 157307 323427
rect 157627 323422 157632 323427
rect 157302 323096 157632 323102
rect 160302 323427 160632 323432
rect 160302 323422 160307 323427
rect 160627 323422 160632 323427
rect 160302 323096 160632 323102
rect 163302 323427 163632 323432
rect 163302 323422 163307 323427
rect 163627 323422 163632 323427
rect 163302 323096 163632 323102
rect 166302 323427 166632 323432
rect 166302 323422 166307 323427
rect 166627 323422 166632 323427
rect 166302 323096 166632 323102
rect 169302 323427 169632 323432
rect 169302 323422 169307 323427
rect 169627 323422 169632 323427
rect 169302 323096 169632 323102
rect 172302 323427 172632 323432
rect 172302 323422 172307 323427
rect 172627 323422 172632 323427
rect 172302 323096 172632 323102
rect 175302 323427 175632 323432
rect 175302 323422 175307 323427
rect 175627 323422 175632 323427
rect 175302 323096 175632 323102
rect 178302 323427 178632 323432
rect 178302 323422 178307 323427
rect 178627 323422 178632 323427
rect 178302 323096 178632 323102
rect 181302 323427 181632 323432
rect 181302 323422 181307 323427
rect 181627 323422 181632 323427
rect 181302 323096 181632 323102
rect 184302 323427 184632 323432
rect 184302 323422 184307 323427
rect 184627 323422 184632 323427
rect 184302 323096 184632 323102
rect 187302 323427 187632 323432
rect 187302 323422 187307 323427
rect 187627 323422 187632 323427
rect 187302 323096 187632 323102
rect 190302 323427 190632 323432
rect 190302 323422 190307 323427
rect 190627 323422 190632 323427
rect 190302 323096 190632 323102
rect 193302 323427 193632 323432
rect 193302 323422 193307 323427
rect 193627 323422 193632 323427
rect 193302 323096 193632 323102
rect 196302 323427 196632 323432
rect 196302 323422 196307 323427
rect 196627 323422 196632 323427
rect 196302 323096 196632 323102
rect 199302 323427 199632 323432
rect 199302 323422 199307 323427
rect 199627 323422 199632 323427
rect 199302 323096 199632 323102
rect 202302 323427 202632 323432
rect 202302 323422 202307 323427
rect 202627 323422 202632 323427
rect 202302 323096 202632 323102
rect 205302 323427 205632 323432
rect 205302 323422 205307 323427
rect 205627 323422 205632 323427
rect 205302 323096 205632 323102
rect 208302 323427 208632 323432
rect 208302 323422 208307 323427
rect 208627 323422 208632 323427
rect 208302 323096 208632 323102
rect 211302 323427 211632 323432
rect 211302 323422 211307 323427
rect 211627 323422 211632 323427
rect 211302 323096 211632 323102
rect 214302 323427 214632 323432
rect 214302 323422 214307 323427
rect 214627 323422 214632 323427
rect 214302 323096 214632 323102
rect 217302 323427 217632 323432
rect 217302 323422 217307 323427
rect 217627 323422 217632 323427
rect 217302 323096 217632 323102
rect 220302 323427 220632 323432
rect 220302 323422 220307 323427
rect 220627 323422 220632 323427
rect 220302 323096 220632 323102
rect 223302 323427 223632 323432
rect 223302 323422 223307 323427
rect 223627 323422 223632 323427
rect 223302 323096 223632 323102
rect 226302 323427 226632 323432
rect 226302 323422 226307 323427
rect 226627 323422 226632 323427
rect 226302 323096 226632 323102
rect 229302 323427 229632 323432
rect 229302 323422 229307 323427
rect 229627 323422 229632 323427
rect 229302 323096 229632 323102
rect 232302 323427 232632 323432
rect 232302 323422 232307 323427
rect 232627 323422 232632 323427
rect 232302 323096 232632 323102
rect 235302 323427 235632 323432
rect 235302 323422 235307 323427
rect 235627 323422 235632 323427
rect 235302 323096 235632 323102
rect 238302 323427 238632 323432
rect 238302 323422 238307 323427
rect 238627 323422 238632 323427
rect 238302 323096 238632 323102
rect 241302 323427 241632 323432
rect 241302 323422 241307 323427
rect 241627 323422 241632 323427
rect 241302 323096 241632 323102
rect 244302 323427 244632 323432
rect 244302 323422 244307 323427
rect 244627 323422 244632 323427
rect 244302 323096 244632 323102
rect 247302 323427 247632 323432
rect 247302 323422 247307 323427
rect 247627 323422 247632 323427
rect 247302 323096 247632 323102
rect 250302 323427 250632 323432
rect 250302 323422 250307 323427
rect 250627 323422 250632 323427
rect 250302 323096 250632 323102
rect 253302 323427 253632 323432
rect 253302 323422 253307 323427
rect 253627 323422 253632 323427
rect 253302 323096 253632 323102
rect 256302 323427 256632 323432
rect 256302 323422 256307 323427
rect 256627 323422 256632 323427
rect 256302 323096 256632 323102
rect 259302 323427 259632 323432
rect 259302 323422 259307 323427
rect 259627 323422 259632 323427
rect 259302 323096 259632 323102
rect 262302 323427 262632 323432
rect 262302 323422 262307 323427
rect 262627 323422 262632 323427
rect 262302 323096 262632 323102
rect 265302 323427 265632 323432
rect 265302 323422 265307 323427
rect 265627 323422 265632 323427
rect 265302 323096 265632 323102
rect 268302 323427 268632 323432
rect 268302 323422 268307 323427
rect 268627 323422 268632 323427
rect 268302 323096 268632 323102
rect 271302 323427 271632 323432
rect 271302 323422 271307 323427
rect 271627 323422 271632 323427
rect 271302 323096 271632 323102
rect 274302 323427 274632 323432
rect 274302 323422 274307 323427
rect 274627 323422 274632 323427
rect 274302 323096 274632 323102
rect 277302 323427 277632 323432
rect 277302 323422 277307 323427
rect 277627 323422 277632 323427
rect 277302 323096 277632 323102
rect 280302 323427 280632 323432
rect 280302 323422 280307 323427
rect 280627 323422 280632 323427
rect 280302 323096 280632 323102
rect 283302 323427 283632 323432
rect 283302 323422 283307 323427
rect 283627 323422 283632 323427
rect 283302 323096 283632 323102
rect 286302 323427 286632 323432
rect 286302 323422 286307 323427
rect 286627 323422 286632 323427
rect 286302 323096 286632 323102
rect 289302 323427 289632 323432
rect 289302 323422 289307 323427
rect 289627 323422 289632 323427
rect 289302 323096 289632 323102
rect 292302 323427 292632 323432
rect 292302 323422 292307 323427
rect 292627 323422 292632 323427
rect 292302 323096 292632 323102
rect 295302 323427 295632 323432
rect 295302 323422 295307 323427
rect 295627 323422 295632 323427
rect 295302 323096 295632 323102
rect 298302 323427 298632 323432
rect 298302 323422 298307 323427
rect 298627 323422 298632 323427
rect 298302 323096 298632 323102
rect 301302 323427 301632 323432
rect 301302 323422 301307 323427
rect 301627 323422 301632 323427
rect 301302 323096 301632 323102
rect 304302 323427 304632 323432
rect 304302 323422 304307 323427
rect 304627 323422 304632 323427
rect 304302 323096 304632 323102
rect 307302 323427 307632 323432
rect 307302 323422 307307 323427
rect 307627 323422 307632 323427
rect 307302 323096 307632 323102
rect 310302 323427 310632 323432
rect 310302 323422 310307 323427
rect 310627 323422 310632 323427
rect 310302 323096 310632 323102
rect 313302 323427 313632 323432
rect 313302 323422 313307 323427
rect 313627 323422 313632 323427
rect 313302 323096 313632 323102
rect 316302 323427 316632 323432
rect 316302 323422 316307 323427
rect 316627 323422 316632 323427
rect 316302 323096 316632 323102
rect 319302 323427 319632 323432
rect 319302 323422 319307 323427
rect 319627 323422 319632 323427
rect 319302 323096 319632 323102
rect 325302 323427 325632 323432
rect 325302 323422 325307 323427
rect 325627 323422 325632 323427
rect 325302 323096 325632 323102
rect 328302 323427 328632 323432
rect 328302 323422 328307 323427
rect 328627 323422 328632 323427
rect 328302 323096 328632 323102
rect 331302 323427 331632 323432
rect 331302 323422 331307 323427
rect 331627 323422 331632 323427
rect 331302 323096 331632 323102
rect 334302 323427 334632 323432
rect 334302 323422 334307 323427
rect 334627 323422 334632 323427
rect 334302 323096 334632 323102
rect 337302 323427 337632 323432
rect 337302 323422 337307 323427
rect 337627 323422 337632 323427
rect 337302 323096 337632 323102
rect 340302 323427 340632 323432
rect 340302 323422 340307 323427
rect 340627 323422 340632 323427
rect 340302 323096 340632 323102
rect 343302 323427 343632 323432
rect 343302 323422 343307 323427
rect 343627 323422 343632 323427
rect 343302 323096 343632 323102
rect 346302 323427 346632 323432
rect 346302 323422 346307 323427
rect 346627 323422 346632 323427
rect 346302 323096 346632 323102
rect 349302 323427 349632 323432
rect 349302 323422 349307 323427
rect 349627 323422 349632 323427
rect 349302 323096 349632 323102
rect 352302 323427 352632 323432
rect 352302 323422 352307 323427
rect 352627 323422 352632 323427
rect 352302 323096 352632 323102
rect 355302 323427 355632 323432
rect 355302 323422 355307 323427
rect 355627 323422 355632 323427
rect 355302 323096 355632 323102
rect 358302 323427 358632 323432
rect 358302 323422 358307 323427
rect 358627 323422 358632 323427
rect 358302 323096 358632 323102
rect 435806 318609 435926 346692
rect 441196 337264 441316 350636
rect 444417 344507 444537 354716
rect 492062 354703 492174 355369
rect 444417 344387 570754 344507
rect 441196 337144 454512 337264
rect 435806 318489 448006 318609
rect 424844 314081 425014 314087
rect 175764 313911 424844 314081
rect 69648 254006 69968 254012
rect 52612 253686 69648 254006
rect 69648 253680 69968 253686
rect 5661 253173 5771 253178
rect 12507 253173 12619 253179
rect 5660 253172 12507 253173
rect 5660 253062 5661 253172
rect 5771 253062 12507 253172
rect 5660 253061 12507 253062
rect 12619 253061 12882 253173
rect 5661 253056 5771 253061
rect 12507 253055 12619 253061
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248959 56028 248964
rect -800 248857 55921 248959
rect 56023 248857 56028 248959
rect -800 248852 56028 248857
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 7127 243720 7217 243726
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 7127 200580 7217 243630
rect 173402 207498 173722 207504
rect 170812 207380 171132 207386
rect 167888 207156 168208 207162
rect 7127 200490 164551 200580
rect 164461 192747 164551 200490
rect 167888 192186 168208 206836
rect 170812 192186 171132 207060
rect 173402 192186 173722 207178
rect 167883 191868 167889 192186
rect 168207 191868 168213 192186
rect 170807 191868 170813 192186
rect 171131 191868 171137 192186
rect 173397 191868 173403 192186
rect 173721 191868 173727 192186
rect 167888 191867 168208 191868
rect 170812 191867 171132 191868
rect 173402 191867 173722 191868
rect 10674 191537 10784 191543
rect 33445 191537 33553 191542
rect 10784 191536 33554 191537
rect 10784 191428 33445 191536
rect 33553 191428 33554 191536
rect 10784 191427 33554 191428
rect 10674 191421 10784 191427
rect 33445 191422 33553 191427
rect 9011 191342 9131 191348
rect 9011 191227 9016 191232
rect 9126 191227 9131 191232
rect 9011 191222 9131 191227
rect 175764 188343 175934 313911
rect 424844 313905 425014 313911
rect 287964 230749 290424 230750
rect 287959 228291 287965 230749
rect 290423 228291 290429 230749
rect 287964 228290 290424 228291
rect 180916 207295 181216 207301
rect 180916 207000 180921 207005
rect 181211 207000 181216 207005
rect 180916 206995 181216 207000
rect 183916 207295 184216 207301
rect 183916 207000 183921 207005
rect 184211 207000 184216 207005
rect 183916 206995 184216 207000
rect 186916 207295 187216 207301
rect 186916 207000 186921 207005
rect 187211 207000 187216 207005
rect 186916 206995 187216 207000
rect 189916 207295 190216 207301
rect 189916 207000 189921 207005
rect 190211 207000 190216 207005
rect 189916 206995 190216 207000
rect 192916 207295 193216 207301
rect 192916 207000 192921 207005
rect 193211 207000 193216 207005
rect 192916 206995 193216 207000
rect 195916 207295 196216 207301
rect 195916 207000 195921 207005
rect 196211 207000 196216 207005
rect 195916 206995 196216 207000
rect 198916 207295 199216 207301
rect 198916 207000 198921 207005
rect 199211 207000 199216 207005
rect 198916 206995 199216 207000
rect 201916 207295 202216 207301
rect 201916 207000 201921 207005
rect 202211 207000 202216 207005
rect 201916 206995 202216 207000
rect 204916 207295 205216 207301
rect 204916 207000 204921 207005
rect 205211 207000 205216 207005
rect 204916 206995 205216 207000
rect 175764 188183 175769 188343
rect 175929 188183 175934 188343
rect 175764 188157 175934 188183
rect 175764 186642 175934 186815
rect 175759 186637 175939 186642
rect 175759 186632 175764 186637
rect 175934 186632 175939 186637
rect 175759 186456 175939 186462
rect 175764 180637 175934 186456
rect 177601 180637 177781 180642
rect 164431 180626 164751 180627
rect 167772 180626 168092 180627
rect 170722 180626 171042 180627
rect 173032 180626 173352 180627
rect 175008 180626 175328 180627
rect 164426 180308 164432 180626
rect 164750 180308 164756 180626
rect 167767 180308 167773 180626
rect 168091 180308 168097 180626
rect 170717 180308 170723 180626
rect 171041 180308 171047 180626
rect 173027 180308 173033 180626
rect 173351 180308 173357 180626
rect 175003 180308 175009 180626
rect 175327 180308 175333 180626
rect 175764 180467 177606 180637
rect 177776 180467 177781 180637
rect 177601 180462 177781 180467
rect 2175 177688 13873 177800
rect -800 176552 13873 177688
rect -800 172888 3527 176552
rect 2175 167688 3527 172888
rect -800 164594 3527 167688
rect 12521 169096 13873 176552
rect 15357 172530 15577 172536
rect 52330 172530 52548 172535
rect 14888 172310 15357 172530
rect 15577 172529 52549 172530
rect 15577 172311 52330 172529
rect 52548 172311 52549 172529
rect 15577 172310 52549 172311
rect 15357 172304 15577 172310
rect 52330 172305 52548 172310
rect 12521 166636 86589 169096
rect 89049 166636 89055 169096
rect 164431 168316 164751 180308
rect 164431 167990 164751 167996
rect 167772 168174 168092 180308
rect 170722 168529 171042 180308
rect 170722 168203 171042 168209
rect 173032 168245 173352 180308
rect 175008 168245 175328 180308
rect 180872 172819 181182 172824
rect 180872 172814 180877 172819
rect 181177 172814 181182 172819
rect 180872 172508 181182 172514
rect 183872 172819 184182 172824
rect 183872 172814 183877 172819
rect 184177 172814 184182 172819
rect 183872 172508 184182 172514
rect 186872 172819 187182 172824
rect 186872 172814 186877 172819
rect 187177 172814 187182 172819
rect 186872 172508 187182 172514
rect 189872 172819 190182 172824
rect 189872 172814 189877 172819
rect 190177 172814 190182 172819
rect 189872 172508 190182 172514
rect 192872 172819 193182 172824
rect 192872 172814 192877 172819
rect 193177 172814 193182 172819
rect 192872 172508 193182 172514
rect 195872 172819 196182 172824
rect 195872 172814 195877 172819
rect 196177 172814 196182 172819
rect 195872 172508 196182 172514
rect 198872 172819 199182 172824
rect 198872 172814 198877 172819
rect 199177 172814 199182 172819
rect 198872 172508 199182 172514
rect 201872 172819 202182 172824
rect 201872 172814 201877 172819
rect 202177 172814 202182 172819
rect 201872 172508 202182 172514
rect 204872 172819 205182 172824
rect 204872 172814 204877 172819
rect 205177 172814 205182 172819
rect 204872 172508 205182 172514
rect 175002 167925 175008 168245
rect 175328 167925 175334 168245
rect 173032 167919 173352 167925
rect 167772 167848 168092 167854
rect 12521 165348 13906 166636
rect 12521 164594 86444 165348
rect -800 162888 86444 164594
rect 88904 162888 88910 165348
rect 13381 154454 15841 162888
rect 13381 151994 86722 154454
rect 89182 151994 89188 154454
rect 13381 147234 15841 151994
rect 13381 144768 15841 144774
rect 13382 136509 15840 136514
rect 13381 136508 86722 136509
rect 13381 134050 13382 136508
rect 15840 134050 86722 136508
rect 13381 134049 86722 134050
rect 89182 134049 89188 136509
rect 13382 134044 15840 134049
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121337 21950 121342
rect -800 121235 21843 121337
rect 21945 121235 21950 121337
rect -800 121230 21950 121235
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 287959 118958 290429 118963
rect 287959 118953 287964 118958
rect 290424 118953 290429 118958
rect 287959 116487 290429 116493
rect 447886 112941 448006 318489
rect 454392 276364 454512 337144
rect 570634 317310 570754 344387
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 570463 317198 584800 317310
rect 570634 316193 570754 317198
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 512453 313652 514829 313764
rect 581256 313652 584800 313764
rect 454392 276244 580683 276364
rect 580563 272888 580683 276244
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 580563 272776 584800 272888
rect 580563 272105 580683 272776
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 512653 269230 514786 269342
rect 582310 269230 584800 269342
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect 573839 217336 573845 222136
rect 578645 217336 578651 222136
rect 573845 204057 578645 217336
rect 573845 199257 574269 204057
rect 579069 199257 579075 204057
rect 573845 196230 579069 199257
rect 502074 193770 502080 196230
rect 504540 193890 584800 196230
rect 502096 191430 502102 193770
rect 504562 191430 584800 193890
rect 573845 186230 578645 191430
rect 502385 183770 502391 186230
rect 504851 183890 584800 186230
rect 502549 181430 502555 183770
rect 505015 181430 584800 183890
rect 573845 167476 578645 181430
rect 573839 162676 573845 167476
rect 578645 162676 578651 167476
rect 582340 149347 584800 151630
rect 501815 146887 501821 149347
rect 504281 146887 513281 149347
rect 576060 146887 584800 149347
rect 582340 146830 584800 146887
rect 582340 139290 584800 141630
rect 502038 136830 502044 139290
rect 504504 136830 513281 139290
rect 576060 136830 584800 139290
rect 447886 112821 571679 112941
rect 571559 92866 571679 112821
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 570398 92754 584800 92866
rect 571559 89505 571679 92754
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect 33622 78124 33722 78129
rect 32898 78120 33627 78124
rect -800 78034 33627 78120
rect 33717 78034 33722 78124
rect -800 78029 33722 78034
rect -800 78008 33701 78029
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 40357 34898
rect 40469 34786 40475 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 46643 13476
rect 46755 13364 46761 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 1849 8748
rect 583520 8636 584800 8748
rect -800 7454 789 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 354 4020
rect 466 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 22111 692011 22219 692119
rect 7013 688089 7331 688093
rect 7013 687779 7017 688089
rect 7017 687779 7327 688089
rect 7327 687779 7331 688089
rect 7013 687775 7331 687779
rect 1920 686005 4378 686009
rect 1920 683555 1924 686005
rect 1924 683555 4374 686005
rect 4374 683555 4378 686005
rect 1920 683551 4378 683555
rect 28682 685548 28750 685552
rect 28682 685488 28686 685548
rect 28686 685488 28746 685548
rect 28746 685488 28750 685548
rect 28682 685484 28750 685488
rect 26807 684464 29267 684469
rect 26807 682004 29262 684464
rect 29262 682004 29267 684464
rect 26807 681999 29267 682004
rect 9017 680857 9125 680861
rect 9017 680757 9021 680857
rect 9021 680757 9121 680857
rect 9121 680757 9125 680857
rect 9017 680753 9125 680757
rect 1920 678110 4378 678114
rect 1920 675660 1924 678110
rect 1924 675660 4374 678110
rect 4374 675660 4378 678110
rect 1920 675656 4378 675660
rect 1920 672888 4378 672892
rect 1920 670438 1924 672888
rect 1924 670438 4374 672888
rect 4374 670438 4378 672888
rect 1920 670434 4378 670438
rect 26515 678115 28975 678120
rect 26515 675655 28970 678115
rect 28970 675655 28975 678115
rect 26515 675650 28975 675655
rect 10675 675031 10783 675139
rect 50826 674488 50936 674598
rect 143668 694385 144068 694390
rect 143668 694000 143673 694385
rect 143673 694000 144063 694385
rect 144063 694000 144068 694385
rect 228439 697491 229477 698529
rect 331192 697349 332128 698285
rect 126037 674486 126145 674594
rect 155830 674103 156210 674108
rect 155830 673738 155835 674103
rect 155835 673738 156205 674103
rect 156205 673738 156210 674103
rect 140627 673664 140632 673729
rect 140632 673664 140702 673729
rect 140702 673664 140707 673729
rect 140627 673659 140707 673664
rect 231034 673684 231352 673996
rect 231034 673678 231038 673684
rect 231038 673678 231348 673684
rect 231348 673678 231352 673684
rect 26348 672893 28808 672898
rect 26348 670433 28803 672893
rect 28803 670433 28808 672893
rect 26348 670428 28808 670433
rect 403010 672740 405470 675200
rect 140633 671130 140701 671134
rect 140633 671070 140637 671130
rect 140637 671070 140697 671130
rect 140697 671070 140701 671130
rect 140633 671066 140701 671070
rect 143668 670346 143673 670731
rect 143673 670346 144063 670731
rect 144063 670346 144068 670731
rect 143668 670341 144068 670346
rect 402810 668426 405270 670886
rect 501550 668426 504010 670886
rect 18915 667760 19235 667765
rect 18915 667440 18920 667760
rect 18920 667440 19235 667760
rect 34054 667755 34372 667759
rect 34054 667445 34058 667755
rect 34058 667445 34368 667755
rect 34368 667445 34372 667755
rect 34054 667441 34372 667445
rect 18915 667435 19235 667440
rect 18915 664760 19235 664765
rect 18915 664440 18920 664760
rect 18920 664440 19235 664760
rect 34054 664755 34372 664759
rect 34054 664445 34058 664755
rect 34058 664445 34368 664755
rect 34368 664445 34372 664755
rect 34054 664441 34372 664445
rect 18915 664435 19235 664440
rect 53664 664723 53982 664727
rect 53664 664413 53668 664723
rect 53668 664413 53978 664723
rect 53978 664413 53982 664723
rect 53664 664409 53982 664413
rect 18820 661990 19140 662310
rect 32571 661991 32889 662309
rect 18915 661760 19235 661765
rect 18915 661440 18920 661760
rect 18920 661440 19235 661760
rect 34054 661755 34372 661759
rect 34054 661445 34058 661755
rect 34058 661445 34368 661755
rect 34368 661445 34372 661755
rect 34054 661441 34372 661445
rect 18915 661435 19235 661440
rect 18820 658990 19140 659310
rect 32571 658991 32889 659309
rect 18915 658760 19235 658765
rect 18915 658440 18920 658760
rect 18920 658440 19235 658760
rect 34054 658755 34372 658759
rect 34054 658445 34058 658755
rect 34058 658445 34368 658755
rect 34368 658445 34372 658755
rect 34054 658441 34372 658445
rect 18915 658435 19235 658440
rect 13652 657326 13972 657331
rect 13652 657006 13967 657326
rect 13967 657006 13972 657326
rect 13652 657001 13972 657006
rect 18820 655990 19140 656310
rect 32571 655991 32889 656309
rect 18915 655760 19235 655765
rect 18915 655440 18920 655760
rect 18920 655440 19235 655760
rect 34054 655755 34372 655759
rect 34054 655445 34058 655755
rect 34058 655445 34368 655755
rect 34368 655445 34372 655755
rect 34054 655441 34372 655445
rect 18915 655435 19235 655440
rect 18820 652990 19140 653310
rect 32571 652991 32889 653309
rect 18915 652760 19235 652765
rect 18915 652440 18920 652760
rect 18920 652440 19235 652760
rect 34054 652755 34372 652759
rect 34054 652445 34058 652755
rect 34058 652445 34368 652755
rect 34368 652445 34372 652755
rect 34054 652441 34372 652445
rect 18915 652435 19235 652440
rect 14835 649252 17295 651712
rect 18820 649990 19140 650310
rect 32571 649991 32889 650309
rect 18915 649760 19235 649765
rect 18915 649440 18920 649760
rect 18920 649440 19235 649760
rect 34054 649755 34372 649759
rect 34054 649445 34058 649755
rect 34058 649445 34368 649755
rect 34368 649445 34372 649755
rect 34054 649441 34372 649445
rect 18915 649435 19235 649440
rect 18820 646990 19140 647310
rect 32571 646991 32889 647309
rect 424845 656024 425013 656028
rect 424845 655864 424849 656024
rect 424849 655864 425009 656024
rect 425009 655864 425013 656024
rect 424845 655860 425013 655864
rect 428429 650409 430889 652869
rect 492826 650141 495284 652599
rect 575238 678818 582000 682402
rect 553289 647541 554147 648399
rect 18915 646760 19235 646765
rect 18915 646440 18920 646760
rect 18920 646440 19235 646760
rect 34054 646755 34372 646759
rect 34054 646445 34058 646755
rect 34058 646445 34368 646755
rect 34368 646445 34372 646755
rect 34054 646441 34372 646445
rect 18915 646435 19235 646440
rect 14754 643842 17214 646302
rect 18820 643990 19140 644310
rect 32571 643991 32889 644309
rect 18915 643760 19235 643765
rect 18915 643440 18920 643760
rect 18920 643440 19235 643760
rect 18915 643435 19235 643440
rect 34054 643755 34372 643759
rect 34054 643445 34058 643755
rect 34058 643445 34368 643755
rect 34368 643445 34372 643755
rect 34054 643441 34372 643445
rect 18820 640990 19140 641310
rect 32571 640991 32889 641309
rect 18915 640760 19235 640765
rect 18915 640440 18920 640760
rect 18920 640440 19235 640760
rect 18915 640435 19235 640440
rect 34054 640755 34372 640759
rect 34054 640445 34058 640755
rect 34058 640445 34368 640755
rect 34368 640445 34372 640755
rect 34054 640441 34372 640445
rect 412602 639784 417402 644584
rect 18820 637990 19140 638310
rect 32571 637991 32889 638309
rect 18915 637760 19235 637765
rect 18915 637440 18920 637760
rect 18920 637440 19235 637760
rect 18915 637435 19235 637440
rect 34054 637755 34372 637759
rect 34054 637445 34058 637755
rect 34058 637445 34368 637755
rect 34368 637445 34372 637755
rect 34054 637441 34372 637445
rect 18820 634990 19140 635310
rect 32571 634991 32889 635309
rect 18915 634760 19235 634765
rect 18915 634440 18920 634760
rect 18920 634440 19235 634760
rect 18915 634435 19235 634440
rect 34054 634755 34372 634759
rect 34054 634445 34058 634755
rect 34058 634445 34368 634755
rect 34368 634445 34372 634755
rect 34054 634441 34372 634445
rect 18820 631990 19140 632310
rect 32571 631991 32889 632309
rect 412469 632244 417269 634584
rect 18915 631760 19235 631765
rect 18915 631440 18920 631760
rect 18920 631440 19235 631760
rect 34054 631755 34372 631759
rect 34054 631445 34058 631755
rect 34058 631445 34368 631755
rect 34368 631445 34372 631755
rect 34054 631441 34372 631445
rect 18915 631435 19235 631440
rect 11334 627835 13792 630293
rect 412468 629784 417269 632244
rect 451369 629784 456169 634584
rect 460694 629784 465494 634584
rect 18915 625760 19235 625765
rect 18915 625440 18920 625760
rect 18920 625440 19235 625760
rect 34054 625755 34372 625759
rect 34054 625445 34058 625755
rect 34058 625445 34368 625755
rect 34368 625445 34372 625755
rect 34054 625441 34372 625445
rect 404762 627989 407222 627994
rect 404762 625529 404767 627989
rect 404767 625529 407222 627989
rect 428430 627984 430888 627988
rect 428430 625534 428434 627984
rect 428434 625534 430884 627984
rect 430884 625534 430888 627984
rect 428430 625530 430888 625534
rect 404762 625524 407222 625529
rect 18915 625435 19235 625440
rect 11078 622087 13833 624842
rect 18820 622990 19140 623310
rect 32571 622991 32889 623309
rect 18915 622760 19235 622765
rect 18915 622440 18920 622760
rect 18920 622440 19235 622760
rect 34054 622755 34372 622759
rect 34054 622445 34058 622755
rect 34058 622445 34368 622755
rect 34368 622445 34372 622755
rect 34054 622441 34372 622445
rect 18915 622435 19235 622440
rect 18820 619990 19140 620310
rect 32571 619991 32889 620309
rect 18915 619760 19235 619765
rect 18915 619440 18920 619760
rect 18920 619440 19235 619760
rect 34054 619755 34372 619759
rect 34054 619445 34058 619755
rect 34058 619445 34368 619755
rect 34368 619445 34372 619755
rect 34054 619441 34372 619445
rect 18915 619435 19235 619440
rect 15232 614713 17987 617468
rect 18820 616990 19140 617310
rect 32571 616991 32889 617309
rect 18915 616760 19235 616765
rect 18915 616440 18920 616760
rect 18920 616440 19235 616760
rect 34054 616755 34372 616759
rect 34054 616445 34058 616755
rect 34058 616445 34368 616755
rect 34368 616445 34372 616755
rect 34054 616441 34372 616445
rect 18915 616435 19235 616440
rect 18820 613990 19140 614310
rect 32571 613991 32889 614309
rect 18915 613760 19235 613765
rect 18915 613440 18920 613760
rect 18920 613440 19235 613760
rect 34054 613755 34372 613759
rect 34054 613445 34058 613755
rect 34058 613445 34368 613755
rect 34368 613445 34372 613755
rect 34054 613441 34372 613445
rect 18915 613435 19235 613440
rect 404902 615819 407362 615824
rect 404902 613359 404907 615819
rect 404907 613359 407362 615819
rect 404902 613354 407362 613359
rect 428430 613360 430888 615818
rect 18820 610990 19140 611310
rect 32571 610991 32889 611309
rect 18915 610760 19235 610765
rect 18915 610440 18920 610760
rect 18920 610440 19235 610760
rect 34054 610755 34372 610759
rect 34054 610445 34058 610755
rect 34058 610445 34368 610755
rect 34368 610445 34372 610755
rect 34054 610441 34372 610445
rect 18915 610435 19235 610440
rect 13717 607375 16472 610130
rect 18820 607990 19140 608310
rect 32571 607991 32889 608309
rect 18915 607760 19235 607765
rect 18915 607440 18920 607760
rect 18920 607440 19235 607760
rect 34054 607755 34372 607759
rect 34054 607445 34058 607755
rect 34058 607445 34368 607755
rect 34368 607445 34372 607755
rect 34054 607441 34372 607445
rect 18915 607435 19235 607440
rect 11078 602850 13833 605645
rect 18820 604990 19140 605310
rect 32571 604991 32889 605309
rect 18915 604760 19235 604765
rect 18915 604440 18920 604760
rect 18920 604440 19235 604760
rect 34054 604755 34372 604759
rect 34054 604445 34058 604755
rect 34058 604445 34368 604755
rect 34368 604445 34372 604755
rect 34054 604441 34372 604445
rect 18915 604435 19235 604440
rect 18820 601990 19140 602310
rect 32571 601991 32889 602309
rect 18915 601760 19235 601765
rect 18915 601440 18920 601760
rect 18920 601440 19235 601760
rect 34054 601755 34372 601759
rect 34054 601445 34058 601755
rect 34058 601445 34368 601755
rect 34368 601445 34372 601755
rect 34054 601441 34372 601445
rect 18915 601435 19235 601440
rect 404413 602180 406873 602185
rect 404413 599720 404418 602180
rect 404418 599720 406873 602180
rect 428430 602175 430888 602179
rect 428430 599725 428434 602175
rect 428434 599725 430884 602175
rect 430884 599725 430888 602175
rect 428430 599721 430888 599725
rect 404413 599715 406873 599720
rect 18820 598990 19140 599310
rect 32571 598991 32889 599309
rect 18915 598760 19235 598765
rect 18915 598440 18920 598760
rect 18920 598440 19235 598760
rect 34054 598755 34372 598759
rect 34054 598445 34058 598755
rect 34058 598445 34368 598755
rect 34368 598445 34372 598755
rect 34054 598441 34372 598445
rect 18915 598435 19235 598440
rect 14987 594555 17742 597310
rect 18820 595990 19140 596310
rect 32571 595991 32889 596309
rect 18915 595760 19235 595765
rect 18915 595440 18920 595760
rect 18920 595440 19235 595760
rect 34054 595755 34372 595759
rect 34054 595445 34058 595755
rect 34058 595445 34368 595755
rect 34368 595445 34372 595755
rect 34054 595441 34372 595445
rect 18915 595435 19235 595440
rect 413053 594404 415511 596862
rect 18820 592990 19140 593310
rect 32571 592991 32889 593309
rect 18915 592760 19235 592765
rect 18915 592440 18920 592760
rect 18920 592440 19235 592760
rect 34054 592755 34372 592759
rect 34054 592445 34058 592755
rect 34058 592445 34368 592755
rect 34368 592445 34372 592755
rect 34054 592441 34372 592445
rect 18915 592435 19235 592440
rect 18820 589990 19140 590310
rect 32571 589991 32889 590309
rect 14577 586732 17332 589487
rect 18915 589760 19235 589765
rect 18915 589440 18920 589760
rect 18920 589440 19235 589760
rect 34054 589755 34372 589759
rect 34054 589445 34058 589755
rect 34058 589445 34368 589755
rect 34368 589445 34372 589755
rect 34054 589441 34372 589445
rect 18915 589435 19235 589440
rect 18820 586990 19140 587310
rect 32571 586991 32889 587309
rect 18915 586760 19235 586765
rect 18915 586440 18920 586760
rect 18920 586440 19235 586760
rect 34054 586755 34372 586759
rect 34054 586445 34058 586755
rect 34058 586445 34368 586755
rect 34368 586445 34372 586755
rect 34054 586441 34372 586445
rect 18915 586435 19235 586440
rect 403713 587353 406173 587358
rect 403713 584893 403718 587353
rect 403718 584893 406173 587353
rect 428430 587348 430888 587352
rect 428430 584898 428434 587348
rect 428434 584898 430884 587348
rect 430884 584898 430888 587348
rect 428430 584894 430888 584898
rect 403713 584888 406173 584893
rect 14536 581284 17291 584039
rect 18820 583990 19140 584310
rect 32571 583991 32889 584309
rect 18915 583760 19235 583765
rect 18915 583440 18920 583760
rect 18920 583440 19235 583760
rect 34054 583755 34372 583759
rect 34054 583445 34058 583755
rect 34058 583445 34368 583755
rect 34368 583445 34372 583755
rect 34054 583441 34372 583445
rect 18915 583435 19235 583440
rect 18820 580990 19140 581310
rect 32571 580991 32889 581309
rect 18915 580760 19235 580765
rect 18915 580440 18920 580760
rect 18920 580440 19235 580760
rect 34054 580755 34372 580759
rect 34054 580445 34058 580755
rect 34058 580445 34368 580755
rect 34368 580445 34372 580755
rect 34054 580441 34372 580445
rect 18915 580435 19235 580440
rect 14577 575836 17332 578591
rect 18820 577990 19140 578310
rect 32571 577991 32889 578309
rect 18915 577760 19235 577765
rect 18915 577440 18920 577760
rect 18920 577440 19235 577760
rect 34054 577755 34372 577759
rect 34054 577445 34058 577755
rect 34058 577445 34368 577755
rect 34368 577445 34372 577755
rect 34054 577441 34372 577445
rect 18915 577435 19235 577440
rect 18820 574990 19140 575310
rect 32571 574991 32889 575309
rect 18915 574760 19235 574765
rect 18915 574440 18920 574760
rect 18920 574440 19235 574760
rect 34054 574755 34372 574759
rect 34054 574445 34058 574755
rect 34058 574445 34368 574755
rect 34368 574445 34372 574755
rect 34054 574441 34372 574445
rect 18915 574435 19235 574440
rect 18820 571990 19140 572310
rect 32571 571991 32889 572309
rect 14946 568832 17701 571587
rect 18915 571760 19235 571765
rect 18915 571440 18920 571760
rect 18920 571440 19235 571760
rect 34054 571755 34372 571759
rect 34054 571445 34058 571755
rect 34058 571445 34368 571755
rect 34368 571445 34372 571755
rect 34054 571441 34372 571445
rect 18915 571435 19235 571440
rect 18820 568990 19140 569310
rect 32571 568991 32889 569309
rect 413175 569040 417975 573840
rect 18915 568760 19235 568765
rect 18915 568440 18920 568760
rect 18920 568440 19235 568760
rect 34054 568755 34372 568759
rect 34054 568445 34058 568755
rect 34058 568445 34368 568755
rect 34368 568445 34372 568755
rect 34054 568441 34372 568445
rect 18915 568435 19235 568440
rect 18820 565990 19140 566310
rect 32571 565991 32889 566309
rect 18915 565760 19235 565765
rect 18915 565440 18920 565760
rect 18920 565440 19235 565760
rect 34054 565755 34372 565759
rect 34054 565445 34058 565755
rect 34058 565445 34368 565755
rect 34368 565445 34372 565755
rect 34054 565441 34372 565445
rect 18915 565435 19235 565440
rect 15150 562115 17905 564870
rect 404348 566278 406808 566283
rect 404348 563818 404353 566278
rect 404353 563818 406808 566278
rect 428430 566273 430888 566277
rect 428430 563823 428434 566273
rect 428434 563823 430884 566273
rect 430884 563823 430888 566273
rect 428430 563819 430888 563823
rect 404348 563813 406808 563818
rect 18820 562990 19140 563310
rect 32571 562991 32889 563309
rect 18915 562760 19235 562765
rect 18915 562440 18920 562760
rect 18920 562440 19235 562760
rect 34054 562755 34372 562759
rect 34054 562445 34058 562755
rect 34058 562445 34368 562755
rect 34368 562445 34372 562755
rect 34054 562441 34372 562445
rect 18915 562435 19235 562440
rect 15355 557978 18110 560733
rect 18820 559990 19140 560310
rect 32571 559991 32889 560309
rect 18915 559760 19235 559765
rect 18915 559440 18920 559760
rect 18920 559440 19235 559760
rect 34054 559755 34372 559759
rect 34054 559445 34058 559755
rect 34058 559445 34368 559755
rect 34368 559445 34372 559755
rect 34054 559441 34372 559445
rect 18915 559435 19235 559440
rect 413355 557385 418155 562185
rect 18820 556990 19140 557310
rect 32571 556991 32889 557309
rect 18915 556760 19235 556765
rect 18915 556440 18920 556760
rect 18920 556440 19235 556760
rect 34054 556755 34372 556759
rect 34054 556445 34058 556755
rect 34058 556445 34368 556755
rect 34368 556445 34372 556755
rect 34054 556441 34372 556445
rect 18915 556435 19235 556440
rect 14659 552079 17414 554834
rect 18820 553990 19140 554310
rect 32571 553991 32889 554309
rect 18915 553760 19235 553765
rect 18915 553440 18920 553760
rect 18920 553440 19235 553760
rect 34054 553755 34372 553759
rect 34054 553445 34058 553755
rect 34058 553445 34368 553755
rect 34368 553445 34372 553755
rect 34054 553441 34372 553445
rect 18915 553435 19235 553440
rect 18820 550990 19140 551310
rect 32571 550991 32889 551309
rect 18915 550760 19235 550765
rect 18915 550440 18920 550760
rect 18920 550440 19235 550760
rect 34054 550755 34372 550759
rect 34054 550445 34058 550755
rect 34058 550445 34368 550755
rect 34368 550445 34372 550755
rect 34054 550441 34372 550445
rect 18915 550435 19235 550440
rect 404422 552465 406882 552470
rect 404422 550005 404427 552465
rect 404427 550005 406882 552465
rect 428430 552460 430888 552464
rect 428430 550010 428434 552460
rect 428434 550010 430884 552460
rect 430884 550010 430888 552460
rect 428430 550006 430888 550010
rect 404422 550000 406882 550005
rect 18820 547990 19140 548310
rect 32571 547991 32889 548309
rect 18915 547760 19235 547765
rect 18915 547440 18920 547760
rect 18920 547440 19235 547760
rect 34054 547755 34372 547759
rect 34054 547445 34058 547755
rect 34058 547445 34368 547755
rect 34368 547445 34372 547755
rect 34054 547441 34372 547445
rect 18915 547435 19235 547440
rect 14946 544666 17701 547421
rect 18820 544990 19140 545310
rect 32571 544991 32889 545309
rect 18915 544760 19235 544765
rect 18915 544440 18920 544760
rect 18920 544440 19235 544760
rect 34054 544755 34372 544759
rect 34054 544445 34058 544755
rect 34058 544445 34368 544755
rect 34368 544445 34372 544755
rect 34054 544441 34372 544445
rect 18915 544435 19235 544440
rect 18820 541990 19140 542310
rect 32571 541991 32889 542309
rect 18915 541760 19235 541765
rect 18915 541440 18920 541760
rect 18920 541440 19235 541760
rect 34054 541755 34372 541759
rect 34054 541445 34058 541755
rect 34058 541445 34368 541755
rect 34368 541445 34372 541755
rect 34054 541441 34372 541445
rect 18915 541435 19235 541440
rect 15724 537989 18479 540744
rect 404128 542841 406588 542846
rect 404128 540381 404133 542841
rect 404133 540381 406588 542841
rect 428430 542836 430888 542840
rect 428430 540386 428434 542836
rect 428434 540386 430884 542836
rect 430884 540386 430888 542836
rect 428430 540382 430888 540386
rect 404128 540376 406588 540381
rect 18820 538990 19140 539310
rect 32571 538991 32889 539309
rect 18915 538760 19235 538765
rect 18915 538440 18920 538760
rect 18920 538440 19235 538760
rect 34054 538755 34372 538759
rect 34054 538445 34058 538755
rect 34058 538445 34368 538755
rect 34368 538445 34372 538755
rect 34054 538441 34372 538445
rect 18915 538435 19235 538440
rect 18820 535990 19140 536310
rect 32571 535991 32889 536309
rect 18915 535760 19235 535765
rect 18915 535440 18920 535760
rect 18920 535440 19235 535760
rect 34054 535755 34372 535759
rect 34054 535445 34058 535755
rect 34058 535445 34368 535755
rect 34368 535445 34372 535755
rect 34054 535441 34372 535445
rect 18915 535435 19235 535440
rect 18820 532990 19140 533310
rect 32571 532991 32889 533309
rect 15314 529879 18069 532634
rect 18915 532760 19235 532765
rect 18915 532440 18920 532760
rect 18920 532440 19235 532760
rect 34054 532755 34372 532759
rect 34054 532445 34058 532755
rect 34058 532445 34368 532755
rect 34368 532445 34372 532755
rect 34054 532441 34372 532445
rect 18915 532435 19235 532440
rect 18820 529990 19140 530310
rect 32571 529991 32889 530309
rect 18915 529760 19235 529765
rect 18915 529440 18920 529760
rect 18920 529440 19235 529760
rect 34054 529755 34372 529759
rect 34054 529445 34058 529755
rect 34058 529445 34368 529755
rect 34368 529445 34372 529755
rect 34054 529441 34372 529445
rect 18915 529435 19235 529440
rect 404128 531893 406588 531898
rect 404128 529433 404133 531893
rect 404133 529433 406588 531893
rect 428430 531888 430888 531892
rect 428430 529438 428434 531888
rect 428434 529438 430884 531888
rect 430884 529438 430888 531888
rect 428430 529434 430888 529438
rect 404128 529428 406588 529433
rect 18820 526990 19140 527310
rect 32571 526991 32889 527309
rect 18915 526760 19235 526765
rect 18915 526440 18920 526760
rect 18920 526440 19235 526760
rect 34054 526755 34372 526759
rect 34054 526445 34058 526755
rect 34058 526445 34368 526755
rect 34368 526445 34372 526755
rect 34054 526441 34372 526445
rect 18915 526435 19235 526440
rect 15437 521441 18192 524196
rect 18820 523990 19140 524310
rect 32571 523991 32889 524309
rect 18915 523760 19235 523765
rect 18915 523440 18920 523760
rect 18920 523440 19235 523760
rect 34054 523755 34372 523759
rect 34054 523445 34058 523755
rect 34058 523445 34368 523755
rect 34368 523445 34372 523755
rect 34054 523441 34372 523445
rect 18915 523435 19235 523440
rect 18820 520990 19140 521310
rect 32571 520991 32889 521309
rect 413053 520820 415511 523278
rect 18915 520760 19235 520765
rect 18915 520440 18920 520760
rect 18920 520440 19235 520760
rect 34054 520755 34372 520759
rect 34054 520445 34058 520755
rect 34058 520445 34368 520755
rect 34368 520445 34372 520755
rect 34054 520441 34372 520445
rect 18915 520435 19235 520440
rect 18820 517990 19140 518310
rect 32571 517991 32889 518309
rect 18915 517760 19235 517765
rect 18915 517440 18920 517760
rect 18920 517440 19235 517760
rect 34054 517755 34372 517759
rect 34054 517445 34058 517755
rect 34058 517445 34368 517755
rect 34368 517445 34372 517755
rect 34054 517441 34372 517445
rect 18915 517435 19235 517440
rect 15355 514110 18110 516865
rect 18820 514990 19140 515310
rect 32571 514991 32889 515309
rect 18820 511990 19140 512310
rect 32571 511991 32889 512309
rect 15232 509235 17987 511990
rect 18915 511760 19235 511765
rect 18915 511440 18920 511760
rect 18920 511440 19235 511760
rect 34054 511755 34372 511759
rect 34054 511445 34058 511755
rect 34058 511445 34368 511755
rect 34368 511445 34372 511755
rect 34054 511441 34372 511445
rect 18915 511435 19235 511440
rect 404174 512943 406634 512948
rect 404174 510483 404179 512943
rect 404179 510483 406634 512943
rect 428430 512938 430888 512942
rect 428430 510488 428434 512938
rect 428434 510488 430884 512938
rect 430884 510488 430888 512938
rect 428430 510484 430888 510488
rect 404174 510478 406634 510483
rect 18820 508990 19140 509310
rect 32571 508991 32889 509309
rect 18915 508760 19235 508765
rect 18915 508440 18920 508760
rect 18920 508440 19235 508760
rect 34054 508755 34372 508759
rect 34054 508445 34058 508755
rect 34058 508445 34368 508755
rect 34368 508445 34372 508755
rect 34054 508441 34372 508445
rect 18915 508435 19235 508440
rect 15642 505549 18397 508304
rect 18820 505990 19140 506310
rect 32571 505991 32889 506309
rect 18915 505760 19235 505765
rect 18915 505440 18920 505760
rect 18920 505440 19235 505760
rect 34054 505755 34372 505759
rect 34054 505445 34058 505755
rect 34058 505445 34368 505755
rect 34368 505445 34372 505755
rect 34054 505441 34372 505445
rect 18915 505435 19235 505440
rect 18820 502990 19140 503310
rect 32571 502991 32889 503309
rect 18915 502760 19235 502765
rect 18915 502440 18920 502760
rect 18920 502440 19235 502760
rect 34054 502755 34372 502759
rect 34054 502445 34058 502755
rect 34058 502445 34368 502755
rect 34368 502445 34372 502755
rect 34054 502441 34372 502445
rect 18915 502435 19235 502440
rect 18820 499990 19140 500310
rect 32571 499991 32889 500309
rect 11078 497132 13833 499927
rect 18915 499760 19235 499765
rect 18915 499440 18920 499760
rect 18920 499440 19235 499760
rect 34054 499755 34372 499759
rect 34054 499445 34058 499755
rect 34058 499445 34368 499755
rect 34368 499445 34372 499755
rect 34054 499441 34372 499445
rect 18915 499435 19235 499440
rect 18820 496990 19140 497310
rect 32571 496991 32889 497309
rect 18915 496760 19235 496765
rect 18915 496440 18920 496760
rect 18920 496440 19235 496760
rect 34054 496755 34372 496759
rect 34054 496445 34058 496755
rect 34058 496445 34368 496755
rect 34368 496445 34372 496755
rect 34054 496441 34372 496445
rect 18915 496435 19235 496440
rect 413053 494836 415511 497294
rect 18820 493990 19140 494310
rect 32571 493991 32889 494309
rect 18915 493760 19235 493765
rect 18915 493440 18920 493760
rect 18920 493440 19235 493760
rect 34054 493755 34372 493759
rect 34054 493445 34058 493755
rect 34058 493445 34368 493755
rect 34368 493445 34372 493755
rect 34054 493441 34372 493445
rect 18915 493435 19235 493440
rect 15273 490148 18028 492903
rect 18820 490990 19140 491310
rect 32571 490991 32889 491309
rect 18915 490760 19235 490765
rect 18915 490440 18920 490760
rect 18920 490440 19235 490760
rect 34054 490755 34372 490759
rect 34054 490445 34058 490755
rect 34058 490445 34368 490755
rect 34368 490445 34372 490755
rect 34054 490441 34372 490445
rect 18915 490435 19235 490440
rect 18820 487990 19140 488310
rect 32571 487991 32889 488309
rect 18915 487760 19235 487765
rect 18915 487440 18920 487760
rect 18920 487440 19235 487760
rect 34054 487755 34372 487759
rect 34054 487445 34058 487755
rect 34058 487445 34368 487755
rect 34368 487445 34372 487755
rect 34054 487441 34372 487445
rect 18915 487435 19235 487440
rect 14495 483430 17250 486185
rect 18820 484990 19140 485310
rect 32571 484991 32889 485309
rect 18915 484760 19235 484765
rect 18915 484440 18920 484760
rect 18920 484440 19235 484760
rect 34054 484755 34372 484759
rect 34054 484445 34058 484755
rect 34058 484445 34368 484755
rect 34368 484445 34372 484755
rect 34054 484441 34372 484445
rect 18915 484435 19235 484440
rect 404455 486407 406915 486412
rect 404455 483947 404460 486407
rect 404460 483947 406915 486407
rect 428430 486402 430888 486406
rect 428430 483952 428434 486402
rect 428434 483952 430884 486402
rect 430884 483952 430888 486402
rect 428430 483948 430888 483952
rect 404455 483942 406915 483947
rect 1920 353274 4378 353278
rect 1920 350824 1924 353274
rect 1924 350824 4374 353274
rect 4374 350824 4378 353274
rect 1920 350820 4378 350824
rect 1920 348745 4378 348749
rect 1920 346295 1924 348745
rect 1924 346295 4374 348745
rect 4374 346295 4378 348745
rect 1920 346291 4378 346295
rect 1920 344235 4378 344239
rect 1920 341785 1924 344235
rect 1924 341785 4374 344235
rect 4374 341785 4378 344235
rect 1920 341781 4378 341785
rect 18820 481990 19140 482310
rect 32571 481991 32889 482309
rect 18915 481760 19235 481765
rect 18915 481440 18920 481760
rect 18920 481440 19235 481760
rect 34054 481755 34372 481759
rect 34054 481445 34058 481755
rect 34058 481445 34368 481755
rect 34368 481445 34372 481755
rect 34054 481441 34372 481445
rect 18915 481435 19235 481440
rect 18820 478990 19140 479310
rect 32571 478991 32889 479309
rect 18915 478760 19235 478765
rect 18915 478440 18920 478760
rect 18920 478440 19235 478760
rect 34054 478755 34372 478759
rect 34054 478445 34058 478755
rect 34058 478445 34368 478755
rect 34368 478445 34372 478755
rect 34054 478441 34372 478445
rect 18915 478435 19235 478440
rect 18820 475990 19140 476310
rect 32571 475991 32889 476309
rect 18915 475760 19235 475765
rect 18915 475440 18920 475760
rect 18920 475440 19235 475760
rect 34054 475755 34372 475759
rect 34054 475445 34058 475755
rect 34058 475445 34368 475755
rect 34368 475445 34372 475755
rect 34054 475441 34372 475445
rect 18915 475435 19235 475440
rect 18820 472990 19140 473310
rect 32571 472991 32889 473309
rect 18915 472760 19235 472765
rect 18915 472440 18920 472760
rect 18920 472440 19235 472760
rect 34054 472755 34372 472759
rect 34054 472445 34058 472755
rect 34058 472445 34368 472755
rect 34368 472445 34372 472755
rect 34054 472441 34372 472445
rect 18915 472435 19235 472440
rect 18820 469990 19140 470310
rect 32571 469991 32889 470309
rect 18915 469760 19235 469765
rect 18915 469440 18920 469760
rect 18920 469440 19235 469760
rect 34054 469755 34372 469759
rect 34054 469445 34058 469755
rect 34058 469445 34368 469755
rect 34368 469445 34372 469755
rect 34054 469441 34372 469445
rect 18915 469435 19235 469440
rect 18820 466990 19140 467310
rect 32571 466991 32889 467309
rect 18915 466760 19235 466765
rect 18915 466440 18920 466760
rect 18920 466440 19235 466760
rect 34054 466755 34372 466759
rect 34054 466445 34058 466755
rect 34058 466445 34368 466755
rect 34368 466445 34372 466755
rect 34054 466441 34372 466445
rect 18915 466435 19235 466440
rect 18820 463990 19140 464310
rect 32571 463991 32889 464309
rect 18915 463760 19235 463765
rect 18915 463440 18920 463760
rect 18920 463440 19235 463760
rect 34054 463755 34372 463759
rect 34054 463445 34058 463755
rect 34058 463445 34368 463755
rect 34368 463445 34372 463755
rect 34054 463441 34372 463445
rect 18915 463435 19235 463440
rect 413053 462872 415511 465330
rect 11078 458587 13833 461424
rect 18820 460990 19140 461310
rect 32571 460991 32889 461309
rect 18915 460760 19235 460765
rect 18915 460440 18920 460760
rect 18920 460440 19235 460760
rect 34054 460755 34372 460759
rect 34054 460445 34058 460755
rect 34058 460445 34368 460755
rect 34368 460445 34372 460755
rect 34054 460441 34372 460445
rect 18915 460435 19235 460440
rect 18820 457990 19140 458310
rect 32571 457991 32889 458309
rect 18915 457760 19235 457765
rect 18915 457440 18920 457760
rect 18920 457440 19235 457760
rect 34054 457755 34372 457759
rect 34054 457445 34058 457755
rect 34058 457445 34368 457755
rect 34368 457445 34372 457755
rect 34054 457441 34372 457445
rect 18915 457435 19235 457440
rect 18820 454990 19140 455310
rect 32571 454991 32889 455309
rect 18915 454760 19235 454765
rect 18915 454440 18920 454760
rect 18920 454440 19235 454760
rect 34054 454755 34372 454759
rect 34054 454445 34058 454755
rect 34058 454445 34368 454755
rect 34368 454445 34372 454755
rect 34054 454441 34372 454445
rect 18915 454435 19235 454440
rect 18820 451990 19140 452310
rect 32571 451991 32889 452309
rect 18915 451760 19235 451765
rect 18915 451440 18920 451760
rect 18920 451440 19235 451760
rect 34054 451755 34372 451759
rect 34054 451445 34058 451755
rect 34058 451445 34368 451755
rect 34368 451445 34372 451755
rect 34054 451441 34372 451445
rect 18915 451435 19235 451440
rect 18820 448990 19140 449310
rect 32571 448991 32889 449309
rect 18915 448760 19235 448765
rect 18915 448440 18920 448760
rect 18920 448440 19235 448760
rect 34054 448755 34372 448759
rect 34054 448445 34058 448755
rect 34058 448445 34368 448755
rect 34368 448445 34372 448755
rect 34054 448441 34372 448445
rect 18915 448435 19235 448440
rect 404476 449962 406936 449967
rect 404476 447502 404481 449962
rect 404481 447502 406936 449962
rect 428430 449957 430888 449961
rect 428430 447507 428434 449957
rect 428434 447507 430884 449957
rect 430884 447507 430888 449957
rect 428430 447503 430888 447507
rect 404476 447497 406936 447502
rect 18820 445990 19140 446310
rect 32571 445991 32889 446309
rect 18915 445760 19235 445765
rect 18915 445440 18920 445760
rect 18920 445440 19235 445760
rect 34054 445755 34372 445759
rect 34054 445445 34058 445755
rect 34058 445445 34368 445755
rect 34368 445445 34372 445755
rect 34054 445441 34372 445445
rect 18915 445435 19235 445440
rect 18820 442990 19140 443310
rect 32571 442991 32889 443309
rect 18915 442760 19235 442765
rect 18915 442440 18920 442760
rect 18920 442440 19235 442760
rect 34054 442755 34372 442759
rect 34054 442445 34058 442755
rect 34058 442445 34368 442755
rect 34368 442445 34372 442755
rect 34054 442441 34372 442445
rect 18915 442435 19235 442440
rect 18820 439990 19140 440310
rect 32571 439991 32889 440309
rect 18915 439760 19235 439765
rect 18915 439440 18920 439760
rect 18920 439440 19235 439760
rect 34054 439755 34372 439759
rect 34054 439445 34058 439755
rect 34058 439445 34368 439755
rect 34368 439445 34372 439755
rect 34054 439441 34372 439445
rect 18915 439435 19235 439440
rect 18820 436990 19140 437310
rect 32571 436991 32889 437309
rect 18915 436760 19235 436765
rect 18915 436440 18920 436760
rect 18920 436440 19235 436760
rect 34054 436755 34372 436759
rect 34054 436445 34058 436755
rect 34058 436445 34368 436755
rect 34368 436445 34372 436755
rect 34054 436441 34372 436445
rect 18915 436435 19235 436440
rect 18820 433990 19140 434310
rect 32571 433991 32889 434309
rect 18915 433760 19235 433765
rect 18915 433440 18920 433760
rect 18920 433440 19235 433760
rect 34054 433755 34372 433759
rect 34054 433445 34058 433755
rect 34058 433445 34368 433755
rect 34368 433445 34372 433755
rect 34054 433441 34372 433445
rect 18915 433435 19235 433440
rect 413053 433439 415511 435897
rect 18820 430990 19140 431310
rect 32571 430991 32889 431309
rect 18915 430760 19235 430765
rect 18915 430440 18920 430760
rect 18920 430440 19235 430760
rect 34054 430755 34372 430759
rect 34054 430445 34058 430755
rect 34058 430445 34368 430755
rect 34368 430445 34372 430755
rect 34054 430441 34372 430445
rect 18915 430435 19235 430440
rect 14457 427174 17212 429929
rect 18820 427990 19140 428310
rect 32571 427991 32889 428309
rect 18915 427760 19235 427765
rect 18915 427440 18920 427760
rect 18920 427440 19235 427760
rect 34054 427755 34372 427759
rect 34054 427445 34058 427755
rect 34058 427445 34368 427755
rect 34368 427445 34372 427755
rect 34054 427441 34372 427445
rect 18915 427435 19235 427440
rect 18820 424990 19140 425310
rect 32571 424991 32889 425309
rect 18915 424760 19235 424765
rect 18915 424440 18920 424760
rect 18920 424440 19235 424760
rect 18915 424435 19235 424440
rect 34054 424755 34372 424759
rect 34054 424445 34058 424755
rect 34058 424445 34368 424755
rect 34368 424445 34372 424755
rect 34054 424441 34372 424445
rect 18820 421990 19140 422310
rect 32571 421991 32889 422309
rect 18915 421760 19235 421765
rect 18915 421440 18920 421760
rect 18920 421440 19235 421760
rect 18915 421435 19235 421440
rect 34054 421755 34372 421759
rect 34054 421445 34058 421755
rect 34058 421445 34368 421755
rect 34368 421445 34372 421755
rect 34054 421441 34372 421445
rect 18820 418990 19140 419310
rect 32571 418991 32889 419309
rect 404808 421579 407268 421584
rect 404808 419119 404813 421579
rect 404813 419119 407268 421579
rect 428430 421574 430888 421578
rect 428430 419124 428434 421574
rect 428434 419124 430884 421574
rect 430884 419124 430888 421574
rect 428430 419120 430888 419124
rect 404808 419114 407268 419119
rect 18915 418760 19235 418765
rect 18915 418440 18920 418760
rect 18920 418440 19235 418760
rect 18915 418435 19235 418440
rect 34054 418755 34372 418759
rect 34054 418445 34058 418755
rect 34058 418445 34368 418755
rect 34368 418445 34372 418755
rect 34054 418441 34372 418445
rect 18820 415990 19140 416310
rect 32571 415991 32889 416309
rect 18915 415760 19235 415765
rect 18915 415440 18920 415760
rect 18920 415440 19235 415760
rect 18915 415435 19235 415440
rect 34054 415755 34372 415759
rect 34054 415445 34058 415755
rect 34058 415445 34368 415755
rect 34368 415445 34372 415755
rect 34054 415441 34372 415445
rect 18820 412990 19140 413310
rect 32571 412991 32889 413309
rect 18915 412760 19235 412765
rect 18915 412440 18920 412760
rect 18920 412440 19235 412760
rect 18915 412435 19235 412440
rect 34054 412755 34372 412759
rect 34054 412445 34058 412755
rect 34058 412445 34368 412755
rect 34368 412445 34372 412755
rect 34054 412441 34372 412445
rect 18820 409990 19140 410310
rect 32571 409991 32889 410309
rect 18915 409760 19235 409765
rect 18915 409440 18920 409760
rect 18920 409440 19235 409760
rect 18915 409435 19235 409440
rect 34054 409755 34372 409759
rect 34054 409445 34058 409755
rect 34058 409445 34368 409755
rect 34368 409445 34372 409755
rect 34054 409441 34372 409445
rect 18820 406990 19140 407310
rect 32571 406991 32889 407309
rect 404574 409691 407034 409696
rect 404574 407231 404579 409691
rect 404579 407231 407034 409691
rect 428430 409686 430888 409690
rect 428430 407236 428434 409686
rect 428434 407236 430884 409686
rect 430884 407236 430888 409686
rect 428430 407232 430888 407236
rect 404574 407226 407034 407231
rect 18915 406760 19235 406765
rect 18915 406440 18920 406760
rect 18920 406440 19235 406760
rect 18915 406435 19235 406440
rect 34054 406755 34372 406759
rect 34054 406445 34058 406755
rect 34058 406445 34368 406755
rect 34368 406445 34372 406755
rect 34054 406441 34372 406445
rect 18820 403990 19140 404310
rect 32571 403991 32889 404309
rect 18915 403760 19235 403765
rect 18915 403440 18920 403760
rect 18920 403440 19235 403760
rect 18915 403435 19235 403440
rect 34054 403755 34372 403759
rect 34054 403445 34058 403755
rect 34058 403445 34368 403755
rect 34368 403445 34372 403755
rect 34054 403441 34372 403445
rect 18820 400990 19140 401310
rect 32571 400991 32889 401309
rect 18820 397990 19140 398310
rect 32571 397991 32889 398309
rect 18915 397760 19235 397765
rect 18915 397440 18920 397760
rect 18920 397440 19235 397760
rect 18915 397435 19235 397440
rect 34054 397755 34372 397759
rect 34054 397445 34058 397755
rect 34058 397445 34368 397755
rect 34368 397445 34372 397755
rect 34054 397441 34372 397445
rect 413053 397336 415511 399794
rect 18820 394990 19140 395310
rect 32571 394991 32889 395309
rect 18915 394760 19235 394765
rect 18915 394440 18920 394760
rect 18920 394440 19235 394760
rect 18915 394435 19235 394440
rect 34054 394755 34372 394759
rect 34054 394445 34058 394755
rect 34058 394445 34368 394755
rect 34368 394445 34372 394755
rect 34054 394441 34372 394445
rect 18820 391990 19140 392310
rect 32571 391991 32889 392309
rect 18915 391760 19235 391765
rect 18915 391440 18920 391760
rect 18920 391440 19235 391760
rect 18915 391435 19235 391440
rect 34054 391755 34372 391759
rect 34054 391445 34058 391755
rect 34058 391445 34368 391755
rect 34368 391445 34372 391755
rect 34054 391441 34372 391445
rect 18820 388990 19140 389310
rect 32571 388991 32889 389309
rect 18915 388760 19235 388765
rect 18915 388440 18920 388760
rect 18920 388440 19235 388760
rect 18915 388435 19235 388440
rect 34054 388755 34372 388759
rect 34054 388445 34058 388755
rect 34058 388445 34368 388755
rect 34368 388445 34372 388755
rect 34054 388441 34372 388445
rect 18820 385990 19140 386310
rect 32571 385991 32889 386309
rect 18915 385760 19235 385765
rect 18915 385440 18920 385760
rect 18920 385440 19235 385760
rect 18915 385435 19235 385440
rect 34054 385755 34372 385759
rect 34054 385445 34058 385755
rect 34058 385445 34368 385755
rect 34368 385445 34372 385755
rect 34054 385441 34372 385445
rect 18820 382990 19140 383310
rect 32571 382991 32889 383309
rect 413053 383309 415511 385767
rect 18915 382760 19235 382765
rect 18915 382440 18920 382760
rect 18920 382440 19235 382760
rect 18915 382435 19235 382440
rect 34054 382755 34372 382759
rect 34054 382445 34058 382755
rect 34058 382445 34368 382755
rect 34368 382445 34372 382755
rect 34054 382441 34372 382445
rect 18820 379990 19140 380310
rect 32571 379991 32889 380309
rect 18915 379760 19235 379765
rect 18915 379440 18920 379760
rect 18920 379440 19235 379760
rect 18915 379435 19235 379440
rect 34054 379755 34372 379759
rect 34054 379445 34058 379755
rect 34058 379445 34368 379755
rect 34368 379445 34372 379755
rect 34054 379441 34372 379445
rect 414103 377762 414393 377767
rect 414103 377472 414388 377762
rect 414388 377472 414393 377762
rect 414103 377467 414393 377472
rect 18820 376990 19140 377310
rect 32571 376991 32889 377309
rect 413995 377075 414285 377080
rect 18915 376760 19235 376765
rect 18915 376440 18920 376760
rect 18920 376440 19235 376760
rect 18915 376435 19235 376440
rect 413995 376785 414280 377075
rect 414280 376785 414285 377075
rect 413995 376780 414285 376785
rect 34054 376755 34372 376759
rect 34054 376445 34058 376755
rect 34058 376445 34368 376755
rect 34368 376445 34372 376755
rect 34054 376441 34372 376445
rect 414248 376208 414538 376213
rect 414248 375918 414533 376208
rect 414533 375918 414538 376208
rect 414248 375913 414538 375918
rect 414031 374653 414321 374658
rect 414031 374363 414316 374653
rect 414316 374363 414321 374653
rect 414031 374358 414321 374363
rect 18820 373990 19140 374310
rect 32571 373991 32889 374309
rect 413999 374054 414289 374059
rect 18915 373760 19235 373765
rect 18915 373440 18920 373760
rect 18920 373440 19235 373760
rect 18915 373435 19235 373440
rect 413999 373764 414284 374054
rect 414284 373764 414289 374054
rect 413999 373759 414289 373764
rect 34054 373755 34372 373759
rect 34054 373445 34058 373755
rect 34058 373445 34368 373755
rect 34368 373445 34372 373755
rect 34054 373441 34372 373445
rect 414357 373194 414647 373199
rect 414357 372904 414642 373194
rect 414642 372904 414647 373194
rect 414357 372899 414647 372904
rect 414250 372477 414540 372482
rect 414250 372187 414535 372477
rect 414535 372187 414540 372477
rect 414250 372182 414540 372187
rect 414357 371832 414647 371837
rect 414357 371542 414642 371832
rect 414642 371542 414647 371832
rect 414357 371537 414647 371542
rect 18820 370990 19140 371310
rect 32571 370991 32889 371309
rect 414781 371295 415071 371300
rect 414781 371005 415066 371295
rect 415066 371005 415071 371295
rect 414781 371000 415071 371005
rect 18915 370760 19235 370765
rect 18915 370440 18920 370760
rect 18920 370440 19235 370760
rect 18915 370435 19235 370440
rect 34054 370755 34372 370759
rect 34054 370445 34058 370755
rect 34058 370445 34368 370755
rect 34368 370445 34372 370755
rect 34054 370441 34372 370445
rect 413777 370704 414067 370709
rect 413777 370414 414062 370704
rect 414062 370414 414067 370704
rect 413777 370409 414067 370414
rect 18820 367990 19140 368310
rect 32571 367991 32889 368309
rect 18915 367760 19235 367765
rect 18915 367440 18920 367760
rect 18920 367440 19235 367760
rect 18915 367435 19235 367440
rect 34054 367755 34372 367759
rect 34054 367445 34058 367755
rect 34058 367445 34368 367755
rect 34368 367445 34372 367755
rect 34054 367441 34372 367445
rect 18820 364990 19140 365310
rect 32571 364991 32889 365309
rect 18915 364760 19235 364765
rect 18915 364440 18920 364760
rect 18920 364440 19235 364760
rect 18915 364435 19235 364440
rect 34054 364755 34372 364759
rect 34054 364445 34058 364755
rect 34058 364445 34368 364755
rect 34368 364445 34372 364755
rect 34054 364441 34372 364445
rect 53819 364409 54137 364727
rect 18820 361990 19140 362310
rect 32571 361991 32889 362309
rect 14741 337916 17496 340671
rect 26655 353279 29115 353284
rect 26655 350819 29110 353279
rect 29110 350819 29115 353279
rect 26655 350814 29115 350819
rect 26581 348750 29041 348755
rect 26581 346290 29036 348750
rect 29036 346290 29041 348750
rect 26581 346285 29041 346290
rect 26581 344240 29041 344245
rect 26581 341780 29036 344240
rect 29036 341780 29041 344240
rect 26581 341775 29041 341780
rect 1920 315910 4378 315914
rect 1920 313460 1924 315910
rect 1924 313460 4374 315910
rect 4374 313460 4378 315910
rect 1920 313456 4378 313460
rect 39941 315915 42401 315920
rect 39941 313455 42396 315915
rect 42396 313455 42401 315915
rect 39941 313450 42401 313455
rect 5660 293269 5772 293381
rect 365000 362051 365170 362221
rect 8382 261315 8462 261320
rect 8382 261250 8387 261315
rect 8387 261250 8457 261315
rect 8457 261250 8462 261315
rect 404520 362175 406980 362180
rect 404520 359715 404525 362175
rect 404525 359715 406980 362175
rect 428430 362170 430888 362174
rect 428430 359720 428434 362170
rect 428434 359720 430884 362170
rect 430884 359720 430888 362170
rect 428430 359716 430888 359720
rect 404520 359710 406980 359715
rect 55308 345751 55626 345755
rect 55308 345441 55312 345751
rect 55312 345441 55622 345751
rect 55622 345441 55626 345751
rect 55308 345437 55626 345441
rect 58308 345751 58626 345755
rect 58308 345441 58312 345751
rect 58312 345441 58622 345751
rect 58622 345441 58626 345751
rect 58308 345437 58626 345441
rect 61308 345751 61626 345755
rect 61308 345441 61312 345751
rect 61312 345441 61622 345751
rect 61622 345441 61626 345751
rect 61308 345437 61626 345441
rect 64308 345751 64626 345755
rect 64308 345441 64312 345751
rect 64312 345441 64622 345751
rect 64622 345441 64626 345751
rect 64308 345437 64626 345441
rect 67308 345751 67626 345755
rect 67308 345441 67312 345751
rect 67312 345441 67622 345751
rect 67622 345441 67626 345751
rect 67308 345437 67626 345441
rect 70308 345751 70626 345755
rect 70308 345441 70312 345751
rect 70312 345441 70622 345751
rect 70622 345441 70626 345751
rect 70308 345437 70626 345441
rect 73308 345751 73626 345755
rect 73308 345441 73312 345751
rect 73312 345441 73622 345751
rect 73622 345441 73626 345751
rect 73308 345437 73626 345441
rect 76308 345751 76626 345755
rect 76308 345441 76312 345751
rect 76312 345441 76622 345751
rect 76622 345441 76626 345751
rect 76308 345437 76626 345441
rect 79308 345751 79626 345755
rect 79308 345441 79312 345751
rect 79312 345441 79622 345751
rect 79622 345441 79626 345751
rect 79308 345437 79626 345441
rect 82308 345751 82626 345755
rect 82308 345441 82312 345751
rect 82312 345441 82622 345751
rect 82622 345441 82626 345751
rect 82308 345437 82626 345441
rect 85308 345751 85626 345755
rect 85308 345441 85312 345751
rect 85312 345441 85622 345751
rect 85622 345441 85626 345751
rect 85308 345437 85626 345441
rect 88308 345751 88626 345755
rect 88308 345441 88312 345751
rect 88312 345441 88622 345751
rect 88622 345441 88626 345751
rect 88308 345437 88626 345441
rect 91308 345751 91626 345755
rect 91308 345441 91312 345751
rect 91312 345441 91622 345751
rect 91622 345441 91626 345751
rect 91308 345437 91626 345441
rect 94308 345751 94626 345755
rect 94308 345441 94312 345751
rect 94312 345441 94622 345751
rect 94622 345441 94626 345751
rect 94308 345437 94626 345441
rect 97308 345751 97626 345755
rect 97308 345441 97312 345751
rect 97312 345441 97622 345751
rect 97622 345441 97626 345751
rect 97308 345437 97626 345441
rect 100308 345751 100626 345755
rect 100308 345441 100312 345751
rect 100312 345441 100622 345751
rect 100622 345441 100626 345751
rect 100308 345437 100626 345441
rect 103308 345751 103626 345755
rect 103308 345441 103312 345751
rect 103312 345441 103622 345751
rect 103622 345441 103626 345751
rect 103308 345437 103626 345441
rect 106308 345751 106626 345755
rect 106308 345441 106312 345751
rect 106312 345441 106622 345751
rect 106622 345441 106626 345751
rect 106308 345437 106626 345441
rect 109308 345751 109626 345755
rect 109308 345441 109312 345751
rect 109312 345441 109622 345751
rect 109622 345441 109626 345751
rect 109308 345437 109626 345441
rect 112308 345751 112626 345755
rect 112308 345441 112312 345751
rect 112312 345441 112622 345751
rect 112622 345441 112626 345751
rect 112308 345437 112626 345441
rect 115308 345751 115626 345755
rect 115308 345441 115312 345751
rect 115312 345441 115622 345751
rect 115622 345441 115626 345751
rect 115308 345437 115626 345441
rect 118308 345751 118626 345755
rect 118308 345441 118312 345751
rect 118312 345441 118622 345751
rect 118622 345441 118626 345751
rect 118308 345437 118626 345441
rect 121308 345751 121626 345755
rect 121308 345441 121312 345751
rect 121312 345441 121622 345751
rect 121622 345441 121626 345751
rect 121308 345437 121626 345441
rect 124308 345751 124626 345755
rect 124308 345441 124312 345751
rect 124312 345441 124622 345751
rect 124622 345441 124626 345751
rect 124308 345437 124626 345441
rect 127308 345751 127626 345755
rect 127308 345441 127312 345751
rect 127312 345441 127622 345751
rect 127622 345441 127626 345751
rect 127308 345437 127626 345441
rect 130308 345751 130626 345755
rect 130308 345441 130312 345751
rect 130312 345441 130622 345751
rect 130622 345441 130626 345751
rect 130308 345437 130626 345441
rect 133308 345751 133626 345755
rect 133308 345441 133312 345751
rect 133312 345441 133622 345751
rect 133622 345441 133626 345751
rect 133308 345437 133626 345441
rect 136308 345751 136626 345755
rect 136308 345441 136312 345751
rect 136312 345441 136622 345751
rect 136622 345441 136626 345751
rect 136308 345437 136626 345441
rect 139308 345751 139626 345755
rect 139308 345441 139312 345751
rect 139312 345441 139622 345751
rect 139622 345441 139626 345751
rect 139308 345437 139626 345441
rect 142308 345751 142626 345755
rect 142308 345441 142312 345751
rect 142312 345441 142622 345751
rect 142622 345441 142626 345751
rect 142308 345437 142626 345441
rect 145308 345751 145626 345755
rect 145308 345441 145312 345751
rect 145312 345441 145622 345751
rect 145622 345441 145626 345751
rect 145308 345437 145626 345441
rect 148308 345751 148626 345755
rect 148308 345441 148312 345751
rect 148312 345441 148622 345751
rect 148622 345441 148626 345751
rect 148308 345437 148626 345441
rect 151308 345751 151626 345755
rect 151308 345441 151312 345751
rect 151312 345441 151622 345751
rect 151622 345441 151626 345751
rect 151308 345437 151626 345441
rect 154308 345751 154626 345755
rect 154308 345441 154312 345751
rect 154312 345441 154622 345751
rect 154622 345441 154626 345751
rect 154308 345437 154626 345441
rect 157308 345751 157626 345755
rect 157308 345441 157312 345751
rect 157312 345441 157622 345751
rect 157622 345441 157626 345751
rect 157308 345437 157626 345441
rect 160308 345751 160626 345755
rect 160308 345441 160312 345751
rect 160312 345441 160622 345751
rect 160622 345441 160626 345751
rect 160308 345437 160626 345441
rect 163308 345751 163626 345755
rect 163308 345441 163312 345751
rect 163312 345441 163622 345751
rect 163622 345441 163626 345751
rect 163308 345437 163626 345441
rect 166308 345751 166626 345755
rect 166308 345441 166312 345751
rect 166312 345441 166622 345751
rect 166622 345441 166626 345751
rect 166308 345437 166626 345441
rect 169308 345751 169626 345755
rect 169308 345441 169312 345751
rect 169312 345441 169622 345751
rect 169622 345441 169626 345751
rect 169308 345437 169626 345441
rect 172308 345751 172626 345755
rect 172308 345441 172312 345751
rect 172312 345441 172622 345751
rect 172622 345441 172626 345751
rect 172308 345437 172626 345441
rect 175308 345751 175626 345755
rect 175308 345441 175312 345751
rect 175312 345441 175622 345751
rect 175622 345441 175626 345751
rect 175308 345437 175626 345441
rect 178308 345751 178626 345755
rect 178308 345441 178312 345751
rect 178312 345441 178622 345751
rect 178622 345441 178626 345751
rect 178308 345437 178626 345441
rect 181308 345751 181626 345755
rect 181308 345441 181312 345751
rect 181312 345441 181622 345751
rect 181622 345441 181626 345751
rect 181308 345437 181626 345441
rect 184308 345751 184626 345755
rect 184308 345441 184312 345751
rect 184312 345441 184622 345751
rect 184622 345441 184626 345751
rect 184308 345437 184626 345441
rect 187308 345751 187626 345755
rect 187308 345441 187312 345751
rect 187312 345441 187622 345751
rect 187622 345441 187626 345751
rect 187308 345437 187626 345441
rect 190308 345751 190626 345755
rect 190308 345441 190312 345751
rect 190312 345441 190622 345751
rect 190622 345441 190626 345751
rect 190308 345437 190626 345441
rect 193308 345751 193626 345755
rect 193308 345441 193312 345751
rect 193312 345441 193622 345751
rect 193622 345441 193626 345751
rect 193308 345437 193626 345441
rect 196308 345751 196626 345755
rect 196308 345441 196312 345751
rect 196312 345441 196622 345751
rect 196622 345441 196626 345751
rect 196308 345437 196626 345441
rect 199308 345751 199626 345755
rect 199308 345441 199312 345751
rect 199312 345441 199622 345751
rect 199622 345441 199626 345751
rect 199308 345437 199626 345441
rect 202308 345751 202626 345755
rect 202308 345441 202312 345751
rect 202312 345441 202622 345751
rect 202622 345441 202626 345751
rect 202308 345437 202626 345441
rect 205308 345751 205626 345755
rect 205308 345441 205312 345751
rect 205312 345441 205622 345751
rect 205622 345441 205626 345751
rect 205308 345437 205626 345441
rect 208308 345751 208626 345755
rect 208308 345441 208312 345751
rect 208312 345441 208622 345751
rect 208622 345441 208626 345751
rect 208308 345437 208626 345441
rect 211308 345751 211626 345755
rect 211308 345441 211312 345751
rect 211312 345441 211622 345751
rect 211622 345441 211626 345751
rect 211308 345437 211626 345441
rect 214308 345751 214626 345755
rect 214308 345441 214312 345751
rect 214312 345441 214622 345751
rect 214622 345441 214626 345751
rect 214308 345437 214626 345441
rect 217308 345751 217626 345755
rect 217308 345441 217312 345751
rect 217312 345441 217622 345751
rect 217622 345441 217626 345751
rect 217308 345437 217626 345441
rect 220308 345751 220626 345755
rect 220308 345441 220312 345751
rect 220312 345441 220622 345751
rect 220622 345441 220626 345751
rect 220308 345437 220626 345441
rect 223308 345751 223626 345755
rect 223308 345441 223312 345751
rect 223312 345441 223622 345751
rect 223622 345441 223626 345751
rect 223308 345437 223626 345441
rect 226308 345751 226626 345755
rect 226308 345441 226312 345751
rect 226312 345441 226622 345751
rect 226622 345441 226626 345751
rect 226308 345437 226626 345441
rect 229308 345751 229626 345755
rect 229308 345441 229312 345751
rect 229312 345441 229622 345751
rect 229622 345441 229626 345751
rect 229308 345437 229626 345441
rect 232308 345751 232626 345755
rect 232308 345441 232312 345751
rect 232312 345441 232622 345751
rect 232622 345441 232626 345751
rect 232308 345437 232626 345441
rect 235308 345751 235626 345755
rect 235308 345441 235312 345751
rect 235312 345441 235622 345751
rect 235622 345441 235626 345751
rect 235308 345437 235626 345441
rect 238308 345751 238626 345755
rect 238308 345441 238312 345751
rect 238312 345441 238622 345751
rect 238622 345441 238626 345751
rect 238308 345437 238626 345441
rect 241308 345751 241626 345755
rect 241308 345441 241312 345751
rect 241312 345441 241622 345751
rect 241622 345441 241626 345751
rect 241308 345437 241626 345441
rect 244308 345751 244626 345755
rect 244308 345441 244312 345751
rect 244312 345441 244622 345751
rect 244622 345441 244626 345751
rect 244308 345437 244626 345441
rect 247308 345751 247626 345755
rect 247308 345441 247312 345751
rect 247312 345441 247622 345751
rect 247622 345441 247626 345751
rect 247308 345437 247626 345441
rect 250308 345751 250626 345755
rect 250308 345441 250312 345751
rect 250312 345441 250622 345751
rect 250622 345441 250626 345751
rect 250308 345437 250626 345441
rect 253308 345751 253626 345755
rect 253308 345441 253312 345751
rect 253312 345441 253622 345751
rect 253622 345441 253626 345751
rect 253308 345437 253626 345441
rect 256308 345751 256626 345755
rect 256308 345441 256312 345751
rect 256312 345441 256622 345751
rect 256622 345441 256626 345751
rect 256308 345437 256626 345441
rect 259308 345751 259626 345755
rect 259308 345441 259312 345751
rect 259312 345441 259622 345751
rect 259622 345441 259626 345751
rect 259308 345437 259626 345441
rect 262308 345751 262626 345755
rect 262308 345441 262312 345751
rect 262312 345441 262622 345751
rect 262622 345441 262626 345751
rect 262308 345437 262626 345441
rect 265308 345751 265626 345755
rect 265308 345441 265312 345751
rect 265312 345441 265622 345751
rect 265622 345441 265626 345751
rect 265308 345437 265626 345441
rect 268308 345751 268626 345755
rect 268308 345441 268312 345751
rect 268312 345441 268622 345751
rect 268622 345441 268626 345751
rect 268308 345437 268626 345441
rect 271308 345751 271626 345755
rect 271308 345441 271312 345751
rect 271312 345441 271622 345751
rect 271622 345441 271626 345751
rect 271308 345437 271626 345441
rect 274308 345751 274626 345755
rect 274308 345441 274312 345751
rect 274312 345441 274622 345751
rect 274622 345441 274626 345751
rect 274308 345437 274626 345441
rect 277308 345751 277626 345755
rect 277308 345441 277312 345751
rect 277312 345441 277622 345751
rect 277622 345441 277626 345751
rect 277308 345437 277626 345441
rect 280308 345751 280626 345755
rect 280308 345441 280312 345751
rect 280312 345441 280622 345751
rect 280622 345441 280626 345751
rect 280308 345437 280626 345441
rect 283308 345751 283626 345755
rect 283308 345441 283312 345751
rect 283312 345441 283622 345751
rect 283622 345441 283626 345751
rect 283308 345437 283626 345441
rect 286308 345751 286626 345755
rect 286308 345441 286312 345751
rect 286312 345441 286622 345751
rect 286622 345441 286626 345751
rect 286308 345437 286626 345441
rect 289308 345751 289626 345755
rect 289308 345441 289312 345751
rect 289312 345441 289622 345751
rect 289622 345441 289626 345751
rect 289308 345437 289626 345441
rect 292308 345751 292626 345755
rect 292308 345441 292312 345751
rect 292312 345441 292622 345751
rect 292622 345441 292626 345751
rect 292308 345437 292626 345441
rect 295308 345751 295626 345755
rect 295308 345441 295312 345751
rect 295312 345441 295622 345751
rect 295622 345441 295626 345751
rect 295308 345437 295626 345441
rect 298308 345751 298626 345755
rect 298308 345441 298312 345751
rect 298312 345441 298622 345751
rect 298622 345441 298626 345751
rect 298308 345437 298626 345441
rect 301308 345751 301626 345755
rect 301308 345441 301312 345751
rect 301312 345441 301622 345751
rect 301622 345441 301626 345751
rect 301308 345437 301626 345441
rect 304308 345751 304626 345755
rect 304308 345441 304312 345751
rect 304312 345441 304622 345751
rect 304622 345441 304626 345751
rect 304308 345437 304626 345441
rect 307308 345751 307626 345755
rect 307308 345441 307312 345751
rect 307312 345441 307622 345751
rect 307622 345441 307626 345751
rect 307308 345437 307626 345441
rect 310308 345751 310626 345755
rect 310308 345441 310312 345751
rect 310312 345441 310622 345751
rect 310622 345441 310626 345751
rect 310308 345437 310626 345441
rect 313308 345751 313626 345755
rect 313308 345441 313312 345751
rect 313312 345441 313622 345751
rect 313622 345441 313626 345751
rect 313308 345437 313626 345441
rect 316308 345751 316626 345755
rect 316308 345441 316312 345751
rect 316312 345441 316622 345751
rect 316622 345441 316626 345751
rect 316308 345437 316626 345441
rect 319308 345751 319626 345755
rect 319308 345441 319312 345751
rect 319312 345441 319622 345751
rect 319622 345441 319626 345751
rect 319308 345437 319626 345441
rect 325308 345751 325626 345755
rect 325308 345441 325312 345751
rect 325312 345441 325622 345751
rect 325622 345441 325626 345751
rect 325308 345437 325626 345441
rect 328308 345751 328626 345755
rect 328308 345441 328312 345751
rect 328312 345441 328622 345751
rect 328622 345441 328626 345751
rect 328308 345437 328626 345441
rect 331308 345751 331626 345755
rect 331308 345441 331312 345751
rect 331312 345441 331622 345751
rect 331622 345441 331626 345751
rect 331308 345437 331626 345441
rect 334308 345751 334626 345755
rect 334308 345441 334312 345751
rect 334312 345441 334622 345751
rect 334622 345441 334626 345751
rect 334308 345437 334626 345441
rect 337308 345751 337626 345755
rect 337308 345441 337312 345751
rect 337312 345441 337622 345751
rect 337622 345441 337626 345751
rect 337308 345437 337626 345441
rect 340308 345751 340626 345755
rect 340308 345441 340312 345751
rect 340312 345441 340622 345751
rect 340622 345441 340626 345751
rect 340308 345437 340626 345441
rect 343308 345751 343626 345755
rect 343308 345441 343312 345751
rect 343312 345441 343622 345751
rect 343622 345441 343626 345751
rect 343308 345437 343626 345441
rect 346308 345751 346626 345755
rect 346308 345441 346312 345751
rect 346312 345441 346622 345751
rect 346622 345441 346626 345751
rect 346308 345437 346626 345441
rect 349308 345751 349626 345755
rect 349308 345441 349312 345751
rect 349312 345441 349622 345751
rect 349622 345441 349626 345751
rect 349308 345437 349626 345441
rect 352308 345751 352626 345755
rect 352308 345441 352312 345751
rect 352312 345441 352622 345751
rect 352622 345441 352626 345751
rect 352308 345437 352626 345441
rect 355308 345751 355626 345755
rect 355308 345441 355312 345751
rect 355312 345441 355622 345751
rect 355622 345441 355626 345751
rect 355308 345437 355626 345441
rect 358308 345751 358626 345755
rect 358308 345441 358312 345751
rect 358312 345441 358622 345751
rect 358622 345441 358626 345751
rect 358308 345437 358626 345441
rect 372486 336904 372786 336909
rect 372486 336604 372781 336904
rect 372781 336604 372786 336904
rect 372486 336599 372786 336604
rect 375486 336904 375786 336909
rect 375486 336604 375781 336904
rect 375781 336604 375786 336904
rect 375486 336599 375786 336604
rect 378486 336904 378786 336909
rect 378486 336604 378781 336904
rect 378781 336604 378786 336904
rect 378486 336599 378786 336604
rect 381486 336904 381786 336909
rect 381486 336604 381781 336904
rect 381781 336604 381786 336904
rect 381486 336599 381786 336604
rect 384486 336904 384786 336909
rect 384486 336604 384781 336904
rect 384781 336604 384786 336904
rect 384486 336599 384786 336604
rect 387486 336904 387786 336909
rect 387486 336604 387781 336904
rect 387781 336604 387786 336904
rect 387486 336599 387786 336604
rect 390486 336904 390786 336909
rect 390486 336604 390781 336904
rect 390781 336604 390786 336904
rect 390486 336599 390786 336604
rect 393486 336904 393786 336909
rect 393486 336604 393781 336904
rect 393781 336604 393786 336904
rect 393486 336599 393786 336604
rect 396486 336904 396786 336909
rect 396486 336604 396781 336904
rect 396781 336604 396786 336904
rect 396486 336599 396786 336604
rect 55302 323107 55307 323422
rect 55307 323107 55627 323422
rect 55627 323107 55632 323422
rect 55302 323102 55632 323107
rect 58302 323107 58307 323422
rect 58307 323107 58627 323422
rect 58627 323107 58632 323422
rect 58302 323102 58632 323107
rect 61302 323107 61307 323422
rect 61307 323107 61627 323422
rect 61627 323107 61632 323422
rect 61302 323102 61632 323107
rect 64302 323107 64307 323422
rect 64307 323107 64627 323422
rect 64627 323107 64632 323422
rect 64302 323102 64632 323107
rect 67302 323107 67307 323422
rect 67307 323107 67627 323422
rect 67627 323107 67632 323422
rect 67302 323102 67632 323107
rect 70302 323107 70307 323422
rect 70307 323107 70627 323422
rect 70627 323107 70632 323422
rect 70302 323102 70632 323107
rect 73302 323107 73307 323422
rect 73307 323107 73627 323422
rect 73627 323107 73632 323422
rect 73302 323102 73632 323107
rect 76302 323107 76307 323422
rect 76307 323107 76627 323422
rect 76627 323107 76632 323422
rect 76302 323102 76632 323107
rect 79302 323107 79307 323422
rect 79307 323107 79627 323422
rect 79627 323107 79632 323422
rect 79302 323102 79632 323107
rect 82302 323107 82307 323422
rect 82307 323107 82627 323422
rect 82627 323107 82632 323422
rect 82302 323102 82632 323107
rect 85302 323107 85307 323422
rect 85307 323107 85627 323422
rect 85627 323107 85632 323422
rect 85302 323102 85632 323107
rect 88302 323107 88307 323422
rect 88307 323107 88627 323422
rect 88627 323107 88632 323422
rect 88302 323102 88632 323107
rect 91302 323107 91307 323422
rect 91307 323107 91627 323422
rect 91627 323107 91632 323422
rect 91302 323102 91632 323107
rect 94302 323107 94307 323422
rect 94307 323107 94627 323422
rect 94627 323107 94632 323422
rect 94302 323102 94632 323107
rect 97302 323107 97307 323422
rect 97307 323107 97627 323422
rect 97627 323107 97632 323422
rect 97302 323102 97632 323107
rect 100302 323107 100307 323422
rect 100307 323107 100627 323422
rect 100627 323107 100632 323422
rect 100302 323102 100632 323107
rect 103302 323107 103307 323422
rect 103307 323107 103627 323422
rect 103627 323107 103632 323422
rect 103302 323102 103632 323107
rect 106302 323107 106307 323422
rect 106307 323107 106627 323422
rect 106627 323107 106632 323422
rect 106302 323102 106632 323107
rect 109302 323107 109307 323422
rect 109307 323107 109627 323422
rect 109627 323107 109632 323422
rect 109302 323102 109632 323107
rect 112302 323107 112307 323422
rect 112307 323107 112627 323422
rect 112627 323107 112632 323422
rect 112302 323102 112632 323107
rect 115302 323107 115307 323422
rect 115307 323107 115627 323422
rect 115627 323107 115632 323422
rect 115302 323102 115632 323107
rect 118302 323107 118307 323422
rect 118307 323107 118627 323422
rect 118627 323107 118632 323422
rect 118302 323102 118632 323107
rect 121302 323107 121307 323422
rect 121307 323107 121627 323422
rect 121627 323107 121632 323422
rect 121302 323102 121632 323107
rect 124302 323107 124307 323422
rect 124307 323107 124627 323422
rect 124627 323107 124632 323422
rect 124302 323102 124632 323107
rect 127302 323107 127307 323422
rect 127307 323107 127627 323422
rect 127627 323107 127632 323422
rect 127302 323102 127632 323107
rect 130302 323107 130307 323422
rect 130307 323107 130627 323422
rect 130627 323107 130632 323422
rect 130302 323102 130632 323107
rect 133302 323107 133307 323422
rect 133307 323107 133627 323422
rect 133627 323107 133632 323422
rect 133302 323102 133632 323107
rect 136302 323107 136307 323422
rect 136307 323107 136627 323422
rect 136627 323107 136632 323422
rect 136302 323102 136632 323107
rect 139302 323107 139307 323422
rect 139307 323107 139627 323422
rect 139627 323107 139632 323422
rect 139302 323102 139632 323107
rect 142302 323107 142307 323422
rect 142307 323107 142627 323422
rect 142627 323107 142632 323422
rect 142302 323102 142632 323107
rect 145302 323107 145307 323422
rect 145307 323107 145627 323422
rect 145627 323107 145632 323422
rect 145302 323102 145632 323107
rect 148302 323107 148307 323422
rect 148307 323107 148627 323422
rect 148627 323107 148632 323422
rect 148302 323102 148632 323107
rect 151302 323107 151307 323422
rect 151307 323107 151627 323422
rect 151627 323107 151632 323422
rect 151302 323102 151632 323107
rect 154302 323107 154307 323422
rect 154307 323107 154627 323422
rect 154627 323107 154632 323422
rect 154302 323102 154632 323107
rect 157302 323107 157307 323422
rect 157307 323107 157627 323422
rect 157627 323107 157632 323422
rect 157302 323102 157632 323107
rect 160302 323107 160307 323422
rect 160307 323107 160627 323422
rect 160627 323107 160632 323422
rect 160302 323102 160632 323107
rect 163302 323107 163307 323422
rect 163307 323107 163627 323422
rect 163627 323107 163632 323422
rect 163302 323102 163632 323107
rect 166302 323107 166307 323422
rect 166307 323107 166627 323422
rect 166627 323107 166632 323422
rect 166302 323102 166632 323107
rect 169302 323107 169307 323422
rect 169307 323107 169627 323422
rect 169627 323107 169632 323422
rect 169302 323102 169632 323107
rect 172302 323107 172307 323422
rect 172307 323107 172627 323422
rect 172627 323107 172632 323422
rect 172302 323102 172632 323107
rect 175302 323107 175307 323422
rect 175307 323107 175627 323422
rect 175627 323107 175632 323422
rect 175302 323102 175632 323107
rect 178302 323107 178307 323422
rect 178307 323107 178627 323422
rect 178627 323107 178632 323422
rect 178302 323102 178632 323107
rect 181302 323107 181307 323422
rect 181307 323107 181627 323422
rect 181627 323107 181632 323422
rect 181302 323102 181632 323107
rect 184302 323107 184307 323422
rect 184307 323107 184627 323422
rect 184627 323107 184632 323422
rect 184302 323102 184632 323107
rect 187302 323107 187307 323422
rect 187307 323107 187627 323422
rect 187627 323107 187632 323422
rect 187302 323102 187632 323107
rect 190302 323107 190307 323422
rect 190307 323107 190627 323422
rect 190627 323107 190632 323422
rect 190302 323102 190632 323107
rect 193302 323107 193307 323422
rect 193307 323107 193627 323422
rect 193627 323107 193632 323422
rect 193302 323102 193632 323107
rect 196302 323107 196307 323422
rect 196307 323107 196627 323422
rect 196627 323107 196632 323422
rect 196302 323102 196632 323107
rect 199302 323107 199307 323422
rect 199307 323107 199627 323422
rect 199627 323107 199632 323422
rect 199302 323102 199632 323107
rect 202302 323107 202307 323422
rect 202307 323107 202627 323422
rect 202627 323107 202632 323422
rect 202302 323102 202632 323107
rect 205302 323107 205307 323422
rect 205307 323107 205627 323422
rect 205627 323107 205632 323422
rect 205302 323102 205632 323107
rect 208302 323107 208307 323422
rect 208307 323107 208627 323422
rect 208627 323107 208632 323422
rect 208302 323102 208632 323107
rect 211302 323107 211307 323422
rect 211307 323107 211627 323422
rect 211627 323107 211632 323422
rect 211302 323102 211632 323107
rect 214302 323107 214307 323422
rect 214307 323107 214627 323422
rect 214627 323107 214632 323422
rect 214302 323102 214632 323107
rect 217302 323107 217307 323422
rect 217307 323107 217627 323422
rect 217627 323107 217632 323422
rect 217302 323102 217632 323107
rect 220302 323107 220307 323422
rect 220307 323107 220627 323422
rect 220627 323107 220632 323422
rect 220302 323102 220632 323107
rect 223302 323107 223307 323422
rect 223307 323107 223627 323422
rect 223627 323107 223632 323422
rect 223302 323102 223632 323107
rect 226302 323107 226307 323422
rect 226307 323107 226627 323422
rect 226627 323107 226632 323422
rect 226302 323102 226632 323107
rect 229302 323107 229307 323422
rect 229307 323107 229627 323422
rect 229627 323107 229632 323422
rect 229302 323102 229632 323107
rect 232302 323107 232307 323422
rect 232307 323107 232627 323422
rect 232627 323107 232632 323422
rect 232302 323102 232632 323107
rect 235302 323107 235307 323422
rect 235307 323107 235627 323422
rect 235627 323107 235632 323422
rect 235302 323102 235632 323107
rect 238302 323107 238307 323422
rect 238307 323107 238627 323422
rect 238627 323107 238632 323422
rect 238302 323102 238632 323107
rect 241302 323107 241307 323422
rect 241307 323107 241627 323422
rect 241627 323107 241632 323422
rect 241302 323102 241632 323107
rect 244302 323107 244307 323422
rect 244307 323107 244627 323422
rect 244627 323107 244632 323422
rect 244302 323102 244632 323107
rect 247302 323107 247307 323422
rect 247307 323107 247627 323422
rect 247627 323107 247632 323422
rect 247302 323102 247632 323107
rect 250302 323107 250307 323422
rect 250307 323107 250627 323422
rect 250627 323107 250632 323422
rect 250302 323102 250632 323107
rect 253302 323107 253307 323422
rect 253307 323107 253627 323422
rect 253627 323107 253632 323422
rect 253302 323102 253632 323107
rect 256302 323107 256307 323422
rect 256307 323107 256627 323422
rect 256627 323107 256632 323422
rect 256302 323102 256632 323107
rect 259302 323107 259307 323422
rect 259307 323107 259627 323422
rect 259627 323107 259632 323422
rect 259302 323102 259632 323107
rect 262302 323107 262307 323422
rect 262307 323107 262627 323422
rect 262627 323107 262632 323422
rect 262302 323102 262632 323107
rect 265302 323107 265307 323422
rect 265307 323107 265627 323422
rect 265627 323107 265632 323422
rect 265302 323102 265632 323107
rect 268302 323107 268307 323422
rect 268307 323107 268627 323422
rect 268627 323107 268632 323422
rect 268302 323102 268632 323107
rect 271302 323107 271307 323422
rect 271307 323107 271627 323422
rect 271627 323107 271632 323422
rect 271302 323102 271632 323107
rect 274302 323107 274307 323422
rect 274307 323107 274627 323422
rect 274627 323107 274632 323422
rect 274302 323102 274632 323107
rect 277302 323107 277307 323422
rect 277307 323107 277627 323422
rect 277627 323107 277632 323422
rect 277302 323102 277632 323107
rect 280302 323107 280307 323422
rect 280307 323107 280627 323422
rect 280627 323107 280632 323422
rect 280302 323102 280632 323107
rect 283302 323107 283307 323422
rect 283307 323107 283627 323422
rect 283627 323107 283632 323422
rect 283302 323102 283632 323107
rect 286302 323107 286307 323422
rect 286307 323107 286627 323422
rect 286627 323107 286632 323422
rect 286302 323102 286632 323107
rect 289302 323107 289307 323422
rect 289307 323107 289627 323422
rect 289627 323107 289632 323422
rect 289302 323102 289632 323107
rect 292302 323107 292307 323422
rect 292307 323107 292627 323422
rect 292627 323107 292632 323422
rect 292302 323102 292632 323107
rect 295302 323107 295307 323422
rect 295307 323107 295627 323422
rect 295627 323107 295632 323422
rect 295302 323102 295632 323107
rect 298302 323107 298307 323422
rect 298307 323107 298627 323422
rect 298627 323107 298632 323422
rect 298302 323102 298632 323107
rect 301302 323107 301307 323422
rect 301307 323107 301627 323422
rect 301627 323107 301632 323422
rect 301302 323102 301632 323107
rect 304302 323107 304307 323422
rect 304307 323107 304627 323422
rect 304627 323107 304632 323422
rect 304302 323102 304632 323107
rect 307302 323107 307307 323422
rect 307307 323107 307627 323422
rect 307627 323107 307632 323422
rect 307302 323102 307632 323107
rect 310302 323107 310307 323422
rect 310307 323107 310627 323422
rect 310627 323107 310632 323422
rect 310302 323102 310632 323107
rect 313302 323107 313307 323422
rect 313307 323107 313627 323422
rect 313627 323107 313632 323422
rect 313302 323102 313632 323107
rect 316302 323107 316307 323422
rect 316307 323107 316627 323422
rect 316627 323107 316632 323422
rect 316302 323102 316632 323107
rect 319302 323107 319307 323422
rect 319307 323107 319627 323422
rect 319627 323107 319632 323422
rect 319302 323102 319632 323107
rect 325302 323107 325307 323422
rect 325307 323107 325627 323422
rect 325627 323107 325632 323422
rect 325302 323102 325632 323107
rect 328302 323107 328307 323422
rect 328307 323107 328627 323422
rect 328627 323107 328632 323422
rect 328302 323102 328632 323107
rect 331302 323107 331307 323422
rect 331307 323107 331627 323422
rect 331627 323107 331632 323422
rect 331302 323102 331632 323107
rect 334302 323107 334307 323422
rect 334307 323107 334627 323422
rect 334627 323107 334632 323422
rect 334302 323102 334632 323107
rect 337302 323107 337307 323422
rect 337307 323107 337627 323422
rect 337627 323107 337632 323422
rect 337302 323102 337632 323107
rect 340302 323107 340307 323422
rect 340307 323107 340627 323422
rect 340627 323107 340632 323422
rect 340302 323102 340632 323107
rect 343302 323107 343307 323422
rect 343307 323107 343627 323422
rect 343627 323107 343632 323422
rect 343302 323102 343632 323107
rect 346302 323107 346307 323422
rect 346307 323107 346627 323422
rect 346627 323107 346632 323422
rect 346302 323102 346632 323107
rect 349302 323107 349307 323422
rect 349307 323107 349627 323422
rect 349627 323107 349632 323422
rect 349302 323102 349632 323107
rect 352302 323107 352307 323422
rect 352307 323107 352627 323422
rect 352627 323107 352632 323422
rect 352302 323102 352632 323107
rect 355302 323107 355307 323422
rect 355307 323107 355627 323422
rect 355627 323107 355632 323422
rect 355302 323102 355632 323107
rect 358302 323107 358307 323422
rect 358307 323107 358627 323422
rect 358627 323107 358632 323422
rect 358302 323102 358632 323107
rect 424844 313911 425014 314081
rect 69648 253686 69968 254006
rect 5661 253062 5771 253172
rect 12507 253061 12619 253173
rect 7127 243630 7217 243720
rect 167888 206836 168208 207156
rect 170812 207060 171132 207380
rect 173402 207178 173722 207498
rect 167889 191868 168207 192186
rect 170813 191868 171131 192186
rect 173403 191868 173721 192186
rect 10674 191427 10784 191537
rect 33445 191428 33553 191536
rect 9011 191337 9131 191342
rect 9011 191232 9016 191337
rect 9016 191232 9126 191337
rect 9126 191232 9131 191337
rect 287965 230745 290423 230749
rect 287965 228295 287969 230745
rect 287969 228295 290419 230745
rect 290419 228295 290423 230745
rect 287965 228291 290423 228295
rect 180916 207290 181216 207295
rect 180916 207005 180921 207290
rect 180921 207005 181211 207290
rect 181211 207005 181216 207290
rect 183916 207290 184216 207295
rect 183916 207005 183921 207290
rect 183921 207005 184211 207290
rect 184211 207005 184216 207290
rect 186916 207290 187216 207295
rect 186916 207005 186921 207290
rect 186921 207005 187211 207290
rect 187211 207005 187216 207290
rect 189916 207290 190216 207295
rect 189916 207005 189921 207290
rect 189921 207005 190211 207290
rect 190211 207005 190216 207290
rect 192916 207290 193216 207295
rect 192916 207005 192921 207290
rect 192921 207005 193211 207290
rect 193211 207005 193216 207290
rect 195916 207290 196216 207295
rect 195916 207005 195921 207290
rect 195921 207005 196211 207290
rect 196211 207005 196216 207290
rect 198916 207290 199216 207295
rect 198916 207005 198921 207290
rect 198921 207005 199211 207290
rect 199211 207005 199216 207290
rect 201916 207290 202216 207295
rect 201916 207005 201921 207290
rect 201921 207005 202211 207290
rect 202211 207005 202216 207290
rect 204916 207290 205216 207295
rect 204916 207005 204921 207290
rect 204921 207005 205211 207290
rect 205211 207005 205216 207290
rect 175759 186467 175764 186632
rect 175764 186467 175934 186632
rect 175934 186467 175939 186632
rect 175759 186462 175939 186467
rect 164432 180308 164750 180626
rect 167773 180308 168091 180626
rect 170723 180308 171041 180626
rect 173033 180308 173351 180626
rect 175009 180308 175327 180626
rect 3527 164594 12521 176552
rect 15357 172310 15577 172530
rect 52330 172311 52548 172529
rect 86589 166636 89049 169096
rect 164431 167996 164751 168316
rect 170722 168209 171042 168529
rect 180872 172519 180877 172814
rect 180877 172519 181177 172814
rect 181177 172519 181182 172814
rect 180872 172514 181182 172519
rect 183872 172519 183877 172814
rect 183877 172519 184177 172814
rect 184177 172519 184182 172814
rect 183872 172514 184182 172519
rect 186872 172519 186877 172814
rect 186877 172519 187177 172814
rect 187177 172519 187182 172814
rect 186872 172514 187182 172519
rect 189872 172519 189877 172814
rect 189877 172519 190177 172814
rect 190177 172519 190182 172814
rect 189872 172514 190182 172519
rect 192872 172519 192877 172814
rect 192877 172519 193177 172814
rect 193177 172519 193182 172814
rect 192872 172514 193182 172519
rect 195872 172519 195877 172814
rect 195877 172519 196177 172814
rect 196177 172519 196182 172814
rect 195872 172514 196182 172519
rect 198872 172519 198877 172814
rect 198877 172519 199177 172814
rect 199177 172519 199182 172814
rect 198872 172514 199182 172519
rect 201872 172519 201877 172814
rect 201877 172519 202177 172814
rect 202177 172519 202182 172814
rect 201872 172514 202182 172519
rect 204872 172519 204877 172814
rect 204877 172519 205177 172814
rect 205177 172519 205182 172814
rect 204872 172514 205182 172519
rect 167772 167854 168092 168174
rect 173032 167925 173352 168245
rect 175008 167925 175328 168245
rect 86444 162888 88904 165348
rect 86722 151994 89182 154454
rect 13381 144774 15841 147234
rect 13382 134050 15840 136508
rect 86722 134049 89182 136509
rect 287959 116498 287964 118953
rect 287964 116498 290424 118953
rect 290424 116498 290429 118953
rect 287959 116493 290429 116498
rect 573845 217336 578645 222136
rect 574269 199257 579069 204057
rect 502080 193890 504540 196230
rect 502080 193770 504562 193890
rect 502102 191430 504562 193770
rect 502391 183890 504851 186230
rect 502391 183770 505015 183890
rect 502555 181430 505015 183770
rect 573845 162676 578645 167476
rect 501821 146887 504281 149347
rect 502044 136830 504504 139290
rect 40357 34786 40469 34898
rect 46643 13364 46755 13476
rect 354 3908 466 4020
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 703788 334294 704800
rect 329294 702300 329837 703788
rect 329590 700672 329837 702300
rect 333913 702300 334294 703788
rect 333913 700672 334190 702300
rect 329590 700390 334190 700672
rect 229190 699708 231180 699960
rect 229190 698530 229597 699708
rect 228350 698529 229597 698530
rect 228350 697491 228439 698529
rect 229477 697552 229597 698529
rect 229477 697491 231180 697552
rect 228350 697490 231180 697491
rect 229190 697460 231180 697490
rect 331191 698285 332129 700390
rect 331191 697349 331192 698285
rect 332128 697349 332129 698285
rect 331191 697042 332129 697349
rect 1919 686009 4379 694260
rect 143667 694000 143668 694001
rect 144068 694000 144069 694001
rect 143667 693999 144069 694000
rect 22110 692119 31923 692120
rect 22110 692011 22111 692119
rect 22219 692011 31923 692119
rect 22110 692010 31923 692011
rect 7012 688093 7332 688094
rect 7012 687775 7013 688093
rect 7331 687775 7332 688093
rect 7012 687774 7332 687775
rect 1919 683551 1920 686009
rect 4378 683551 4379 686009
rect 1919 678114 4379 683551
rect 1919 675656 1920 678114
rect 4378 675656 4379 678114
rect 1919 672892 4379 675656
rect 1919 670434 1920 672892
rect 4378 670434 4379 672892
rect 1919 353278 4379 670434
rect 1919 350820 1920 353278
rect 4378 350820 4379 353278
rect 1919 348749 4379 350820
rect 1919 346291 1920 348749
rect 4378 346291 4379 348749
rect 1919 344239 4379 346291
rect 1919 341781 1920 344239
rect 4378 341781 4379 344239
rect 1919 315914 4379 341781
rect 1919 313456 1920 315914
rect 4378 313456 4379 315914
rect 1919 177800 4379 313456
rect 8387 685552 28751 685553
rect 8387 685484 28682 685552
rect 28750 685484 28751 685552
rect 8387 685483 28751 685484
rect 5659 293381 5773 293382
rect 5659 293269 5660 293381
rect 5772 293269 5773 293381
rect 5659 293268 5773 293269
rect 5660 253172 5772 293268
rect 8387 261321 8457 685483
rect 26806 684469 26808 684470
rect 26806 681999 26807 684469
rect 26806 681998 26808 681999
rect 9016 680861 9126 680862
rect 9016 680753 9017 680861
rect 9125 680753 9126 680861
rect 8381 261320 8463 261321
rect 8381 261250 8382 261320
rect 8462 261250 8463 261320
rect 8381 261249 8463 261250
rect 5660 253062 5661 253172
rect 5771 253062 5772 253172
rect 5660 253061 5772 253062
rect 9016 191343 9126 680753
rect 26514 678120 26516 678121
rect 26514 675650 26515 678120
rect 26514 675649 26516 675650
rect 10674 675139 10784 675140
rect 10674 675031 10675 675139
rect 10783 675031 10784 675139
rect 10674 191538 10784 675031
rect 26347 672898 26349 672899
rect 26347 670428 26348 672898
rect 26347 670427 26349 670428
rect 19234 667765 19236 667766
rect 19235 667435 19236 667765
rect 19234 667434 19236 667435
rect 19234 664765 19236 664766
rect 19235 664435 19236 664765
rect 19234 664434 19236 664435
rect 19139 662310 19141 662311
rect 19140 661990 19141 662310
rect 19139 661989 19141 661990
rect 19234 661765 19236 661766
rect 19235 661435 19236 661765
rect 19234 661434 19236 661435
rect 19139 659310 19141 659311
rect 19140 658990 19141 659310
rect 19139 658989 19141 658990
rect 19234 658765 19236 658766
rect 19235 658435 19236 658765
rect 19234 658434 19236 658435
rect 13651 657331 13973 657332
rect 13651 657001 13652 657331
rect 13972 657001 13973 657331
rect 13651 657000 13973 657001
rect 19139 656310 19141 656311
rect 19140 655990 19141 656310
rect 19139 655989 19141 655990
rect 19234 655765 19236 655766
rect 19235 655435 19236 655765
rect 19234 655434 19236 655435
rect 19139 653310 19141 653311
rect 19140 652990 19141 653310
rect 19139 652989 19141 652990
rect 19234 652765 19236 652766
rect 19235 652435 19236 652765
rect 19234 652434 19236 652435
rect 19139 650310 19141 650311
rect 19140 649990 19141 650310
rect 19139 649989 19141 649990
rect 19234 649765 19236 649766
rect 19235 649435 19236 649765
rect 19234 649434 19236 649435
rect 19139 647310 19141 647311
rect 19140 646990 19141 647310
rect 19139 646989 19141 646990
rect 19234 646765 19236 646766
rect 19235 646435 19236 646765
rect 19234 646434 19236 646435
rect 19139 644310 19141 644311
rect 19140 643990 19141 644310
rect 19139 643989 19141 643990
rect 19234 643765 19236 643766
rect 19235 643435 19236 643765
rect 19234 643434 19236 643435
rect 19139 641310 19141 641311
rect 19140 640990 19141 641310
rect 19139 640989 19141 640990
rect 19234 640765 19236 640766
rect 19235 640435 19236 640765
rect 19234 640434 19236 640435
rect 19139 638310 19141 638311
rect 19140 637990 19141 638310
rect 19139 637989 19141 637990
rect 19234 637765 19236 637766
rect 19235 637435 19236 637765
rect 19234 637434 19236 637435
rect 19139 635310 19141 635311
rect 19140 634990 19141 635310
rect 19139 634989 19141 634990
rect 19234 634765 19236 634766
rect 19235 634435 19236 634765
rect 19234 634434 19236 634435
rect 19139 632310 19141 632311
rect 19140 631990 19141 632310
rect 19139 631989 19141 631990
rect 19234 631765 19236 631766
rect 19235 631435 19236 631765
rect 19234 631434 19236 631435
rect 11333 630293 13793 630294
rect 11333 627835 11334 630293
rect 13792 627835 13793 630293
rect 11333 627834 13793 627835
rect 19234 625765 19236 625766
rect 19235 625435 19236 625765
rect 19234 625434 19236 625435
rect 11077 624842 11079 624843
rect 11077 622087 11078 624842
rect 19139 623310 19141 623311
rect 19140 622990 19141 623310
rect 19139 622989 19141 622990
rect 19234 622765 19236 622766
rect 19235 622435 19236 622765
rect 19234 622434 19236 622435
rect 11077 622086 11079 622087
rect 19139 620310 19141 620311
rect 19140 619990 19141 620310
rect 19139 619989 19141 619990
rect 19234 619765 19236 619766
rect 19235 619435 19236 619765
rect 19234 619434 19236 619435
rect 19139 617310 19141 617311
rect 19140 616990 19141 617310
rect 19139 616989 19141 616990
rect 19234 616765 19236 616766
rect 19235 616435 19236 616765
rect 19234 616434 19236 616435
rect 15231 614713 15232 614714
rect 17987 614713 17988 614714
rect 15231 614712 17988 614713
rect 19139 614310 19141 614311
rect 19140 613990 19141 614310
rect 19139 613989 19141 613990
rect 19234 613765 19236 613766
rect 19235 613435 19236 613765
rect 19234 613434 19236 613435
rect 19139 611310 19141 611311
rect 19140 610990 19141 611310
rect 19139 610989 19141 610990
rect 19234 610765 19236 610766
rect 19235 610435 19236 610765
rect 19234 610434 19236 610435
rect 19139 608310 19141 608311
rect 19140 607990 19141 608310
rect 19139 607989 19141 607990
rect 19234 607765 19236 607766
rect 19235 607435 19236 607765
rect 19234 607434 19236 607435
rect 11077 605645 11079 605646
rect 11077 602850 11078 605645
rect 19139 605310 19141 605311
rect 19140 604990 19141 605310
rect 19139 604989 19141 604990
rect 19234 604765 19236 604766
rect 19235 604435 19236 604765
rect 19234 604434 19236 604435
rect 11077 602849 11079 602850
rect 19139 602310 19141 602311
rect 19140 601990 19141 602310
rect 19139 601989 19141 601990
rect 19234 601765 19236 601766
rect 19235 601435 19236 601765
rect 19234 601434 19236 601435
rect 19139 599310 19141 599311
rect 19140 598990 19141 599310
rect 19139 598989 19141 598990
rect 19234 598765 19236 598766
rect 19235 598435 19236 598765
rect 19234 598434 19236 598435
rect 19139 596310 19141 596311
rect 19140 595990 19141 596310
rect 19139 595989 19141 595990
rect 19234 595765 19236 595766
rect 19235 595435 19236 595765
rect 19234 595434 19236 595435
rect 19139 593310 19141 593311
rect 19140 592990 19141 593310
rect 19139 592989 19141 592990
rect 19234 592765 19236 592766
rect 19235 592435 19236 592765
rect 19234 592434 19236 592435
rect 19139 590310 19141 590311
rect 19140 589990 19141 590310
rect 19139 589989 19141 589990
rect 19234 589765 19236 589766
rect 19235 589435 19236 589765
rect 19234 589434 19236 589435
rect 19139 587310 19141 587311
rect 19140 586990 19141 587310
rect 19139 586989 19141 586990
rect 19234 586765 19236 586766
rect 19235 586435 19236 586765
rect 19234 586434 19236 586435
rect 19139 584310 19141 584311
rect 19140 583990 19141 584310
rect 19139 583989 19141 583990
rect 19234 583765 19236 583766
rect 19235 583435 19236 583765
rect 19234 583434 19236 583435
rect 19139 581310 19141 581311
rect 19140 580990 19141 581310
rect 19139 580989 19141 580990
rect 19234 580765 19236 580766
rect 19235 580435 19236 580765
rect 19234 580434 19236 580435
rect 19139 578310 19141 578311
rect 19140 577990 19141 578310
rect 19139 577989 19141 577990
rect 19234 577765 19236 577766
rect 19235 577435 19236 577765
rect 19234 577434 19236 577435
rect 19139 575310 19141 575311
rect 19140 574990 19141 575310
rect 19139 574989 19141 574990
rect 19234 574765 19236 574766
rect 19235 574435 19236 574765
rect 19234 574434 19236 574435
rect 19139 572310 19141 572311
rect 19140 571990 19141 572310
rect 19139 571989 19141 571990
rect 19234 571765 19236 571766
rect 19235 571435 19236 571765
rect 19234 571434 19236 571435
rect 19139 569310 19141 569311
rect 19140 568990 19141 569310
rect 19139 568989 19141 568990
rect 19234 568765 19236 568766
rect 19235 568435 19236 568765
rect 19234 568434 19236 568435
rect 19139 566310 19141 566311
rect 19140 565990 19141 566310
rect 19139 565989 19141 565990
rect 19234 565765 19236 565766
rect 19235 565435 19236 565765
rect 19234 565434 19236 565435
rect 19139 563310 19141 563311
rect 19140 562990 19141 563310
rect 19139 562989 19141 562990
rect 19234 562765 19236 562766
rect 19235 562435 19236 562765
rect 19234 562434 19236 562435
rect 19139 560310 19141 560311
rect 19140 559990 19141 560310
rect 19139 559989 19141 559990
rect 19234 559765 19236 559766
rect 19235 559435 19236 559765
rect 19234 559434 19236 559435
rect 19139 557310 19141 557311
rect 19140 556990 19141 557310
rect 19139 556989 19141 556990
rect 19234 556765 19236 556766
rect 19235 556435 19236 556765
rect 19234 556434 19236 556435
rect 17413 554834 17415 554835
rect 17414 552079 17415 554834
rect 19139 554310 19141 554311
rect 19140 553990 19141 554310
rect 19139 553989 19141 553990
rect 19234 553765 19236 553766
rect 19235 553435 19236 553765
rect 19234 553434 19236 553435
rect 17413 552078 17415 552079
rect 19139 551310 19141 551311
rect 19140 550990 19141 551310
rect 19139 550989 19141 550990
rect 19234 550765 19236 550766
rect 19235 550435 19236 550765
rect 19234 550434 19236 550435
rect 19139 548310 19141 548311
rect 19140 547990 19141 548310
rect 19139 547989 19141 547990
rect 19234 547765 19236 547766
rect 19235 547435 19236 547765
rect 19234 547434 19236 547435
rect 19139 545310 19141 545311
rect 19140 544990 19141 545310
rect 19139 544989 19141 544990
rect 19234 544765 19236 544766
rect 19235 544435 19236 544765
rect 19234 544434 19236 544435
rect 19139 542310 19141 542311
rect 19140 541990 19141 542310
rect 19139 541989 19141 541990
rect 19234 541765 19236 541766
rect 19235 541435 19236 541765
rect 19234 541434 19236 541435
rect 19139 539310 19141 539311
rect 19140 538990 19141 539310
rect 19139 538989 19141 538990
rect 19234 538765 19236 538766
rect 19235 538435 19236 538765
rect 19234 538434 19236 538435
rect 19139 536310 19141 536311
rect 19140 535990 19141 536310
rect 19139 535989 19141 535990
rect 19234 535765 19236 535766
rect 19235 535435 19236 535765
rect 19234 535434 19236 535435
rect 19139 533310 19141 533311
rect 19140 532990 19141 533310
rect 19139 532989 19141 532990
rect 19234 532765 19236 532766
rect 19235 532435 19236 532765
rect 19234 532434 19236 532435
rect 19139 530310 19141 530311
rect 19140 529990 19141 530310
rect 19139 529989 19141 529990
rect 19234 529765 19236 529766
rect 19235 529435 19236 529765
rect 19234 529434 19236 529435
rect 19139 527310 19141 527311
rect 19140 526990 19141 527310
rect 19139 526989 19141 526990
rect 19234 526765 19236 526766
rect 19235 526435 19236 526765
rect 19234 526434 19236 526435
rect 19139 524310 19141 524311
rect 19140 523990 19141 524310
rect 19139 523989 19141 523990
rect 19234 523765 19236 523766
rect 19235 523435 19236 523765
rect 19234 523434 19236 523435
rect 19139 521310 19141 521311
rect 19140 520990 19141 521310
rect 19139 520989 19141 520990
rect 19234 520765 19236 520766
rect 19235 520435 19236 520765
rect 19234 520434 19236 520435
rect 19139 518310 19141 518311
rect 19140 517990 19141 518310
rect 19139 517989 19141 517990
rect 19234 517765 19236 517766
rect 19235 517435 19236 517765
rect 19234 517434 19236 517435
rect 19139 515310 19141 515311
rect 19140 514990 19141 515310
rect 19139 514989 19141 514990
rect 19139 512310 19141 512311
rect 19140 511990 19141 512310
rect 19139 511989 19141 511990
rect 19234 511765 19236 511766
rect 19235 511435 19236 511765
rect 19234 511434 19236 511435
rect 19139 509310 19141 509311
rect 19140 508990 19141 509310
rect 19139 508989 19141 508990
rect 19234 508765 19236 508766
rect 19235 508435 19236 508765
rect 19234 508434 19236 508435
rect 18396 508304 18398 508305
rect 18397 505549 18398 508304
rect 19139 506310 19141 506311
rect 19140 505990 19141 506310
rect 19139 505989 19141 505990
rect 18396 505548 18398 505549
rect 19234 505765 19236 505766
rect 19235 505435 19236 505765
rect 19234 505434 19236 505435
rect 19139 503310 19141 503311
rect 19140 502990 19141 503310
rect 19139 502989 19141 502990
rect 19234 502765 19236 502766
rect 19235 502435 19236 502765
rect 19234 502434 19236 502435
rect 19139 500310 19141 500311
rect 19140 499990 19141 500310
rect 19139 499989 19141 499990
rect 11077 499927 11079 499928
rect 11077 497132 11078 499927
rect 19234 499765 19236 499766
rect 19235 499435 19236 499765
rect 19234 499434 19236 499435
rect 11077 497131 11079 497132
rect 19139 497310 19141 497311
rect 19140 496990 19141 497310
rect 19139 496989 19141 496990
rect 19234 496765 19236 496766
rect 19235 496435 19236 496765
rect 19234 496434 19236 496435
rect 19139 494310 19141 494311
rect 19140 493990 19141 494310
rect 19139 493989 19141 493990
rect 19234 493765 19236 493766
rect 19235 493435 19236 493765
rect 19234 493434 19236 493435
rect 19139 491310 19141 491311
rect 19140 490990 19141 491310
rect 19139 490989 19141 490990
rect 19234 490765 19236 490766
rect 19235 490435 19236 490765
rect 19234 490434 19236 490435
rect 19139 488310 19141 488311
rect 19140 487990 19141 488310
rect 19139 487989 19141 487990
rect 19234 487765 19236 487766
rect 19235 487435 19236 487765
rect 19234 487434 19236 487435
rect 19139 485310 19141 485311
rect 19140 484990 19141 485310
rect 19139 484989 19141 484990
rect 19234 484765 19236 484766
rect 19235 484435 19236 484765
rect 19234 484434 19236 484435
rect 19139 482310 19141 482311
rect 19140 481990 19141 482310
rect 19139 481989 19141 481990
rect 19234 481765 19236 481766
rect 19235 481435 19236 481765
rect 19234 481434 19236 481435
rect 19139 479310 19141 479311
rect 19140 478990 19141 479310
rect 19139 478989 19141 478990
rect 19234 478765 19236 478766
rect 19235 478435 19236 478765
rect 19234 478434 19236 478435
rect 19139 476310 19141 476311
rect 19140 475990 19141 476310
rect 19139 475989 19141 475990
rect 19234 475765 19236 475766
rect 19235 475435 19236 475765
rect 19234 475434 19236 475435
rect 19139 473310 19141 473311
rect 19140 472990 19141 473310
rect 19139 472989 19141 472990
rect 19234 472765 19236 472766
rect 19235 472435 19236 472765
rect 19234 472434 19236 472435
rect 19139 470310 19141 470311
rect 19140 469990 19141 470310
rect 19139 469989 19141 469990
rect 19234 469765 19236 469766
rect 19235 469435 19236 469765
rect 19234 469434 19236 469435
rect 19139 467310 19141 467311
rect 19140 466990 19141 467310
rect 19139 466989 19141 466990
rect 19234 466765 19236 466766
rect 19235 466435 19236 466765
rect 19234 466434 19236 466435
rect 19139 464310 19141 464311
rect 19140 463990 19141 464310
rect 19139 463989 19141 463990
rect 19234 463765 19236 463766
rect 19235 463435 19236 463765
rect 19234 463434 19236 463435
rect 11077 461424 13834 461425
rect 11077 458587 11078 461424
rect 13833 461383 13834 461424
rect 13833 458628 14868 461383
rect 19139 461310 19141 461311
rect 19140 460990 19141 461310
rect 19139 460989 19141 460990
rect 19234 460765 19236 460766
rect 19235 460435 19236 460765
rect 19234 460434 19236 460435
rect 13833 458587 13834 458628
rect 11077 458586 13834 458587
rect 19139 458310 19141 458311
rect 19140 457990 19141 458310
rect 19139 457989 19141 457990
rect 19234 457765 19236 457766
rect 19235 457435 19236 457765
rect 19234 457434 19236 457435
rect 19139 455310 19141 455311
rect 19140 454990 19141 455310
rect 19139 454989 19141 454990
rect 19234 454765 19236 454766
rect 19235 454435 19236 454765
rect 19234 454434 19236 454435
rect 19139 452310 19141 452311
rect 19140 451990 19141 452310
rect 19139 451989 19141 451990
rect 19234 451765 19236 451766
rect 19235 451435 19236 451765
rect 19234 451434 19236 451435
rect 19139 449310 19141 449311
rect 19140 448990 19141 449310
rect 19139 448989 19141 448990
rect 19234 448765 19236 448766
rect 19235 448435 19236 448765
rect 19234 448434 19236 448435
rect 19139 446310 19141 446311
rect 19140 445990 19141 446310
rect 19139 445989 19141 445990
rect 19234 445765 19236 445766
rect 19235 445435 19236 445765
rect 19234 445434 19236 445435
rect 19139 443310 19141 443311
rect 19140 442990 19141 443310
rect 19139 442989 19141 442990
rect 19234 442765 19236 442766
rect 19235 442435 19236 442765
rect 19234 442434 19236 442435
rect 19139 440310 19141 440311
rect 19140 439990 19141 440310
rect 19139 439989 19141 439990
rect 19234 439765 19236 439766
rect 19235 439435 19236 439765
rect 19234 439434 19236 439435
rect 19139 437310 19141 437311
rect 19140 436990 19141 437310
rect 19139 436989 19141 436990
rect 19234 436765 19236 436766
rect 19235 436435 19236 436765
rect 19234 436434 19236 436435
rect 19139 434310 19141 434311
rect 19140 433990 19141 434310
rect 19139 433989 19141 433990
rect 19234 433765 19236 433766
rect 19235 433435 19236 433765
rect 19234 433434 19236 433435
rect 19139 431310 19141 431311
rect 19140 430990 19141 431310
rect 19139 430989 19141 430990
rect 19234 430765 19236 430766
rect 19235 430435 19236 430765
rect 19234 430434 19236 430435
rect 19139 428310 19141 428311
rect 19140 427990 19141 428310
rect 19139 427989 19141 427990
rect 19234 427765 19236 427766
rect 19235 427435 19236 427765
rect 19234 427434 19236 427435
rect 19139 425310 19141 425311
rect 19140 424990 19141 425310
rect 19139 424989 19141 424990
rect 19234 424765 19236 424766
rect 19235 424435 19236 424765
rect 19234 424434 19236 424435
rect 19139 422310 19141 422311
rect 19140 421990 19141 422310
rect 19139 421989 19141 421990
rect 19234 421765 19236 421766
rect 19235 421435 19236 421765
rect 19234 421434 19236 421435
rect 19139 419310 19141 419311
rect 19140 418990 19141 419310
rect 19139 418989 19141 418990
rect 19234 418765 19236 418766
rect 19235 418435 19236 418765
rect 19234 418434 19236 418435
rect 19139 416310 19141 416311
rect 19140 415990 19141 416310
rect 19139 415989 19141 415990
rect 19234 415765 19236 415766
rect 19235 415435 19236 415765
rect 19234 415434 19236 415435
rect 19139 413310 19141 413311
rect 19140 412990 19141 413310
rect 19139 412989 19141 412990
rect 19234 412765 19236 412766
rect 19235 412435 19236 412765
rect 19234 412434 19236 412435
rect 19139 410310 19141 410311
rect 19140 409990 19141 410310
rect 19139 409989 19141 409990
rect 19234 409765 19236 409766
rect 19235 409435 19236 409765
rect 19234 409434 19236 409435
rect 19139 407310 19141 407311
rect 19140 406990 19141 407310
rect 19139 406989 19141 406990
rect 19234 406765 19236 406766
rect 19235 406435 19236 406765
rect 19234 406434 19236 406435
rect 19139 404310 19141 404311
rect 19140 403990 19141 404310
rect 19139 403989 19141 403990
rect 19234 403765 19236 403766
rect 19235 403435 19236 403765
rect 19234 403434 19236 403435
rect 19139 401310 19141 401311
rect 19140 400990 19141 401310
rect 19139 400989 19141 400990
rect 19139 398310 19141 398311
rect 19140 397990 19141 398310
rect 19139 397989 19141 397990
rect 19234 397765 19236 397766
rect 19235 397435 19236 397765
rect 19234 397434 19236 397435
rect 19139 395310 19141 395311
rect 19140 394990 19141 395310
rect 19139 394989 19141 394990
rect 19234 394765 19236 394766
rect 19235 394435 19236 394765
rect 19234 394434 19236 394435
rect 19139 392310 19141 392311
rect 19140 391990 19141 392310
rect 19139 391989 19141 391990
rect 19234 391765 19236 391766
rect 19235 391435 19236 391765
rect 19234 391434 19236 391435
rect 19139 389310 19141 389311
rect 19140 388990 19141 389310
rect 19139 388989 19141 388990
rect 19234 388765 19236 388766
rect 19235 388435 19236 388765
rect 19234 388434 19236 388435
rect 19139 386310 19141 386311
rect 19140 385990 19141 386310
rect 19139 385989 19141 385990
rect 19234 385765 19236 385766
rect 19235 385435 19236 385765
rect 19234 385434 19236 385435
rect 19139 383310 19141 383311
rect 19140 382990 19141 383310
rect 19139 382989 19141 382990
rect 19234 382765 19236 382766
rect 19235 382435 19236 382765
rect 19234 382434 19236 382435
rect 19139 380310 19141 380311
rect 19140 379990 19141 380310
rect 19139 379989 19141 379990
rect 19234 379765 19236 379766
rect 19235 379435 19236 379765
rect 19234 379434 19236 379435
rect 19139 377310 19141 377311
rect 19140 376990 19141 377310
rect 19139 376989 19141 376990
rect 19234 376765 19236 376766
rect 19235 376435 19236 376765
rect 19234 376434 19236 376435
rect 19139 374310 19141 374311
rect 19140 373990 19141 374310
rect 19139 373989 19141 373990
rect 19234 373765 19236 373766
rect 19235 373435 19236 373765
rect 19234 373434 19236 373435
rect 19139 371310 19141 371311
rect 19140 370990 19141 371310
rect 19139 370989 19141 370990
rect 19234 370765 19236 370766
rect 19235 370435 19236 370765
rect 19234 370434 19236 370435
rect 19139 368310 19141 368311
rect 19140 367990 19141 368310
rect 19139 367989 19141 367990
rect 19234 367765 19236 367766
rect 19235 367435 19236 367765
rect 19234 367434 19236 367435
rect 19139 365310 19141 365311
rect 19140 364990 19141 365310
rect 19139 364989 19141 364990
rect 19234 364765 19236 364766
rect 19235 364435 19236 364765
rect 19234 364434 19236 364435
rect 19139 362310 19141 362311
rect 19140 361990 19141 362310
rect 19139 361989 19141 361990
rect 31813 358331 31923 692010
rect 50825 674598 50937 674599
rect 50825 674595 50826 674598
rect 46878 674488 50826 674595
rect 50936 674595 50937 674598
rect 50936 674594 126146 674595
rect 50936 674488 126037 674594
rect 46878 674486 126037 674488
rect 126145 674486 126146 674594
rect 46878 674485 126146 674486
rect 46878 670057 46988 674485
rect 155835 674109 156205 682425
rect 574553 682650 577887 682687
rect 574553 682402 582200 682650
rect 574553 678818 575238 682402
rect 582000 678818 582200 682402
rect 574553 678570 582200 678818
rect 405469 675200 405471 675201
rect 155829 674108 156211 674109
rect 155829 673738 155830 674108
rect 156210 673738 156211 674108
rect 155829 673737 156211 673738
rect 231033 673996 231353 673997
rect 140626 673729 140708 673730
rect 140626 673659 140627 673729
rect 140707 673659 140708 673729
rect 231033 673678 231034 673996
rect 231352 673678 231353 673996
rect 231033 673677 231353 673678
rect 140626 673658 140708 673659
rect 140632 671134 140702 673658
rect 405470 672740 405471 675200
rect 405469 672739 405471 672740
rect 140632 671066 140633 671134
rect 140701 671066 140702 671134
rect 140632 671065 140702 671066
rect 402809 670886 405271 670887
rect 402809 670885 402810 670886
rect 405270 670885 405271 670886
rect 143667 670731 144069 670732
rect 143667 670730 143668 670731
rect 144068 670730 144069 670731
rect 501549 670886 504011 670887
rect 501549 670885 501550 670886
rect 504010 670885 504011 670886
rect 34053 667759 34373 667760
rect 34053 667441 34054 667759
rect 34372 667441 34373 667759
rect 34053 667440 34373 667441
rect 358691 666311 403637 666631
rect 408464 665164 409289 666667
rect 574553 665164 577887 678570
rect 34053 664759 34373 664760
rect 34053 664441 34054 664759
rect 34372 664441 34373 664759
rect 34053 664440 34373 664441
rect 53663 664727 53983 664728
rect 53663 664409 53664 664727
rect 53982 664409 53983 664727
rect 53663 664408 53983 664409
rect 358691 663311 403637 663631
rect 32570 662309 51843 662310
rect 32570 661991 32571 662309
rect 32889 662286 51843 662309
rect 32889 662014 51547 662286
rect 51819 662014 51843 662286
rect 32889 661991 51843 662014
rect 32570 661990 51843 661991
rect 408150 661830 577887 665164
rect 34053 661759 34373 661760
rect 34053 661441 34054 661759
rect 34372 661441 34373 661759
rect 34053 661440 34373 661441
rect 358691 660311 403637 660631
rect 32570 659309 51843 659310
rect 32570 658991 32571 659309
rect 32889 659286 51843 659309
rect 32889 659014 51547 659286
rect 51819 659014 51843 659286
rect 32889 658991 51843 659014
rect 32570 658990 51843 658991
rect 34053 658759 34373 658760
rect 34053 658441 34054 658759
rect 34372 658441 34373 658759
rect 34053 658440 34373 658441
rect 358691 657311 403637 657631
rect 32570 656309 51843 656310
rect 32570 655991 32571 656309
rect 32889 656286 51843 656309
rect 32889 656014 51547 656286
rect 51819 656014 51843 656286
rect 32889 655991 51843 656014
rect 32570 655990 51843 655991
rect 34053 655759 34373 655760
rect 34053 655441 34054 655759
rect 34372 655441 34373 655759
rect 34053 655440 34373 655441
rect 358691 654311 403637 654631
rect 32570 653309 51843 653310
rect 32570 652991 32571 653309
rect 32889 653286 51843 653309
rect 32889 653014 51547 653286
rect 51819 653014 51843 653286
rect 32889 652991 51843 653014
rect 32570 652990 51843 652991
rect 34053 652759 34373 652760
rect 34053 652441 34054 652759
rect 34372 652441 34373 652759
rect 34053 652440 34373 652441
rect 358691 651311 403637 651631
rect 32570 650309 51843 650310
rect 32570 649991 32571 650309
rect 32889 650286 51843 650309
rect 32889 650014 51547 650286
rect 51819 650014 51843 650286
rect 32889 649991 51843 650014
rect 32570 649990 51843 649991
rect 34053 649759 34373 649760
rect 34053 649441 34054 649759
rect 34372 649441 34373 649759
rect 34053 649440 34373 649441
rect 358691 648311 403637 648631
rect 32570 647309 51843 647310
rect 32570 646991 32571 647309
rect 32889 647286 51843 647309
rect 32889 647014 51547 647286
rect 51819 647014 51843 647286
rect 32889 646991 51843 647014
rect 32570 646990 51843 646991
rect 34053 646759 34373 646760
rect 34053 646441 34054 646759
rect 34372 646441 34373 646759
rect 34053 646440 34373 646441
rect 358691 645311 403637 645631
rect 32570 644309 51843 644310
rect 32570 643991 32571 644309
rect 32889 644286 51843 644309
rect 32889 644014 51547 644286
rect 51819 644014 51843 644286
rect 32889 643991 51843 644014
rect 32570 643990 51843 643991
rect 34053 643759 34373 643760
rect 34053 643441 34054 643759
rect 34372 643441 34373 643759
rect 34053 643440 34373 643441
rect 358691 642311 403637 642631
rect 32570 641309 51843 641310
rect 32570 640991 32571 641309
rect 32889 641286 51843 641309
rect 32889 641014 51547 641286
rect 51819 641014 51843 641286
rect 32889 640991 51843 641014
rect 32570 640990 51843 640991
rect 34053 640759 34373 640760
rect 34053 640441 34054 640759
rect 34372 640441 34373 640759
rect 34053 640440 34373 640441
rect 358691 639311 403637 639631
rect 32570 638309 51843 638310
rect 32570 637991 32571 638309
rect 32889 638286 51843 638309
rect 32889 638014 51547 638286
rect 51819 638014 51843 638286
rect 32889 637991 51843 638014
rect 32570 637990 51843 637991
rect 34053 637759 34373 637760
rect 34053 637441 34054 637759
rect 34372 637441 34373 637759
rect 34053 637440 34373 637441
rect 358691 636311 403637 636631
rect 32570 635309 51843 635310
rect 32570 634991 32571 635309
rect 32889 635286 51843 635309
rect 32889 635014 51547 635286
rect 51819 635014 51843 635286
rect 32889 634991 51843 635014
rect 32570 634990 51843 634991
rect 34053 634759 34373 634760
rect 34053 634441 34054 634759
rect 34372 634441 34373 634759
rect 34053 634440 34373 634441
rect 358691 633311 403637 633631
rect 32570 632309 51843 632310
rect 32570 631991 32571 632309
rect 32889 632286 51843 632309
rect 32889 632014 51547 632286
rect 51819 632014 51843 632286
rect 32889 631991 51843 632014
rect 32570 631990 51843 631991
rect 34053 631759 34373 631760
rect 34053 631441 34054 631759
rect 34372 631441 34373 631759
rect 34053 631440 34373 631441
rect 358691 630311 403637 630631
rect 407221 627994 407223 627995
rect 358691 627311 403637 627631
rect 34053 625759 34373 625760
rect 34053 625441 34054 625759
rect 34372 625441 34373 625759
rect 407222 625524 407223 627994
rect 407221 625523 407223 625524
rect 34053 625440 34373 625441
rect 358691 624311 403637 624631
rect 32570 623309 51843 623310
rect 32570 622991 32571 623309
rect 32889 623286 51843 623309
rect 32889 623014 51547 623286
rect 51819 623014 51843 623286
rect 32889 622991 51843 623014
rect 32570 622990 51843 622991
rect 34053 622759 34373 622760
rect 34053 622441 34054 622759
rect 34372 622441 34373 622759
rect 34053 622440 34373 622441
rect 358691 621311 403637 621631
rect 32570 620309 51843 620310
rect 32570 619991 32571 620309
rect 32889 620286 51843 620309
rect 32889 620014 51547 620286
rect 51819 620014 51843 620286
rect 32889 619991 51843 620014
rect 32570 619990 51843 619991
rect 34053 619759 34373 619760
rect 34053 619441 34054 619759
rect 34372 619441 34373 619759
rect 34053 619440 34373 619441
rect 358691 618311 403637 618631
rect 32570 617309 51843 617310
rect 32570 616991 32571 617309
rect 32889 617286 51843 617309
rect 32889 617014 51547 617286
rect 51819 617014 51843 617286
rect 32889 616991 51843 617014
rect 32570 616990 51843 616991
rect 34053 616759 34373 616760
rect 34053 616441 34054 616759
rect 34372 616441 34373 616759
rect 34053 616440 34373 616441
rect 407361 615824 407363 615825
rect 358691 615311 403637 615631
rect 32570 614309 51843 614310
rect 32570 613991 32571 614309
rect 32889 614286 51843 614309
rect 32889 614014 51547 614286
rect 51819 614014 51843 614286
rect 32889 613991 51843 614014
rect 32570 613990 51843 613991
rect 34053 613759 34373 613760
rect 34053 613441 34054 613759
rect 34372 613441 34373 613759
rect 34053 613440 34373 613441
rect 407362 613354 407363 615824
rect 407361 613353 407363 613354
rect 358691 612311 403637 612631
rect 32570 611309 51843 611310
rect 32570 610991 32571 611309
rect 32889 611286 51843 611309
rect 32889 611014 51547 611286
rect 51819 611014 51843 611286
rect 32889 610991 51843 611014
rect 32570 610990 51843 610991
rect 34053 610759 34373 610760
rect 34053 610441 34054 610759
rect 34372 610441 34373 610759
rect 34053 610440 34373 610441
rect 358691 609311 403637 609631
rect 32570 608309 51843 608310
rect 32570 607991 32571 608309
rect 32889 608286 51843 608309
rect 32889 608014 51547 608286
rect 51819 608014 51843 608286
rect 32889 607991 51843 608014
rect 32570 607990 51843 607991
rect 34053 607759 34373 607760
rect 34053 607441 34054 607759
rect 34372 607441 34373 607759
rect 34053 607440 34373 607441
rect 358691 606311 403637 606631
rect 32570 605309 51843 605310
rect 32570 604991 32571 605309
rect 32889 605286 51843 605309
rect 32889 605014 51547 605286
rect 51819 605014 51843 605286
rect 32889 604991 51843 605014
rect 32570 604990 51843 604991
rect 34053 604759 34373 604760
rect 34053 604441 34054 604759
rect 34372 604441 34373 604759
rect 34053 604440 34373 604441
rect 358691 603311 403637 603631
rect 32570 602309 51843 602310
rect 32570 601991 32571 602309
rect 32889 602286 51843 602309
rect 32889 602014 51547 602286
rect 51819 602014 51843 602286
rect 32889 601991 51843 602014
rect 32570 601990 51843 601991
rect 406872 602185 406874 602186
rect 34053 601759 34373 601760
rect 34053 601441 34054 601759
rect 34372 601441 34373 601759
rect 34053 601440 34373 601441
rect 358691 600311 403637 600631
rect 406873 599715 406874 602185
rect 406872 599714 406874 599715
rect 32570 599309 51843 599310
rect 32570 598991 32571 599309
rect 32889 599286 51843 599309
rect 32889 599014 51547 599286
rect 51819 599014 51843 599286
rect 32889 598991 51843 599014
rect 32570 598990 51843 598991
rect 34053 598759 34373 598760
rect 34053 598441 34054 598759
rect 34372 598441 34373 598759
rect 34053 598440 34373 598441
rect 358691 597311 403637 597631
rect 32570 596309 51843 596310
rect 32570 595991 32571 596309
rect 32889 596286 51843 596309
rect 32889 596014 51547 596286
rect 51819 596014 51843 596286
rect 32889 595991 51843 596014
rect 32570 595990 51843 595991
rect 34053 595759 34373 595760
rect 34053 595441 34054 595759
rect 34372 595441 34373 595759
rect 34053 595440 34373 595441
rect 358691 594311 403637 594631
rect 32570 593309 51843 593310
rect 32570 592991 32571 593309
rect 32889 593286 51843 593309
rect 32889 593014 51547 593286
rect 51819 593014 51843 593286
rect 32889 592991 51843 593014
rect 32570 592990 51843 592991
rect 34053 592759 34373 592760
rect 34053 592441 34054 592759
rect 34372 592441 34373 592759
rect 34053 592440 34373 592441
rect 358691 591311 403637 591631
rect 32570 590309 51843 590310
rect 32570 589991 32571 590309
rect 32889 590286 51843 590309
rect 32889 590014 51547 590286
rect 51819 590014 51843 590286
rect 32889 589991 51843 590014
rect 32570 589990 51843 589991
rect 34053 589759 34373 589760
rect 34053 589441 34054 589759
rect 34372 589441 34373 589759
rect 34053 589440 34373 589441
rect 358691 588311 403637 588631
rect 406172 587358 406174 587359
rect 32570 587309 51843 587310
rect 32570 586991 32571 587309
rect 32889 587286 51843 587309
rect 32889 587014 51547 587286
rect 51819 587014 51843 587286
rect 32889 586991 51843 587014
rect 32570 586990 51843 586991
rect 34053 586759 34373 586760
rect 34053 586441 34054 586759
rect 34372 586441 34373 586759
rect 34053 586440 34373 586441
rect 358691 585311 403637 585631
rect 406173 584888 406174 587358
rect 406172 584887 406174 584888
rect 32570 584309 51843 584310
rect 32570 583991 32571 584309
rect 32889 584286 51843 584309
rect 32889 584014 51547 584286
rect 51819 584014 51843 584286
rect 32889 583991 51843 584014
rect 32570 583990 51843 583991
rect 34053 583759 34373 583760
rect 34053 583441 34054 583759
rect 34372 583441 34373 583759
rect 34053 583440 34373 583441
rect 358691 582311 403637 582631
rect 32570 581309 51843 581310
rect 32570 580991 32571 581309
rect 32889 581286 51843 581309
rect 32889 581014 51547 581286
rect 51819 581014 51843 581286
rect 32889 580991 51843 581014
rect 32570 580990 51843 580991
rect 34053 580759 34373 580760
rect 34053 580441 34054 580759
rect 34372 580441 34373 580759
rect 34053 580440 34373 580441
rect 358691 579311 403637 579631
rect 32570 578309 51843 578310
rect 32570 577991 32571 578309
rect 32889 578286 51843 578309
rect 32889 578014 51547 578286
rect 51819 578014 51843 578286
rect 32889 577991 51843 578014
rect 32570 577990 51843 577991
rect 34053 577759 34373 577760
rect 34053 577441 34054 577759
rect 34372 577441 34373 577759
rect 34053 577440 34373 577441
rect 358691 576311 403637 576631
rect 32570 575309 51843 575310
rect 32570 574991 32571 575309
rect 32889 575286 51843 575309
rect 32889 575014 51547 575286
rect 51819 575014 51843 575286
rect 32889 574991 51843 575014
rect 32570 574990 51843 574991
rect 34053 574759 34373 574760
rect 34053 574441 34054 574759
rect 34372 574441 34373 574759
rect 34053 574440 34373 574441
rect 358691 573311 403637 573631
rect 32570 572309 51843 572310
rect 32570 571991 32571 572309
rect 32889 572286 51843 572309
rect 32889 572014 51547 572286
rect 51819 572014 51843 572286
rect 32889 571991 51843 572014
rect 32570 571990 51843 571991
rect 34053 571759 34373 571760
rect 34053 571441 34054 571759
rect 34372 571441 34373 571759
rect 34053 571440 34373 571441
rect 358691 570311 403637 570631
rect 32570 569309 51843 569310
rect 32570 568991 32571 569309
rect 32889 569286 51843 569309
rect 32889 569014 51547 569286
rect 51819 569014 51843 569286
rect 32889 568991 51843 569014
rect 32570 568990 51843 568991
rect 34053 568759 34373 568760
rect 34053 568441 34054 568759
rect 34372 568441 34373 568759
rect 34053 568440 34373 568441
rect 358691 567311 403637 567631
rect 32570 566309 51843 566310
rect 32570 565991 32571 566309
rect 32889 566286 51843 566309
rect 32889 566014 51547 566286
rect 51819 566014 51843 566286
rect 32889 565991 51843 566014
rect 32570 565990 51843 565991
rect 406807 566283 406809 566284
rect 34053 565759 34373 565760
rect 34053 565441 34054 565759
rect 34372 565441 34373 565759
rect 34053 565440 34373 565441
rect 358691 564311 403637 564631
rect 406808 563813 406809 566283
rect 406807 563812 406809 563813
rect 32570 563309 51843 563310
rect 32570 562991 32571 563309
rect 32889 563286 51843 563309
rect 32889 563014 51547 563286
rect 51819 563014 51843 563286
rect 32889 562991 51843 563014
rect 32570 562990 51843 562991
rect 34053 562759 34373 562760
rect 34053 562441 34054 562759
rect 34372 562441 34373 562759
rect 34053 562440 34373 562441
rect 358691 561311 403637 561631
rect 32570 560309 51843 560310
rect 32570 559991 32571 560309
rect 32889 560286 51843 560309
rect 32889 560014 51547 560286
rect 51819 560014 51843 560286
rect 32889 559991 51843 560014
rect 32570 559990 51843 559991
rect 34053 559759 34373 559760
rect 34053 559441 34054 559759
rect 34372 559441 34373 559759
rect 34053 559440 34373 559441
rect 358691 558311 403637 558631
rect 32570 557309 51843 557310
rect 32570 556991 32571 557309
rect 32889 557286 51843 557309
rect 32889 557014 51547 557286
rect 51819 557014 51843 557286
rect 32889 556991 51843 557014
rect 32570 556990 51843 556991
rect 34053 556759 34373 556760
rect 34053 556441 34054 556759
rect 34372 556441 34373 556759
rect 34053 556440 34373 556441
rect 358691 555311 403637 555631
rect 32570 554309 51843 554310
rect 32570 553991 32571 554309
rect 32889 554286 51843 554309
rect 32889 554014 51547 554286
rect 51819 554014 51843 554286
rect 32889 553991 51843 554014
rect 32570 553990 51843 553991
rect 34053 553759 34373 553760
rect 34053 553441 34054 553759
rect 34372 553441 34373 553759
rect 34053 553440 34373 553441
rect 358691 552311 403637 552631
rect 406881 552470 406883 552471
rect 32570 551309 51843 551310
rect 32570 550991 32571 551309
rect 32889 551286 51843 551309
rect 32889 551014 51547 551286
rect 51819 551014 51843 551286
rect 32889 550991 51843 551014
rect 32570 550990 51843 550991
rect 34053 550759 34373 550760
rect 34053 550441 34054 550759
rect 34372 550441 34373 550759
rect 34053 550440 34373 550441
rect 406882 550000 406883 552470
rect 406881 549999 406883 550000
rect 358691 549311 403637 549631
rect 32570 548309 51843 548310
rect 32570 547991 32571 548309
rect 32889 548286 51843 548309
rect 32889 548014 51547 548286
rect 51819 548014 51843 548286
rect 32889 547991 51843 548014
rect 32570 547990 51843 547991
rect 34053 547759 34373 547760
rect 34053 547441 34054 547759
rect 34372 547441 34373 547759
rect 34053 547440 34373 547441
rect 358691 546311 403637 546631
rect 32570 545309 51843 545310
rect 32570 544991 32571 545309
rect 32889 545286 51843 545309
rect 32889 545014 51547 545286
rect 51819 545014 51843 545286
rect 32889 544991 51843 545014
rect 32570 544990 51843 544991
rect 34053 544759 34373 544760
rect 34053 544441 34054 544759
rect 34372 544441 34373 544759
rect 34053 544440 34373 544441
rect 358691 543311 403637 543631
rect 406587 542846 406589 542847
rect 32570 542309 51843 542310
rect 32570 541991 32571 542309
rect 32889 542286 51843 542309
rect 32889 542014 51547 542286
rect 51819 542014 51843 542286
rect 32889 541991 51843 542014
rect 32570 541990 51843 541991
rect 34053 541759 34373 541760
rect 34053 541441 34054 541759
rect 34372 541441 34373 541759
rect 34053 541440 34373 541441
rect 358691 540311 403637 540631
rect 406588 540376 406589 542846
rect 406587 540375 406589 540376
rect 32570 539309 51843 539310
rect 32570 538991 32571 539309
rect 32889 539286 51843 539309
rect 32889 539014 51547 539286
rect 51819 539014 51843 539286
rect 32889 538991 51843 539014
rect 32570 538990 51843 538991
rect 34053 538759 34373 538760
rect 34053 538441 34054 538759
rect 34372 538441 34373 538759
rect 34053 538440 34373 538441
rect 358691 537311 403637 537631
rect 32570 536309 51843 536310
rect 32570 535991 32571 536309
rect 32889 536286 51843 536309
rect 32889 536014 51547 536286
rect 51819 536014 51843 536286
rect 32889 535991 51843 536014
rect 32570 535990 51843 535991
rect 34053 535759 34373 535760
rect 34053 535441 34054 535759
rect 34372 535441 34373 535759
rect 34053 535440 34373 535441
rect 358691 534311 403637 534631
rect 32570 533309 51843 533310
rect 32570 532991 32571 533309
rect 32889 533286 51843 533309
rect 32889 533014 51547 533286
rect 51819 533014 51843 533286
rect 32889 532991 51843 533014
rect 32570 532990 51843 532991
rect 34053 532759 34373 532760
rect 34053 532441 34054 532759
rect 34372 532441 34373 532759
rect 34053 532440 34373 532441
rect 406587 531898 406589 531899
rect 358691 531311 403637 531631
rect 32570 530309 51843 530310
rect 32570 529991 32571 530309
rect 32889 530286 51843 530309
rect 32889 530014 51547 530286
rect 51819 530014 51843 530286
rect 32889 529991 51843 530014
rect 32570 529990 51843 529991
rect 34053 529759 34373 529760
rect 34053 529441 34054 529759
rect 34372 529441 34373 529759
rect 34053 529440 34373 529441
rect 406588 529428 406589 531898
rect 406587 529427 406589 529428
rect 358691 528311 403637 528631
rect 32570 527309 51843 527310
rect 32570 526991 32571 527309
rect 32889 527286 51843 527309
rect 32889 527014 51547 527286
rect 51819 527014 51843 527286
rect 32889 526991 51843 527014
rect 32570 526990 51843 526991
rect 34053 526759 34373 526760
rect 34053 526441 34054 526759
rect 34372 526441 34373 526759
rect 34053 526440 34373 526441
rect 358691 525311 403637 525631
rect 32570 524309 51843 524310
rect 32570 523991 32571 524309
rect 32889 524286 51843 524309
rect 32889 524014 51547 524286
rect 51819 524014 51843 524286
rect 32889 523991 51843 524014
rect 32570 523990 51843 523991
rect 34053 523759 34373 523760
rect 34053 523441 34054 523759
rect 34372 523441 34373 523759
rect 34053 523440 34373 523441
rect 358691 522311 403637 522631
rect 32570 521309 51843 521310
rect 32570 520991 32571 521309
rect 32889 521286 51843 521309
rect 32889 521014 51547 521286
rect 51819 521014 51843 521286
rect 32889 520991 51843 521014
rect 32570 520990 51843 520991
rect 34053 520759 34373 520760
rect 34053 520441 34054 520759
rect 34372 520441 34373 520759
rect 34053 520440 34373 520441
rect 358691 519311 403637 519631
rect 32570 518309 51843 518310
rect 32570 517991 32571 518309
rect 32889 518286 51843 518309
rect 32889 518014 51547 518286
rect 51819 518014 51843 518286
rect 32889 517991 51843 518014
rect 32570 517990 51843 517991
rect 34053 517759 34373 517760
rect 34053 517441 34054 517759
rect 34372 517441 34373 517759
rect 34053 517440 34373 517441
rect 358691 516311 403637 516631
rect 32570 515309 51843 515310
rect 32570 514991 32571 515309
rect 32889 515286 51843 515309
rect 32889 515014 51547 515286
rect 51819 515014 51843 515286
rect 32889 514991 51843 515014
rect 32570 514990 51843 514991
rect 358691 513311 403637 513631
rect 406633 512948 406635 512949
rect 32570 512309 51843 512310
rect 32570 511991 32571 512309
rect 32889 512286 51843 512309
rect 32889 512014 51547 512286
rect 51819 512014 51843 512286
rect 32889 511991 51843 512014
rect 32570 511990 51843 511991
rect 34053 511759 34373 511760
rect 34053 511441 34054 511759
rect 34372 511441 34373 511759
rect 34053 511440 34373 511441
rect 358691 510311 403637 510631
rect 406634 510478 406635 512948
rect 406633 510477 406635 510478
rect 32570 509309 51843 509310
rect 32570 508991 32571 509309
rect 32889 509286 51843 509309
rect 32889 509014 51547 509286
rect 51819 509014 51843 509286
rect 32889 508991 51843 509014
rect 32570 508990 51843 508991
rect 34053 508759 34373 508760
rect 34053 508441 34054 508759
rect 34372 508441 34373 508759
rect 34053 508440 34373 508441
rect 358691 507311 403637 507631
rect 32570 506309 51843 506310
rect 32570 505991 32571 506309
rect 32889 506286 51843 506309
rect 32889 506014 51547 506286
rect 51819 506014 51843 506286
rect 32889 505991 51843 506014
rect 32570 505990 51843 505991
rect 34053 505759 34373 505760
rect 34053 505441 34054 505759
rect 34372 505441 34373 505759
rect 34053 505440 34373 505441
rect 358691 504311 403637 504631
rect 32570 503309 51843 503310
rect 32570 502991 32571 503309
rect 32889 503286 51843 503309
rect 32889 503014 51547 503286
rect 51819 503014 51843 503286
rect 32889 502991 51843 503014
rect 32570 502990 51843 502991
rect 34053 502759 34373 502760
rect 34053 502441 34054 502759
rect 34372 502441 34373 502759
rect 34053 502440 34373 502441
rect 358691 501311 403637 501631
rect 32570 500309 51843 500310
rect 32570 499991 32571 500309
rect 32889 500286 51843 500309
rect 32889 500014 51547 500286
rect 51819 500014 51843 500286
rect 32889 499991 51843 500014
rect 32570 499990 51843 499991
rect 34053 499759 34373 499760
rect 34053 499441 34054 499759
rect 34372 499441 34373 499759
rect 34053 499440 34373 499441
rect 358691 498311 403637 498631
rect 32570 497309 51843 497310
rect 32570 496991 32571 497309
rect 32889 497286 51843 497309
rect 32889 497014 51547 497286
rect 51819 497014 51843 497286
rect 32889 496991 51843 497014
rect 32570 496990 51843 496991
rect 34053 496759 34373 496760
rect 34053 496441 34054 496759
rect 34372 496441 34373 496759
rect 34053 496440 34373 496441
rect 358691 495311 403637 495631
rect 32570 494309 51843 494310
rect 32570 493991 32571 494309
rect 32889 494286 51843 494309
rect 32889 494014 51547 494286
rect 51819 494014 51843 494286
rect 32889 493991 51843 494014
rect 32570 493990 51843 493991
rect 34053 493759 34373 493760
rect 34053 493441 34054 493759
rect 34372 493441 34373 493759
rect 34053 493440 34373 493441
rect 358691 492311 403637 492631
rect 32570 491309 51843 491310
rect 32570 490991 32571 491309
rect 32889 491286 51843 491309
rect 32889 491014 51547 491286
rect 51819 491014 51843 491286
rect 32889 490991 51843 491014
rect 32570 490990 51843 490991
rect 34053 490759 34373 490760
rect 34053 490441 34054 490759
rect 34372 490441 34373 490759
rect 34053 490440 34373 490441
rect 358691 489311 403637 489631
rect 32570 488309 51843 488310
rect 32570 487991 32571 488309
rect 32889 488286 51843 488309
rect 32889 488014 51547 488286
rect 51819 488014 51843 488286
rect 32889 487991 51843 488014
rect 32570 487990 51843 487991
rect 34053 487759 34373 487760
rect 34053 487441 34054 487759
rect 34372 487441 34373 487759
rect 34053 487440 34373 487441
rect 358691 486311 403637 486631
rect 406914 486412 406916 486413
rect 32570 485309 51843 485310
rect 32570 484991 32571 485309
rect 32889 485286 51843 485309
rect 32889 485014 51547 485286
rect 51819 485014 51843 485286
rect 32889 484991 51843 485014
rect 32570 484990 51843 484991
rect 34053 484759 34373 484760
rect 34053 484441 34054 484759
rect 34372 484441 34373 484759
rect 34053 484440 34373 484441
rect 406915 483942 406916 486412
rect 406914 483941 406916 483942
rect 358691 483311 403637 483631
rect 32570 482309 51843 482310
rect 32570 481991 32571 482309
rect 32889 482286 51843 482309
rect 32889 482014 51547 482286
rect 51819 482014 51843 482286
rect 32889 481991 51843 482014
rect 32570 481990 51843 481991
rect 34053 481759 34373 481760
rect 34053 481441 34054 481759
rect 34372 481441 34373 481759
rect 34053 481440 34373 481441
rect 358691 480311 403637 480631
rect 32570 479309 51843 479310
rect 32570 478991 32571 479309
rect 32889 479286 51843 479309
rect 32889 479014 51547 479286
rect 51819 479014 51843 479286
rect 32889 478991 51843 479014
rect 32570 478990 51843 478991
rect 34053 478759 34373 478760
rect 34053 478441 34054 478759
rect 34372 478441 34373 478759
rect 34053 478440 34373 478441
rect 358691 477311 403637 477631
rect 32570 476309 51843 476310
rect 32570 475991 32571 476309
rect 32889 476286 51843 476309
rect 32889 476014 51547 476286
rect 51819 476014 51843 476286
rect 32889 475991 51843 476014
rect 32570 475990 51843 475991
rect 34053 475759 34373 475760
rect 34053 475441 34054 475759
rect 34372 475441 34373 475759
rect 34053 475440 34373 475441
rect 358691 474311 403637 474631
rect 32570 473309 51843 473310
rect 32570 472991 32571 473309
rect 32889 473286 51843 473309
rect 32889 473014 51547 473286
rect 51819 473014 51843 473286
rect 32889 472991 51843 473014
rect 32570 472990 51843 472991
rect 34053 472759 34373 472760
rect 34053 472441 34054 472759
rect 34372 472441 34373 472759
rect 34053 472440 34373 472441
rect 358691 471311 403637 471631
rect 32570 470309 51843 470310
rect 32570 469991 32571 470309
rect 32889 470286 51843 470309
rect 32889 470014 51547 470286
rect 51819 470014 51843 470286
rect 32889 469991 51843 470014
rect 32570 469990 51843 469991
rect 34053 469759 34373 469760
rect 34053 469441 34054 469759
rect 34372 469441 34373 469759
rect 34053 469440 34373 469441
rect 358691 468311 403637 468631
rect 32570 467309 51843 467310
rect 32570 466991 32571 467309
rect 32889 467286 51843 467309
rect 32889 467014 51547 467286
rect 51819 467014 51843 467286
rect 32889 466991 51843 467014
rect 32570 466990 51843 466991
rect 34053 466759 34373 466760
rect 34053 466441 34054 466759
rect 34372 466441 34373 466759
rect 34053 466440 34373 466441
rect 358691 465311 403637 465631
rect 32570 464309 51843 464310
rect 32570 463991 32571 464309
rect 32889 464286 51843 464309
rect 32889 464014 51547 464286
rect 51819 464014 51843 464286
rect 32889 463991 51843 464014
rect 32570 463990 51843 463991
rect 34053 463759 34373 463760
rect 34053 463441 34054 463759
rect 34372 463441 34373 463759
rect 34053 463440 34373 463441
rect 358691 462311 403637 462631
rect 32570 461309 51843 461310
rect 32570 460991 32571 461309
rect 32889 461286 51843 461309
rect 32889 461014 51547 461286
rect 51819 461014 51843 461286
rect 32889 460991 51843 461014
rect 32570 460990 51843 460991
rect 34053 460759 34373 460760
rect 34053 460441 34054 460759
rect 34372 460441 34373 460759
rect 34053 460440 34373 460441
rect 358691 459311 403637 459631
rect 32570 458309 51843 458310
rect 32570 457991 32571 458309
rect 32889 458286 51843 458309
rect 32889 458014 51547 458286
rect 51819 458014 51843 458286
rect 32889 457991 51843 458014
rect 32570 457990 51843 457991
rect 34053 457759 34373 457760
rect 34053 457441 34054 457759
rect 34372 457441 34373 457759
rect 34053 457440 34373 457441
rect 358691 456311 403637 456631
rect 32570 455309 51843 455310
rect 32570 454991 32571 455309
rect 32889 455286 51843 455309
rect 32889 455014 51547 455286
rect 51819 455014 51843 455286
rect 32889 454991 51843 455014
rect 32570 454990 51843 454991
rect 34053 454759 34373 454760
rect 34053 454441 34054 454759
rect 34372 454441 34373 454759
rect 34053 454440 34373 454441
rect 358691 453311 403637 453631
rect 32570 452309 51843 452310
rect 32570 451991 32571 452309
rect 32889 452286 51843 452309
rect 32889 452014 51547 452286
rect 51819 452014 51843 452286
rect 32889 451991 51843 452014
rect 32570 451990 51843 451991
rect 34053 451759 34373 451760
rect 34053 451441 34054 451759
rect 34372 451441 34373 451759
rect 34053 451440 34373 451441
rect 358691 450311 403637 450631
rect 406935 449967 406937 449968
rect 32570 449309 51843 449310
rect 32570 448991 32571 449309
rect 32889 449286 51843 449309
rect 32889 449014 51547 449286
rect 51819 449014 51843 449286
rect 32889 448991 51843 449014
rect 32570 448990 51843 448991
rect 34053 448759 34373 448760
rect 34053 448441 34054 448759
rect 34372 448441 34373 448759
rect 34053 448440 34373 448441
rect 358691 447311 403637 447631
rect 406936 447497 406937 449967
rect 406935 447496 406937 447497
rect 32570 446309 51843 446310
rect 32570 445991 32571 446309
rect 32889 446286 51843 446309
rect 32889 446014 51547 446286
rect 51819 446014 51843 446286
rect 32889 445991 51843 446014
rect 32570 445990 51843 445991
rect 34053 445759 34373 445760
rect 34053 445441 34054 445759
rect 34372 445441 34373 445759
rect 34053 445440 34373 445441
rect 358691 444311 403637 444631
rect 32570 443309 51843 443310
rect 32570 442991 32571 443309
rect 32889 443286 51843 443309
rect 32889 443014 51547 443286
rect 51819 443014 51843 443286
rect 32889 442991 51843 443014
rect 32570 442990 51843 442991
rect 34053 442759 34373 442760
rect 34053 442441 34054 442759
rect 34372 442441 34373 442759
rect 34053 442440 34373 442441
rect 358691 441311 403637 441631
rect 32570 440309 51843 440310
rect 32570 439991 32571 440309
rect 32889 440286 51843 440309
rect 32889 440014 51547 440286
rect 51819 440014 51843 440286
rect 32889 439991 51843 440014
rect 32570 439990 51843 439991
rect 34053 439759 34373 439760
rect 34053 439441 34054 439759
rect 34372 439441 34373 439759
rect 34053 439440 34373 439441
rect 358691 438311 403637 438631
rect 32570 437309 51843 437310
rect 32570 436991 32571 437309
rect 32889 437286 51843 437309
rect 32889 437014 51547 437286
rect 51819 437014 51843 437286
rect 32889 436991 51843 437014
rect 32570 436990 51843 436991
rect 34053 436759 34373 436760
rect 34053 436441 34054 436759
rect 34372 436441 34373 436759
rect 34053 436440 34373 436441
rect 358691 435311 403637 435631
rect 32570 434309 51843 434310
rect 32570 433991 32571 434309
rect 32889 434286 51843 434309
rect 32889 434014 51547 434286
rect 51819 434014 51843 434286
rect 32889 433991 51843 434014
rect 32570 433990 51843 433991
rect 34053 433759 34373 433760
rect 34053 433441 34054 433759
rect 34372 433441 34373 433759
rect 34053 433440 34373 433441
rect 358691 432311 403637 432631
rect 32570 431309 51843 431310
rect 32570 430991 32571 431309
rect 32889 431286 51843 431309
rect 32889 431014 51547 431286
rect 51819 431014 51843 431286
rect 32889 430991 51843 431014
rect 32570 430990 51843 430991
rect 34053 430759 34373 430760
rect 34053 430441 34054 430759
rect 34372 430441 34373 430759
rect 34053 430440 34373 430441
rect 358691 429311 403637 429631
rect 32570 428309 51843 428310
rect 32570 427991 32571 428309
rect 32889 428286 51843 428309
rect 32889 428014 51547 428286
rect 51819 428014 51843 428286
rect 32889 427991 51843 428014
rect 32570 427990 51843 427991
rect 34053 427759 34373 427760
rect 34053 427441 34054 427759
rect 34372 427441 34373 427759
rect 34053 427440 34373 427441
rect 358691 426311 403637 426631
rect 32570 425309 51843 425310
rect 32570 424991 32571 425309
rect 32889 425286 51843 425309
rect 32889 425014 51547 425286
rect 51819 425014 51843 425286
rect 32889 424991 51843 425014
rect 32570 424990 51843 424991
rect 34053 424759 34373 424760
rect 34053 424441 34054 424759
rect 34372 424441 34373 424759
rect 34053 424440 34373 424441
rect 358691 423311 403637 423631
rect 32570 422309 51843 422310
rect 32570 421991 32571 422309
rect 32889 422286 51843 422309
rect 32889 422014 51547 422286
rect 51819 422014 51843 422286
rect 32889 421991 51843 422014
rect 32570 421990 51843 421991
rect 34053 421759 34373 421760
rect 34053 421441 34054 421759
rect 34372 421441 34373 421759
rect 34053 421440 34373 421441
rect 407267 421584 407269 421585
rect 358691 420311 403637 420631
rect 32570 419309 51843 419310
rect 32570 418991 32571 419309
rect 32889 419286 51843 419309
rect 32889 419014 51547 419286
rect 51819 419014 51843 419286
rect 407268 419114 407269 421584
rect 407267 419113 407269 419114
rect 32889 418991 51843 419014
rect 32570 418990 51843 418991
rect 34053 418759 34373 418760
rect 34053 418441 34054 418759
rect 34372 418441 34373 418759
rect 34053 418440 34373 418441
rect 358691 417311 403637 417631
rect 32570 416309 51843 416310
rect 32570 415991 32571 416309
rect 32889 416286 51843 416309
rect 32889 416014 51547 416286
rect 51819 416014 51843 416286
rect 32889 415991 51843 416014
rect 32570 415990 51843 415991
rect 34053 415759 34373 415760
rect 34053 415441 34054 415759
rect 34372 415441 34373 415759
rect 34053 415440 34373 415441
rect 358691 414311 403637 414631
rect 32570 413309 51843 413310
rect 32570 412991 32571 413309
rect 32889 413286 51843 413309
rect 32889 413014 51547 413286
rect 51819 413014 51843 413286
rect 32889 412991 51843 413014
rect 32570 412990 51843 412991
rect 34053 412759 34373 412760
rect 34053 412441 34054 412759
rect 34372 412441 34373 412759
rect 34053 412440 34373 412441
rect 358691 411311 403637 411631
rect 32570 410309 51843 410310
rect 32570 409991 32571 410309
rect 32889 410286 51843 410309
rect 32889 410014 51547 410286
rect 51819 410014 51843 410286
rect 32889 409991 51843 410014
rect 32570 409990 51843 409991
rect 34053 409759 34373 409760
rect 34053 409441 34054 409759
rect 34372 409441 34373 409759
rect 34053 409440 34373 409441
rect 407033 409696 407035 409697
rect 358691 408311 403637 408631
rect 32570 407309 51843 407310
rect 32570 406991 32571 407309
rect 32889 407286 51843 407309
rect 32889 407014 51547 407286
rect 51819 407014 51843 407286
rect 407034 407226 407035 409696
rect 407033 407225 407035 407226
rect 32889 406991 51843 407014
rect 32570 406990 51843 406991
rect 34053 406759 34373 406760
rect 34053 406441 34054 406759
rect 34372 406441 34373 406759
rect 34053 406440 34373 406441
rect 358691 405311 403637 405631
rect 32570 404309 51843 404310
rect 32570 403991 32571 404309
rect 32889 404286 51843 404309
rect 32889 404014 51547 404286
rect 51819 404014 51843 404286
rect 32889 403991 51843 404014
rect 32570 403990 51843 403991
rect 34053 403759 34373 403760
rect 34053 403441 34054 403759
rect 34372 403441 34373 403759
rect 34053 403440 34373 403441
rect 358691 402311 403637 402631
rect 32570 401309 51843 401310
rect 32570 400991 32571 401309
rect 32889 401286 51843 401309
rect 32889 401014 51547 401286
rect 51819 401014 51843 401286
rect 32889 400991 51843 401014
rect 32570 400990 51843 400991
rect 358691 399311 403637 399631
rect 32570 398309 51843 398310
rect 32570 397991 32571 398309
rect 32889 398286 51843 398309
rect 32889 398014 51547 398286
rect 51819 398014 51843 398286
rect 32889 397991 51843 398014
rect 32570 397990 51843 397991
rect 34053 397759 34373 397760
rect 34053 397441 34054 397759
rect 34372 397441 34373 397759
rect 34053 397440 34373 397441
rect 358691 396311 403637 396631
rect 32570 395309 51843 395310
rect 32570 394991 32571 395309
rect 32889 395286 51843 395309
rect 32889 395014 51547 395286
rect 51819 395014 51843 395286
rect 32889 394991 51843 395014
rect 32570 394990 51843 394991
rect 34053 394759 34373 394760
rect 34053 394441 34054 394759
rect 34372 394441 34373 394759
rect 34053 394440 34373 394441
rect 358691 393311 403637 393631
rect 32570 392309 51843 392310
rect 32570 391991 32571 392309
rect 32889 392286 51843 392309
rect 32889 392014 51547 392286
rect 51819 392014 51843 392286
rect 32889 391991 51843 392014
rect 32570 391990 51843 391991
rect 34053 391759 34373 391760
rect 34053 391441 34054 391759
rect 34372 391441 34373 391759
rect 34053 391440 34373 391441
rect 358691 390311 403637 390631
rect 32570 389309 51843 389310
rect 32570 388991 32571 389309
rect 32889 389286 51843 389309
rect 32889 389014 51547 389286
rect 51819 389014 51843 389286
rect 32889 388991 51843 389014
rect 32570 388990 51843 388991
rect 34053 388759 34373 388760
rect 34053 388441 34054 388759
rect 34372 388441 34373 388759
rect 34053 388440 34373 388441
rect 358691 387311 403637 387631
rect 32570 386309 51843 386310
rect 32570 385991 32571 386309
rect 32889 386286 51843 386309
rect 32889 386014 51547 386286
rect 51819 386014 51843 386286
rect 32889 385991 51843 386014
rect 32570 385990 51843 385991
rect 34053 385759 34373 385760
rect 34053 385441 34054 385759
rect 34372 385441 34373 385759
rect 34053 385440 34373 385441
rect 358691 384311 403637 384631
rect 32570 383309 51843 383310
rect 32570 382991 32571 383309
rect 32889 383286 51843 383309
rect 32889 383014 51547 383286
rect 51819 383014 51843 383286
rect 32889 382991 51843 383014
rect 32570 382990 51843 382991
rect 34053 382759 34373 382760
rect 34053 382441 34054 382759
rect 34372 382441 34373 382759
rect 34053 382440 34373 382441
rect 358691 381311 403637 381631
rect 32570 380309 51843 380310
rect 32570 379991 32571 380309
rect 32889 380286 51843 380309
rect 32889 380014 51547 380286
rect 51819 380014 51843 380286
rect 32889 379991 51843 380014
rect 32570 379990 51843 379991
rect 34053 379759 34373 379760
rect 34053 379441 34054 379759
rect 34372 379441 34373 379759
rect 34053 379440 34373 379441
rect 358691 378311 403637 378631
rect 32570 377309 51843 377310
rect 32570 376991 32571 377309
rect 32889 377286 51843 377309
rect 32889 377014 51547 377286
rect 51819 377014 51843 377286
rect 32889 376991 51843 377014
rect 32570 376990 51843 376991
rect 34053 376759 34373 376760
rect 34053 376441 34054 376759
rect 34372 376441 34373 376759
rect 34053 376440 34373 376441
rect 358395 375607 403637 375631
rect 358395 375335 358419 375607
rect 358691 375335 403637 375607
rect 358395 375311 403637 375335
rect 32570 374309 51843 374310
rect 32570 373991 32571 374309
rect 32889 374286 51843 374309
rect 32889 374014 51547 374286
rect 51819 374014 51843 374286
rect 32889 373991 51843 374014
rect 32570 373990 51843 373991
rect 34053 373759 34373 373760
rect 34053 373441 34054 373759
rect 34372 373441 34373 373759
rect 34053 373440 34373 373441
rect 32570 371309 51843 371310
rect 32570 370991 32571 371309
rect 32889 371286 51843 371309
rect 32889 371014 51547 371286
rect 51819 371014 51843 371286
rect 32889 370991 51843 371014
rect 32570 370990 51843 370991
rect 34053 370759 34373 370760
rect 34053 370441 34054 370759
rect 34372 370441 34373 370759
rect 34053 370440 34373 370441
rect 32570 368309 51843 368310
rect 32570 367991 32571 368309
rect 32889 368286 51843 368309
rect 32889 368014 51547 368286
rect 51819 368014 51843 368286
rect 32889 367991 51843 368014
rect 32570 367990 51843 367991
rect 34053 367759 34373 367760
rect 34053 367441 34054 367759
rect 34372 367441 34373 367759
rect 34053 367440 34373 367441
rect 408464 367222 409289 661830
rect 424844 656028 425014 656029
rect 424844 655860 424845 656028
rect 425013 655860 425014 656028
rect 417401 644584 417403 644585
rect 417402 639784 417403 644584
rect 417401 639783 417403 639784
rect 417268 634584 417270 634585
rect 417269 629784 417270 634584
rect 417268 629783 417270 629784
rect 413052 596862 415512 596863
rect 413052 594404 413053 596862
rect 415511 594404 415512 596862
rect 413052 594403 415512 594404
rect 413052 523278 415512 523279
rect 413052 520820 413053 523278
rect 415511 520820 415512 523278
rect 413052 520819 415512 520820
rect 413052 497294 415512 497295
rect 413052 494836 413053 497294
rect 415511 494836 415512 497294
rect 413052 494835 415512 494836
rect 413052 465330 415512 465331
rect 413052 462872 413053 465330
rect 415511 462872 415512 465330
rect 413052 462871 415512 462872
rect 413052 435897 415512 435898
rect 413052 433439 413053 435897
rect 415511 433439 415512 435897
rect 413052 433438 415512 433439
rect 413052 399794 415512 399795
rect 413052 397336 413053 399794
rect 415511 397336 415512 399794
rect 413052 397335 415512 397336
rect 413052 385767 415512 385768
rect 413052 383309 413053 385767
rect 415511 383309 415512 385767
rect 413052 383308 415512 383309
rect 395276 366397 409289 367222
rect 32570 365309 51843 365310
rect 32570 364991 32571 365309
rect 32889 365286 51843 365309
rect 32889 365014 51547 365286
rect 51819 365014 51843 365286
rect 32889 364991 51843 365014
rect 32570 364990 51843 364991
rect 34053 364759 34373 364760
rect 34053 364441 34054 364759
rect 34372 364441 34373 364759
rect 34053 364440 34373 364441
rect 53818 364727 54138 364728
rect 53818 364409 53819 364727
rect 54137 364409 54138 364727
rect 53818 364408 54138 364409
rect 32570 362309 51843 362310
rect 32570 361991 32571 362309
rect 32889 362286 51843 362309
rect 32889 362014 51547 362286
rect 51819 362014 51843 362286
rect 32889 361991 51843 362014
rect 32570 361990 51843 361991
rect 406979 362180 406981 362181
rect 406980 359710 406981 362180
rect 406979 359709 406981 359710
rect 45905 358331 46015 358342
rect 31813 358221 50244 358331
rect 26654 353284 26656 353285
rect 26654 350814 26655 353284
rect 26654 350813 26656 350814
rect 26580 348755 26582 348756
rect 26580 346285 26581 348755
rect 26580 346284 26582 346285
rect 26580 344245 26582 344246
rect 26580 341775 26581 344245
rect 26580 341774 26582 341775
rect 45905 333339 46015 358221
rect 55307 345755 55627 345756
rect 55307 345437 55308 345755
rect 55626 345437 55627 345755
rect 55307 345436 55627 345437
rect 58307 345755 58627 345756
rect 58307 345437 58308 345755
rect 58626 345437 58627 345755
rect 58307 345436 58627 345437
rect 61307 345755 61627 345756
rect 61307 345437 61308 345755
rect 61626 345437 61627 345755
rect 61307 345436 61627 345437
rect 64307 345755 64627 345756
rect 64307 345437 64308 345755
rect 64626 345437 64627 345755
rect 64307 345436 64627 345437
rect 67307 345755 67627 345756
rect 67307 345437 67308 345755
rect 67626 345437 67627 345755
rect 67307 345436 67627 345437
rect 70307 345755 70627 345756
rect 70307 345437 70308 345755
rect 70626 345437 70627 345755
rect 70307 345436 70627 345437
rect 73307 345755 73627 345756
rect 73307 345437 73308 345755
rect 73626 345437 73627 345755
rect 73307 345436 73627 345437
rect 76307 345755 76627 345756
rect 76307 345437 76308 345755
rect 76626 345437 76627 345755
rect 76307 345436 76627 345437
rect 79307 345755 79627 345756
rect 79307 345437 79308 345755
rect 79626 345437 79627 345755
rect 79307 345436 79627 345437
rect 82307 345755 82627 345756
rect 82307 345437 82308 345755
rect 82626 345437 82627 345755
rect 82307 345436 82627 345437
rect 85307 345755 85627 345756
rect 85307 345437 85308 345755
rect 85626 345437 85627 345755
rect 85307 345436 85627 345437
rect 88307 345755 88627 345756
rect 88307 345437 88308 345755
rect 88626 345437 88627 345755
rect 88307 345436 88627 345437
rect 91307 345755 91627 345756
rect 91307 345437 91308 345755
rect 91626 345437 91627 345755
rect 91307 345436 91627 345437
rect 94307 345755 94627 345756
rect 94307 345437 94308 345755
rect 94626 345437 94627 345755
rect 94307 345436 94627 345437
rect 97307 345755 97627 345756
rect 97307 345437 97308 345755
rect 97626 345437 97627 345755
rect 97307 345436 97627 345437
rect 100307 345755 100627 345756
rect 100307 345437 100308 345755
rect 100626 345437 100627 345755
rect 100307 345436 100627 345437
rect 103307 345755 103627 345756
rect 103307 345437 103308 345755
rect 103626 345437 103627 345755
rect 103307 345436 103627 345437
rect 106307 345755 106627 345756
rect 106307 345437 106308 345755
rect 106626 345437 106627 345755
rect 106307 345436 106627 345437
rect 109307 345755 109627 345756
rect 109307 345437 109308 345755
rect 109626 345437 109627 345755
rect 109307 345436 109627 345437
rect 112307 345755 112627 345756
rect 112307 345437 112308 345755
rect 112626 345437 112627 345755
rect 112307 345436 112627 345437
rect 115307 345755 115627 345756
rect 115307 345437 115308 345755
rect 115626 345437 115627 345755
rect 115307 345436 115627 345437
rect 118307 345755 118627 345756
rect 118307 345437 118308 345755
rect 118626 345437 118627 345755
rect 118307 345436 118627 345437
rect 121307 345755 121627 345756
rect 121307 345437 121308 345755
rect 121626 345437 121627 345755
rect 121307 345436 121627 345437
rect 124307 345755 124627 345756
rect 124307 345437 124308 345755
rect 124626 345437 124627 345755
rect 124307 345436 124627 345437
rect 127307 345755 127627 345756
rect 127307 345437 127308 345755
rect 127626 345437 127627 345755
rect 127307 345436 127627 345437
rect 130307 345755 130627 345756
rect 130307 345437 130308 345755
rect 130626 345437 130627 345755
rect 130307 345436 130627 345437
rect 133307 345755 133627 345756
rect 133307 345437 133308 345755
rect 133626 345437 133627 345755
rect 133307 345436 133627 345437
rect 136307 345755 136627 345756
rect 136307 345437 136308 345755
rect 136626 345437 136627 345755
rect 136307 345436 136627 345437
rect 139307 345755 139627 345756
rect 139307 345437 139308 345755
rect 139626 345437 139627 345755
rect 139307 345436 139627 345437
rect 142307 345755 142627 345756
rect 142307 345437 142308 345755
rect 142626 345437 142627 345755
rect 142307 345436 142627 345437
rect 145307 345755 145627 345756
rect 145307 345437 145308 345755
rect 145626 345437 145627 345755
rect 145307 345436 145627 345437
rect 148307 345755 148627 345756
rect 148307 345437 148308 345755
rect 148626 345437 148627 345755
rect 148307 345436 148627 345437
rect 151307 345755 151627 345756
rect 151307 345437 151308 345755
rect 151626 345437 151627 345755
rect 151307 345436 151627 345437
rect 154307 345755 154627 345756
rect 154307 345437 154308 345755
rect 154626 345437 154627 345755
rect 154307 345436 154627 345437
rect 157307 345755 157627 345756
rect 157307 345437 157308 345755
rect 157626 345437 157627 345755
rect 157307 345436 157627 345437
rect 160307 345755 160627 345756
rect 160307 345437 160308 345755
rect 160626 345437 160627 345755
rect 160307 345436 160627 345437
rect 163307 345755 163627 345756
rect 163307 345437 163308 345755
rect 163626 345437 163627 345755
rect 163307 345436 163627 345437
rect 166307 345755 166627 345756
rect 166307 345437 166308 345755
rect 166626 345437 166627 345755
rect 166307 345436 166627 345437
rect 169307 345755 169627 345756
rect 169307 345437 169308 345755
rect 169626 345437 169627 345755
rect 169307 345436 169627 345437
rect 172307 345755 172627 345756
rect 172307 345437 172308 345755
rect 172626 345437 172627 345755
rect 172307 345436 172627 345437
rect 175307 345755 175627 345756
rect 175307 345437 175308 345755
rect 175626 345437 175627 345755
rect 175307 345436 175627 345437
rect 178307 345755 178627 345756
rect 178307 345437 178308 345755
rect 178626 345437 178627 345755
rect 178307 345436 178627 345437
rect 181307 345755 181627 345756
rect 181307 345437 181308 345755
rect 181626 345437 181627 345755
rect 181307 345436 181627 345437
rect 184307 345755 184627 345756
rect 184307 345437 184308 345755
rect 184626 345437 184627 345755
rect 184307 345436 184627 345437
rect 187307 345755 187627 345756
rect 187307 345437 187308 345755
rect 187626 345437 187627 345755
rect 187307 345436 187627 345437
rect 190307 345755 190627 345756
rect 190307 345437 190308 345755
rect 190626 345437 190627 345755
rect 190307 345436 190627 345437
rect 193307 345755 193627 345756
rect 193307 345437 193308 345755
rect 193626 345437 193627 345755
rect 193307 345436 193627 345437
rect 196307 345755 196627 345756
rect 196307 345437 196308 345755
rect 196626 345437 196627 345755
rect 196307 345436 196627 345437
rect 199307 345755 199627 345756
rect 199307 345437 199308 345755
rect 199626 345437 199627 345755
rect 199307 345436 199627 345437
rect 202307 345755 202627 345756
rect 202307 345437 202308 345755
rect 202626 345437 202627 345755
rect 202307 345436 202627 345437
rect 205307 345755 205627 345756
rect 205307 345437 205308 345755
rect 205626 345437 205627 345755
rect 205307 345436 205627 345437
rect 208307 345755 208627 345756
rect 208307 345437 208308 345755
rect 208626 345437 208627 345755
rect 208307 345436 208627 345437
rect 211307 345755 211627 345756
rect 211307 345437 211308 345755
rect 211626 345437 211627 345755
rect 211307 345436 211627 345437
rect 214307 345755 214627 345756
rect 214307 345437 214308 345755
rect 214626 345437 214627 345755
rect 214307 345436 214627 345437
rect 217307 345755 217627 345756
rect 217307 345437 217308 345755
rect 217626 345437 217627 345755
rect 217307 345436 217627 345437
rect 220307 345755 220627 345756
rect 220307 345437 220308 345755
rect 220626 345437 220627 345755
rect 220307 345436 220627 345437
rect 223307 345755 223627 345756
rect 223307 345437 223308 345755
rect 223626 345437 223627 345755
rect 223307 345436 223627 345437
rect 226307 345755 226627 345756
rect 226307 345437 226308 345755
rect 226626 345437 226627 345755
rect 226307 345436 226627 345437
rect 229307 345755 229627 345756
rect 229307 345437 229308 345755
rect 229626 345437 229627 345755
rect 229307 345436 229627 345437
rect 232307 345755 232627 345756
rect 232307 345437 232308 345755
rect 232626 345437 232627 345755
rect 232307 345436 232627 345437
rect 235307 345755 235627 345756
rect 235307 345437 235308 345755
rect 235626 345437 235627 345755
rect 235307 345436 235627 345437
rect 238307 345755 238627 345756
rect 238307 345437 238308 345755
rect 238626 345437 238627 345755
rect 238307 345436 238627 345437
rect 241307 345755 241627 345756
rect 241307 345437 241308 345755
rect 241626 345437 241627 345755
rect 241307 345436 241627 345437
rect 244307 345755 244627 345756
rect 244307 345437 244308 345755
rect 244626 345437 244627 345755
rect 244307 345436 244627 345437
rect 247307 345755 247627 345756
rect 247307 345437 247308 345755
rect 247626 345437 247627 345755
rect 247307 345436 247627 345437
rect 250307 345755 250627 345756
rect 250307 345437 250308 345755
rect 250626 345437 250627 345755
rect 250307 345436 250627 345437
rect 253307 345755 253627 345756
rect 253307 345437 253308 345755
rect 253626 345437 253627 345755
rect 253307 345436 253627 345437
rect 256307 345755 256627 345756
rect 256307 345437 256308 345755
rect 256626 345437 256627 345755
rect 256307 345436 256627 345437
rect 259307 345755 259627 345756
rect 259307 345437 259308 345755
rect 259626 345437 259627 345755
rect 259307 345436 259627 345437
rect 262307 345755 262627 345756
rect 262307 345437 262308 345755
rect 262626 345437 262627 345755
rect 262307 345436 262627 345437
rect 265307 345755 265627 345756
rect 265307 345437 265308 345755
rect 265626 345437 265627 345755
rect 265307 345436 265627 345437
rect 268307 345755 268627 345756
rect 268307 345437 268308 345755
rect 268626 345437 268627 345755
rect 268307 345436 268627 345437
rect 271307 345755 271627 345756
rect 271307 345437 271308 345755
rect 271626 345437 271627 345755
rect 271307 345436 271627 345437
rect 274307 345755 274627 345756
rect 274307 345437 274308 345755
rect 274626 345437 274627 345755
rect 274307 345436 274627 345437
rect 277307 345755 277627 345756
rect 277307 345437 277308 345755
rect 277626 345437 277627 345755
rect 277307 345436 277627 345437
rect 280307 345755 280627 345756
rect 280307 345437 280308 345755
rect 280626 345437 280627 345755
rect 280307 345436 280627 345437
rect 283307 345755 283627 345756
rect 283307 345437 283308 345755
rect 283626 345437 283627 345755
rect 283307 345436 283627 345437
rect 286307 345755 286627 345756
rect 286307 345437 286308 345755
rect 286626 345437 286627 345755
rect 286307 345436 286627 345437
rect 289307 345755 289627 345756
rect 289307 345437 289308 345755
rect 289626 345437 289627 345755
rect 289307 345436 289627 345437
rect 292307 345755 292627 345756
rect 292307 345437 292308 345755
rect 292626 345437 292627 345755
rect 292307 345436 292627 345437
rect 295307 345755 295627 345756
rect 295307 345437 295308 345755
rect 295626 345437 295627 345755
rect 295307 345436 295627 345437
rect 298307 345755 298627 345756
rect 298307 345437 298308 345755
rect 298626 345437 298627 345755
rect 298307 345436 298627 345437
rect 301307 345755 301627 345756
rect 301307 345437 301308 345755
rect 301626 345437 301627 345755
rect 301307 345436 301627 345437
rect 304307 345755 304627 345756
rect 304307 345437 304308 345755
rect 304626 345437 304627 345755
rect 304307 345436 304627 345437
rect 307307 345755 307627 345756
rect 307307 345437 307308 345755
rect 307626 345437 307627 345755
rect 307307 345436 307627 345437
rect 310307 345755 310627 345756
rect 310307 345437 310308 345755
rect 310626 345437 310627 345755
rect 310307 345436 310627 345437
rect 313307 345755 313627 345756
rect 313307 345437 313308 345755
rect 313626 345437 313627 345755
rect 313307 345436 313627 345437
rect 316307 345755 316627 345756
rect 316307 345437 316308 345755
rect 316626 345437 316627 345755
rect 316307 345436 316627 345437
rect 319307 345755 319627 345756
rect 319307 345437 319308 345755
rect 319626 345437 319627 345755
rect 319307 345436 319627 345437
rect 325307 345755 325627 345756
rect 325307 345437 325308 345755
rect 325626 345437 325627 345755
rect 325307 345436 325627 345437
rect 328307 345755 328627 345756
rect 328307 345437 328308 345755
rect 328626 345437 328627 345755
rect 328307 345436 328627 345437
rect 331307 345755 331627 345756
rect 331307 345437 331308 345755
rect 331626 345437 331627 345755
rect 331307 345436 331627 345437
rect 334307 345755 334627 345756
rect 334307 345437 334308 345755
rect 334626 345437 334627 345755
rect 334307 345436 334627 345437
rect 337307 345755 337627 345756
rect 337307 345437 337308 345755
rect 337626 345437 337627 345755
rect 337307 345436 337627 345437
rect 340307 345755 340627 345756
rect 340307 345437 340308 345755
rect 340626 345437 340627 345755
rect 340307 345436 340627 345437
rect 343307 345755 343627 345756
rect 343307 345437 343308 345755
rect 343626 345437 343627 345755
rect 343307 345436 343627 345437
rect 346307 345755 346627 345756
rect 346307 345437 346308 345755
rect 346626 345437 346627 345755
rect 346307 345436 346627 345437
rect 349307 345755 349627 345756
rect 349307 345437 349308 345755
rect 349626 345437 349627 345755
rect 349307 345436 349627 345437
rect 352307 345755 352627 345756
rect 352307 345437 352308 345755
rect 352626 345437 352627 345755
rect 352307 345436 352627 345437
rect 355307 345755 355627 345756
rect 355307 345437 355308 345755
rect 355626 345437 355627 345755
rect 355307 345436 355627 345437
rect 358307 345755 358627 345756
rect 358307 345437 358308 345755
rect 358626 345437 358627 345755
rect 358307 345436 358627 345437
rect 29741 333229 46015 333339
rect 12506 253173 12620 253174
rect 12506 253061 12507 253173
rect 12619 253061 12620 253173
rect 12506 253060 12620 253061
rect 12507 201638 12619 253060
rect 15357 201638 15577 201898
rect 12507 201526 15843 201638
rect 10673 191537 10785 191538
rect 10673 191427 10674 191537
rect 10784 191427 10785 191537
rect 10673 191426 10785 191427
rect 9010 191342 9132 191343
rect 9010 191232 9011 191342
rect 9131 191232 9132 191342
rect 9010 191231 9132 191232
rect 1919 176552 13873 177800
rect 1919 164695 3527 176552
rect 2175 164594 3527 164695
rect 12521 164594 13873 176552
rect 15357 172531 15577 201526
rect 29741 179969 29851 333229
rect 55301 323422 55633 323423
rect 55301 323421 55302 323422
rect 55632 323421 55633 323422
rect 58301 323422 58633 323423
rect 58301 323421 58302 323422
rect 58632 323421 58633 323422
rect 61301 323422 61633 323423
rect 61301 323421 61302 323422
rect 61632 323421 61633 323422
rect 64301 323422 64633 323423
rect 64301 323421 64302 323422
rect 64632 323421 64633 323422
rect 67301 323422 67633 323423
rect 67301 323421 67302 323422
rect 67632 323421 67633 323422
rect 70301 323422 70633 323423
rect 70301 323421 70302 323422
rect 70632 323421 70633 323422
rect 73301 323422 73633 323423
rect 73301 323421 73302 323422
rect 73632 323421 73633 323422
rect 76301 323422 76633 323423
rect 76301 323421 76302 323422
rect 76632 323421 76633 323422
rect 79301 323422 79633 323423
rect 79301 323421 79302 323422
rect 79632 323421 79633 323422
rect 82301 323422 82633 323423
rect 82301 323421 82302 323422
rect 82632 323421 82633 323422
rect 85301 323422 85633 323423
rect 85301 323421 85302 323422
rect 85632 323421 85633 323422
rect 88301 323422 88633 323423
rect 88301 323421 88302 323422
rect 88632 323421 88633 323422
rect 91301 323422 91633 323423
rect 91301 323421 91302 323422
rect 91632 323421 91633 323422
rect 94301 323422 94633 323423
rect 94301 323421 94302 323422
rect 94632 323421 94633 323422
rect 97301 323422 97633 323423
rect 97301 323421 97302 323422
rect 97632 323421 97633 323422
rect 100301 323422 100633 323423
rect 100301 323421 100302 323422
rect 100632 323421 100633 323422
rect 103301 323422 103633 323423
rect 103301 323421 103302 323422
rect 103632 323421 103633 323422
rect 106301 323422 106633 323423
rect 106301 323421 106302 323422
rect 106632 323421 106633 323422
rect 109301 323422 109633 323423
rect 109301 323421 109302 323422
rect 109632 323421 109633 323422
rect 112301 323422 112633 323423
rect 112301 323421 112302 323422
rect 112632 323421 112633 323422
rect 115301 323422 115633 323423
rect 115301 323421 115302 323422
rect 115632 323421 115633 323422
rect 118301 323422 118633 323423
rect 118301 323421 118302 323422
rect 118632 323421 118633 323422
rect 121301 323422 121633 323423
rect 121301 323421 121302 323422
rect 121632 323421 121633 323422
rect 124301 323422 124633 323423
rect 124301 323421 124302 323422
rect 124632 323421 124633 323422
rect 127301 323422 127633 323423
rect 127301 323421 127302 323422
rect 127632 323421 127633 323422
rect 130301 323422 130633 323423
rect 130301 323421 130302 323422
rect 130632 323421 130633 323422
rect 133301 323422 133633 323423
rect 133301 323421 133302 323422
rect 133632 323421 133633 323422
rect 136301 323422 136633 323423
rect 136301 323421 136302 323422
rect 136632 323421 136633 323422
rect 139301 323422 139633 323423
rect 139301 323421 139302 323422
rect 139632 323421 139633 323422
rect 142301 323422 142633 323423
rect 142301 323421 142302 323422
rect 142632 323421 142633 323422
rect 145301 323422 145633 323423
rect 145301 323421 145302 323422
rect 145632 323421 145633 323422
rect 148301 323422 148633 323423
rect 148301 323421 148302 323422
rect 148632 323421 148633 323422
rect 151301 323422 151633 323423
rect 151301 323421 151302 323422
rect 151632 323421 151633 323422
rect 154301 323422 154633 323423
rect 154301 323421 154302 323422
rect 154632 323421 154633 323422
rect 157301 323422 157633 323423
rect 157301 323421 157302 323422
rect 157632 323421 157633 323422
rect 160301 323422 160633 323423
rect 160301 323421 160302 323422
rect 160632 323421 160633 323422
rect 163301 323422 163633 323423
rect 163301 323421 163302 323422
rect 163632 323421 163633 323422
rect 166301 323422 166633 323423
rect 166301 323421 166302 323422
rect 166632 323421 166633 323422
rect 169301 323422 169633 323423
rect 169301 323421 169302 323422
rect 169632 323421 169633 323422
rect 172301 323422 172633 323423
rect 172301 323421 172302 323422
rect 172632 323421 172633 323422
rect 175301 323422 175633 323423
rect 175301 323421 175302 323422
rect 175632 323421 175633 323422
rect 178301 323422 178633 323423
rect 178301 323421 178302 323422
rect 178632 323421 178633 323422
rect 181301 323422 181633 323423
rect 181301 323421 181302 323422
rect 181632 323421 181633 323422
rect 184301 323422 184633 323423
rect 184301 323421 184302 323422
rect 184632 323421 184633 323422
rect 187301 323422 187633 323423
rect 187301 323421 187302 323422
rect 187632 323421 187633 323422
rect 190301 323422 190633 323423
rect 190301 323421 190302 323422
rect 190632 323421 190633 323422
rect 193301 323422 193633 323423
rect 193301 323421 193302 323422
rect 193632 323421 193633 323422
rect 196301 323422 196633 323423
rect 196301 323421 196302 323422
rect 196632 323421 196633 323422
rect 199301 323422 199633 323423
rect 199301 323421 199302 323422
rect 199632 323421 199633 323422
rect 202301 323422 202633 323423
rect 202301 323421 202302 323422
rect 202632 323421 202633 323422
rect 205301 323422 205633 323423
rect 205301 323421 205302 323422
rect 205632 323421 205633 323422
rect 208301 323422 208633 323423
rect 208301 323421 208302 323422
rect 208632 323421 208633 323422
rect 211301 323422 211633 323423
rect 211301 323421 211302 323422
rect 211632 323421 211633 323422
rect 214301 323422 214633 323423
rect 214301 323421 214302 323422
rect 214632 323421 214633 323422
rect 217301 323422 217633 323423
rect 217301 323421 217302 323422
rect 217632 323421 217633 323422
rect 220301 323422 220633 323423
rect 220301 323421 220302 323422
rect 220632 323421 220633 323422
rect 223301 323422 223633 323423
rect 223301 323421 223302 323422
rect 223632 323421 223633 323422
rect 226301 323422 226633 323423
rect 226301 323421 226302 323422
rect 226632 323421 226633 323422
rect 229301 323422 229633 323423
rect 229301 323421 229302 323422
rect 229632 323421 229633 323422
rect 232301 323422 232633 323423
rect 232301 323421 232302 323422
rect 232632 323421 232633 323422
rect 235301 323422 235633 323423
rect 235301 323421 235302 323422
rect 235632 323421 235633 323422
rect 238301 323422 238633 323423
rect 238301 323421 238302 323422
rect 238632 323421 238633 323422
rect 241301 323422 241633 323423
rect 241301 323421 241302 323422
rect 241632 323421 241633 323422
rect 244301 323422 244633 323423
rect 244301 323421 244302 323422
rect 244632 323421 244633 323422
rect 247301 323422 247633 323423
rect 247301 323421 247302 323422
rect 247632 323421 247633 323422
rect 250301 323422 250633 323423
rect 250301 323421 250302 323422
rect 250632 323421 250633 323422
rect 253301 323422 253633 323423
rect 253301 323421 253302 323422
rect 253632 323421 253633 323422
rect 256301 323422 256633 323423
rect 256301 323421 256302 323422
rect 256632 323421 256633 323422
rect 259301 323422 259633 323423
rect 259301 323421 259302 323422
rect 259632 323421 259633 323422
rect 262301 323422 262633 323423
rect 262301 323421 262302 323422
rect 262632 323421 262633 323422
rect 265301 323422 265633 323423
rect 265301 323421 265302 323422
rect 265632 323421 265633 323422
rect 268301 323422 268633 323423
rect 268301 323421 268302 323422
rect 268632 323421 268633 323422
rect 271301 323422 271633 323423
rect 271301 323421 271302 323422
rect 271632 323421 271633 323422
rect 274301 323422 274633 323423
rect 274301 323421 274302 323422
rect 274632 323421 274633 323422
rect 277301 323422 277633 323423
rect 277301 323421 277302 323422
rect 277632 323421 277633 323422
rect 280301 323422 280633 323423
rect 280301 323421 280302 323422
rect 280632 323421 280633 323422
rect 283301 323422 283633 323423
rect 283301 323421 283302 323422
rect 283632 323421 283633 323422
rect 286301 323422 286633 323423
rect 286301 323421 286302 323422
rect 286632 323421 286633 323422
rect 289301 323422 289633 323423
rect 289301 323421 289302 323422
rect 289632 323421 289633 323422
rect 292301 323422 292633 323423
rect 292301 323421 292302 323422
rect 292632 323421 292633 323422
rect 295301 323422 295633 323423
rect 295301 323421 295302 323422
rect 295632 323421 295633 323422
rect 298301 323422 298633 323423
rect 298301 323421 298302 323422
rect 298632 323421 298633 323422
rect 301301 323422 301633 323423
rect 301301 323421 301302 323422
rect 301632 323421 301633 323422
rect 304301 323422 304633 323423
rect 304301 323421 304302 323422
rect 304632 323421 304633 323422
rect 307301 323422 307633 323423
rect 307301 323421 307302 323422
rect 307632 323421 307633 323422
rect 310301 323422 310633 323423
rect 310301 323421 310302 323422
rect 310632 323421 310633 323422
rect 313301 323422 313633 323423
rect 313301 323421 313302 323422
rect 313632 323421 313633 323422
rect 316301 323422 316633 323423
rect 316301 323421 316302 323422
rect 316632 323421 316633 323422
rect 319301 323422 319633 323423
rect 319301 323421 319302 323422
rect 319632 323421 319633 323422
rect 325301 323422 325633 323423
rect 325301 323421 325302 323422
rect 325632 323421 325633 323422
rect 328301 323422 328633 323423
rect 328301 323421 328302 323422
rect 328632 323421 328633 323422
rect 331301 323422 331633 323423
rect 331301 323421 331302 323422
rect 331632 323421 331633 323422
rect 334301 323422 334633 323423
rect 334301 323421 334302 323422
rect 334632 323421 334633 323422
rect 337301 323422 337633 323423
rect 337301 323421 337302 323422
rect 337632 323421 337633 323422
rect 340301 323422 340633 323423
rect 340301 323421 340302 323422
rect 340632 323421 340633 323422
rect 343301 323422 343633 323423
rect 343301 323421 343302 323422
rect 343632 323421 343633 323422
rect 346301 323422 346633 323423
rect 346301 323421 346302 323422
rect 346632 323421 346633 323422
rect 349301 323422 349633 323423
rect 349301 323421 349302 323422
rect 349632 323421 349633 323422
rect 352301 323422 352633 323423
rect 352301 323421 352302 323422
rect 352632 323421 352633 323422
rect 355301 323422 355633 323423
rect 355301 323421 355302 323422
rect 355632 323421 355633 323422
rect 358301 323422 358633 323423
rect 358301 323421 358302 323422
rect 358632 323421 358633 323422
rect 39940 315920 39942 315921
rect 39940 313450 39941 315920
rect 39940 313449 39942 313450
rect 97424 315891 99884 315915
rect 97424 313479 97448 315891
rect 99860 313479 99884 315891
rect 69647 254006 69969 254007
rect 69647 253686 69648 254006
rect 69968 253686 69969 254006
rect 69647 253685 69969 253686
rect 69648 214521 69968 253685
rect 97424 230750 99884 313479
rect 120117 315891 122577 315915
rect 120117 313479 120141 315891
rect 122553 313479 122577 315891
rect 120117 230750 122577 313479
rect 143536 315891 145996 315915
rect 143536 313479 143560 315891
rect 145972 313479 145996 315891
rect 424844 314082 425014 655860
rect 428428 652869 430890 652870
rect 428428 650409 428429 652869
rect 430889 650409 430890 652869
rect 428428 650408 430890 650409
rect 492825 652599 495285 652600
rect 428429 627988 430889 650408
rect 492825 650141 492826 652599
rect 495284 650141 495285 652599
rect 451368 634584 456170 634585
rect 451368 634583 451369 634584
rect 456169 634583 456170 634584
rect 460693 634584 465495 634585
rect 460693 634583 460694 634584
rect 465494 634583 465495 634584
rect 428429 625530 428430 627988
rect 430888 625530 430889 627988
rect 428429 615818 430889 625530
rect 428429 613360 428430 615818
rect 430888 613360 430889 615818
rect 428429 602179 430889 613360
rect 428429 599721 428430 602179
rect 430888 599721 430889 602179
rect 428429 587352 430889 599721
rect 428429 584894 428430 587352
rect 430888 584894 430889 587352
rect 428429 566277 430889 584894
rect 428429 563819 428430 566277
rect 430888 563819 430889 566277
rect 428429 552464 430889 563819
rect 428429 550006 428430 552464
rect 430888 550006 430889 552464
rect 428429 542840 430889 550006
rect 428429 540382 428430 542840
rect 430888 540382 430889 542840
rect 428429 531892 430889 540382
rect 428429 529434 428430 531892
rect 430888 529434 430889 531892
rect 428429 512942 430889 529434
rect 428429 510484 428430 512942
rect 430888 510484 430889 512942
rect 428429 486406 430889 510484
rect 428429 483948 428430 486406
rect 430888 483948 430889 486406
rect 428429 449961 430889 483948
rect 428429 447503 428430 449961
rect 430888 447503 430889 449961
rect 428429 421578 430889 447503
rect 428429 419120 428430 421578
rect 430888 419120 430889 421578
rect 428429 409690 430889 419120
rect 428429 407232 428430 409690
rect 430888 407232 430889 409690
rect 428429 362174 430889 407232
rect 428429 359716 428430 362174
rect 430888 359716 430889 362174
rect 424843 314081 425015 314082
rect 424843 313911 424844 314081
rect 425014 313911 425015 314081
rect 424843 313910 425015 313911
rect 143536 230750 145996 313479
rect 428429 294486 430889 359716
rect 492825 230750 495285 650141
rect 86876 230749 495285 230750
rect 86876 230726 287965 230749
rect 89288 228314 287965 230726
rect 86876 228291 287965 228314
rect 290423 228291 495285 230749
rect 86876 228290 495285 228291
rect 512860 648399 554148 648400
rect 512860 647541 553289 648399
rect 554147 647541 554148 648399
rect 512860 647540 554148 647541
rect 69648 214201 142794 214521
rect 142474 198586 142794 214201
rect 156541 203679 158303 228290
rect 173401 207178 173402 207179
rect 173722 207178 173723 207179
rect 173401 207177 173723 207178
rect 170811 207060 170812 207061
rect 171132 207060 171133 207061
rect 170811 207059 171133 207060
rect 167887 206836 167888 206837
rect 168208 206836 168209 206837
rect 167887 206835 168209 206836
rect 156541 201965 156565 203679
rect 158279 201965 158303 203679
rect 156541 201941 158303 201965
rect 141920 198033 143271 198586
rect 141920 197761 142258 198033
rect 142530 197761 143271 198033
rect 141920 197302 143271 197761
rect 89090 196007 157941 196031
rect 89090 194293 156203 196007
rect 157917 194293 157941 196007
rect 89090 194269 157941 194293
rect 163189 192163 163509 205508
rect 174310 203679 176072 228290
rect 174310 201965 174334 203679
rect 176048 201965 176072 203679
rect 174310 201941 176072 201965
rect 178419 203679 180181 228290
rect 178419 201965 178443 203679
rect 180157 201965 180181 203679
rect 178419 201941 180181 201965
rect 190957 203679 192719 228290
rect 190957 201965 190981 203679
rect 192695 201965 192719 203679
rect 190957 201941 192719 201965
rect 207499 203679 209261 228290
rect 207499 201965 207523 203679
rect 209237 201965 209261 203679
rect 207499 201941 209261 201965
rect 504539 196230 504541 196231
rect 504540 193891 504541 196230
rect 504561 193890 504563 193891
rect 163189 191891 163213 192163
rect 163485 191891 163509 192163
rect 163189 191867 163509 191891
rect 167888 192186 168208 192187
rect 167888 191868 167889 192186
rect 168207 191868 168208 192186
rect 167888 191867 168208 191868
rect 170812 192186 171132 192187
rect 170812 191868 170813 192186
rect 171131 191868 171132 192186
rect 170812 191867 171132 191868
rect 173402 192186 173722 192187
rect 173402 191868 173403 192186
rect 173721 191868 173722 192186
rect 173402 191867 173722 191868
rect 33444 191536 162771 191537
rect 33444 191428 33445 191536
rect 33553 191428 162771 191536
rect 504562 191430 504563 193890
rect 504561 191429 504563 191430
rect 33444 191427 162771 191428
rect 142554 191013 164013 191037
rect 142554 190741 163717 191013
rect 163989 190741 164013 191013
rect 142554 190717 164013 190741
rect 153047 188975 163131 188999
rect 153047 188703 162835 188975
rect 163107 188703 163131 188975
rect 153047 188679 163131 188703
rect 512860 188567 513720 647540
rect 578644 222136 578646 222137
rect 578645 217336 578646 222136
rect 578644 217335 578646 217336
rect 579068 204057 579070 204058
rect 579069 199257 579070 204057
rect 579068 199256 579070 199257
rect 205113 187707 513720 188567
rect 175758 186632 175940 186633
rect 175758 186462 175759 186632
rect 175939 186462 175940 186632
rect 175758 186461 175940 186462
rect 504850 186230 504852 186231
rect 153080 185822 163131 185846
rect 153080 185550 162835 185822
rect 163107 185550 163131 185822
rect 153080 185526 163131 185550
rect 504851 183891 504852 186230
rect 505014 183890 505016 183891
rect 152814 183130 163131 183154
rect 152814 182858 162835 183130
rect 163107 182858 163131 183130
rect 152814 182834 163131 182858
rect 505015 181430 505016 183890
rect 505014 181429 505016 181430
rect 153039 180603 163161 180627
rect 153039 180331 162865 180603
rect 163137 180331 163161 180603
rect 153039 180307 163161 180331
rect 164431 180626 164751 180627
rect 164431 180308 164432 180626
rect 164750 180308 164751 180626
rect 164431 180307 164751 180308
rect 165181 179969 165291 180956
rect 29741 179859 165291 179969
rect 165881 178039 166101 181051
rect 167772 180626 168092 180627
rect 167772 180308 167773 180626
rect 168091 180308 168092 180626
rect 167772 180307 168092 180308
rect 40276 177819 166101 178039
rect 15356 172530 15578 172531
rect 15356 172310 15357 172530
rect 15577 172310 15578 172530
rect 15356 172309 15578 172310
rect 2175 163346 13873 164594
rect 13380 147234 15842 147235
rect 13380 144774 13381 147234
rect 15841 144774 15842 147234
rect 13380 144773 15842 144774
rect 13381 136508 15841 144773
rect 13381 134050 13382 136508
rect 15840 134050 15841 136508
rect 13381 124806 15841 134050
rect 13381 103327 15841 122346
rect 40276 34898 40496 177819
rect 168881 176521 169101 181111
rect 170722 180626 171042 180627
rect 170722 180308 170723 180626
rect 171041 180308 171042 180626
rect 170722 180307 171042 180308
rect 40276 34786 40357 34898
rect 40469 34786 40496 34898
rect 40276 34595 40496 34786
rect 46533 176301 169101 176521
rect 46533 13477 46753 176301
rect 171881 175537 172101 181117
rect 173032 180626 173352 180627
rect 173032 180308 173033 180626
rect 173351 180308 173352 180626
rect 173032 180307 173352 180308
rect 175008 180626 175328 180627
rect 175008 180308 175009 180626
rect 175327 180308 175328 180626
rect 175008 180307 175328 180308
rect 52329 175317 172101 175537
rect 52329 172529 52549 175317
rect 52329 172311 52330 172529
rect 52548 172311 52549 172529
rect 52329 171265 52549 172311
rect 156179 173279 157941 173303
rect 156179 171565 156203 173279
rect 157917 171565 157941 173279
rect 86588 169096 86590 169097
rect 86588 166636 86589 169096
rect 86588 166635 86590 166636
rect 86443 165348 86445 165349
rect 86443 162888 86444 165348
rect 86443 162887 86445 162888
rect 86721 154454 86723 154455
rect 86721 151994 86722 154454
rect 86721 151993 86723 151994
rect 86721 136509 86723 136510
rect 86721 134049 86722 136509
rect 86721 134048 86723 134049
rect 156179 117757 157941 171565
rect 162512 173046 164274 173070
rect 162512 171332 162536 173046
rect 164250 171332 164274 173046
rect 162512 117457 164274 171332
rect 177697 173046 179459 173070
rect 177697 171332 177721 173046
rect 179435 171332 179459 173046
rect 196479 173046 198241 173070
rect 170721 168529 171043 168530
rect 170721 168528 170722 168529
rect 171042 168528 171043 168529
rect 164430 168316 164752 168317
rect 164430 168315 164431 168316
rect 164751 168315 164752 168316
rect 173031 168245 173353 168246
rect 173031 168244 173032 168245
rect 173352 168244 173353 168245
rect 167771 168174 168093 168175
rect 167771 168173 167772 168174
rect 168092 168173 168093 168174
rect 175007 168245 175009 168246
rect 175007 167925 175008 168245
rect 175007 167924 175009 167925
rect 177697 117058 179459 171332
rect 196479 171332 196503 173046
rect 198217 171332 198241 173046
rect 207668 173046 209430 173070
rect 196479 117457 198241 171332
rect 196479 114996 198241 115695
rect 207668 171332 207692 173046
rect 209406 171332 209430 173046
rect 207668 117557 209430 171332
rect 578644 167476 578646 167477
rect 578645 162676 578646 167476
rect 578644 162675 578646 162676
rect 504280 149347 504282 149348
rect 504281 146887 504282 149347
rect 504280 146886 504282 146887
rect 504503 139290 504505 139291
rect 504504 136830 504505 139290
rect 504503 136829 504505 136830
rect 287958 118953 290430 118954
rect 287958 118952 287959 118953
rect 290429 118952 290430 118953
rect 207668 115495 209430 115795
rect 46533 13476 46756 13477
rect 46533 13364 46643 13476
rect 46755 13364 46756 13476
rect 46533 13363 46756 13364
rect 46533 12024 46753 13363
rect 353 4020 467 4021
rect 353 3908 354 4020
rect 466 3908 467 4020
rect 353 3907 467 3908
<< via4 >>
rect 329837 700672 333913 703788
rect 229597 697552 231180 699708
rect 143667 694390 144069 694391
rect 143667 694001 143668 694390
rect 143668 694001 144068 694390
rect 144068 694001 144069 694390
rect 7036 687798 7308 688070
rect 26808 684469 29268 684470
rect 26808 681999 29267 684469
rect 29267 681999 29268 684469
rect 26808 681998 29268 681999
rect 7012 243720 7332 243835
rect 7012 243630 7127 243720
rect 7127 243630 7217 243720
rect 7217 243630 7332 243720
rect 7012 243515 7332 243630
rect 26516 678120 28976 678121
rect 26516 675650 28975 678120
rect 28975 675650 28976 678120
rect 26516 675649 28976 675650
rect 26349 672898 28809 672899
rect 26349 670428 28808 672898
rect 28808 670428 28809 672898
rect 26349 670427 28809 670428
rect 18914 667765 19234 667766
rect 18914 667435 18915 667765
rect 18915 667435 19234 667765
rect 18914 667434 19234 667435
rect 18914 664765 19234 664766
rect 18914 664435 18915 664765
rect 18915 664435 19234 664765
rect 18914 664434 19234 664435
rect 18819 662310 19139 662311
rect 18819 661990 18820 662310
rect 18820 661990 19139 662310
rect 18819 661989 19139 661990
rect 18914 661765 19234 661766
rect 18914 661435 18915 661765
rect 18915 661435 19234 661765
rect 18914 661434 19234 661435
rect 18819 659310 19139 659311
rect 18819 658990 18820 659310
rect 18820 658990 19139 659310
rect 18819 658989 19139 658990
rect 18914 658765 19234 658766
rect 18914 658435 18915 658765
rect 18915 658435 19234 658765
rect 18914 658434 19234 658435
rect 18819 656310 19139 656311
rect 18819 655990 18820 656310
rect 18820 655990 19139 656310
rect 18819 655989 19139 655990
rect 18914 655765 19234 655766
rect 18914 655435 18915 655765
rect 18915 655435 19234 655765
rect 18914 655434 19234 655435
rect 18819 653310 19139 653311
rect 18819 652990 18820 653310
rect 18820 652990 19139 653310
rect 18819 652989 19139 652990
rect 18914 652765 19234 652766
rect 18914 652435 18915 652765
rect 18915 652435 19234 652765
rect 18914 652434 19234 652435
rect 14834 651712 17296 651713
rect 14834 649252 14835 651712
rect 14835 649252 17295 651712
rect 17295 649252 17296 651712
rect 18819 650310 19139 650311
rect 18819 649990 18820 650310
rect 18820 649990 19139 650310
rect 18819 649989 19139 649990
rect 18914 649765 19234 649766
rect 18914 649435 18915 649765
rect 18915 649435 19234 649765
rect 18914 649434 19234 649435
rect 14834 649251 17296 649252
rect 18819 647310 19139 647311
rect 18819 646990 18820 647310
rect 18820 646990 19139 647310
rect 18819 646989 19139 646990
rect 18914 646765 19234 646766
rect 18914 646435 18915 646765
rect 18915 646435 19234 646765
rect 18914 646434 19234 646435
rect 14753 646302 17215 646303
rect 14753 643842 14754 646302
rect 14754 643842 17214 646302
rect 17214 643842 17215 646302
rect 18819 644310 19139 644311
rect 18819 643990 18820 644310
rect 18820 643990 19139 644310
rect 18819 643989 19139 643990
rect 14753 643841 17215 643842
rect 18914 643765 19234 643766
rect 18914 643435 18915 643765
rect 18915 643435 19234 643765
rect 18914 643434 19234 643435
rect 18819 641310 19139 641311
rect 18819 640990 18820 641310
rect 18820 640990 19139 641310
rect 18819 640989 19139 640990
rect 18914 640765 19234 640766
rect 18914 640435 18915 640765
rect 18915 640435 19234 640765
rect 18914 640434 19234 640435
rect 18819 638310 19139 638311
rect 18819 637990 18820 638310
rect 18820 637990 19139 638310
rect 18819 637989 19139 637990
rect 18914 637765 19234 637766
rect 18914 637435 18915 637765
rect 18915 637435 19234 637765
rect 18914 637434 19234 637435
rect 18819 635310 19139 635311
rect 18819 634990 18820 635310
rect 18820 634990 19139 635310
rect 18819 634989 19139 634990
rect 18914 634765 19234 634766
rect 18914 634435 18915 634765
rect 18915 634435 19234 634765
rect 18914 634434 19234 634435
rect 18819 632310 19139 632311
rect 18819 631990 18820 632310
rect 18820 631990 19139 632310
rect 18819 631989 19139 631990
rect 18914 631765 19234 631766
rect 18914 631435 18915 631765
rect 18915 631435 19234 631765
rect 18914 631434 19234 631435
rect 11357 627858 13769 630270
rect 18914 625765 19234 625766
rect 18914 625435 18915 625765
rect 18915 625435 19234 625765
rect 18914 625434 19234 625435
rect 11079 624842 13834 624843
rect 11079 622087 13833 624842
rect 13833 622087 13834 624842
rect 18819 623310 19139 623311
rect 18819 622990 18820 623310
rect 18820 622990 19139 623310
rect 18819 622989 19139 622990
rect 18914 622765 19234 622766
rect 18914 622435 18915 622765
rect 18915 622435 19234 622765
rect 18914 622434 19234 622435
rect 11079 622086 13834 622087
rect 18819 620310 19139 620311
rect 18819 619990 18820 620310
rect 18820 619990 19139 620310
rect 18819 619989 19139 619990
rect 18914 619765 19234 619766
rect 18914 619435 18915 619765
rect 18915 619435 19234 619765
rect 18914 619434 19234 619435
rect 15231 617468 17988 617469
rect 15231 614714 15232 617468
rect 15232 614714 17987 617468
rect 17987 614714 17988 617468
rect 18819 617310 19139 617311
rect 18819 616990 18820 617310
rect 18820 616990 19139 617310
rect 18819 616989 19139 616990
rect 18914 616765 19234 616766
rect 18914 616435 18915 616765
rect 18915 616435 19234 616765
rect 18914 616434 19234 616435
rect 18819 614310 19139 614311
rect 18819 613990 18820 614310
rect 18820 613990 19139 614310
rect 18819 613989 19139 613990
rect 18914 613765 19234 613766
rect 18914 613435 18915 613765
rect 18915 613435 19234 613765
rect 18914 613434 19234 613435
rect 18819 611310 19139 611311
rect 18819 610990 18820 611310
rect 18820 610990 19139 611310
rect 18819 610989 19139 610990
rect 18914 610765 19234 610766
rect 18914 610435 18915 610765
rect 18915 610435 19234 610765
rect 18914 610434 19234 610435
rect 13716 610130 16473 610131
rect 13716 607375 13717 610130
rect 13717 607375 16472 610130
rect 16472 607375 16473 610130
rect 18819 608310 19139 608311
rect 18819 607990 18820 608310
rect 18820 607990 19139 608310
rect 18819 607989 19139 607990
rect 18914 607765 19234 607766
rect 18914 607435 18915 607765
rect 18915 607435 19234 607765
rect 18914 607434 19234 607435
rect 13716 607374 16473 607375
rect 11079 605645 13834 605646
rect 11079 602850 13833 605645
rect 13833 602850 13834 605645
rect 18819 605310 19139 605311
rect 18819 604990 18820 605310
rect 18820 604990 19139 605310
rect 18819 604989 19139 604990
rect 18914 604765 19234 604766
rect 18914 604435 18915 604765
rect 18915 604435 19234 604765
rect 18914 604434 19234 604435
rect 11079 602849 13834 602850
rect 18819 602310 19139 602311
rect 18819 601990 18820 602310
rect 18820 601990 19139 602310
rect 18819 601989 19139 601990
rect 18914 601765 19234 601766
rect 18914 601435 18915 601765
rect 18915 601435 19234 601765
rect 18914 601434 19234 601435
rect 18819 599310 19139 599311
rect 18819 598990 18820 599310
rect 18820 598990 19139 599310
rect 18819 598989 19139 598990
rect 18914 598765 19234 598766
rect 18914 598435 18915 598765
rect 18915 598435 19234 598765
rect 18914 598434 19234 598435
rect 14986 597310 17743 597311
rect 14986 594555 14987 597310
rect 14987 594555 17742 597310
rect 17742 594555 17743 597310
rect 18819 596310 19139 596311
rect 18819 595990 18820 596310
rect 18820 595990 19139 596310
rect 18819 595989 19139 595990
rect 18914 595765 19234 595766
rect 18914 595435 18915 595765
rect 18915 595435 19234 595765
rect 18914 595434 19234 595435
rect 14986 594554 17743 594555
rect 18819 593310 19139 593311
rect 18819 592990 18820 593310
rect 18820 592990 19139 593310
rect 18819 592989 19139 592990
rect 18914 592765 19234 592766
rect 18914 592435 18915 592765
rect 18915 592435 19234 592765
rect 18914 592434 19234 592435
rect 18819 590310 19139 590311
rect 18819 589990 18820 590310
rect 18820 589990 19139 590310
rect 18819 589989 19139 589990
rect 18914 589765 19234 589766
rect 14576 589487 17333 589488
rect 14576 586732 14577 589487
rect 14577 586732 17332 589487
rect 17332 586732 17333 589487
rect 18914 589435 18915 589765
rect 18915 589435 19234 589765
rect 18914 589434 19234 589435
rect 18819 587310 19139 587311
rect 18819 586990 18820 587310
rect 18820 586990 19139 587310
rect 18819 586989 19139 586990
rect 14576 586731 17333 586732
rect 18914 586765 19234 586766
rect 18914 586435 18915 586765
rect 18915 586435 19234 586765
rect 18914 586434 19234 586435
rect 18819 584310 19139 584311
rect 14535 584039 17292 584040
rect 14535 581284 14536 584039
rect 14536 581284 17291 584039
rect 17291 581284 17292 584039
rect 18819 583990 18820 584310
rect 18820 583990 19139 584310
rect 18819 583989 19139 583990
rect 18914 583765 19234 583766
rect 18914 583435 18915 583765
rect 18915 583435 19234 583765
rect 18914 583434 19234 583435
rect 14535 581283 17292 581284
rect 18819 581310 19139 581311
rect 18819 580990 18820 581310
rect 18820 580990 19139 581310
rect 18819 580989 19139 580990
rect 18914 580765 19234 580766
rect 18914 580435 18915 580765
rect 18915 580435 19234 580765
rect 18914 580434 19234 580435
rect 14576 578591 17333 578592
rect 14576 575836 14577 578591
rect 14577 575836 17332 578591
rect 17332 575836 17333 578591
rect 18819 578310 19139 578311
rect 18819 577990 18820 578310
rect 18820 577990 19139 578310
rect 18819 577989 19139 577990
rect 18914 577765 19234 577766
rect 18914 577435 18915 577765
rect 18915 577435 19234 577765
rect 18914 577434 19234 577435
rect 14576 575835 17333 575836
rect 18819 575310 19139 575311
rect 18819 574990 18820 575310
rect 18820 574990 19139 575310
rect 18819 574989 19139 574990
rect 18914 574765 19234 574766
rect 18914 574435 18915 574765
rect 18915 574435 19234 574765
rect 18914 574434 19234 574435
rect 18819 572310 19139 572311
rect 18819 571990 18820 572310
rect 18820 571990 19139 572310
rect 18819 571989 19139 571990
rect 18914 571765 19234 571766
rect 14945 571587 17702 571588
rect 14945 568832 14946 571587
rect 14946 568832 17701 571587
rect 17701 568832 17702 571587
rect 18914 571435 18915 571765
rect 18915 571435 19234 571765
rect 18914 571434 19234 571435
rect 18819 569310 19139 569311
rect 18819 568990 18820 569310
rect 18820 568990 19139 569310
rect 18819 568989 19139 568990
rect 14945 568831 17702 568832
rect 18914 568765 19234 568766
rect 18914 568435 18915 568765
rect 18915 568435 19234 568765
rect 18914 568434 19234 568435
rect 18819 566310 19139 566311
rect 18819 565990 18820 566310
rect 18820 565990 19139 566310
rect 18819 565989 19139 565990
rect 18914 565765 19234 565766
rect 18914 565435 18915 565765
rect 18915 565435 19234 565765
rect 18914 565434 19234 565435
rect 15149 564870 17906 564871
rect 15149 562115 15150 564870
rect 15150 562115 17905 564870
rect 17905 562115 17906 564870
rect 18819 563310 19139 563311
rect 18819 562990 18820 563310
rect 18820 562990 19139 563310
rect 18819 562989 19139 562990
rect 18914 562765 19234 562766
rect 18914 562435 18915 562765
rect 18915 562435 19234 562765
rect 18914 562434 19234 562435
rect 15149 562114 17906 562115
rect 15354 560733 18111 560734
rect 15354 557978 15355 560733
rect 15355 557978 18110 560733
rect 18110 557978 18111 560733
rect 18819 560310 19139 560311
rect 18819 559990 18820 560310
rect 18820 559990 19139 560310
rect 18819 559989 19139 559990
rect 18914 559765 19234 559766
rect 18914 559435 18915 559765
rect 18915 559435 19234 559765
rect 18914 559434 19234 559435
rect 15354 557977 18111 557978
rect 18819 557310 19139 557311
rect 18819 556990 18820 557310
rect 18820 556990 19139 557310
rect 18819 556989 19139 556990
rect 18914 556765 19234 556766
rect 18914 556435 18915 556765
rect 18915 556435 19234 556765
rect 18914 556434 19234 556435
rect 14658 554834 17413 554835
rect 14658 552079 14659 554834
rect 14659 552079 17413 554834
rect 18819 554310 19139 554311
rect 18819 553990 18820 554310
rect 18820 553990 19139 554310
rect 18819 553989 19139 553990
rect 18914 553765 19234 553766
rect 18914 553435 18915 553765
rect 18915 553435 19234 553765
rect 18914 553434 19234 553435
rect 14658 552078 17413 552079
rect 18819 551310 19139 551311
rect 18819 550990 18820 551310
rect 18820 550990 19139 551310
rect 18819 550989 19139 550990
rect 18914 550765 19234 550766
rect 18914 550435 18915 550765
rect 18915 550435 19234 550765
rect 18914 550434 19234 550435
rect 18819 548310 19139 548311
rect 18819 547990 18820 548310
rect 18820 547990 19139 548310
rect 18819 547989 19139 547990
rect 18914 547765 19234 547766
rect 18914 547435 18915 547765
rect 18915 547435 19234 547765
rect 18914 547434 19234 547435
rect 14945 547421 17702 547422
rect 14945 544666 14946 547421
rect 14946 544666 17701 547421
rect 17701 544666 17702 547421
rect 18819 545310 19139 545311
rect 18819 544990 18820 545310
rect 18820 544990 19139 545310
rect 18819 544989 19139 544990
rect 14945 544665 17702 544666
rect 18914 544765 19234 544766
rect 18914 544435 18915 544765
rect 18915 544435 19234 544765
rect 18914 544434 19234 544435
rect 18819 542310 19139 542311
rect 18819 541990 18820 542310
rect 18820 541990 19139 542310
rect 18819 541989 19139 541990
rect 18914 541765 19234 541766
rect 18914 541435 18915 541765
rect 18915 541435 19234 541765
rect 18914 541434 19234 541435
rect 15723 540744 18480 540745
rect 15723 537989 15724 540744
rect 15724 537989 18479 540744
rect 18479 537989 18480 540744
rect 18819 539310 19139 539311
rect 18819 538990 18820 539310
rect 18820 538990 19139 539310
rect 18819 538989 19139 538990
rect 18914 538765 19234 538766
rect 18914 538435 18915 538765
rect 18915 538435 19234 538765
rect 18914 538434 19234 538435
rect 15723 537988 18480 537989
rect 18819 536310 19139 536311
rect 18819 535990 18820 536310
rect 18820 535990 19139 536310
rect 18819 535989 19139 535990
rect 18914 535765 19234 535766
rect 18914 535435 18915 535765
rect 18915 535435 19234 535765
rect 18914 535434 19234 535435
rect 18819 533310 19139 533311
rect 18819 532990 18820 533310
rect 18820 532990 19139 533310
rect 18819 532989 19139 532990
rect 18914 532765 19234 532766
rect 15313 532634 18070 532635
rect 15313 529879 15314 532634
rect 15314 529879 18069 532634
rect 18069 529879 18070 532634
rect 18914 532435 18915 532765
rect 18915 532435 19234 532765
rect 18914 532434 19234 532435
rect 18819 530310 19139 530311
rect 18819 529990 18820 530310
rect 18820 529990 19139 530310
rect 18819 529989 19139 529990
rect 15313 529878 18070 529879
rect 18914 529765 19234 529766
rect 18914 529435 18915 529765
rect 18915 529435 19234 529765
rect 18914 529434 19234 529435
rect 18819 527310 19139 527311
rect 18819 526990 18820 527310
rect 18820 526990 19139 527310
rect 18819 526989 19139 526990
rect 18914 526765 19234 526766
rect 18914 526435 18915 526765
rect 18915 526435 19234 526765
rect 18914 526434 19234 526435
rect 18819 524310 19139 524311
rect 15436 524196 18193 524197
rect 15436 521441 15437 524196
rect 15437 521441 18192 524196
rect 18192 521441 18193 524196
rect 18819 523990 18820 524310
rect 18820 523990 19139 524310
rect 18819 523989 19139 523990
rect 18914 523765 19234 523766
rect 18914 523435 18915 523765
rect 18915 523435 19234 523765
rect 18914 523434 19234 523435
rect 15436 521440 18193 521441
rect 18819 521310 19139 521311
rect 18819 520990 18820 521310
rect 18820 520990 19139 521310
rect 18819 520989 19139 520990
rect 18914 520765 19234 520766
rect 18914 520435 18915 520765
rect 18915 520435 19234 520765
rect 18914 520434 19234 520435
rect 18819 518310 19139 518311
rect 18819 517990 18820 518310
rect 18820 517990 19139 518310
rect 18819 517989 19139 517990
rect 18914 517765 19234 517766
rect 18914 517435 18915 517765
rect 18915 517435 19234 517765
rect 18914 517434 19234 517435
rect 15354 516865 18111 516866
rect 15354 514110 15355 516865
rect 15355 514110 18110 516865
rect 18110 514110 18111 516865
rect 18819 515310 19139 515311
rect 18819 514990 18820 515310
rect 18820 514990 19139 515310
rect 18819 514989 19139 514990
rect 15354 514109 18111 514110
rect 18819 512310 19139 512311
rect 15231 511990 17988 511991
rect 15231 509235 15232 511990
rect 15232 509235 17987 511990
rect 17987 509235 17988 511990
rect 18819 511990 18820 512310
rect 18820 511990 19139 512310
rect 18819 511989 19139 511990
rect 18914 511765 19234 511766
rect 18914 511435 18915 511765
rect 18915 511435 19234 511765
rect 18914 511434 19234 511435
rect 15231 509234 17988 509235
rect 18819 509310 19139 509311
rect 18819 508990 18820 509310
rect 18820 508990 19139 509310
rect 18819 508989 19139 508990
rect 18914 508765 19234 508766
rect 18914 508435 18915 508765
rect 18915 508435 19234 508765
rect 18914 508434 19234 508435
rect 15641 508304 18396 508305
rect 15641 505549 15642 508304
rect 15642 505549 18396 508304
rect 18819 506310 19139 506311
rect 18819 505990 18820 506310
rect 18820 505990 19139 506310
rect 18819 505989 19139 505990
rect 15641 505548 18396 505549
rect 18914 505765 19234 505766
rect 18914 505435 18915 505765
rect 18915 505435 19234 505765
rect 18914 505434 19234 505435
rect 18819 503310 19139 503311
rect 18819 502990 18820 503310
rect 18820 502990 19139 503310
rect 18819 502989 19139 502990
rect 18914 502765 19234 502766
rect 18914 502435 18915 502765
rect 18915 502435 19234 502765
rect 18914 502434 19234 502435
rect 18819 500310 19139 500311
rect 18819 499990 18820 500310
rect 18820 499990 19139 500310
rect 18819 499989 19139 499990
rect 11079 499927 13834 499928
rect 11079 497132 13833 499927
rect 13833 497132 13834 499927
rect 18914 499765 19234 499766
rect 18914 499435 18915 499765
rect 18915 499435 19234 499765
rect 18914 499434 19234 499435
rect 11079 497131 13834 497132
rect 18819 497310 19139 497311
rect 18819 496990 18820 497310
rect 18820 496990 19139 497310
rect 18819 496989 19139 496990
rect 18914 496765 19234 496766
rect 18914 496435 18915 496765
rect 18915 496435 19234 496765
rect 18914 496434 19234 496435
rect 18819 494310 19139 494311
rect 18819 493990 18820 494310
rect 18820 493990 19139 494310
rect 18819 493989 19139 493990
rect 18914 493765 19234 493766
rect 18914 493435 18915 493765
rect 18915 493435 19234 493765
rect 18914 493434 19234 493435
rect 15272 492903 18029 492904
rect 15272 490148 15273 492903
rect 15273 490148 18028 492903
rect 18028 490148 18029 492903
rect 18819 491310 19139 491311
rect 18819 490990 18820 491310
rect 18820 490990 19139 491310
rect 18819 490989 19139 490990
rect 18914 490765 19234 490766
rect 18914 490435 18915 490765
rect 18915 490435 19234 490765
rect 18914 490434 19234 490435
rect 15272 490147 18029 490148
rect 18819 488310 19139 488311
rect 18819 487990 18820 488310
rect 18820 487990 19139 488310
rect 18819 487989 19139 487990
rect 18914 487765 19234 487766
rect 18914 487435 18915 487765
rect 18915 487435 19234 487765
rect 18914 487434 19234 487435
rect 14494 486185 17251 486186
rect 14494 483430 14495 486185
rect 14495 483430 17250 486185
rect 17250 483430 17251 486185
rect 18819 485310 19139 485311
rect 18819 484990 18820 485310
rect 18820 484990 19139 485310
rect 18819 484989 19139 484990
rect 18914 484765 19234 484766
rect 18914 484435 18915 484765
rect 18915 484435 19234 484765
rect 18914 484434 19234 484435
rect 14494 483429 17251 483430
rect 18819 482310 19139 482311
rect 18819 481990 18820 482310
rect 18820 481990 19139 482310
rect 18819 481989 19139 481990
rect 18914 481765 19234 481766
rect 18914 481435 18915 481765
rect 18915 481435 19234 481765
rect 18914 481434 19234 481435
rect 18819 479310 19139 479311
rect 18819 478990 18820 479310
rect 18820 478990 19139 479310
rect 18819 478989 19139 478990
rect 18914 478765 19234 478766
rect 18914 478435 18915 478765
rect 18915 478435 19234 478765
rect 18914 478434 19234 478435
rect 18819 476310 19139 476311
rect 18819 475990 18820 476310
rect 18820 475990 19139 476310
rect 18819 475989 19139 475990
rect 18914 475765 19234 475766
rect 18914 475435 18915 475765
rect 18915 475435 19234 475765
rect 18914 475434 19234 475435
rect 18819 473310 19139 473311
rect 18819 472990 18820 473310
rect 18820 472990 19139 473310
rect 18819 472989 19139 472990
rect 18914 472765 19234 472766
rect 18914 472435 18915 472765
rect 18915 472435 19234 472765
rect 18914 472434 19234 472435
rect 18819 470310 19139 470311
rect 18819 469990 18820 470310
rect 18820 469990 19139 470310
rect 18819 469989 19139 469990
rect 18914 469765 19234 469766
rect 18914 469435 18915 469765
rect 18915 469435 19234 469765
rect 18914 469434 19234 469435
rect 18819 467310 19139 467311
rect 18819 466990 18820 467310
rect 18820 466990 19139 467310
rect 18819 466989 19139 466990
rect 18914 466765 19234 466766
rect 18914 466435 18915 466765
rect 18915 466435 19234 466765
rect 18914 466434 19234 466435
rect 18819 464310 19139 464311
rect 18819 463990 18820 464310
rect 18820 463990 19139 464310
rect 18819 463989 19139 463990
rect 18914 463765 19234 463766
rect 18914 463435 18915 463765
rect 18915 463435 19234 463765
rect 18914 463434 19234 463435
rect 14868 458628 17623 461383
rect 18819 461310 19139 461311
rect 18819 460990 18820 461310
rect 18820 460990 19139 461310
rect 18819 460989 19139 460990
rect 18914 460765 19234 460766
rect 18914 460435 18915 460765
rect 18915 460435 19234 460765
rect 18914 460434 19234 460435
rect 18819 458310 19139 458311
rect 18819 457990 18820 458310
rect 18820 457990 19139 458310
rect 18819 457989 19139 457990
rect 18914 457765 19234 457766
rect 18914 457435 18915 457765
rect 18915 457435 19234 457765
rect 18914 457434 19234 457435
rect 18819 455310 19139 455311
rect 18819 454990 18820 455310
rect 18820 454990 19139 455310
rect 18819 454989 19139 454990
rect 18914 454765 19234 454766
rect 18914 454435 18915 454765
rect 18915 454435 19234 454765
rect 18914 454434 19234 454435
rect 18819 452310 19139 452311
rect 18819 451990 18820 452310
rect 18820 451990 19139 452310
rect 18819 451989 19139 451990
rect 18914 451765 19234 451766
rect 18914 451435 18915 451765
rect 18915 451435 19234 451765
rect 18914 451434 19234 451435
rect 18819 449310 19139 449311
rect 18819 448990 18820 449310
rect 18820 448990 19139 449310
rect 18819 448989 19139 448990
rect 18914 448765 19234 448766
rect 18914 448435 18915 448765
rect 18915 448435 19234 448765
rect 18914 448434 19234 448435
rect 18819 446310 19139 446311
rect 18819 445990 18820 446310
rect 18820 445990 19139 446310
rect 18819 445989 19139 445990
rect 18914 445765 19234 445766
rect 18914 445435 18915 445765
rect 18915 445435 19234 445765
rect 18914 445434 19234 445435
rect 18819 443310 19139 443311
rect 18819 442990 18820 443310
rect 18820 442990 19139 443310
rect 18819 442989 19139 442990
rect 18914 442765 19234 442766
rect 18914 442435 18915 442765
rect 18915 442435 19234 442765
rect 18914 442434 19234 442435
rect 18819 440310 19139 440311
rect 18819 439990 18820 440310
rect 18820 439990 19139 440310
rect 18819 439989 19139 439990
rect 18914 439765 19234 439766
rect 18914 439435 18915 439765
rect 18915 439435 19234 439765
rect 18914 439434 19234 439435
rect 18819 437310 19139 437311
rect 18819 436990 18820 437310
rect 18820 436990 19139 437310
rect 18819 436989 19139 436990
rect 18914 436765 19234 436766
rect 18914 436435 18915 436765
rect 18915 436435 19234 436765
rect 18914 436434 19234 436435
rect 18819 434310 19139 434311
rect 18819 433990 18820 434310
rect 18820 433990 19139 434310
rect 18819 433989 19139 433990
rect 18914 433765 19234 433766
rect 18914 433435 18915 433765
rect 18915 433435 19234 433765
rect 18914 433434 19234 433435
rect 18819 431310 19139 431311
rect 18819 430990 18820 431310
rect 18820 430990 19139 431310
rect 18819 430989 19139 430990
rect 18914 430765 19234 430766
rect 18914 430435 18915 430765
rect 18915 430435 19234 430765
rect 18914 430434 19234 430435
rect 14456 429929 17213 429930
rect 14456 427174 14457 429929
rect 14457 427174 17212 429929
rect 17212 427174 17213 429929
rect 18819 428310 19139 428311
rect 18819 427990 18820 428310
rect 18820 427990 19139 428310
rect 18819 427989 19139 427990
rect 18914 427765 19234 427766
rect 18914 427435 18915 427765
rect 18915 427435 19234 427765
rect 18914 427434 19234 427435
rect 14456 427173 17213 427174
rect 18819 425310 19139 425311
rect 18819 424990 18820 425310
rect 18820 424990 19139 425310
rect 18819 424989 19139 424990
rect 18914 424765 19234 424766
rect 18914 424435 18915 424765
rect 18915 424435 19234 424765
rect 18914 424434 19234 424435
rect 18819 422310 19139 422311
rect 18819 421990 18820 422310
rect 18820 421990 19139 422310
rect 18819 421989 19139 421990
rect 18914 421765 19234 421766
rect 18914 421435 18915 421765
rect 18915 421435 19234 421765
rect 18914 421434 19234 421435
rect 18819 419310 19139 419311
rect 18819 418990 18820 419310
rect 18820 418990 19139 419310
rect 18819 418989 19139 418990
rect 18914 418765 19234 418766
rect 18914 418435 18915 418765
rect 18915 418435 19234 418765
rect 18914 418434 19234 418435
rect 18819 416310 19139 416311
rect 18819 415990 18820 416310
rect 18820 415990 19139 416310
rect 18819 415989 19139 415990
rect 18914 415765 19234 415766
rect 18914 415435 18915 415765
rect 18915 415435 19234 415765
rect 18914 415434 19234 415435
rect 18819 413310 19139 413311
rect 18819 412990 18820 413310
rect 18820 412990 19139 413310
rect 18819 412989 19139 412990
rect 18914 412765 19234 412766
rect 18914 412435 18915 412765
rect 18915 412435 19234 412765
rect 18914 412434 19234 412435
rect 18819 410310 19139 410311
rect 18819 409990 18820 410310
rect 18820 409990 19139 410310
rect 18819 409989 19139 409990
rect 18914 409765 19234 409766
rect 18914 409435 18915 409765
rect 18915 409435 19234 409765
rect 18914 409434 19234 409435
rect 18819 407310 19139 407311
rect 18819 406990 18820 407310
rect 18820 406990 19139 407310
rect 18819 406989 19139 406990
rect 18914 406765 19234 406766
rect 18914 406435 18915 406765
rect 18915 406435 19234 406765
rect 18914 406434 19234 406435
rect 18819 404310 19139 404311
rect 18819 403990 18820 404310
rect 18820 403990 19139 404310
rect 18819 403989 19139 403990
rect 18914 403765 19234 403766
rect 18914 403435 18915 403765
rect 18915 403435 19234 403765
rect 18914 403434 19234 403435
rect 18819 401310 19139 401311
rect 18819 400990 18820 401310
rect 18820 400990 19139 401310
rect 18819 400989 19139 400990
rect 18819 398310 19139 398311
rect 18819 397990 18820 398310
rect 18820 397990 19139 398310
rect 18819 397989 19139 397990
rect 18914 397765 19234 397766
rect 18914 397435 18915 397765
rect 18915 397435 19234 397765
rect 18914 397434 19234 397435
rect 18819 395310 19139 395311
rect 18819 394990 18820 395310
rect 18820 394990 19139 395310
rect 18819 394989 19139 394990
rect 18914 394765 19234 394766
rect 18914 394435 18915 394765
rect 18915 394435 19234 394765
rect 18914 394434 19234 394435
rect 18819 392310 19139 392311
rect 18819 391990 18820 392310
rect 18820 391990 19139 392310
rect 18819 391989 19139 391990
rect 18914 391765 19234 391766
rect 18914 391435 18915 391765
rect 18915 391435 19234 391765
rect 18914 391434 19234 391435
rect 18819 389310 19139 389311
rect 18819 388990 18820 389310
rect 18820 388990 19139 389310
rect 18819 388989 19139 388990
rect 18914 388765 19234 388766
rect 18914 388435 18915 388765
rect 18915 388435 19234 388765
rect 18914 388434 19234 388435
rect 18819 386310 19139 386311
rect 18819 385990 18820 386310
rect 18820 385990 19139 386310
rect 18819 385989 19139 385990
rect 18914 385765 19234 385766
rect 18914 385435 18915 385765
rect 18915 385435 19234 385765
rect 18914 385434 19234 385435
rect 18819 383310 19139 383311
rect 18819 382990 18820 383310
rect 18820 382990 19139 383310
rect 18819 382989 19139 382990
rect 18914 382765 19234 382766
rect 18914 382435 18915 382765
rect 18915 382435 19234 382765
rect 18914 382434 19234 382435
rect 18819 380310 19139 380311
rect 18819 379990 18820 380310
rect 18820 379990 19139 380310
rect 18819 379989 19139 379990
rect 18914 379765 19234 379766
rect 18914 379435 18915 379765
rect 18915 379435 19234 379765
rect 18914 379434 19234 379435
rect 18819 377310 19139 377311
rect 18819 376990 18820 377310
rect 18820 376990 19139 377310
rect 18819 376989 19139 376990
rect 18914 376765 19234 376766
rect 18914 376435 18915 376765
rect 18915 376435 19234 376765
rect 18914 376434 19234 376435
rect 18819 374310 19139 374311
rect 18819 373990 18820 374310
rect 18820 373990 19139 374310
rect 18819 373989 19139 373990
rect 18914 373765 19234 373766
rect 18914 373435 18915 373765
rect 18915 373435 19234 373765
rect 18914 373434 19234 373435
rect 18819 371310 19139 371311
rect 18819 370990 18820 371310
rect 18820 370990 19139 371310
rect 18819 370989 19139 370990
rect 18914 370765 19234 370766
rect 18914 370435 18915 370765
rect 18915 370435 19234 370765
rect 18914 370434 19234 370435
rect 18819 368310 19139 368311
rect 18819 367990 18820 368310
rect 18820 367990 19139 368310
rect 18819 367989 19139 367990
rect 18914 367765 19234 367766
rect 18914 367435 18915 367765
rect 18915 367435 19234 367765
rect 18914 367434 19234 367435
rect 18819 365310 19139 365311
rect 18819 364990 18820 365310
rect 18820 364990 19139 365310
rect 18819 364989 19139 364990
rect 18914 364765 19234 364766
rect 18914 364435 18915 364765
rect 18915 364435 19234 364765
rect 18914 364434 19234 364435
rect 18819 362310 19139 362311
rect 18819 361990 18820 362310
rect 18820 361990 19139 362310
rect 18819 361989 19139 361990
rect 155835 682425 156205 682795
rect 402985 675200 405469 675201
rect 231057 673701 231329 673973
rect 402985 672740 403010 675200
rect 403010 672740 405469 675200
rect 402985 672739 405469 672740
rect 143667 670341 143668 670730
rect 143668 670341 144068 670730
rect 144068 670341 144069 670730
rect 143667 670340 144069 670341
rect 402809 668426 402810 670885
rect 402810 668426 405270 670885
rect 405270 668426 405271 670885
rect 402809 668425 405271 668426
rect 501549 668426 501550 670885
rect 501550 668426 504010 670885
rect 504010 668426 504011 670885
rect 501549 668425 504011 668426
rect 34077 667464 34349 667736
rect 358419 666335 358691 666607
rect 403637 666311 403981 666631
rect 34077 664464 34349 664736
rect 53687 664432 53959 664704
rect 358419 663335 358691 663607
rect 403637 663311 403981 663631
rect 51547 662014 51819 662286
rect 34077 661464 34349 661736
rect 358419 660335 358691 660607
rect 403637 660311 403981 660631
rect 51547 659014 51819 659286
rect 34077 658464 34349 658736
rect 358419 657335 358691 657607
rect 403637 657311 403981 657631
rect 51547 656014 51819 656286
rect 34077 655464 34349 655736
rect 358419 654335 358691 654607
rect 403637 654311 403981 654631
rect 51547 653014 51819 653286
rect 34077 652464 34349 652736
rect 358419 651335 358691 651607
rect 403637 651311 403981 651631
rect 51547 650014 51819 650286
rect 34077 649464 34349 649736
rect 358419 648335 358691 648607
rect 403637 648311 403981 648631
rect 51547 647014 51819 647286
rect 34077 646464 34349 646736
rect 358419 645335 358691 645607
rect 403637 645311 403981 645631
rect 51547 644014 51819 644286
rect 34077 643464 34349 643736
rect 358419 642335 358691 642607
rect 403637 642311 403981 642631
rect 51547 641014 51819 641286
rect 34077 640464 34349 640736
rect 358419 639335 358691 639607
rect 403637 639311 403981 639631
rect 51547 638014 51819 638286
rect 34077 637464 34349 637736
rect 358419 636335 358691 636607
rect 403637 636311 403981 636631
rect 51547 635014 51819 635286
rect 34077 634464 34349 634736
rect 358419 633335 358691 633607
rect 403637 633311 403981 633631
rect 51547 632014 51819 632286
rect 34077 631464 34349 631736
rect 358419 630335 358691 630607
rect 403637 630311 403981 630631
rect 404761 627994 407221 627995
rect 358419 627335 358691 627607
rect 403637 627311 403981 627631
rect 34077 625464 34349 625736
rect 404761 625524 404762 627994
rect 404762 625524 407221 627994
rect 404761 625523 407221 625524
rect 358419 624335 358691 624607
rect 403637 624311 403981 624631
rect 51547 623014 51819 623286
rect 34077 622464 34349 622736
rect 358419 621335 358691 621607
rect 403637 621311 403981 621631
rect 51547 620014 51819 620286
rect 34077 619464 34349 619736
rect 358419 618335 358691 618607
rect 403637 618311 403981 618631
rect 51547 617014 51819 617286
rect 34077 616464 34349 616736
rect 404901 615824 407361 615825
rect 358419 615335 358691 615607
rect 403637 615311 403981 615631
rect 51547 614014 51819 614286
rect 34077 613464 34349 613736
rect 404901 613354 404902 615824
rect 404902 613354 407361 615824
rect 404901 613353 407361 613354
rect 358419 612335 358691 612607
rect 403637 612311 403981 612631
rect 51547 611014 51819 611286
rect 34077 610464 34349 610736
rect 358419 609335 358691 609607
rect 403637 609311 403981 609631
rect 51547 608014 51819 608286
rect 34077 607464 34349 607736
rect 358419 606335 358691 606607
rect 403637 606311 403981 606631
rect 51547 605014 51819 605286
rect 34077 604464 34349 604736
rect 358419 603335 358691 603607
rect 403637 603311 403981 603631
rect 51547 602014 51819 602286
rect 404412 602185 406872 602186
rect 34077 601464 34349 601736
rect 358419 600335 358691 600607
rect 403637 600311 403981 600631
rect 404412 599715 404413 602185
rect 404413 599715 406872 602185
rect 404412 599714 406872 599715
rect 51547 599014 51819 599286
rect 34077 598464 34349 598736
rect 358419 597335 358691 597607
rect 403637 597311 403981 597631
rect 51547 596014 51819 596286
rect 34077 595464 34349 595736
rect 358419 594335 358691 594607
rect 403637 594311 403981 594631
rect 51547 593014 51819 593286
rect 34077 592464 34349 592736
rect 358419 591335 358691 591607
rect 403637 591311 403981 591631
rect 51547 590014 51819 590286
rect 34077 589464 34349 589736
rect 358419 588335 358691 588607
rect 403637 588311 403981 588631
rect 403712 587358 406172 587359
rect 51547 587014 51819 587286
rect 34077 586464 34349 586736
rect 403712 585631 403713 587358
rect 358419 585335 358691 585607
rect 403637 585311 403713 585631
rect 403712 584888 403713 585311
rect 403713 584888 406172 587358
rect 403712 584887 406172 584888
rect 51547 584014 51819 584286
rect 34077 583464 34349 583736
rect 358419 582335 358691 582607
rect 403637 582311 403981 582631
rect 51547 581014 51819 581286
rect 34077 580464 34349 580736
rect 358419 579335 358691 579607
rect 403637 579311 403981 579631
rect 51547 578014 51819 578286
rect 34077 577464 34349 577736
rect 358419 576335 358691 576607
rect 403637 576311 403981 576631
rect 51547 575014 51819 575286
rect 34077 574464 34349 574736
rect 358419 573335 358691 573607
rect 403637 573311 403981 573631
rect 51547 572014 51819 572286
rect 34077 571464 34349 571736
rect 358419 570335 358691 570607
rect 403637 570311 403981 570631
rect 51547 569014 51819 569286
rect 34077 568464 34349 568736
rect 358419 567335 358691 567607
rect 403637 567311 403981 567631
rect 51547 566014 51819 566286
rect 404347 566283 406807 566284
rect 34077 565464 34349 565736
rect 358419 564335 358691 564607
rect 403637 564311 403981 564631
rect 404347 563813 404348 566283
rect 404348 563813 406807 566283
rect 404347 563812 406807 563813
rect 51547 563014 51819 563286
rect 34077 562464 34349 562736
rect 358419 561335 358691 561607
rect 403637 561311 403981 561631
rect 51547 560014 51819 560286
rect 34077 559464 34349 559736
rect 358419 558335 358691 558607
rect 403637 558311 403981 558631
rect 51547 557014 51819 557286
rect 34077 556464 34349 556736
rect 358419 555335 358691 555607
rect 403637 555311 403981 555631
rect 51547 554014 51819 554286
rect 34077 553464 34349 553736
rect 358419 552335 358691 552607
rect 403637 552311 403981 552631
rect 404421 552470 406881 552471
rect 51547 551014 51819 551286
rect 34077 550464 34349 550736
rect 404421 550000 404422 552470
rect 404422 550000 406881 552470
rect 404421 549999 406881 550000
rect 358419 549335 358691 549607
rect 403637 549311 403981 549631
rect 51547 548014 51819 548286
rect 34077 547464 34349 547736
rect 358419 546335 358691 546607
rect 403637 546311 403981 546631
rect 51547 545014 51819 545286
rect 34077 544464 34349 544736
rect 358419 543335 358691 543607
rect 403637 543311 403981 543631
rect 404127 542846 406587 542847
rect 51547 542014 51819 542286
rect 34077 541464 34349 541736
rect 358419 540335 358691 540607
rect 403637 540311 403981 540631
rect 404127 540376 404128 542846
rect 404128 540376 406587 542846
rect 404127 540375 406587 540376
rect 51547 539014 51819 539286
rect 34077 538464 34349 538736
rect 358419 537335 358691 537607
rect 403637 537311 403981 537631
rect 51547 536014 51819 536286
rect 34077 535464 34349 535736
rect 358419 534335 358691 534607
rect 403637 534311 403981 534631
rect 51547 533014 51819 533286
rect 34077 532464 34349 532736
rect 404127 531898 406587 531899
rect 358419 531335 358691 531607
rect 403637 531311 403981 531631
rect 51547 530014 51819 530286
rect 34077 529464 34349 529736
rect 404127 529428 404128 531898
rect 404128 529428 406587 531898
rect 404127 529427 406587 529428
rect 358419 528335 358691 528607
rect 403637 528311 403981 528631
rect 51547 527014 51819 527286
rect 34077 526464 34349 526736
rect 358419 525335 358691 525607
rect 403637 525311 403981 525631
rect 51547 524014 51819 524286
rect 34077 523464 34349 523736
rect 358419 522335 358691 522607
rect 403637 522311 403981 522631
rect 51547 521014 51819 521286
rect 34077 520464 34349 520736
rect 358419 519335 358691 519607
rect 403637 519311 403981 519631
rect 51547 518014 51819 518286
rect 34077 517464 34349 517736
rect 358419 516335 358691 516607
rect 403637 516311 403981 516631
rect 51547 515014 51819 515286
rect 358419 513335 358691 513607
rect 403637 513311 403981 513631
rect 404173 512948 406633 512949
rect 51547 512014 51819 512286
rect 34077 511464 34349 511736
rect 358419 510335 358691 510607
rect 403637 510311 403981 510631
rect 404173 510478 404174 512948
rect 404174 510478 406633 512948
rect 404173 510477 406633 510478
rect 51547 509014 51819 509286
rect 34077 508464 34349 508736
rect 358419 507335 358691 507607
rect 403637 507311 403981 507631
rect 51547 506014 51819 506286
rect 34077 505464 34349 505736
rect 358419 504335 358691 504607
rect 403637 504311 403981 504631
rect 51547 503014 51819 503286
rect 34077 502464 34349 502736
rect 358419 501335 358691 501607
rect 403637 501311 403981 501631
rect 51547 500014 51819 500286
rect 34077 499464 34349 499736
rect 358419 498335 358691 498607
rect 403637 498311 403981 498631
rect 51547 497014 51819 497286
rect 34077 496464 34349 496736
rect 358419 495335 358691 495607
rect 403637 495311 403981 495631
rect 51547 494014 51819 494286
rect 34077 493464 34349 493736
rect 358419 492335 358691 492607
rect 403637 492311 403981 492631
rect 51547 491014 51819 491286
rect 34077 490464 34349 490736
rect 358419 489335 358691 489607
rect 403637 489311 403981 489631
rect 51547 488014 51819 488286
rect 34077 487464 34349 487736
rect 358419 486335 358691 486607
rect 403637 486311 403981 486631
rect 404454 486412 406914 486413
rect 51547 485014 51819 485286
rect 34077 484464 34349 484736
rect 404454 483942 404455 486412
rect 404455 483942 406914 486412
rect 404454 483941 406914 483942
rect 358419 483335 358691 483607
rect 403637 483311 403981 483631
rect 51547 482014 51819 482286
rect 34077 481464 34349 481736
rect 358419 480335 358691 480607
rect 403637 480311 403981 480631
rect 51547 479014 51819 479286
rect 34077 478464 34349 478736
rect 358419 477335 358691 477607
rect 403637 477311 403981 477631
rect 51547 476014 51819 476286
rect 34077 475464 34349 475736
rect 358419 474335 358691 474607
rect 403637 474311 403981 474631
rect 51547 473014 51819 473286
rect 34077 472464 34349 472736
rect 358419 471335 358691 471607
rect 403637 471311 403981 471631
rect 51547 470014 51819 470286
rect 34077 469464 34349 469736
rect 358419 468335 358691 468607
rect 403637 468311 403981 468631
rect 51547 467014 51819 467286
rect 34077 466464 34349 466736
rect 358419 465335 358691 465607
rect 403637 465311 403981 465631
rect 51547 464014 51819 464286
rect 34077 463464 34349 463736
rect 358419 462335 358691 462607
rect 403637 462311 403981 462631
rect 51547 461014 51819 461286
rect 34077 460464 34349 460736
rect 358419 459335 358691 459607
rect 403637 459311 403981 459631
rect 51547 458014 51819 458286
rect 34077 457464 34349 457736
rect 358419 456335 358691 456607
rect 403637 456311 403981 456631
rect 51547 455014 51819 455286
rect 34077 454464 34349 454736
rect 358419 453335 358691 453607
rect 403637 453311 403981 453631
rect 51547 452014 51819 452286
rect 34077 451464 34349 451736
rect 358419 450335 358691 450607
rect 403637 450311 403981 450631
rect 404475 449967 406935 449968
rect 51547 449014 51819 449286
rect 34077 448464 34349 448736
rect 358419 447335 358691 447607
rect 403637 447311 403981 447631
rect 404475 447497 404476 449967
rect 404476 447497 406935 449967
rect 404475 447496 406935 447497
rect 51547 446014 51819 446286
rect 34077 445464 34349 445736
rect 358419 444335 358691 444607
rect 403637 444311 403981 444631
rect 51547 443014 51819 443286
rect 34077 442464 34349 442736
rect 358419 441335 358691 441607
rect 403637 441311 403981 441631
rect 51547 440014 51819 440286
rect 34077 439464 34349 439736
rect 358419 438335 358691 438607
rect 403637 438311 403981 438631
rect 51547 437014 51819 437286
rect 34077 436464 34349 436736
rect 358419 435335 358691 435607
rect 403637 435311 403981 435631
rect 51547 434014 51819 434286
rect 34077 433464 34349 433736
rect 358419 432335 358691 432607
rect 403637 432311 403981 432631
rect 51547 431014 51819 431286
rect 34077 430464 34349 430736
rect 358419 429335 358691 429607
rect 403637 429311 403981 429631
rect 51547 428014 51819 428286
rect 34077 427464 34349 427736
rect 358419 426335 358691 426607
rect 403637 426311 403981 426631
rect 51547 425014 51819 425286
rect 34077 424464 34349 424736
rect 358419 423335 358691 423607
rect 403637 423311 403981 423631
rect 51547 422014 51819 422286
rect 34077 421464 34349 421736
rect 404807 421584 407267 421585
rect 358419 420335 358691 420607
rect 403637 420311 403981 420631
rect 51547 419014 51819 419286
rect 404807 419114 404808 421584
rect 404808 419114 407267 421584
rect 404807 419113 407267 419114
rect 34077 418464 34349 418736
rect 358419 417335 358691 417607
rect 403637 417311 403981 417631
rect 51547 416014 51819 416286
rect 34077 415464 34349 415736
rect 358419 414335 358691 414607
rect 403637 414311 403981 414631
rect 51547 413014 51819 413286
rect 34077 412464 34349 412736
rect 358419 411335 358691 411607
rect 403637 411311 403981 411631
rect 51547 410014 51819 410286
rect 34077 409464 34349 409736
rect 404573 409696 407033 409697
rect 358419 408335 358691 408607
rect 403637 408311 403981 408631
rect 51547 407014 51819 407286
rect 404573 407226 404574 409696
rect 404574 407226 407033 409696
rect 404573 407225 407033 407226
rect 34077 406464 34349 406736
rect 358419 405335 358691 405607
rect 403637 405311 403981 405631
rect 51547 404014 51819 404286
rect 34077 403464 34349 403736
rect 358419 402335 358691 402607
rect 403637 402311 403981 402631
rect 51547 401014 51819 401286
rect 358419 399335 358691 399607
rect 403637 399311 403981 399631
rect 51547 398014 51819 398286
rect 34077 397464 34349 397736
rect 358419 396335 358691 396607
rect 403637 396311 403981 396631
rect 51547 395014 51819 395286
rect 34077 394464 34349 394736
rect 358419 393335 358691 393607
rect 403637 393311 403981 393631
rect 51547 392014 51819 392286
rect 34077 391464 34349 391736
rect 358419 390335 358691 390607
rect 403637 390311 403981 390631
rect 51547 389014 51819 389286
rect 34077 388464 34349 388736
rect 358419 387335 358691 387607
rect 403637 387311 403981 387631
rect 51547 386014 51819 386286
rect 34077 385464 34349 385736
rect 358419 384335 358691 384607
rect 403637 384311 403981 384631
rect 51547 383014 51819 383286
rect 34077 382464 34349 382736
rect 358419 381335 358691 381607
rect 403637 381311 403981 381631
rect 51547 380014 51819 380286
rect 34077 379464 34349 379736
rect 358419 378335 358691 378607
rect 403637 378311 403981 378631
rect 51547 377014 51819 377286
rect 34077 376464 34349 376736
rect 358419 375335 358691 375607
rect 403637 375311 403981 375631
rect 51547 374014 51819 374286
rect 34077 373464 34349 373736
rect 51547 371014 51819 371286
rect 34077 370464 34349 370736
rect 51547 368014 51819 368286
rect 34077 367464 34349 367736
rect 412601 644584 417401 644585
rect 412601 639784 412602 644584
rect 412602 639784 417401 644584
rect 412601 639783 417401 639784
rect 412468 634584 417268 634585
rect 412468 632245 412469 634584
rect 412467 632244 412469 632245
rect 412469 632244 417268 634584
rect 412467 629784 412468 632244
rect 412468 629784 417268 632244
rect 412467 629783 417268 629784
rect 413076 594427 415488 596839
rect 413174 573840 417976 573841
rect 413174 569040 413175 573840
rect 413175 569040 417975 573840
rect 417975 569040 417976 573840
rect 413174 569039 417976 569040
rect 413354 562185 418156 562186
rect 413354 557385 413355 562185
rect 413355 557385 418155 562185
rect 418155 557385 418156 562185
rect 413354 557384 418156 557385
rect 413076 520843 415488 523255
rect 413076 494859 415488 497271
rect 413076 462895 415488 465307
rect 413076 433462 415488 435874
rect 413076 397359 415488 399771
rect 413076 383332 415488 385744
rect 414088 377767 414408 377777
rect 414088 377467 414103 377767
rect 414103 377467 414393 377767
rect 414393 377467 414408 377767
rect 414088 377457 414408 377467
rect 413980 377080 414300 377090
rect 413980 376780 413995 377080
rect 413995 376780 414285 377080
rect 414285 376780 414300 377080
rect 413980 376770 414300 376780
rect 414233 376213 414553 376223
rect 414233 375913 414248 376213
rect 414248 375913 414538 376213
rect 414538 375913 414553 376213
rect 414233 375903 414553 375913
rect 414016 374658 414336 374668
rect 414016 374358 414031 374658
rect 414031 374358 414321 374658
rect 414321 374358 414336 374658
rect 414016 374348 414336 374358
rect 413984 374059 414304 374069
rect 413984 373759 413999 374059
rect 413999 373759 414289 374059
rect 414289 373759 414304 374059
rect 413984 373749 414304 373759
rect 414342 373199 414662 373209
rect 414342 372899 414357 373199
rect 414357 372899 414647 373199
rect 414647 372899 414662 373199
rect 414342 372889 414662 372899
rect 414235 372482 414555 372492
rect 414235 372182 414250 372482
rect 414250 372182 414540 372482
rect 414540 372182 414555 372482
rect 414235 372172 414555 372182
rect 414342 371837 414662 371847
rect 414342 371537 414357 371837
rect 414357 371537 414647 371837
rect 414647 371537 414662 371837
rect 414342 371527 414662 371537
rect 414766 371300 415086 371310
rect 414766 371000 414781 371300
rect 414781 371000 415071 371300
rect 415071 371000 415086 371300
rect 414766 370990 415086 371000
rect 413762 370709 414082 370719
rect 413762 370409 413777 370709
rect 413777 370409 414067 370709
rect 414067 370409 414082 370709
rect 413762 370399 414082 370409
rect 51547 365014 51819 365286
rect 34077 364464 34349 364736
rect 53842 364432 54114 364704
rect 51547 362014 51819 362286
rect 364925 362221 365245 362296
rect 364925 362051 365000 362221
rect 365000 362051 365170 362221
rect 365170 362051 365245 362221
rect 364925 361976 365245 362051
rect 404519 362180 406979 362181
rect 404519 359710 404520 362180
rect 404520 359710 406979 362180
rect 404519 359709 406979 359710
rect 26656 353284 29116 353285
rect 26656 350814 29115 353284
rect 29115 350814 29116 353284
rect 26656 350813 29116 350814
rect 26582 348755 29042 348756
rect 26582 346285 29041 348755
rect 29041 346285 29042 348755
rect 26582 346284 29042 346285
rect 26582 344245 29042 344246
rect 26582 341775 29041 344245
rect 29041 341775 29042 344245
rect 26582 341774 29042 341775
rect 14740 340671 17497 340672
rect 14740 337916 14741 340671
rect 14741 337916 17496 340671
rect 17496 337916 17497 340671
rect 14740 337915 17497 337916
rect 55331 345460 55603 345732
rect 58331 345460 58603 345732
rect 61331 345460 61603 345732
rect 64331 345460 64603 345732
rect 67331 345460 67603 345732
rect 70331 345460 70603 345732
rect 73331 345460 73603 345732
rect 76331 345460 76603 345732
rect 79331 345460 79603 345732
rect 82331 345460 82603 345732
rect 85331 345460 85603 345732
rect 88331 345460 88603 345732
rect 91331 345460 91603 345732
rect 94331 345460 94603 345732
rect 97331 345460 97603 345732
rect 100331 345460 100603 345732
rect 103331 345460 103603 345732
rect 106331 345460 106603 345732
rect 109331 345460 109603 345732
rect 112331 345460 112603 345732
rect 115331 345460 115603 345732
rect 118331 345460 118603 345732
rect 121331 345460 121603 345732
rect 124331 345460 124603 345732
rect 127331 345460 127603 345732
rect 130331 345460 130603 345732
rect 133331 345460 133603 345732
rect 136331 345460 136603 345732
rect 139331 345460 139603 345732
rect 142331 345460 142603 345732
rect 145331 345460 145603 345732
rect 148331 345460 148603 345732
rect 151331 345460 151603 345732
rect 154331 345460 154603 345732
rect 157331 345460 157603 345732
rect 160331 345460 160603 345732
rect 163331 345460 163603 345732
rect 166331 345460 166603 345732
rect 169331 345460 169603 345732
rect 172331 345460 172603 345732
rect 175331 345460 175603 345732
rect 178331 345460 178603 345732
rect 181331 345460 181603 345732
rect 184331 345460 184603 345732
rect 187331 345460 187603 345732
rect 190331 345460 190603 345732
rect 193331 345460 193603 345732
rect 196331 345460 196603 345732
rect 199331 345460 199603 345732
rect 202331 345460 202603 345732
rect 205331 345460 205603 345732
rect 208331 345460 208603 345732
rect 211331 345460 211603 345732
rect 214331 345460 214603 345732
rect 217331 345460 217603 345732
rect 220331 345460 220603 345732
rect 223331 345460 223603 345732
rect 226331 345460 226603 345732
rect 229331 345460 229603 345732
rect 232331 345460 232603 345732
rect 235331 345460 235603 345732
rect 238331 345460 238603 345732
rect 241331 345460 241603 345732
rect 244331 345460 244603 345732
rect 247331 345460 247603 345732
rect 250331 345460 250603 345732
rect 253331 345460 253603 345732
rect 256331 345460 256603 345732
rect 259331 345460 259603 345732
rect 262331 345460 262603 345732
rect 265331 345460 265603 345732
rect 268331 345460 268603 345732
rect 271331 345460 271603 345732
rect 274331 345460 274603 345732
rect 277331 345460 277603 345732
rect 280331 345460 280603 345732
rect 283331 345460 283603 345732
rect 286331 345460 286603 345732
rect 289331 345460 289603 345732
rect 292331 345460 292603 345732
rect 295331 345460 295603 345732
rect 298331 345460 298603 345732
rect 301331 345460 301603 345732
rect 304331 345460 304603 345732
rect 307331 345460 307603 345732
rect 310331 345460 310603 345732
rect 313331 345460 313603 345732
rect 316331 345460 316603 345732
rect 319331 345460 319603 345732
rect 325331 345460 325603 345732
rect 328331 345460 328603 345732
rect 331331 345460 331603 345732
rect 334331 345460 334603 345732
rect 337331 345460 337603 345732
rect 340331 345460 340603 345732
rect 343331 345460 343603 345732
rect 346331 345460 346603 345732
rect 349331 345460 349603 345732
rect 352331 345460 352603 345732
rect 355331 345460 355603 345732
rect 358331 345460 358603 345732
rect 372476 336909 372796 336914
rect 372476 336599 372486 336909
rect 372486 336599 372786 336909
rect 372786 336599 372796 336909
rect 372476 336594 372796 336599
rect 375476 336909 375796 336914
rect 375476 336599 375486 336909
rect 375486 336599 375786 336909
rect 375786 336599 375796 336909
rect 375476 336594 375796 336599
rect 378476 336909 378796 336914
rect 378476 336599 378486 336909
rect 378486 336599 378786 336909
rect 378786 336599 378796 336909
rect 378476 336594 378796 336599
rect 381476 336909 381796 336914
rect 381476 336599 381486 336909
rect 381486 336599 381786 336909
rect 381786 336599 381796 336909
rect 381476 336594 381796 336599
rect 384476 336909 384796 336914
rect 384476 336599 384486 336909
rect 384486 336599 384786 336909
rect 384786 336599 384796 336909
rect 384476 336594 384796 336599
rect 387476 336909 387796 336914
rect 387476 336599 387486 336909
rect 387486 336599 387786 336909
rect 387786 336599 387796 336909
rect 387476 336594 387796 336599
rect 390476 336909 390796 336914
rect 390476 336599 390486 336909
rect 390486 336599 390786 336909
rect 390786 336599 390796 336909
rect 390476 336594 390796 336599
rect 393476 336909 393796 336914
rect 393476 336599 393486 336909
rect 393486 336599 393786 336909
rect 393786 336599 393796 336909
rect 393476 336594 393796 336599
rect 396476 336909 396796 336914
rect 396476 336599 396486 336909
rect 396486 336599 396786 336909
rect 396786 336599 396796 336909
rect 396476 336594 396796 336599
rect 55301 323102 55302 323421
rect 55302 323102 55632 323421
rect 55632 323102 55633 323421
rect 55301 323101 55633 323102
rect 58301 323102 58302 323421
rect 58302 323102 58632 323421
rect 58632 323102 58633 323421
rect 58301 323101 58633 323102
rect 61301 323102 61302 323421
rect 61302 323102 61632 323421
rect 61632 323102 61633 323421
rect 61301 323101 61633 323102
rect 64301 323102 64302 323421
rect 64302 323102 64632 323421
rect 64632 323102 64633 323421
rect 64301 323101 64633 323102
rect 67301 323102 67302 323421
rect 67302 323102 67632 323421
rect 67632 323102 67633 323421
rect 67301 323101 67633 323102
rect 70301 323102 70302 323421
rect 70302 323102 70632 323421
rect 70632 323102 70633 323421
rect 70301 323101 70633 323102
rect 73301 323102 73302 323421
rect 73302 323102 73632 323421
rect 73632 323102 73633 323421
rect 73301 323101 73633 323102
rect 76301 323102 76302 323421
rect 76302 323102 76632 323421
rect 76632 323102 76633 323421
rect 76301 323101 76633 323102
rect 79301 323102 79302 323421
rect 79302 323102 79632 323421
rect 79632 323102 79633 323421
rect 79301 323101 79633 323102
rect 82301 323102 82302 323421
rect 82302 323102 82632 323421
rect 82632 323102 82633 323421
rect 82301 323101 82633 323102
rect 85301 323102 85302 323421
rect 85302 323102 85632 323421
rect 85632 323102 85633 323421
rect 85301 323101 85633 323102
rect 88301 323102 88302 323421
rect 88302 323102 88632 323421
rect 88632 323102 88633 323421
rect 88301 323101 88633 323102
rect 91301 323102 91302 323421
rect 91302 323102 91632 323421
rect 91632 323102 91633 323421
rect 91301 323101 91633 323102
rect 94301 323102 94302 323421
rect 94302 323102 94632 323421
rect 94632 323102 94633 323421
rect 94301 323101 94633 323102
rect 97301 323102 97302 323421
rect 97302 323102 97632 323421
rect 97632 323102 97633 323421
rect 97301 323101 97633 323102
rect 100301 323102 100302 323421
rect 100302 323102 100632 323421
rect 100632 323102 100633 323421
rect 100301 323101 100633 323102
rect 103301 323102 103302 323421
rect 103302 323102 103632 323421
rect 103632 323102 103633 323421
rect 103301 323101 103633 323102
rect 106301 323102 106302 323421
rect 106302 323102 106632 323421
rect 106632 323102 106633 323421
rect 106301 323101 106633 323102
rect 109301 323102 109302 323421
rect 109302 323102 109632 323421
rect 109632 323102 109633 323421
rect 109301 323101 109633 323102
rect 112301 323102 112302 323421
rect 112302 323102 112632 323421
rect 112632 323102 112633 323421
rect 112301 323101 112633 323102
rect 115301 323102 115302 323421
rect 115302 323102 115632 323421
rect 115632 323102 115633 323421
rect 115301 323101 115633 323102
rect 118301 323102 118302 323421
rect 118302 323102 118632 323421
rect 118632 323102 118633 323421
rect 118301 323101 118633 323102
rect 121301 323102 121302 323421
rect 121302 323102 121632 323421
rect 121632 323102 121633 323421
rect 121301 323101 121633 323102
rect 124301 323102 124302 323421
rect 124302 323102 124632 323421
rect 124632 323102 124633 323421
rect 124301 323101 124633 323102
rect 127301 323102 127302 323421
rect 127302 323102 127632 323421
rect 127632 323102 127633 323421
rect 127301 323101 127633 323102
rect 130301 323102 130302 323421
rect 130302 323102 130632 323421
rect 130632 323102 130633 323421
rect 130301 323101 130633 323102
rect 133301 323102 133302 323421
rect 133302 323102 133632 323421
rect 133632 323102 133633 323421
rect 133301 323101 133633 323102
rect 136301 323102 136302 323421
rect 136302 323102 136632 323421
rect 136632 323102 136633 323421
rect 136301 323101 136633 323102
rect 139301 323102 139302 323421
rect 139302 323102 139632 323421
rect 139632 323102 139633 323421
rect 139301 323101 139633 323102
rect 142301 323102 142302 323421
rect 142302 323102 142632 323421
rect 142632 323102 142633 323421
rect 142301 323101 142633 323102
rect 145301 323102 145302 323421
rect 145302 323102 145632 323421
rect 145632 323102 145633 323421
rect 145301 323101 145633 323102
rect 148301 323102 148302 323421
rect 148302 323102 148632 323421
rect 148632 323102 148633 323421
rect 148301 323101 148633 323102
rect 151301 323102 151302 323421
rect 151302 323102 151632 323421
rect 151632 323102 151633 323421
rect 151301 323101 151633 323102
rect 154301 323102 154302 323421
rect 154302 323102 154632 323421
rect 154632 323102 154633 323421
rect 154301 323101 154633 323102
rect 157301 323102 157302 323421
rect 157302 323102 157632 323421
rect 157632 323102 157633 323421
rect 157301 323101 157633 323102
rect 160301 323102 160302 323421
rect 160302 323102 160632 323421
rect 160632 323102 160633 323421
rect 160301 323101 160633 323102
rect 163301 323102 163302 323421
rect 163302 323102 163632 323421
rect 163632 323102 163633 323421
rect 163301 323101 163633 323102
rect 166301 323102 166302 323421
rect 166302 323102 166632 323421
rect 166632 323102 166633 323421
rect 166301 323101 166633 323102
rect 169301 323102 169302 323421
rect 169302 323102 169632 323421
rect 169632 323102 169633 323421
rect 169301 323101 169633 323102
rect 172301 323102 172302 323421
rect 172302 323102 172632 323421
rect 172632 323102 172633 323421
rect 172301 323101 172633 323102
rect 175301 323102 175302 323421
rect 175302 323102 175632 323421
rect 175632 323102 175633 323421
rect 175301 323101 175633 323102
rect 178301 323102 178302 323421
rect 178302 323102 178632 323421
rect 178632 323102 178633 323421
rect 178301 323101 178633 323102
rect 181301 323102 181302 323421
rect 181302 323102 181632 323421
rect 181632 323102 181633 323421
rect 181301 323101 181633 323102
rect 184301 323102 184302 323421
rect 184302 323102 184632 323421
rect 184632 323102 184633 323421
rect 184301 323101 184633 323102
rect 187301 323102 187302 323421
rect 187302 323102 187632 323421
rect 187632 323102 187633 323421
rect 187301 323101 187633 323102
rect 190301 323102 190302 323421
rect 190302 323102 190632 323421
rect 190632 323102 190633 323421
rect 190301 323101 190633 323102
rect 193301 323102 193302 323421
rect 193302 323102 193632 323421
rect 193632 323102 193633 323421
rect 193301 323101 193633 323102
rect 196301 323102 196302 323421
rect 196302 323102 196632 323421
rect 196632 323102 196633 323421
rect 196301 323101 196633 323102
rect 199301 323102 199302 323421
rect 199302 323102 199632 323421
rect 199632 323102 199633 323421
rect 199301 323101 199633 323102
rect 202301 323102 202302 323421
rect 202302 323102 202632 323421
rect 202632 323102 202633 323421
rect 202301 323101 202633 323102
rect 205301 323102 205302 323421
rect 205302 323102 205632 323421
rect 205632 323102 205633 323421
rect 205301 323101 205633 323102
rect 208301 323102 208302 323421
rect 208302 323102 208632 323421
rect 208632 323102 208633 323421
rect 208301 323101 208633 323102
rect 211301 323102 211302 323421
rect 211302 323102 211632 323421
rect 211632 323102 211633 323421
rect 211301 323101 211633 323102
rect 214301 323102 214302 323421
rect 214302 323102 214632 323421
rect 214632 323102 214633 323421
rect 214301 323101 214633 323102
rect 217301 323102 217302 323421
rect 217302 323102 217632 323421
rect 217632 323102 217633 323421
rect 217301 323101 217633 323102
rect 220301 323102 220302 323421
rect 220302 323102 220632 323421
rect 220632 323102 220633 323421
rect 220301 323101 220633 323102
rect 223301 323102 223302 323421
rect 223302 323102 223632 323421
rect 223632 323102 223633 323421
rect 223301 323101 223633 323102
rect 226301 323102 226302 323421
rect 226302 323102 226632 323421
rect 226632 323102 226633 323421
rect 226301 323101 226633 323102
rect 228301 323101 228633 323421
rect 229301 323102 229302 323421
rect 229302 323102 229632 323421
rect 229632 323102 229633 323421
rect 229301 323101 229633 323102
rect 232301 323102 232302 323421
rect 232302 323102 232632 323421
rect 232632 323102 232633 323421
rect 232301 323101 232633 323102
rect 235301 323102 235302 323421
rect 235302 323102 235632 323421
rect 235632 323102 235633 323421
rect 235301 323101 235633 323102
rect 238301 323102 238302 323421
rect 238302 323102 238632 323421
rect 238632 323102 238633 323421
rect 238301 323101 238633 323102
rect 241301 323102 241302 323421
rect 241302 323102 241632 323421
rect 241632 323102 241633 323421
rect 241301 323101 241633 323102
rect 244301 323102 244302 323421
rect 244302 323102 244632 323421
rect 244632 323102 244633 323421
rect 244301 323101 244633 323102
rect 247301 323102 247302 323421
rect 247302 323102 247632 323421
rect 247632 323102 247633 323421
rect 247301 323101 247633 323102
rect 250301 323102 250302 323421
rect 250302 323102 250632 323421
rect 250632 323102 250633 323421
rect 250301 323101 250633 323102
rect 253301 323102 253302 323421
rect 253302 323102 253632 323421
rect 253632 323102 253633 323421
rect 253301 323101 253633 323102
rect 256301 323102 256302 323421
rect 256302 323102 256632 323421
rect 256632 323102 256633 323421
rect 256301 323101 256633 323102
rect 258301 323101 258633 323421
rect 259301 323102 259302 323421
rect 259302 323102 259632 323421
rect 259632 323102 259633 323421
rect 259301 323101 259633 323102
rect 262301 323102 262302 323421
rect 262302 323102 262632 323421
rect 262632 323102 262633 323421
rect 262301 323101 262633 323102
rect 265301 323102 265302 323421
rect 265302 323102 265632 323421
rect 265632 323102 265633 323421
rect 265301 323101 265633 323102
rect 268301 323102 268302 323421
rect 268302 323102 268632 323421
rect 268632 323102 268633 323421
rect 268301 323101 268633 323102
rect 269301 323101 269633 323421
rect 271301 323102 271302 323421
rect 271302 323102 271632 323421
rect 271632 323102 271633 323421
rect 271301 323101 271633 323102
rect 274301 323102 274302 323421
rect 274302 323102 274632 323421
rect 274632 323102 274633 323421
rect 274301 323101 274633 323102
rect 277301 323102 277302 323421
rect 277302 323102 277632 323421
rect 277632 323102 277633 323421
rect 277301 323101 277633 323102
rect 278301 323101 278633 323421
rect 279301 323101 279633 323421
rect 280301 323102 280302 323421
rect 280302 323102 280632 323421
rect 280632 323102 280633 323421
rect 280301 323101 280633 323102
rect 283301 323102 283302 323421
rect 283302 323102 283632 323421
rect 283632 323102 283633 323421
rect 283301 323101 283633 323102
rect 286301 323102 286302 323421
rect 286302 323102 286632 323421
rect 286632 323102 286633 323421
rect 286301 323101 286633 323102
rect 288301 323101 288633 323421
rect 289301 323102 289302 323421
rect 289302 323102 289632 323421
rect 289632 323102 289633 323421
rect 289301 323101 289633 323102
rect 292301 323102 292302 323421
rect 292302 323102 292632 323421
rect 292632 323102 292633 323421
rect 292301 323101 292633 323102
rect 295301 323102 295302 323421
rect 295302 323102 295632 323421
rect 295632 323102 295633 323421
rect 295301 323101 295633 323102
rect 298301 323102 298302 323421
rect 298302 323102 298632 323421
rect 298632 323102 298633 323421
rect 298301 323101 298633 323102
rect 299301 323101 299633 323421
rect 301301 323102 301302 323421
rect 301302 323102 301632 323421
rect 301632 323102 301633 323421
rect 301301 323101 301633 323102
rect 304301 323102 304302 323421
rect 304302 323102 304632 323421
rect 304632 323102 304633 323421
rect 304301 323101 304633 323102
rect 307301 323102 307302 323421
rect 307302 323102 307632 323421
rect 307632 323102 307633 323421
rect 307301 323101 307633 323102
rect 310301 323102 310302 323421
rect 310302 323102 310632 323421
rect 310632 323102 310633 323421
rect 310301 323101 310633 323102
rect 313301 323102 313302 323421
rect 313302 323102 313632 323421
rect 313632 323102 313633 323421
rect 313301 323101 313633 323102
rect 316301 323102 316302 323421
rect 316302 323102 316632 323421
rect 316632 323102 316633 323421
rect 316301 323101 316633 323102
rect 318301 323101 318633 323421
rect 319301 323102 319302 323421
rect 319302 323102 319632 323421
rect 319632 323102 319633 323421
rect 319301 323101 319633 323102
rect 325301 323102 325302 323421
rect 325302 323102 325632 323421
rect 325632 323102 325633 323421
rect 325301 323101 325633 323102
rect 328301 323102 328302 323421
rect 328302 323102 328632 323421
rect 328632 323102 328633 323421
rect 328301 323101 328633 323102
rect 329301 323101 329633 323421
rect 331301 323102 331302 323421
rect 331302 323102 331632 323421
rect 331632 323102 331633 323421
rect 331301 323101 331633 323102
rect 334301 323102 334302 323421
rect 334302 323102 334632 323421
rect 334632 323102 334633 323421
rect 334301 323101 334633 323102
rect 337301 323102 337302 323421
rect 337302 323102 337632 323421
rect 337632 323102 337633 323421
rect 337301 323101 337633 323102
rect 338301 323101 338633 323421
rect 339301 323101 339633 323421
rect 340301 323102 340302 323421
rect 340302 323102 340632 323421
rect 340632 323102 340633 323421
rect 340301 323101 340633 323102
rect 343301 323102 343302 323421
rect 343302 323102 343632 323421
rect 343632 323102 343633 323421
rect 343301 323101 343633 323102
rect 346301 323102 346302 323421
rect 346302 323102 346632 323421
rect 346632 323102 346633 323421
rect 346301 323101 346633 323102
rect 348301 323101 348633 323421
rect 349301 323102 349302 323421
rect 349302 323102 349632 323421
rect 349632 323102 349633 323421
rect 349301 323101 349633 323102
rect 352301 323102 352302 323421
rect 352302 323102 352632 323421
rect 352632 323102 352633 323421
rect 352301 323101 352633 323102
rect 355301 323102 355302 323421
rect 355302 323102 355632 323421
rect 355632 323102 355633 323421
rect 355301 323101 355633 323102
rect 358301 323102 358302 323421
rect 358302 323102 358632 323421
rect 358632 323102 358633 323421
rect 358301 323101 358633 323102
rect 39942 315920 42402 315921
rect 39942 313450 42401 315920
rect 42401 313450 42402 315920
rect 39942 313449 42402 313450
rect 97448 313479 99860 315891
rect 120141 313479 122553 315891
rect 143560 313479 145972 315891
rect 451368 629784 451369 634583
rect 451369 629784 456169 634583
rect 456169 629784 456170 634583
rect 451368 629783 456170 629784
rect 460693 629784 460694 634583
rect 460694 629784 465494 634583
rect 465494 629784 465495 634583
rect 460693 629783 465495 629784
rect 86876 228314 89288 230726
rect 173401 207498 173723 207499
rect 170811 207380 171133 207381
rect 167887 207156 168209 207157
rect 167887 206837 167888 207156
rect 167888 206837 168208 207156
rect 168208 206837 168209 207156
rect 170811 207061 170812 207380
rect 170812 207061 171132 207380
rect 171132 207061 171133 207380
rect 173401 207179 173402 207498
rect 173402 207179 173722 207498
rect 173722 207179 173723 207498
rect 156565 201965 158279 203679
rect 163189 205508 163509 205828
rect 142258 197761 142530 198033
rect 87328 194269 89090 196031
rect 156203 194293 157917 196007
rect 176811 207061 177133 207381
rect 174334 201965 176048 203679
rect 180906 207295 181226 207310
rect 180906 207005 180916 207295
rect 180916 207005 181216 207295
rect 181216 207005 181226 207295
rect 182811 207061 183133 207381
rect 183906 207295 184226 207310
rect 180906 206990 181226 207005
rect 183906 207005 183916 207295
rect 183916 207005 184216 207295
rect 184216 207005 184226 207295
rect 183906 206990 184226 207005
rect 186906 207295 187226 207310
rect 186906 207005 186916 207295
rect 186916 207005 187216 207295
rect 187216 207005 187226 207295
rect 186906 206990 187226 207005
rect 189906 207295 190226 207310
rect 189906 207005 189916 207295
rect 189916 207005 190216 207295
rect 190216 207005 190226 207295
rect 189906 206990 190226 207005
rect 178443 201965 180157 203679
rect 192906 207295 193226 207310
rect 192906 207005 192916 207295
rect 192916 207005 193216 207295
rect 193216 207005 193226 207295
rect 192906 206990 193226 207005
rect 195906 207295 196226 207310
rect 195906 207005 195916 207295
rect 195916 207005 196216 207295
rect 196216 207005 196226 207295
rect 195906 206990 196226 207005
rect 198906 207295 199226 207310
rect 198906 207005 198916 207295
rect 198916 207005 199216 207295
rect 199216 207005 199226 207295
rect 198906 206990 199226 207005
rect 201906 207295 202226 207310
rect 201906 207005 201916 207295
rect 201916 207005 202216 207295
rect 202216 207005 202226 207295
rect 201906 206990 202226 207005
rect 204906 207295 205226 207310
rect 204906 207005 204916 207295
rect 204916 207005 205216 207295
rect 205216 207005 205226 207295
rect 204906 206990 205226 207005
rect 190981 201965 192695 203679
rect 207523 201965 209237 203679
rect 502079 196230 504539 196231
rect 502079 193770 502080 196230
rect 502080 193891 504539 196230
rect 502080 193890 504540 193891
rect 504540 193890 504561 193891
rect 502080 193770 504561 193890
rect 502079 193769 502102 193770
rect 163213 191891 163485 192163
rect 167912 191891 168184 192163
rect 170836 191891 171108 192163
rect 173426 191891 173698 192163
rect 502101 191430 502102 193769
rect 502102 191430 504561 193770
rect 502101 191429 504561 191430
rect 142234 190717 142554 191037
rect 163717 190741 163989 191013
rect 152727 188679 153047 188999
rect 162835 188703 163107 188975
rect 573844 222136 578644 222137
rect 573844 217336 573845 222136
rect 573845 217336 578644 222136
rect 573844 217335 578644 217336
rect 574268 204057 579068 204058
rect 574268 199257 574269 204057
rect 574269 199257 579068 204057
rect 574268 199256 579068 199257
rect 502390 186230 504850 186231
rect 152760 185526 153080 185846
rect 162835 185550 163107 185822
rect 502390 183770 502391 186230
rect 502391 183891 504850 186230
rect 502391 183890 504851 183891
rect 504851 183890 505014 183891
rect 502391 183770 505014 183890
rect 502390 183769 502555 183770
rect 152494 182834 152814 183154
rect 162835 182858 163107 183130
rect 502554 181430 502555 183769
rect 502555 181430 505014 183770
rect 502554 181429 505014 181430
rect 152719 180307 153039 180627
rect 162865 180331 163137 180603
rect 164455 180331 164727 180603
rect 167796 180331 168068 180603
rect 13381 122346 15841 124806
rect 170746 180331 171018 180603
rect 173056 180331 173328 180603
rect 175032 180331 175304 180603
rect 156203 171565 157917 173279
rect 86590 169096 89050 169097
rect 86590 166636 89049 169096
rect 89049 166636 89050 169096
rect 86590 166635 89050 166636
rect 86445 165348 88905 165349
rect 86445 162888 88904 165348
rect 88904 162888 88905 165348
rect 86445 162887 88905 162888
rect 86723 154454 89183 154455
rect 86723 151994 89182 154454
rect 89182 151994 89183 154454
rect 86723 151993 89183 151994
rect 86723 136509 89183 136510
rect 86723 134049 89182 136509
rect 89182 134049 89183 136509
rect 86723 134048 89183 134049
rect 156179 115995 157941 117757
rect 162536 171332 164250 173046
rect 177721 171332 179435 173046
rect 180867 172814 181187 172824
rect 180867 172514 180872 172814
rect 180872 172514 181182 172814
rect 181182 172514 181187 172814
rect 180867 172504 181187 172514
rect 183867 172814 184187 172824
rect 183867 172514 183872 172814
rect 183872 172514 184182 172814
rect 184182 172514 184187 172814
rect 183867 172504 184187 172514
rect 186867 172814 187187 172824
rect 186867 172514 186872 172814
rect 186872 172514 187182 172814
rect 187182 172514 187187 172814
rect 186867 172504 187187 172514
rect 189867 172814 190187 172824
rect 189867 172514 189872 172814
rect 189872 172514 190182 172814
rect 190182 172514 190187 172814
rect 189867 172504 190187 172514
rect 192867 172814 193187 172824
rect 192867 172514 192872 172814
rect 192872 172514 193182 172814
rect 193182 172514 193187 172814
rect 192867 172504 193187 172514
rect 195867 172814 196187 172824
rect 195867 172514 195872 172814
rect 195872 172514 196182 172814
rect 196182 172514 196187 172814
rect 195867 172504 196187 172514
rect 164430 167996 164431 168315
rect 164431 167996 164751 168315
rect 164751 167996 164752 168315
rect 170721 168209 170722 168528
rect 170722 168209 171042 168528
rect 171042 168209 171043 168528
rect 170721 168208 171043 168209
rect 164430 167995 164752 167996
rect 167771 167854 167772 168173
rect 167772 167854 168092 168173
rect 168092 167854 168093 168173
rect 173031 167925 173032 168244
rect 173032 167925 173352 168244
rect 173352 167925 173353 168244
rect 173031 167924 173353 167925
rect 175009 168245 175329 168246
rect 175009 167925 175328 168245
rect 175328 167925 175329 168245
rect 175009 167924 175329 167925
rect 167771 167853 168093 167854
rect 162512 115695 164274 117457
rect 177697 115296 179459 117058
rect 196503 171332 198217 173046
rect 198867 172814 199187 172824
rect 198867 172514 198872 172814
rect 198872 172514 199182 172814
rect 199182 172514 199187 172814
rect 198867 172504 199187 172514
rect 201867 172814 202187 172824
rect 201867 172514 201872 172814
rect 201872 172514 202182 172814
rect 202182 172514 202187 172814
rect 201867 172504 202187 172514
rect 204867 172814 205187 172824
rect 204867 172514 204872 172814
rect 204872 172514 205182 172814
rect 205182 172514 205187 172814
rect 204867 172504 205187 172514
rect 196479 115695 198241 117457
rect 207692 171332 209406 173046
rect 573844 167476 578644 167477
rect 573844 162676 573845 167476
rect 573845 162676 578644 167476
rect 573844 162675 578644 162676
rect 501820 149347 504280 149348
rect 501820 146887 501821 149347
rect 501821 146887 504280 149347
rect 501820 146886 504280 146887
rect 502043 139290 504503 139291
rect 502043 136830 502044 139290
rect 502044 136830 504503 139290
rect 502043 136829 504503 136830
rect 207668 115795 209430 117557
rect 287958 116493 287959 118952
rect 287959 116493 290429 118952
rect 290429 116493 290430 118952
rect 287958 116492 290430 116493
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 703788 334294 704800
rect 329294 702300 329837 703788
rect 229160 699708 231660 702300
rect 329590 700672 329837 702300
rect 333913 702300 334294 703788
rect 333913 700672 334230 702300
rect 329590 700360 334230 700672
rect 229160 697552 229597 699708
rect 231180 697552 231660 699708
rect 229160 697490 231660 697552
rect 16414 694935 416859 695062
rect 14675 694391 416859 694935
rect 14675 694001 143667 694391
rect 144069 694001 416859 694391
rect 14675 692602 416859 694001
rect 7012 688070 7332 688094
rect 7012 687798 7036 688070
rect 7308 687798 7332 688070
rect 7012 243859 7332 687798
rect 14675 667766 20482 692602
rect 26624 684495 405609 684501
rect 26624 684470 407019 684495
rect 26624 681998 26808 684470
rect 29268 682795 407019 684470
rect 29268 682425 155835 682795
rect 156205 682425 407019 682795
rect 29268 682041 407019 682425
rect 29268 681998 29292 682041
rect 26624 681974 29292 681998
rect 26624 678145 29084 681974
rect 230913 679619 374371 679939
rect 26492 678121 29084 678145
rect 26492 675649 26516 678121
rect 28976 675649 29084 678121
rect 26492 675625 29084 675649
rect 26624 672923 29084 675625
rect 231033 673973 231353 679619
rect 374051 676649 374371 679619
rect 373871 676329 376329 676649
rect 231033 673701 231057 673973
rect 231329 673701 231353 673973
rect 231033 673677 231353 673701
rect 26325 672899 29084 672923
rect 26325 670427 26349 672899
rect 28809 670427 29084 672899
rect 26325 670403 29084 670427
rect 14675 667434 18914 667766
rect 19234 667434 20482 667766
rect 14675 664766 20482 667434
rect 14675 664434 18914 664766
rect 19234 664434 20482 664766
rect 14675 662311 20482 664434
rect 14675 661989 18819 662311
rect 19139 661989 20482 662311
rect 14675 661766 20482 661989
rect 14675 661434 18914 661766
rect 19234 661434 20482 661766
rect 14675 659311 20482 661434
rect 14675 658989 18819 659311
rect 19139 658989 20482 659311
rect 14675 658766 20482 658989
rect 14675 658434 18914 658766
rect 19234 658434 20482 658766
rect 14675 656311 20482 658434
rect 14675 655989 18819 656311
rect 19139 655989 20482 656311
rect 14675 655766 20482 655989
rect 14675 655434 18914 655766
rect 19234 655434 20482 655766
rect 14675 653311 20482 655434
rect 14675 652989 18819 653311
rect 19139 652989 20482 653311
rect 14675 652766 20482 652989
rect 14675 652434 18914 652766
rect 19234 652434 20482 652766
rect 14675 651713 20482 652434
rect 14675 649251 14834 651713
rect 17296 650311 20482 651713
rect 17296 649989 18819 650311
rect 19139 649989 20482 650311
rect 17296 649766 20482 649989
rect 17296 649434 18914 649766
rect 19234 649434 20482 649766
rect 17296 649251 20482 649434
rect 14675 647311 20482 649251
rect 14675 646989 18819 647311
rect 19139 646989 20482 647311
rect 14675 646766 20482 646989
rect 14675 646434 18914 646766
rect 19234 646434 20482 646766
rect 14675 646303 20482 646434
rect 14675 643841 14753 646303
rect 17215 644311 20482 646303
rect 17215 643989 18819 644311
rect 19139 643989 20482 644311
rect 17215 643841 20482 643989
rect 14675 643766 20482 643841
rect 14675 643434 18914 643766
rect 19234 643434 20482 643766
rect 14675 641311 20482 643434
rect 14675 640989 18819 641311
rect 19139 640989 20482 641311
rect 14675 640766 20482 640989
rect 14675 640434 18914 640766
rect 19234 640434 20482 640766
rect 14675 638311 20482 640434
rect 14675 637989 18819 638311
rect 19139 637989 20482 638311
rect 14675 637766 20482 637989
rect 14675 637434 18914 637766
rect 19234 637434 20482 637766
rect 14675 635311 20482 637434
rect 14675 634989 18819 635311
rect 19139 634989 20482 635311
rect 14675 634766 20482 634989
rect 14675 634434 18914 634766
rect 19234 634434 20482 634766
rect 14675 632311 20482 634434
rect 14675 631989 18819 632311
rect 19139 631989 20482 632311
rect 14675 631766 20482 631989
rect 14675 631434 18914 631766
rect 19234 631434 20482 631766
rect 14675 630294 20482 631434
rect 11333 630270 20482 630294
rect 11333 627858 11357 630270
rect 13769 627858 20482 630270
rect 11333 627834 20482 627858
rect 14675 625766 20482 627834
rect 14675 625434 18914 625766
rect 19234 625434 20482 625766
rect 11055 624843 13858 624867
rect 11055 622086 11079 624843
rect 13834 624842 13858 624843
rect 14675 624842 20482 625434
rect 13834 623311 20482 624842
rect 13834 622989 18819 623311
rect 19139 622989 20482 623311
rect 13834 622766 20482 622989
rect 13834 622434 18914 622766
rect 19234 622434 20482 622766
rect 13834 622087 20482 622434
rect 13834 622086 13858 622087
rect 11055 622062 13858 622086
rect 14675 620311 20482 622087
rect 14675 619989 18819 620311
rect 19139 619989 20482 620311
rect 14675 619766 20482 619989
rect 14675 619434 18914 619766
rect 19234 619434 20482 619766
rect 14675 617469 20482 619434
rect 14675 614714 15231 617469
rect 17988 617311 20482 617469
rect 17988 616989 18819 617311
rect 19139 616989 20482 617311
rect 17988 616766 20482 616989
rect 17988 616434 18914 616766
rect 19234 616434 20482 616766
rect 17988 614714 20482 616434
rect 14675 614311 20482 614714
rect 14675 613989 18819 614311
rect 19139 613989 20482 614311
rect 14675 613766 20482 613989
rect 14675 613434 18914 613766
rect 19234 613434 20482 613766
rect 14675 611311 20482 613434
rect 14675 610989 18819 611311
rect 19139 610989 20482 611311
rect 14675 610766 20482 610989
rect 14675 610434 18914 610766
rect 19234 610434 20482 610766
rect 14675 610155 20482 610434
rect 13692 610131 20482 610155
rect 13692 607374 13716 610131
rect 16473 608311 20482 610131
rect 16473 607989 18819 608311
rect 19139 607989 20482 608311
rect 16473 607766 20482 607989
rect 16473 607434 18914 607766
rect 19234 607434 20482 607766
rect 16473 607374 20482 607434
rect 13692 607350 20482 607374
rect 11055 605646 13858 605670
rect 11055 602849 11079 605646
rect 13834 605625 13858 605646
rect 14675 605625 20482 607350
rect 13834 605311 20482 605625
rect 13834 604989 18819 605311
rect 19139 604989 20482 605311
rect 13834 604766 20482 604989
rect 13834 604434 18914 604766
rect 19234 604434 20482 604766
rect 13834 602870 20482 604434
rect 13834 602849 13858 602870
rect 11055 602825 13858 602849
rect 14675 602311 20482 602870
rect 14675 601989 18819 602311
rect 19139 601989 20482 602311
rect 14675 601766 20482 601989
rect 14675 601434 18914 601766
rect 19234 601434 20482 601766
rect 14675 599311 20482 601434
rect 14675 598989 18819 599311
rect 19139 598989 20482 599311
rect 14675 598766 20482 598989
rect 14675 598434 18914 598766
rect 19234 598434 20482 598766
rect 14675 597311 20482 598434
rect 14675 594554 14986 597311
rect 17743 596311 20482 597311
rect 17743 595989 18819 596311
rect 19139 595989 20482 596311
rect 17743 595766 20482 595989
rect 17743 595434 18914 595766
rect 19234 595434 20482 595766
rect 17743 594554 20482 595434
rect 14675 593311 20482 594554
rect 14675 592989 18819 593311
rect 19139 592989 20482 593311
rect 14675 592766 20482 592989
rect 14675 592434 18914 592766
rect 19234 592434 20482 592766
rect 14675 590311 20482 592434
rect 14675 589989 18819 590311
rect 19139 589989 20482 590311
rect 14675 589766 20482 589989
rect 14675 589512 18914 589766
rect 14552 589488 18914 589512
rect 14552 586731 14576 589488
rect 17333 589434 18914 589488
rect 19234 589434 20482 589766
rect 17333 587311 20482 589434
rect 17333 586989 18819 587311
rect 19139 586989 20482 587311
rect 17333 586766 20482 586989
rect 17333 586731 18914 586766
rect 14552 586707 18914 586731
rect 14675 586434 18914 586707
rect 19234 586434 20482 586766
rect 14675 584311 20482 586434
rect 14675 584064 18819 584311
rect 14511 584040 18819 584064
rect 14511 581283 14535 584040
rect 17292 583989 18819 584040
rect 19139 583989 20482 584311
rect 17292 583766 20482 583989
rect 17292 583434 18914 583766
rect 19234 583434 20482 583766
rect 17292 581311 20482 583434
rect 17292 581283 18819 581311
rect 14511 581259 18819 581283
rect 14675 580989 18819 581259
rect 19139 580989 20482 581311
rect 14675 580766 20482 580989
rect 14675 580434 18914 580766
rect 19234 580434 20482 580766
rect 14675 578616 20482 580434
rect 14552 578592 20482 578616
rect 14552 575835 14576 578592
rect 17333 578311 20482 578592
rect 17333 577989 18819 578311
rect 19139 577989 20482 578311
rect 17333 577766 20482 577989
rect 17333 577434 18914 577766
rect 19234 577434 20482 577766
rect 17333 575835 20482 577434
rect 14552 575811 20482 575835
rect 14675 575311 20482 575811
rect 14675 574989 18819 575311
rect 19139 574989 20482 575311
rect 14675 574766 20482 574989
rect 14675 574434 18914 574766
rect 19234 574434 20482 574766
rect 14675 572311 20482 574434
rect 14675 571989 18819 572311
rect 19139 571989 20482 572311
rect 14675 571766 20482 571989
rect 14675 571588 18914 571766
rect 14675 568831 14945 571588
rect 17702 571434 18914 571588
rect 19234 571434 20482 571766
rect 17702 569311 20482 571434
rect 17702 568989 18819 569311
rect 19139 568989 20482 569311
rect 17702 568831 20482 568989
rect 14675 568766 20482 568831
rect 14675 568434 18914 568766
rect 19234 568434 20482 568766
rect 14675 566311 20482 568434
rect 14675 565989 18819 566311
rect 19139 565989 20482 566311
rect 14675 565766 20482 565989
rect 14675 565434 18914 565766
rect 19234 565434 20482 565766
rect 14675 564871 20482 565434
rect 14675 562114 15149 564871
rect 17906 563311 20482 564871
rect 17906 562989 18819 563311
rect 19139 562989 20482 563311
rect 17906 562766 20482 562989
rect 17906 562434 18914 562766
rect 19234 562434 20482 562766
rect 17906 562114 20482 562434
rect 14675 560734 20482 562114
rect 14675 557977 15354 560734
rect 18111 560311 20482 560734
rect 18111 559989 18819 560311
rect 19139 559989 20482 560311
rect 18111 559766 20482 559989
rect 18111 559434 18914 559766
rect 19234 559434 20482 559766
rect 18111 557977 20482 559434
rect 14675 557311 20482 557977
rect 14675 556989 18819 557311
rect 19139 556989 20482 557311
rect 14675 556766 20482 556989
rect 14675 556434 18914 556766
rect 19234 556434 20482 556766
rect 14675 554859 20482 556434
rect 14634 554835 20482 554859
rect 14634 552078 14658 554835
rect 17413 554311 20482 554835
rect 17413 553989 18819 554311
rect 19139 553989 20482 554311
rect 17413 553766 20482 553989
rect 17413 553434 18914 553766
rect 19234 553434 20482 553766
rect 17413 552078 20482 553434
rect 14634 552054 20482 552078
rect 14675 551311 20482 552054
rect 14675 550989 18819 551311
rect 19139 550989 20482 551311
rect 14675 550766 20482 550989
rect 14675 550434 18914 550766
rect 19234 550434 20482 550766
rect 14675 548311 20482 550434
rect 14675 547989 18819 548311
rect 19139 547989 20482 548311
rect 14675 547766 20482 547989
rect 14675 547434 18914 547766
rect 19234 547434 20482 547766
rect 14675 547422 20482 547434
rect 14675 544665 14945 547422
rect 17702 545311 20482 547422
rect 17702 544989 18819 545311
rect 19139 544989 20482 545311
rect 17702 544766 20482 544989
rect 17702 544665 18914 544766
rect 14675 544434 18914 544665
rect 19234 544434 20482 544766
rect 14675 542311 20482 544434
rect 14675 541989 18819 542311
rect 19139 541989 20482 542311
rect 14675 541766 20482 541989
rect 14675 541434 18914 541766
rect 19234 541434 20482 541766
rect 14675 540745 20482 541434
rect 14675 537988 15723 540745
rect 18480 539311 20482 540745
rect 18480 538989 18819 539311
rect 19139 538989 20482 539311
rect 18480 538766 20482 538989
rect 18480 538434 18914 538766
rect 19234 538434 20482 538766
rect 18480 537988 20482 538434
rect 14675 536311 20482 537988
rect 14675 535989 18819 536311
rect 19139 535989 20482 536311
rect 14675 535766 20482 535989
rect 14675 535434 18914 535766
rect 19234 535434 20482 535766
rect 14675 533311 20482 535434
rect 14675 532989 18819 533311
rect 19139 532989 20482 533311
rect 14675 532766 20482 532989
rect 14675 532635 18914 532766
rect 14675 529878 15313 532635
rect 18070 532434 18914 532635
rect 19234 532434 20482 532766
rect 18070 530311 20482 532434
rect 18070 529989 18819 530311
rect 19139 529989 20482 530311
rect 18070 529878 20482 529989
rect 14675 529766 20482 529878
rect 14675 529434 18914 529766
rect 19234 529434 20482 529766
rect 14675 527311 20482 529434
rect 14675 526989 18819 527311
rect 19139 526989 20482 527311
rect 14675 526766 20482 526989
rect 14675 526434 18914 526766
rect 19234 526434 20482 526766
rect 14675 524311 20482 526434
rect 14675 524197 18819 524311
rect 14675 521440 15436 524197
rect 18193 523989 18819 524197
rect 19139 523989 20482 524311
rect 18193 523766 20482 523989
rect 18193 523434 18914 523766
rect 19234 523434 20482 523766
rect 18193 521440 20482 523434
rect 14675 521311 20482 521440
rect 14675 520989 18819 521311
rect 19139 520989 20482 521311
rect 14675 520766 20482 520989
rect 14675 520434 18914 520766
rect 19234 520434 20482 520766
rect 14675 518311 20482 520434
rect 14675 517989 18819 518311
rect 19139 517989 20482 518311
rect 14675 517766 20482 517989
rect 14675 517434 18914 517766
rect 19234 517434 20482 517766
rect 14675 516866 20482 517434
rect 14675 514109 15354 516866
rect 18111 515311 20482 516866
rect 18111 514989 18819 515311
rect 19139 514989 20482 515311
rect 18111 514109 20482 514989
rect 14675 512311 20482 514109
rect 14675 511991 18819 512311
rect 14675 509234 15231 511991
rect 17988 511989 18819 511991
rect 19139 511989 20482 512311
rect 17988 511766 20482 511989
rect 17988 511434 18914 511766
rect 19234 511434 20482 511766
rect 17988 509311 20482 511434
rect 17988 509234 18819 509311
rect 14675 508989 18819 509234
rect 19139 508989 20482 509311
rect 14675 508766 20482 508989
rect 14675 508434 18914 508766
rect 19234 508434 20482 508766
rect 14675 508305 20482 508434
rect 14675 505548 15641 508305
rect 18396 506311 20482 508305
rect 18396 505989 18819 506311
rect 19139 505989 20482 506311
rect 18396 505766 20482 505989
rect 18396 505548 18914 505766
rect 14675 505434 18914 505548
rect 19234 505434 20482 505766
rect 14675 503311 20482 505434
rect 14675 502989 18819 503311
rect 19139 502989 20482 503311
rect 14675 502766 20482 502989
rect 14675 502434 18914 502766
rect 19234 502434 20482 502766
rect 14675 500311 20482 502434
rect 14675 499989 18819 500311
rect 19139 499989 20482 500311
rect 11055 499928 13858 499952
rect 11055 497131 11079 499928
rect 13834 499907 13858 499928
rect 14675 499907 20482 499989
rect 13834 499766 20482 499907
rect 13834 499434 18914 499766
rect 19234 499434 20482 499766
rect 13834 497311 20482 499434
rect 13834 497152 18819 497311
rect 13834 497131 13858 497152
rect 11055 497107 13858 497131
rect 14675 496989 18819 497152
rect 19139 496989 20482 497311
rect 14675 496766 20482 496989
rect 14675 496434 18914 496766
rect 19234 496434 20482 496766
rect 14675 494311 20482 496434
rect 14675 493989 18819 494311
rect 19139 493989 20482 494311
rect 14675 493766 20482 493989
rect 14675 493434 18914 493766
rect 19234 493434 20482 493766
rect 14675 492904 20482 493434
rect 14675 490147 15272 492904
rect 18029 491311 20482 492904
rect 18029 490989 18819 491311
rect 19139 490989 20482 491311
rect 18029 490766 20482 490989
rect 18029 490434 18914 490766
rect 19234 490434 20482 490766
rect 18029 490147 20482 490434
rect 14675 488311 20482 490147
rect 14675 487989 18819 488311
rect 19139 487989 20482 488311
rect 14675 487766 20482 487989
rect 14675 487434 18914 487766
rect 19234 487434 20482 487766
rect 14675 486210 20482 487434
rect 14470 486186 20482 486210
rect 14470 483429 14494 486186
rect 17251 485311 20482 486186
rect 17251 484989 18819 485311
rect 19139 484989 20482 485311
rect 17251 484766 20482 484989
rect 17251 484434 18914 484766
rect 19234 484434 20482 484766
rect 17251 483429 20482 484434
rect 14470 483405 20482 483429
rect 14675 482311 20482 483405
rect 14675 481989 18819 482311
rect 19139 481989 20482 482311
rect 14675 481766 20482 481989
rect 14675 481434 18914 481766
rect 19234 481434 20482 481766
rect 14675 479311 20482 481434
rect 14675 478989 18819 479311
rect 19139 478989 20482 479311
rect 14675 478766 20482 478989
rect 14675 478434 18914 478766
rect 19234 478434 20482 478766
rect 14675 476311 20482 478434
rect 14675 475989 18819 476311
rect 19139 475989 20482 476311
rect 14675 475766 20482 475989
rect 14675 475434 18914 475766
rect 19234 475434 20482 475766
rect 14675 473311 20482 475434
rect 14675 472989 18819 473311
rect 19139 472989 20482 473311
rect 14675 472766 20482 472989
rect 14675 472434 18914 472766
rect 19234 472434 20482 472766
rect 14675 470311 20482 472434
rect 14675 469989 18819 470311
rect 19139 469989 20482 470311
rect 14675 469766 20482 469989
rect 14675 469434 18914 469766
rect 19234 469434 20482 469766
rect 14675 467311 20482 469434
rect 14675 466989 18819 467311
rect 19139 466989 20482 467311
rect 14675 466766 20482 466989
rect 14675 466434 18914 466766
rect 19234 466434 20482 466766
rect 14675 464311 20482 466434
rect 14675 463989 18819 464311
rect 19139 463989 20482 464311
rect 14675 463766 20482 463989
rect 14675 463434 18914 463766
rect 19234 463434 20482 463766
rect 14675 461383 20482 463434
rect 14675 458628 14868 461383
rect 17623 461311 20482 461383
rect 17623 460989 18819 461311
rect 19139 460989 20482 461311
rect 17623 460766 20482 460989
rect 17623 460434 18914 460766
rect 19234 460434 20482 460766
rect 17623 458628 20482 460434
rect 14675 458311 20482 458628
rect 14675 457989 18819 458311
rect 19139 457989 20482 458311
rect 14675 457766 20482 457989
rect 14675 457434 18914 457766
rect 19234 457434 20482 457766
rect 14675 455311 20482 457434
rect 14675 454989 18819 455311
rect 19139 454989 20482 455311
rect 14675 454766 20482 454989
rect 14675 454434 18914 454766
rect 19234 454434 20482 454766
rect 14675 452311 20482 454434
rect 14675 451989 18819 452311
rect 19139 451989 20482 452311
rect 14675 451766 20482 451989
rect 14675 451434 18914 451766
rect 19234 451434 20482 451766
rect 14675 449311 20482 451434
rect 14675 448989 18819 449311
rect 19139 448989 20482 449311
rect 14675 448766 20482 448989
rect 14675 448434 18914 448766
rect 19234 448434 20482 448766
rect 14675 446311 20482 448434
rect 14675 445989 18819 446311
rect 19139 445989 20482 446311
rect 14675 445766 20482 445989
rect 14675 445434 18914 445766
rect 19234 445434 20482 445766
rect 14675 443311 20482 445434
rect 14675 442989 18819 443311
rect 19139 442989 20482 443311
rect 14675 442766 20482 442989
rect 14675 442434 18914 442766
rect 19234 442434 20482 442766
rect 14675 440311 20482 442434
rect 14675 439989 18819 440311
rect 19139 439989 20482 440311
rect 14675 439766 20482 439989
rect 14675 439434 18914 439766
rect 19234 439434 20482 439766
rect 14675 437311 20482 439434
rect 14675 436989 18819 437311
rect 19139 436989 20482 437311
rect 14675 436766 20482 436989
rect 14675 436434 18914 436766
rect 19234 436434 20482 436766
rect 14675 434311 20482 436434
rect 14675 433989 18819 434311
rect 19139 433989 20482 434311
rect 14675 433766 20482 433989
rect 14675 433434 18914 433766
rect 19234 433434 20482 433766
rect 14675 431311 20482 433434
rect 14675 430989 18819 431311
rect 19139 430989 20482 431311
rect 14675 430766 20482 430989
rect 14675 430434 18914 430766
rect 19234 430434 20482 430766
rect 14675 429954 20482 430434
rect 14432 429930 20482 429954
rect 14432 427173 14456 429930
rect 17213 428311 20482 429930
rect 17213 427989 18819 428311
rect 19139 427989 20482 428311
rect 17213 427766 20482 427989
rect 17213 427434 18914 427766
rect 19234 427434 20482 427766
rect 17213 427173 20482 427434
rect 14432 427149 20482 427173
rect 14675 425311 20482 427149
rect 14675 424989 18819 425311
rect 19139 424989 20482 425311
rect 14675 424766 20482 424989
rect 14675 424434 18914 424766
rect 19234 424434 20482 424766
rect 14675 422311 20482 424434
rect 14675 421989 18819 422311
rect 19139 421989 20482 422311
rect 14675 421766 20482 421989
rect 14675 421434 18914 421766
rect 19234 421434 20482 421766
rect 14675 419311 20482 421434
rect 14675 418989 18819 419311
rect 19139 418989 20482 419311
rect 14675 418766 20482 418989
rect 14675 418434 18914 418766
rect 19234 418434 20482 418766
rect 14675 416311 20482 418434
rect 14675 415989 18819 416311
rect 19139 415989 20482 416311
rect 14675 415766 20482 415989
rect 14675 415434 18914 415766
rect 19234 415434 20482 415766
rect 14675 413311 20482 415434
rect 14675 412989 18819 413311
rect 19139 412989 20482 413311
rect 14675 412766 20482 412989
rect 14675 412434 18914 412766
rect 19234 412434 20482 412766
rect 14675 410311 20482 412434
rect 14675 409989 18819 410311
rect 19139 409989 20482 410311
rect 14675 409766 20482 409989
rect 14675 409434 18914 409766
rect 19234 409434 20482 409766
rect 14675 407311 20482 409434
rect 14675 406989 18819 407311
rect 19139 406989 20482 407311
rect 14675 406766 20482 406989
rect 14675 406434 18914 406766
rect 19234 406434 20482 406766
rect 14675 404311 20482 406434
rect 14675 403989 18819 404311
rect 19139 403989 20482 404311
rect 14675 403766 20482 403989
rect 14675 403434 18914 403766
rect 19234 403434 20482 403766
rect 14675 401311 20482 403434
rect 14675 400989 18819 401311
rect 19139 400989 20482 401311
rect 14675 398311 20482 400989
rect 14675 397989 18819 398311
rect 19139 397989 20482 398311
rect 14675 397766 20482 397989
rect 14675 397434 18914 397766
rect 19234 397434 20482 397766
rect 14675 395311 20482 397434
rect 14675 394989 18819 395311
rect 19139 394989 20482 395311
rect 14675 394766 20482 394989
rect 14675 394434 18914 394766
rect 19234 394434 20482 394766
rect 14675 392311 20482 394434
rect 14675 391989 18819 392311
rect 19139 391989 20482 392311
rect 14675 391766 20482 391989
rect 14675 391434 18914 391766
rect 19234 391434 20482 391766
rect 14675 389311 20482 391434
rect 14675 388989 18819 389311
rect 19139 388989 20482 389311
rect 14675 388766 20482 388989
rect 14675 388434 18914 388766
rect 19234 388434 20482 388766
rect 14675 386311 20482 388434
rect 14675 385989 18819 386311
rect 19139 385989 20482 386311
rect 14675 385766 20482 385989
rect 14675 385434 18914 385766
rect 19234 385434 20482 385766
rect 14675 383311 20482 385434
rect 14675 382989 18819 383311
rect 19139 382989 20482 383311
rect 14675 382766 20482 382989
rect 14675 382434 18914 382766
rect 19234 382434 20482 382766
rect 14675 380311 20482 382434
rect 14675 379989 18819 380311
rect 19139 379989 20482 380311
rect 14675 379766 20482 379989
rect 14675 379434 18914 379766
rect 19234 379434 20482 379766
rect 14675 377311 20482 379434
rect 14675 376989 18819 377311
rect 19139 376989 20482 377311
rect 14675 376766 20482 376989
rect 14675 376434 18914 376766
rect 19234 376434 20482 376766
rect 14675 374311 20482 376434
rect 14675 373989 18819 374311
rect 19139 373989 20482 374311
rect 14675 373766 20482 373989
rect 14675 373434 18914 373766
rect 19234 373434 20482 373766
rect 14675 371311 20482 373434
rect 14675 370989 18819 371311
rect 19139 370989 20482 371311
rect 14675 370766 20482 370989
rect 14675 370434 18914 370766
rect 19234 370434 20482 370766
rect 14675 368311 20482 370434
rect 14675 367989 18819 368311
rect 19139 367989 20482 368311
rect 14675 367766 20482 367989
rect 14675 367434 18914 367766
rect 19234 367434 20482 367766
rect 14675 365311 20482 367434
rect 14675 364989 18819 365311
rect 19139 364989 20482 365311
rect 14675 364766 20482 364989
rect 14675 364434 18914 364766
rect 19234 364434 20482 364766
rect 14675 362311 20482 364434
rect 14675 361989 18819 362311
rect 19139 361989 20482 362311
rect 14675 340672 20482 361989
rect 26624 666911 29084 670403
rect 143643 670730 144093 670754
rect 143643 670340 143667 670730
rect 144069 670340 144093 670730
rect 143643 670316 144093 670340
rect 34053 667736 34373 667760
rect 34053 667464 34077 667736
rect 34349 667464 34373 667736
rect 34053 667440 34373 667464
rect 26624 666591 33713 666911
rect 26624 663911 29084 666591
rect 34053 664736 34373 664760
rect 34053 664464 34077 664736
rect 34349 664464 34373 664736
rect 34053 664440 34373 664464
rect 53663 664704 54897 664728
rect 53663 664432 53687 664704
rect 53959 664432 54897 664704
rect 53663 664408 54897 664432
rect 26624 663591 33713 663911
rect 26624 660911 29084 663591
rect 51523 662286 51843 662310
rect 51523 662014 51547 662286
rect 51819 662014 51843 662286
rect 51523 661990 51843 662014
rect 34053 661736 34373 661760
rect 34053 661464 34077 661736
rect 34349 661464 34373 661736
rect 34053 661440 34373 661464
rect 26624 660591 33713 660911
rect 26624 657911 29084 660591
rect 51523 659286 51843 659310
rect 51523 659014 51547 659286
rect 51819 659014 51843 659286
rect 51523 658990 51843 659014
rect 34053 658736 34373 658760
rect 34053 658464 34077 658736
rect 34349 658464 34373 658736
rect 34053 658440 34373 658464
rect 26624 657591 33713 657911
rect 26624 654911 29084 657591
rect 51523 656286 51843 656310
rect 51523 656014 51547 656286
rect 51819 656014 51843 656286
rect 51523 655990 51843 656014
rect 34053 655736 34373 655760
rect 34053 655464 34077 655736
rect 34349 655464 34373 655736
rect 34053 655440 34373 655464
rect 374051 655260 374371 676329
rect 402810 675201 407019 682041
rect 402810 672739 402985 675201
rect 405469 672739 407019 675201
rect 402810 670909 407019 672739
rect 402785 670885 407019 670909
rect 402785 668425 402809 670885
rect 405271 668425 407019 670885
rect 402785 668401 407019 668425
rect 362730 654940 374371 655260
rect 402810 666631 407019 668401
rect 402810 666311 403637 666631
rect 403981 666311 407019 666631
rect 402810 663631 407019 666311
rect 402810 663311 403637 663631
rect 403981 663311 407019 663631
rect 402810 660631 407019 663311
rect 402810 660311 403637 660631
rect 403981 660311 407019 660631
rect 402810 657631 407019 660311
rect 402810 657311 403637 657631
rect 403981 657311 407019 657631
rect 26624 654591 33713 654911
rect 26624 651911 29084 654591
rect 51523 653286 51843 653310
rect 51523 653014 51547 653286
rect 51819 653014 51843 653286
rect 51523 652990 51843 653014
rect 34053 652736 34373 652760
rect 34053 652464 34077 652736
rect 34349 652464 34373 652736
rect 34053 652440 34373 652464
rect 26624 651591 33713 651911
rect 26624 648911 29084 651591
rect 51523 650286 51843 650310
rect 51523 650014 51547 650286
rect 51819 650014 51843 650286
rect 51523 649990 51843 650014
rect 34053 649736 34373 649760
rect 34053 649464 34077 649736
rect 34349 649464 34373 649736
rect 34053 649440 34373 649464
rect 26624 648591 33713 648911
rect 26624 645911 29084 648591
rect 51523 647286 51843 647310
rect 51523 647014 51547 647286
rect 51819 647014 51843 647286
rect 51523 646990 51843 647014
rect 34053 646736 34373 646760
rect 34053 646464 34077 646736
rect 34349 646464 34373 646736
rect 34053 646440 34373 646464
rect 26624 645591 33713 645911
rect 26624 642911 29084 645591
rect 51523 644286 51843 644310
rect 51523 644014 51547 644286
rect 51819 644014 51843 644286
rect 51523 643990 51843 644014
rect 34053 643736 34373 643760
rect 34053 643464 34077 643736
rect 34349 643464 34373 643736
rect 34053 643440 34373 643464
rect 26624 642591 33713 642911
rect 26624 639911 29084 642591
rect 51523 641286 51843 641310
rect 51523 641014 51547 641286
rect 51819 641014 51843 641286
rect 51523 640990 51843 641014
rect 34053 640736 34373 640760
rect 34053 640464 34077 640736
rect 34349 640464 34373 640736
rect 34053 640440 34373 640464
rect 26624 639591 33713 639911
rect 26624 636911 29084 639591
rect 51523 638286 51843 638310
rect 51523 638014 51547 638286
rect 51819 638014 51843 638286
rect 51523 637990 51843 638014
rect 34053 637736 34373 637760
rect 34053 637464 34077 637736
rect 34349 637464 34373 637736
rect 34053 637440 34373 637464
rect 26624 636591 33713 636911
rect 26624 633911 29084 636591
rect 51523 635286 51843 635310
rect 51523 635014 51547 635286
rect 51819 635014 51843 635286
rect 51523 634990 51843 635014
rect 34053 634736 34373 634760
rect 34053 634464 34077 634736
rect 34349 634464 34373 634736
rect 34053 634440 34373 634464
rect 26624 633591 33713 633911
rect 26624 630911 29084 633591
rect 51523 632286 51843 632310
rect 51523 632014 51547 632286
rect 51819 632014 51843 632286
rect 51523 631990 51843 632014
rect 34053 631736 34373 631760
rect 34053 631464 34077 631736
rect 34349 631464 34373 631736
rect 34053 631440 34373 631464
rect 26624 630591 33713 630911
rect 26624 627911 29084 630591
rect 26624 627591 33713 627911
rect 26624 624911 29084 627591
rect 34053 625736 34373 625760
rect 34053 625464 34077 625736
rect 34349 625464 34373 625736
rect 34053 625440 34373 625464
rect 26624 624591 33713 624911
rect 26624 621911 29084 624591
rect 51523 623286 51843 623310
rect 51523 623014 51547 623286
rect 51819 623014 51843 623286
rect 51523 622990 51843 623014
rect 34053 622736 34373 622760
rect 34053 622464 34077 622736
rect 34349 622464 34373 622736
rect 34053 622440 34373 622464
rect 26624 621591 33713 621911
rect 26624 618911 29084 621591
rect 51523 620286 51843 620310
rect 51523 620014 51547 620286
rect 51819 620014 51843 620286
rect 51523 619990 51843 620014
rect 34053 619736 34373 619760
rect 34053 619464 34077 619736
rect 34349 619464 34373 619736
rect 34053 619440 34373 619464
rect 26624 618591 33713 618911
rect 26624 615911 29084 618591
rect 51523 617286 51843 617310
rect 51523 617014 51547 617286
rect 51819 617014 51843 617286
rect 51523 616990 51843 617014
rect 34053 616736 34373 616760
rect 34053 616464 34077 616736
rect 34349 616464 34373 616736
rect 34053 616440 34373 616464
rect 26624 615591 33713 615911
rect 26624 612911 29084 615591
rect 51523 614286 51843 614310
rect 51523 614014 51547 614286
rect 51819 614014 51843 614286
rect 51523 613990 51843 614014
rect 34053 613736 34373 613760
rect 34053 613464 34077 613736
rect 34349 613464 34373 613736
rect 34053 613440 34373 613464
rect 26624 612591 33713 612911
rect 26624 609911 29084 612591
rect 51523 611286 51843 611310
rect 51523 611014 51547 611286
rect 51819 611014 51843 611286
rect 51523 610990 51843 611014
rect 34053 610736 34373 610760
rect 34053 610464 34077 610736
rect 34349 610464 34373 610736
rect 34053 610440 34373 610464
rect 26624 609591 33713 609911
rect 26624 606911 29084 609591
rect 51523 608286 51843 608310
rect 51523 608014 51547 608286
rect 51819 608014 51843 608286
rect 51523 607990 51843 608014
rect 34053 607736 34373 607760
rect 34053 607464 34077 607736
rect 34349 607464 34373 607736
rect 34053 607440 34373 607464
rect 26624 606591 33713 606911
rect 26624 603911 29084 606591
rect 51523 605286 51843 605310
rect 51523 605014 51547 605286
rect 51819 605014 51843 605286
rect 51523 604990 51843 605014
rect 34053 604736 34373 604760
rect 34053 604464 34077 604736
rect 34349 604464 34373 604736
rect 34053 604440 34373 604464
rect 26624 603591 33713 603911
rect 26624 600911 29084 603591
rect 51523 602286 51843 602310
rect 51523 602014 51547 602286
rect 51819 602014 51843 602286
rect 51523 601990 51843 602014
rect 34053 601736 34373 601760
rect 34053 601464 34077 601736
rect 34349 601464 34373 601736
rect 34053 601440 34373 601464
rect 26624 600591 33713 600911
rect 26624 597911 29084 600591
rect 51523 599286 51843 599310
rect 51523 599014 51547 599286
rect 51819 599014 51843 599286
rect 51523 598990 51843 599014
rect 34053 598736 34373 598760
rect 34053 598464 34077 598736
rect 34349 598464 34373 598736
rect 34053 598440 34373 598464
rect 26624 597591 33713 597911
rect 26624 594911 29084 597591
rect 51523 596286 51843 596310
rect 51523 596014 51547 596286
rect 51819 596014 51843 596286
rect 51523 595990 51843 596014
rect 34053 595736 34373 595760
rect 34053 595464 34077 595736
rect 34349 595464 34373 595736
rect 34053 595440 34373 595464
rect 26624 594591 33713 594911
rect 26624 591911 29084 594591
rect 51523 593286 51843 593310
rect 51523 593014 51547 593286
rect 51819 593014 51843 593286
rect 51523 592990 51843 593014
rect 34053 592736 34373 592760
rect 34053 592464 34077 592736
rect 34349 592464 34373 592736
rect 34053 592440 34373 592464
rect 26624 591591 33713 591911
rect 26624 588911 29084 591591
rect 51523 590286 51843 590310
rect 51523 590014 51547 590286
rect 51819 590014 51843 590286
rect 51523 589990 51843 590014
rect 34053 589736 34373 589760
rect 34053 589464 34077 589736
rect 34349 589464 34373 589736
rect 34053 589440 34373 589464
rect 26624 588591 33713 588911
rect 26624 585911 29084 588591
rect 51523 587286 51843 587310
rect 51523 587014 51547 587286
rect 51819 587014 51843 587286
rect 51523 586990 51843 587014
rect 34053 586736 34373 586760
rect 34053 586464 34077 586736
rect 34349 586464 34373 586736
rect 34053 586440 34373 586464
rect 26624 585591 33713 585911
rect 26624 582911 29084 585591
rect 51523 584286 51843 584310
rect 51523 584014 51547 584286
rect 51819 584014 51843 584286
rect 51523 583990 51843 584014
rect 34053 583736 34373 583760
rect 34053 583464 34077 583736
rect 34349 583464 34373 583736
rect 34053 583440 34373 583464
rect 26624 582591 33713 582911
rect 26624 579911 29084 582591
rect 51523 581286 51843 581310
rect 51523 581014 51547 581286
rect 51819 581014 51843 581286
rect 51523 580990 51843 581014
rect 34053 580736 34373 580760
rect 34053 580464 34077 580736
rect 34349 580464 34373 580736
rect 34053 580440 34373 580464
rect 26624 579591 33713 579911
rect 26624 576911 29084 579591
rect 51523 578286 51843 578310
rect 51523 578014 51547 578286
rect 51819 578014 51843 578286
rect 51523 577990 51843 578014
rect 34053 577736 34373 577760
rect 34053 577464 34077 577736
rect 34349 577464 34373 577736
rect 34053 577440 34373 577464
rect 26624 576591 33713 576911
rect 26624 573911 29084 576591
rect 51523 575286 51843 575310
rect 51523 575014 51547 575286
rect 51819 575014 51843 575286
rect 51523 574990 51843 575014
rect 34053 574736 34373 574760
rect 34053 574464 34077 574736
rect 34349 574464 34373 574736
rect 34053 574440 34373 574464
rect 26624 573591 33713 573911
rect 26624 570911 29084 573591
rect 51523 572286 51843 572310
rect 51523 572014 51547 572286
rect 51819 572014 51843 572286
rect 51523 571990 51843 572014
rect 34053 571736 34373 571760
rect 34053 571464 34077 571736
rect 34349 571464 34373 571736
rect 34053 571440 34373 571464
rect 26624 570591 33713 570911
rect 26624 567911 29084 570591
rect 51523 569286 51843 569310
rect 51523 569014 51547 569286
rect 51819 569014 51843 569286
rect 51523 568990 51843 569014
rect 34053 568736 34373 568760
rect 34053 568464 34077 568736
rect 34349 568464 34373 568736
rect 34053 568440 34373 568464
rect 26624 567591 33713 567911
rect 26624 564911 29084 567591
rect 51523 566286 51843 566310
rect 51523 566014 51547 566286
rect 51819 566014 51843 566286
rect 51523 565990 51843 566014
rect 34053 565736 34373 565760
rect 34053 565464 34077 565736
rect 34349 565464 34373 565736
rect 34053 565440 34373 565464
rect 26624 564591 33713 564911
rect 26624 561911 29084 564591
rect 51523 563286 51843 563310
rect 51523 563014 51547 563286
rect 51819 563014 51843 563286
rect 51523 562990 51843 563014
rect 34053 562736 34373 562760
rect 34053 562464 34077 562736
rect 34349 562464 34373 562736
rect 34053 562440 34373 562464
rect 26624 561591 33713 561911
rect 26624 558911 29084 561591
rect 51523 560286 51843 560310
rect 51523 560014 51547 560286
rect 51819 560014 51843 560286
rect 51523 559990 51843 560014
rect 34053 559736 34373 559760
rect 34053 559464 34077 559736
rect 34349 559464 34373 559736
rect 34053 559440 34373 559464
rect 26624 558591 33713 558911
rect 26624 555911 29084 558591
rect 51523 557286 51843 557310
rect 51523 557014 51547 557286
rect 51819 557014 51843 557286
rect 51523 556990 51843 557014
rect 34053 556736 34373 556760
rect 34053 556464 34077 556736
rect 34349 556464 34373 556736
rect 34053 556440 34373 556464
rect 26624 555591 33713 555911
rect 26624 552911 29084 555591
rect 51523 554286 51843 554310
rect 51523 554014 51547 554286
rect 51819 554014 51843 554286
rect 51523 553990 51843 554014
rect 34053 553736 34373 553760
rect 34053 553464 34077 553736
rect 34349 553464 34373 553736
rect 34053 553440 34373 553464
rect 26624 552591 33713 552911
rect 26624 549911 29084 552591
rect 51523 551286 51843 551310
rect 51523 551014 51547 551286
rect 51819 551014 51843 551286
rect 51523 550990 51843 551014
rect 34053 550736 34373 550760
rect 34053 550464 34077 550736
rect 34349 550464 34373 550736
rect 34053 550440 34373 550464
rect 26624 549591 33713 549911
rect 26624 546911 29084 549591
rect 51523 548286 51843 548310
rect 51523 548014 51547 548286
rect 51819 548014 51843 548286
rect 51523 547990 51843 548014
rect 34053 547736 34373 547760
rect 34053 547464 34077 547736
rect 34349 547464 34373 547736
rect 34053 547440 34373 547464
rect 26624 546591 33713 546911
rect 26624 543911 29084 546591
rect 51523 545286 51843 545310
rect 51523 545014 51547 545286
rect 51819 545014 51843 545286
rect 51523 544990 51843 545014
rect 34053 544736 34373 544760
rect 34053 544464 34077 544736
rect 34349 544464 34373 544736
rect 34053 544440 34373 544464
rect 26624 543591 33713 543911
rect 26624 540911 29084 543591
rect 51523 542286 51843 542310
rect 51523 542014 51547 542286
rect 51819 542014 51843 542286
rect 51523 541990 51843 542014
rect 34053 541736 34373 541760
rect 34053 541464 34077 541736
rect 34349 541464 34373 541736
rect 34053 541440 34373 541464
rect 26624 540591 33713 540911
rect 26624 537911 29084 540591
rect 51523 539286 51843 539310
rect 51523 539014 51547 539286
rect 51819 539014 51843 539286
rect 51523 538990 51843 539014
rect 34053 538736 34373 538760
rect 34053 538464 34077 538736
rect 34349 538464 34373 538736
rect 34053 538440 34373 538464
rect 26624 537591 33713 537911
rect 26624 534911 29084 537591
rect 51523 536286 51843 536310
rect 51523 536014 51547 536286
rect 51819 536014 51843 536286
rect 51523 535990 51843 536014
rect 34053 535736 34373 535760
rect 34053 535464 34077 535736
rect 34349 535464 34373 535736
rect 34053 535440 34373 535464
rect 26624 534591 33713 534911
rect 26624 531911 29084 534591
rect 51523 533286 51843 533310
rect 51523 533014 51547 533286
rect 51819 533014 51843 533286
rect 51523 532990 51843 533014
rect 34053 532736 34373 532760
rect 34053 532464 34077 532736
rect 34349 532464 34373 532736
rect 34053 532440 34373 532464
rect 26624 531591 33713 531911
rect 26624 528911 29084 531591
rect 51523 530286 51843 530310
rect 51523 530014 51547 530286
rect 51819 530014 51843 530286
rect 51523 529990 51843 530014
rect 34053 529736 34373 529760
rect 34053 529464 34077 529736
rect 34349 529464 34373 529736
rect 34053 529440 34373 529464
rect 26624 528591 33713 528911
rect 26624 525911 29084 528591
rect 51523 527286 51843 527310
rect 51523 527014 51547 527286
rect 51819 527014 51843 527286
rect 51523 526990 51843 527014
rect 34053 526736 34373 526760
rect 34053 526464 34077 526736
rect 34349 526464 34373 526736
rect 34053 526440 34373 526464
rect 26624 525591 33713 525911
rect 26624 522911 29084 525591
rect 51523 524286 51843 524310
rect 51523 524014 51547 524286
rect 51819 524014 51843 524286
rect 51523 523990 51843 524014
rect 34053 523736 34373 523760
rect 34053 523464 34077 523736
rect 34349 523464 34373 523736
rect 34053 523440 34373 523464
rect 26624 522591 33713 522911
rect 26624 519911 29084 522591
rect 51523 521286 51843 521310
rect 51523 521014 51547 521286
rect 51819 521014 51843 521286
rect 51523 520990 51843 521014
rect 34053 520736 34373 520760
rect 34053 520464 34077 520736
rect 34349 520464 34373 520736
rect 34053 520440 34373 520464
rect 26624 519591 33713 519911
rect 26624 516911 29084 519591
rect 51523 518286 51843 518310
rect 51523 518014 51547 518286
rect 51819 518014 51843 518286
rect 51523 517990 51843 518014
rect 34053 517736 34373 517760
rect 34053 517464 34077 517736
rect 34349 517464 34373 517736
rect 34053 517440 34373 517464
rect 26624 516591 33713 516911
rect 26624 513911 29084 516591
rect 51523 515286 51843 515310
rect 51523 515014 51547 515286
rect 51819 515014 51843 515286
rect 51523 514990 51843 515014
rect 26624 513591 33713 513911
rect 26624 510911 29084 513591
rect 51523 512286 51843 512310
rect 51523 512014 51547 512286
rect 51819 512014 51843 512286
rect 51523 511990 51843 512014
rect 34053 511736 34373 511760
rect 34053 511464 34077 511736
rect 34349 511464 34373 511736
rect 34053 511440 34373 511464
rect 26624 510591 33713 510911
rect 26624 507911 29084 510591
rect 51523 509286 51843 509310
rect 51523 509014 51547 509286
rect 51819 509014 51843 509286
rect 51523 508990 51843 509014
rect 34053 508736 34373 508760
rect 34053 508464 34077 508736
rect 34349 508464 34373 508736
rect 34053 508440 34373 508464
rect 26624 507591 33713 507911
rect 26624 504911 29084 507591
rect 51523 506286 51843 506310
rect 51523 506014 51547 506286
rect 51819 506014 51843 506286
rect 51523 505990 51843 506014
rect 34053 505736 34373 505760
rect 34053 505464 34077 505736
rect 34349 505464 34373 505736
rect 34053 505440 34373 505464
rect 26624 504591 33713 504911
rect 26624 501911 29084 504591
rect 51523 503286 51843 503310
rect 51523 503014 51547 503286
rect 51819 503014 51843 503286
rect 51523 502990 51843 503014
rect 34053 502736 34373 502760
rect 34053 502464 34077 502736
rect 34349 502464 34373 502736
rect 34053 502440 34373 502464
rect 26624 501591 33713 501911
rect 26624 498911 29084 501591
rect 51523 500286 51843 500310
rect 51523 500014 51547 500286
rect 51819 500014 51843 500286
rect 51523 499990 51843 500014
rect 34053 499736 34373 499760
rect 34053 499464 34077 499736
rect 34349 499464 34373 499736
rect 34053 499440 34373 499464
rect 26624 498591 33713 498911
rect 26624 495911 29084 498591
rect 51523 497286 51843 497310
rect 51523 497014 51547 497286
rect 51819 497014 51843 497286
rect 51523 496990 51843 497014
rect 34053 496736 34373 496760
rect 34053 496464 34077 496736
rect 34349 496464 34373 496736
rect 34053 496440 34373 496464
rect 26624 495591 33713 495911
rect 26624 492911 29084 495591
rect 51523 494286 51843 494310
rect 51523 494014 51547 494286
rect 51819 494014 51843 494286
rect 51523 493990 51843 494014
rect 34053 493736 34373 493760
rect 34053 493464 34077 493736
rect 34349 493464 34373 493736
rect 34053 493440 34373 493464
rect 26624 492591 33713 492911
rect 26624 489911 29084 492591
rect 51523 491286 51843 491310
rect 51523 491014 51547 491286
rect 51819 491014 51843 491286
rect 51523 490990 51843 491014
rect 34053 490736 34373 490760
rect 34053 490464 34077 490736
rect 34349 490464 34373 490736
rect 34053 490440 34373 490464
rect 26624 489591 33713 489911
rect 26624 486911 29084 489591
rect 51523 488286 51843 488310
rect 51523 488014 51547 488286
rect 51819 488014 51843 488286
rect 51523 487990 51843 488014
rect 34053 487736 34373 487760
rect 34053 487464 34077 487736
rect 34349 487464 34373 487736
rect 34053 487440 34373 487464
rect 26624 486591 33713 486911
rect 26624 483911 29084 486591
rect 51523 485286 51843 485310
rect 51523 485014 51547 485286
rect 51819 485014 51843 485286
rect 51523 484990 51843 485014
rect 34053 484736 34373 484760
rect 34053 484464 34077 484736
rect 34349 484464 34373 484736
rect 34053 484440 34373 484464
rect 26624 483591 33713 483911
rect 26624 480911 29084 483591
rect 51523 482286 51843 482310
rect 51523 482014 51547 482286
rect 51819 482014 51843 482286
rect 51523 481990 51843 482014
rect 34053 481736 34373 481760
rect 34053 481464 34077 481736
rect 34349 481464 34373 481736
rect 34053 481440 34373 481464
rect 26624 480591 33713 480911
rect 26624 477911 29084 480591
rect 51523 479286 51843 479310
rect 51523 479014 51547 479286
rect 51819 479014 51843 479286
rect 51523 478990 51843 479014
rect 34053 478736 34373 478760
rect 34053 478464 34077 478736
rect 34349 478464 34373 478736
rect 34053 478440 34373 478464
rect 26624 477591 33713 477911
rect 26624 474911 29084 477591
rect 51523 476286 51843 476310
rect 51523 476014 51547 476286
rect 51819 476014 51843 476286
rect 51523 475990 51843 476014
rect 34053 475736 34373 475760
rect 34053 475464 34077 475736
rect 34349 475464 34373 475736
rect 34053 475440 34373 475464
rect 26624 474591 33713 474911
rect 26624 471911 29084 474591
rect 51523 473286 51843 473310
rect 51523 473014 51547 473286
rect 51819 473014 51843 473286
rect 51523 472990 51843 473014
rect 34053 472736 34373 472760
rect 34053 472464 34077 472736
rect 34349 472464 34373 472736
rect 34053 472440 34373 472464
rect 26624 471591 33713 471911
rect 26624 468911 29084 471591
rect 51523 470286 51843 470310
rect 51523 470014 51547 470286
rect 51819 470014 51843 470286
rect 51523 469990 51843 470014
rect 34053 469736 34373 469760
rect 34053 469464 34077 469736
rect 34349 469464 34373 469736
rect 34053 469440 34373 469464
rect 26624 468591 33713 468911
rect 26624 465911 29084 468591
rect 51523 467286 51843 467310
rect 51523 467014 51547 467286
rect 51819 467014 51843 467286
rect 51523 466990 51843 467014
rect 34053 466736 34373 466760
rect 34053 466464 34077 466736
rect 34349 466464 34373 466736
rect 34053 466440 34373 466464
rect 26624 465591 33713 465911
rect 26624 462911 29084 465591
rect 51523 464286 51843 464310
rect 51523 464014 51547 464286
rect 51819 464014 51843 464286
rect 51523 463990 51843 464014
rect 34053 463736 34373 463760
rect 34053 463464 34077 463736
rect 34349 463464 34373 463736
rect 34053 463440 34373 463464
rect 26624 462591 33713 462911
rect 26624 459911 29084 462591
rect 51523 461286 51843 461310
rect 51523 461014 51547 461286
rect 51819 461014 51843 461286
rect 51523 460990 51843 461014
rect 34053 460736 34373 460760
rect 34053 460464 34077 460736
rect 34349 460464 34373 460736
rect 34053 460440 34373 460464
rect 26624 459591 33713 459911
rect 26624 456911 29084 459591
rect 51523 458286 51843 458310
rect 51523 458014 51547 458286
rect 51819 458014 51843 458286
rect 51523 457990 51843 458014
rect 34053 457736 34373 457760
rect 34053 457464 34077 457736
rect 34349 457464 34373 457736
rect 34053 457440 34373 457464
rect 26624 456591 33713 456911
rect 26624 453911 29084 456591
rect 51523 455286 51843 455310
rect 51523 455014 51547 455286
rect 51819 455014 51843 455286
rect 51523 454990 51843 455014
rect 34053 454736 34373 454760
rect 34053 454464 34077 454736
rect 34349 454464 34373 454736
rect 34053 454440 34373 454464
rect 26624 453591 33713 453911
rect 26624 450911 29084 453591
rect 51523 452286 51843 452310
rect 51523 452014 51547 452286
rect 51819 452014 51843 452286
rect 51523 451990 51843 452014
rect 34053 451736 34373 451760
rect 34053 451464 34077 451736
rect 34349 451464 34373 451736
rect 34053 451440 34373 451464
rect 26624 450591 33713 450911
rect 26624 447911 29084 450591
rect 51523 449286 51843 449310
rect 51523 449014 51547 449286
rect 51819 449014 51843 449286
rect 51523 448990 51843 449014
rect 34053 448736 34373 448760
rect 34053 448464 34077 448736
rect 34349 448464 34373 448736
rect 34053 448440 34373 448464
rect 26624 447591 33713 447911
rect 26624 444911 29084 447591
rect 51523 446286 51843 446310
rect 51523 446014 51547 446286
rect 51819 446014 51843 446286
rect 51523 445990 51843 446014
rect 34053 445736 34373 445760
rect 34053 445464 34077 445736
rect 34349 445464 34373 445736
rect 34053 445440 34373 445464
rect 26624 444591 33713 444911
rect 26624 441911 29084 444591
rect 51523 443286 51843 443310
rect 51523 443014 51547 443286
rect 51819 443014 51843 443286
rect 51523 442990 51843 443014
rect 34053 442736 34373 442760
rect 34053 442464 34077 442736
rect 34349 442464 34373 442736
rect 34053 442440 34373 442464
rect 26624 441591 33713 441911
rect 26624 438911 29084 441591
rect 51523 440286 51843 440310
rect 51523 440014 51547 440286
rect 51819 440014 51843 440286
rect 51523 439990 51843 440014
rect 34053 439736 34373 439760
rect 34053 439464 34077 439736
rect 34349 439464 34373 439736
rect 34053 439440 34373 439464
rect 26624 438591 33713 438911
rect 26624 435911 29084 438591
rect 51523 437286 51843 437310
rect 51523 437014 51547 437286
rect 51819 437014 51843 437286
rect 51523 436990 51843 437014
rect 34053 436736 34373 436760
rect 34053 436464 34077 436736
rect 34349 436464 34373 436736
rect 34053 436440 34373 436464
rect 26624 435591 33713 435911
rect 26624 432911 29084 435591
rect 51523 434286 51843 434310
rect 51523 434014 51547 434286
rect 51819 434014 51843 434286
rect 51523 433990 51843 434014
rect 34053 433736 34373 433760
rect 34053 433464 34077 433736
rect 34349 433464 34373 433736
rect 34053 433440 34373 433464
rect 26624 432591 33713 432911
rect 26624 429911 29084 432591
rect 51523 431286 51843 431310
rect 51523 431014 51547 431286
rect 51819 431014 51843 431286
rect 51523 430990 51843 431014
rect 34053 430736 34373 430760
rect 34053 430464 34077 430736
rect 34349 430464 34373 430736
rect 34053 430440 34373 430464
rect 26624 429591 33713 429911
rect 26624 426911 29084 429591
rect 51523 428286 51843 428310
rect 51523 428014 51547 428286
rect 51819 428014 51843 428286
rect 51523 427990 51843 428014
rect 34053 427736 34373 427760
rect 34053 427464 34077 427736
rect 34349 427464 34373 427736
rect 34053 427440 34373 427464
rect 26624 426591 33713 426911
rect 26624 423911 29084 426591
rect 51523 425286 51843 425310
rect 51523 425014 51547 425286
rect 51819 425014 51843 425286
rect 51523 424990 51843 425014
rect 34053 424736 34373 424760
rect 34053 424464 34077 424736
rect 34349 424464 34373 424736
rect 34053 424440 34373 424464
rect 26624 423591 33713 423911
rect 26624 420911 29084 423591
rect 51523 422286 51843 422310
rect 51523 422014 51547 422286
rect 51819 422014 51843 422286
rect 51523 421990 51843 422014
rect 34053 421736 34373 421760
rect 34053 421464 34077 421736
rect 34349 421464 34373 421736
rect 34053 421440 34373 421464
rect 26624 420591 33713 420911
rect 26624 417911 29084 420591
rect 51523 419286 51843 419310
rect 51523 419014 51547 419286
rect 51819 419014 51843 419286
rect 51523 418990 51843 419014
rect 34053 418736 34373 418760
rect 34053 418464 34077 418736
rect 34349 418464 34373 418736
rect 34053 418440 34373 418464
rect 26624 417591 33713 417911
rect 26624 414911 29084 417591
rect 51523 416286 51843 416310
rect 51523 416014 51547 416286
rect 51819 416014 51843 416286
rect 51523 415990 51843 416014
rect 34053 415736 34373 415760
rect 34053 415464 34077 415736
rect 34349 415464 34373 415736
rect 34053 415440 34373 415464
rect 26624 414591 33713 414911
rect 26624 411911 29084 414591
rect 51523 413286 51843 413310
rect 51523 413014 51547 413286
rect 51819 413014 51843 413286
rect 51523 412990 51843 413014
rect 34053 412736 34373 412760
rect 34053 412464 34077 412736
rect 34349 412464 34373 412736
rect 34053 412440 34373 412464
rect 26624 411591 33713 411911
rect 26624 408911 29084 411591
rect 51523 410286 51843 410310
rect 51523 410014 51547 410286
rect 51819 410014 51843 410286
rect 51523 409990 51843 410014
rect 34053 409736 34373 409760
rect 34053 409464 34077 409736
rect 34349 409464 34373 409736
rect 34053 409440 34373 409464
rect 26624 408591 33713 408911
rect 26624 405911 29084 408591
rect 51523 407286 51843 407310
rect 51523 407014 51547 407286
rect 51819 407014 51843 407286
rect 51523 406990 51843 407014
rect 34053 406736 34373 406760
rect 34053 406464 34077 406736
rect 34349 406464 34373 406736
rect 34053 406440 34373 406464
rect 26624 405591 33713 405911
rect 26624 402911 29084 405591
rect 51523 404286 51843 404310
rect 51523 404014 51547 404286
rect 51819 404014 51843 404286
rect 51523 403990 51843 404014
rect 34053 403736 34373 403760
rect 34053 403464 34077 403736
rect 34349 403464 34373 403736
rect 34053 403440 34373 403464
rect 26624 402591 33713 402911
rect 26624 399911 29084 402591
rect 51523 401286 51843 401310
rect 51523 401014 51547 401286
rect 51819 401014 51843 401286
rect 51523 400990 51843 401014
rect 26624 399591 33713 399911
rect 26624 396911 29084 399591
rect 51523 398286 51843 398310
rect 51523 398014 51547 398286
rect 51819 398014 51843 398286
rect 51523 397990 51843 398014
rect 34053 397736 34373 397760
rect 34053 397464 34077 397736
rect 34349 397464 34373 397736
rect 34053 397440 34373 397464
rect 26624 396591 33713 396911
rect 26624 393911 29084 396591
rect 51523 395286 51843 395310
rect 51523 395014 51547 395286
rect 51819 395014 51843 395286
rect 51523 394990 51843 395014
rect 34053 394736 34373 394760
rect 34053 394464 34077 394736
rect 34349 394464 34373 394736
rect 34053 394440 34373 394464
rect 26624 393591 33713 393911
rect 26624 390911 29084 393591
rect 51523 392286 51843 392310
rect 51523 392014 51547 392286
rect 51819 392014 51843 392286
rect 51523 391990 51843 392014
rect 34053 391736 34373 391760
rect 34053 391464 34077 391736
rect 34349 391464 34373 391736
rect 34053 391440 34373 391464
rect 26624 390591 33713 390911
rect 26624 387911 29084 390591
rect 51523 389286 51843 389310
rect 51523 389014 51547 389286
rect 51819 389014 51843 389286
rect 51523 388990 51843 389014
rect 34053 388736 34373 388760
rect 34053 388464 34077 388736
rect 34349 388464 34373 388736
rect 34053 388440 34373 388464
rect 26624 387591 33713 387911
rect 26624 384911 29084 387591
rect 51523 386286 51843 386310
rect 51523 386014 51547 386286
rect 51819 386014 51843 386286
rect 51523 385990 51843 386014
rect 34053 385736 34373 385760
rect 34053 385464 34077 385736
rect 34349 385464 34373 385736
rect 34053 385440 34373 385464
rect 26624 384591 33713 384911
rect 26624 381911 29084 384591
rect 51523 383286 51843 383310
rect 51523 383014 51547 383286
rect 51819 383014 51843 383286
rect 51523 382990 51843 383014
rect 34053 382736 34373 382760
rect 34053 382464 34077 382736
rect 34349 382464 34373 382736
rect 34053 382440 34373 382464
rect 26624 381591 33713 381911
rect 26624 378911 29084 381591
rect 51523 380286 51843 380310
rect 51523 380014 51547 380286
rect 51819 380014 51843 380286
rect 51523 379990 51843 380014
rect 34053 379736 34373 379760
rect 34053 379464 34077 379736
rect 34349 379464 34373 379736
rect 34053 379440 34373 379464
rect 26624 378591 33713 378911
rect 26624 375911 29084 378591
rect 51523 377286 51843 377310
rect 51523 377014 51547 377286
rect 51819 377014 51843 377286
rect 51523 376990 51843 377014
rect 34053 376736 34373 376760
rect 34053 376464 34077 376736
rect 34349 376464 34373 376736
rect 34053 376440 34373 376464
rect 26624 375591 33713 375911
rect 358395 375607 358715 375631
rect 26624 372911 29084 375591
rect 358395 375335 358419 375607
rect 358691 375335 358715 375607
rect 358395 375311 358715 375335
rect 51523 374286 51843 374310
rect 51523 374014 51547 374286
rect 51819 374014 51843 374286
rect 51523 373990 51843 374014
rect 34053 373736 34373 373760
rect 34053 373464 34077 373736
rect 34349 373464 34373 373736
rect 34053 373440 34373 373464
rect 26624 372591 33713 372911
rect 26624 369911 29084 372591
rect 51523 371286 51843 371310
rect 51523 371014 51547 371286
rect 51819 371014 51843 371286
rect 51523 370990 51843 371014
rect 34053 370736 34373 370760
rect 34053 370464 34077 370736
rect 34349 370464 34373 370736
rect 34053 370440 34373 370464
rect 26624 369591 33713 369911
rect 26624 366911 29084 369591
rect 51523 368286 51843 368310
rect 51523 368014 51547 368286
rect 51819 368014 51843 368286
rect 51523 367990 51843 368014
rect 34053 367736 34373 367760
rect 34053 367464 34077 367736
rect 34349 367464 34373 367736
rect 34053 367440 34373 367464
rect 26624 366591 33713 366911
rect 26624 363911 29084 366591
rect 362730 366160 363050 654940
rect 402810 654631 407019 657311
rect 402810 654311 403637 654631
rect 403981 654311 407019 654631
rect 402810 651631 407019 654311
rect 402810 651311 403637 651631
rect 403981 651311 407019 651631
rect 402810 648631 407019 651311
rect 402810 648311 403637 648631
rect 403981 648311 407019 648631
rect 402810 645631 407019 648311
rect 402810 645311 403637 645631
rect 403981 645311 407019 645631
rect 402810 642631 407019 645311
rect 413052 644609 415512 692602
rect 501525 670885 504035 670909
rect 501525 668425 501549 670885
rect 504011 668425 504035 670885
rect 501525 668401 504035 668425
rect 402810 642311 403637 642631
rect 403981 642311 407019 642631
rect 402810 639631 407019 642311
rect 412577 644585 417425 644609
rect 412577 639783 412601 644585
rect 417401 639783 417425 644585
rect 412577 639759 417425 639783
rect 402810 639311 403637 639631
rect 403981 639311 407019 639631
rect 402810 636631 407019 639311
rect 402810 636311 403637 636631
rect 403981 636311 407019 636631
rect 402810 633631 407019 636311
rect 413052 634609 415512 639759
rect 402810 633311 403637 633631
rect 403981 633311 407019 633631
rect 402810 630631 407019 633311
rect 412444 634585 417292 634609
rect 412444 632269 412468 634585
rect 402810 630311 403637 630631
rect 403981 630311 407019 630631
rect 402810 628019 407019 630311
rect 412443 632245 412468 632269
rect 412443 629783 412467 632245
rect 417268 629783 417292 634585
rect 412443 629759 417292 629783
rect 451344 634583 456194 634607
rect 451344 629783 451368 634583
rect 456170 629783 456194 634583
rect 451344 629759 456194 629783
rect 460669 634583 465519 634607
rect 460669 629783 460693 634583
rect 465495 629783 465519 634583
rect 460669 629759 465519 629783
rect 402810 627995 407245 628019
rect 402810 627631 404761 627995
rect 402810 627311 403637 627631
rect 403981 627311 404761 627631
rect 402810 625523 404761 627311
rect 407221 625523 407245 627995
rect 402810 625499 407245 625523
rect 402810 624631 407019 625499
rect 402810 624311 403637 624631
rect 403981 624311 407019 624631
rect 402810 621631 407019 624311
rect 402810 621311 403637 621631
rect 403981 621311 407019 621631
rect 402810 618631 407019 621311
rect 402810 618311 403637 618631
rect 403981 618311 407019 618631
rect 402810 615849 407019 618311
rect 402810 615825 407385 615849
rect 402810 615631 404901 615825
rect 402810 615311 403637 615631
rect 403981 615311 404901 615631
rect 402810 613353 404901 615311
rect 407361 613353 407385 615825
rect 402810 613329 407385 613353
rect 402810 612631 407019 613329
rect 402810 612311 403637 612631
rect 403981 612311 407019 612631
rect 402810 609631 407019 612311
rect 402810 609311 403637 609631
rect 403981 609311 407019 609631
rect 402810 606631 407019 609311
rect 402810 606311 403637 606631
rect 403981 606311 407019 606631
rect 402810 603631 407019 606311
rect 402810 603311 403637 603631
rect 403981 603311 407019 603631
rect 402810 602186 407019 603311
rect 402810 600631 404412 602186
rect 402810 600311 403637 600631
rect 403981 600311 404412 600631
rect 402810 599714 404412 600311
rect 406872 599714 407019 602186
rect 402810 597631 407019 599714
rect 402810 597311 403637 597631
rect 403981 597311 407019 597631
rect 402810 594631 407019 597311
rect 402810 594311 403637 594631
rect 403981 594311 407019 594631
rect 402810 591631 407019 594311
rect 402810 591311 403637 591631
rect 403981 591311 407019 591631
rect 402810 588631 407019 591311
rect 402810 588311 403637 588631
rect 403981 588311 407019 588631
rect 402810 587359 407019 588311
rect 402810 585631 403712 587359
rect 402810 585311 403637 585631
rect 402810 584887 403712 585311
rect 406172 584887 407019 587359
rect 402810 582631 407019 584887
rect 402810 582311 403637 582631
rect 403981 582311 407019 582631
rect 402810 579631 407019 582311
rect 402810 579311 403637 579631
rect 403981 579311 407019 579631
rect 402810 576631 407019 579311
rect 402810 576311 403637 576631
rect 403981 576311 407019 576631
rect 402810 573631 407019 576311
rect 402810 573311 403637 573631
rect 403981 573311 407019 573631
rect 402810 570631 407019 573311
rect 402810 570311 403637 570631
rect 403981 570311 407019 570631
rect 402810 567631 407019 570311
rect 402810 567311 403637 567631
rect 403981 567311 407019 567631
rect 402810 566284 407019 567311
rect 402810 564631 404347 566284
rect 402810 564311 403637 564631
rect 403981 564311 404347 564631
rect 402810 563812 404347 564311
rect 406807 563812 407019 566284
rect 402810 561631 407019 563812
rect 402810 561311 403637 561631
rect 403981 561311 407019 561631
rect 402810 558631 407019 561311
rect 402810 558311 403637 558631
rect 403981 558311 407019 558631
rect 402810 555631 407019 558311
rect 402810 555311 403637 555631
rect 403981 555311 407019 555631
rect 402810 552631 407019 555311
rect 402810 552311 403637 552631
rect 403981 552471 407019 552631
rect 403981 552311 404421 552471
rect 402810 549999 404421 552311
rect 406881 549999 407019 552471
rect 402810 549631 407019 549999
rect 402810 549311 403637 549631
rect 403981 549311 407019 549631
rect 402810 546631 407019 549311
rect 402810 546311 403637 546631
rect 403981 546311 407019 546631
rect 402810 543631 407019 546311
rect 402810 543311 403637 543631
rect 403981 543311 407019 543631
rect 402810 542847 407019 543311
rect 402810 540631 404127 542847
rect 402810 540311 403637 540631
rect 403981 540375 404127 540631
rect 406587 540375 407019 542847
rect 403981 540311 407019 540375
rect 402810 537631 407019 540311
rect 402810 537311 403637 537631
rect 403981 537311 407019 537631
rect 402810 534631 407019 537311
rect 402810 534311 403637 534631
rect 403981 534311 407019 534631
rect 402810 531899 407019 534311
rect 402810 531631 404127 531899
rect 402810 531311 403637 531631
rect 403981 531311 404127 531631
rect 402810 529427 404127 531311
rect 406587 529427 407019 531899
rect 402810 528631 407019 529427
rect 402810 528311 403637 528631
rect 403981 528311 407019 528631
rect 402810 525631 407019 528311
rect 402810 525311 403637 525631
rect 403981 525311 407019 525631
rect 402810 522631 407019 525311
rect 402810 522311 403637 522631
rect 403981 522311 407019 522631
rect 402810 519631 407019 522311
rect 402810 519311 403637 519631
rect 403981 519311 407019 519631
rect 402810 516631 407019 519311
rect 402810 516311 403637 516631
rect 403981 516311 407019 516631
rect 402810 513631 407019 516311
rect 402810 513311 403637 513631
rect 403981 513311 407019 513631
rect 402810 512949 407019 513311
rect 402810 510631 404173 512949
rect 402810 510311 403637 510631
rect 403981 510477 404173 510631
rect 406633 510477 407019 512949
rect 403981 510311 407019 510477
rect 402810 507631 407019 510311
rect 402810 507311 403637 507631
rect 403981 507311 407019 507631
rect 402810 504631 407019 507311
rect 402810 504311 403637 504631
rect 403981 504311 407019 504631
rect 402810 501631 407019 504311
rect 402810 501311 403637 501631
rect 403981 501311 407019 501631
rect 402810 498631 407019 501311
rect 402810 498311 403637 498631
rect 403981 498311 407019 498631
rect 402810 495631 407019 498311
rect 402810 495311 403637 495631
rect 403981 495311 407019 495631
rect 402810 492631 407019 495311
rect 402810 492311 403637 492631
rect 403981 492311 407019 492631
rect 402810 489631 407019 492311
rect 402810 489311 403637 489631
rect 403981 489311 407019 489631
rect 402810 486631 407019 489311
rect 402810 486311 403637 486631
rect 403981 486413 407019 486631
rect 403981 486311 404454 486413
rect 402810 483941 404454 486311
rect 406914 483941 407019 486413
rect 402810 483631 407019 483941
rect 402810 483311 403637 483631
rect 403981 483311 407019 483631
rect 402810 480631 407019 483311
rect 402810 480311 403637 480631
rect 403981 480311 407019 480631
rect 402810 477631 407019 480311
rect 402810 477311 403637 477631
rect 403981 477311 407019 477631
rect 402810 474631 407019 477311
rect 402810 474311 403637 474631
rect 403981 474311 407019 474631
rect 402810 471631 407019 474311
rect 402810 471311 403637 471631
rect 403981 471311 407019 471631
rect 402810 468631 407019 471311
rect 402810 468311 403637 468631
rect 403981 468311 407019 468631
rect 402810 465631 407019 468311
rect 402810 465311 403637 465631
rect 403981 465311 407019 465631
rect 402810 462631 407019 465311
rect 402810 462311 403637 462631
rect 403981 462311 407019 462631
rect 402810 459631 407019 462311
rect 402810 459311 403637 459631
rect 403981 459311 407019 459631
rect 402810 456631 407019 459311
rect 402810 456311 403637 456631
rect 403981 456311 407019 456631
rect 402810 453631 407019 456311
rect 402810 453311 403637 453631
rect 403981 453311 407019 453631
rect 402810 450631 407019 453311
rect 402810 450311 403637 450631
rect 403981 450311 407019 450631
rect 402810 449968 407019 450311
rect 402810 447631 404475 449968
rect 402810 447311 403637 447631
rect 403981 447496 404475 447631
rect 406935 447496 407019 449968
rect 403981 447311 407019 447496
rect 402810 444631 407019 447311
rect 402810 444311 403637 444631
rect 403981 444311 407019 444631
rect 402810 441631 407019 444311
rect 402810 441311 403637 441631
rect 403981 441311 407019 441631
rect 402810 438631 407019 441311
rect 402810 438311 403637 438631
rect 403981 438311 407019 438631
rect 402810 435631 407019 438311
rect 402810 435311 403637 435631
rect 403981 435311 407019 435631
rect 402810 432631 407019 435311
rect 402810 432311 403637 432631
rect 403981 432311 407019 432631
rect 402810 429631 407019 432311
rect 402810 429311 403637 429631
rect 403981 429311 407019 429631
rect 402810 426631 407019 429311
rect 402810 426311 403637 426631
rect 403981 426311 407019 426631
rect 402810 423631 407019 426311
rect 402810 423311 403637 423631
rect 403981 423311 407019 423631
rect 402810 421609 407019 423311
rect 413052 596839 415512 629759
rect 413052 594427 413076 596839
rect 415488 594427 415512 596839
rect 413052 573865 415512 594427
rect 413052 573841 418000 573865
rect 413052 569039 413174 573841
rect 417976 569039 418000 573841
rect 413052 569015 418000 569039
rect 413052 562210 415512 569015
rect 413052 562186 418180 562210
rect 413052 557384 413354 562186
rect 418156 557384 418180 562186
rect 413052 557360 418180 557384
rect 413052 523255 415512 557360
rect 413052 520843 413076 523255
rect 415488 520843 415512 523255
rect 413052 497271 415512 520843
rect 413052 494859 413076 497271
rect 415488 494859 415512 497271
rect 413052 465307 415512 494859
rect 413052 462895 413076 465307
rect 415488 462895 415512 465307
rect 413052 435874 415512 462895
rect 413052 433462 413076 435874
rect 415488 433462 415512 435874
rect 402810 421585 407291 421609
rect 402810 420631 404807 421585
rect 402810 420311 403637 420631
rect 403981 420311 404807 420631
rect 402810 419113 404807 420311
rect 407267 419113 407291 421585
rect 402810 419089 407291 419113
rect 402810 417631 407019 419089
rect 402810 417311 403637 417631
rect 403981 417311 407019 417631
rect 402810 414631 407019 417311
rect 402810 414311 403637 414631
rect 403981 414311 407019 414631
rect 402810 411631 407019 414311
rect 402810 411311 403637 411631
rect 403981 411311 407019 411631
rect 402810 409721 407019 411311
rect 402810 409697 407057 409721
rect 402810 408631 404573 409697
rect 402810 408311 403637 408631
rect 403981 408311 404573 408631
rect 402810 407225 404573 408311
rect 407033 407225 407057 409697
rect 402810 407201 407057 407225
rect 402810 405631 407019 407201
rect 402810 405311 403637 405631
rect 403981 405311 407019 405631
rect 402810 402631 407019 405311
rect 402810 402311 403637 402631
rect 403981 402311 407019 402631
rect 402810 399631 407019 402311
rect 402810 399311 403637 399631
rect 403981 399311 407019 399631
rect 402810 396631 407019 399311
rect 402810 396311 403637 396631
rect 403981 396311 407019 396631
rect 402810 393631 407019 396311
rect 402810 393311 403637 393631
rect 403981 393311 407019 393631
rect 402810 390631 407019 393311
rect 402810 390311 403637 390631
rect 403981 390311 407019 390631
rect 402810 387631 407019 390311
rect 402810 387311 403637 387631
rect 403981 387311 407019 387631
rect 402810 384631 407019 387311
rect 402810 384311 403637 384631
rect 403981 384311 407019 384631
rect 402810 381631 407019 384311
rect 402810 381311 403637 381631
rect 403981 381311 407019 381631
rect 402810 378631 407019 381311
rect 402810 378311 403637 378631
rect 403981 378311 407019 378631
rect 402810 375631 407019 378311
rect 402810 375311 403637 375631
rect 403981 375311 407019 375631
rect 362730 365840 365245 366160
rect 51523 365286 51843 365310
rect 51523 365014 51547 365286
rect 51819 365014 51843 365286
rect 51523 364990 51843 365014
rect 34053 364736 34373 364760
rect 34053 364464 34077 364736
rect 34349 364464 34373 364736
rect 34053 364440 34373 364464
rect 53818 364704 56737 364728
rect 53818 364432 53842 364704
rect 54114 364432 56737 364704
rect 53818 364408 56737 364432
rect 26624 363591 33713 363911
rect 26624 360911 29084 363591
rect 364925 362320 365245 365840
rect 51523 362286 51843 362310
rect 51523 362014 51547 362286
rect 51819 362014 51843 362286
rect 51523 361990 51843 362014
rect 364901 362296 365269 362320
rect 364901 361976 364925 362296
rect 365245 361976 365269 362296
rect 364901 361952 365269 361976
rect 402810 362181 407019 375311
rect 26624 360591 33713 360911
rect 26624 353309 29084 360591
rect 402810 359709 404519 362181
rect 406979 359709 407019 362181
rect 26624 353285 29140 353309
rect 26624 350813 26656 353285
rect 29116 350813 29140 353285
rect 26624 350789 29140 350813
rect 26624 348780 29084 350789
rect 26558 348756 29084 348780
rect 26558 346284 26582 348756
rect 29042 346284 29084 348756
rect 26558 346260 29084 346284
rect 26624 344270 29084 346260
rect 55307 345732 55627 345756
rect 55307 345460 55331 345732
rect 55603 345460 55627 345732
rect 55307 345436 55627 345460
rect 58307 345732 58627 345756
rect 58307 345460 58331 345732
rect 58603 345460 58627 345732
rect 58307 345436 58627 345460
rect 61307 345732 61627 345756
rect 61307 345460 61331 345732
rect 61603 345460 61627 345732
rect 61307 345436 61627 345460
rect 64307 345732 64627 345756
rect 64307 345460 64331 345732
rect 64603 345460 64627 345732
rect 64307 345436 64627 345460
rect 67307 345732 67627 345756
rect 67307 345460 67331 345732
rect 67603 345460 67627 345732
rect 67307 345436 67627 345460
rect 70307 345732 70627 345756
rect 70307 345460 70331 345732
rect 70603 345460 70627 345732
rect 70307 345436 70627 345460
rect 73307 345732 73627 345756
rect 73307 345460 73331 345732
rect 73603 345460 73627 345732
rect 73307 345436 73627 345460
rect 76307 345732 76627 345756
rect 76307 345460 76331 345732
rect 76603 345460 76627 345732
rect 76307 345436 76627 345460
rect 79307 345732 79627 345756
rect 79307 345460 79331 345732
rect 79603 345460 79627 345732
rect 79307 345436 79627 345460
rect 82307 345732 82627 345756
rect 82307 345460 82331 345732
rect 82603 345460 82627 345732
rect 82307 345436 82627 345460
rect 85307 345732 85627 345756
rect 85307 345460 85331 345732
rect 85603 345460 85627 345732
rect 85307 345436 85627 345460
rect 88307 345732 88627 345756
rect 88307 345460 88331 345732
rect 88603 345460 88627 345732
rect 88307 345436 88627 345460
rect 91307 345732 91627 345756
rect 91307 345460 91331 345732
rect 91603 345460 91627 345732
rect 91307 345436 91627 345460
rect 94307 345732 94627 345756
rect 94307 345460 94331 345732
rect 94603 345460 94627 345732
rect 94307 345436 94627 345460
rect 97307 345732 97627 345756
rect 97307 345460 97331 345732
rect 97603 345460 97627 345732
rect 97307 345436 97627 345460
rect 100307 345732 100627 345756
rect 100307 345460 100331 345732
rect 100603 345460 100627 345732
rect 100307 345436 100627 345460
rect 103307 345732 103627 345756
rect 103307 345460 103331 345732
rect 103603 345460 103627 345732
rect 103307 345436 103627 345460
rect 106307 345732 106627 345756
rect 106307 345460 106331 345732
rect 106603 345460 106627 345732
rect 106307 345436 106627 345460
rect 109307 345732 109627 345756
rect 109307 345460 109331 345732
rect 109603 345460 109627 345732
rect 109307 345436 109627 345460
rect 112307 345732 112627 345756
rect 112307 345460 112331 345732
rect 112603 345460 112627 345732
rect 112307 345436 112627 345460
rect 115307 345732 115627 345756
rect 115307 345460 115331 345732
rect 115603 345460 115627 345732
rect 115307 345436 115627 345460
rect 118307 345732 118627 345756
rect 118307 345460 118331 345732
rect 118603 345460 118627 345732
rect 118307 345436 118627 345460
rect 121307 345732 121627 345756
rect 121307 345460 121331 345732
rect 121603 345460 121627 345732
rect 121307 345436 121627 345460
rect 124307 345732 124627 345756
rect 124307 345460 124331 345732
rect 124603 345460 124627 345732
rect 124307 345436 124627 345460
rect 127307 345732 127627 345756
rect 127307 345460 127331 345732
rect 127603 345460 127627 345732
rect 127307 345436 127627 345460
rect 130307 345732 130627 345756
rect 130307 345460 130331 345732
rect 130603 345460 130627 345732
rect 130307 345436 130627 345460
rect 133307 345732 133627 345756
rect 133307 345460 133331 345732
rect 133603 345460 133627 345732
rect 133307 345436 133627 345460
rect 136307 345732 136627 345756
rect 136307 345460 136331 345732
rect 136603 345460 136627 345732
rect 136307 345436 136627 345460
rect 139307 345732 139627 345756
rect 139307 345460 139331 345732
rect 139603 345460 139627 345732
rect 139307 345436 139627 345460
rect 142307 345732 142627 345756
rect 142307 345460 142331 345732
rect 142603 345460 142627 345732
rect 142307 345436 142627 345460
rect 145307 345732 145627 345756
rect 145307 345460 145331 345732
rect 145603 345460 145627 345732
rect 145307 345436 145627 345460
rect 148307 345732 148627 345756
rect 148307 345460 148331 345732
rect 148603 345460 148627 345732
rect 148307 345436 148627 345460
rect 151307 345732 151627 345756
rect 151307 345460 151331 345732
rect 151603 345460 151627 345732
rect 151307 345436 151627 345460
rect 154307 345732 154627 345756
rect 154307 345460 154331 345732
rect 154603 345460 154627 345732
rect 154307 345436 154627 345460
rect 157307 345732 157627 345756
rect 157307 345460 157331 345732
rect 157603 345460 157627 345732
rect 157307 345436 157627 345460
rect 160307 345732 160627 345756
rect 160307 345460 160331 345732
rect 160603 345460 160627 345732
rect 160307 345436 160627 345460
rect 163307 345732 163627 345756
rect 163307 345460 163331 345732
rect 163603 345460 163627 345732
rect 163307 345436 163627 345460
rect 166307 345732 166627 345756
rect 166307 345460 166331 345732
rect 166603 345460 166627 345732
rect 166307 345436 166627 345460
rect 169307 345732 169627 345756
rect 169307 345460 169331 345732
rect 169603 345460 169627 345732
rect 169307 345436 169627 345460
rect 172307 345732 172627 345756
rect 172307 345460 172331 345732
rect 172603 345460 172627 345732
rect 172307 345436 172627 345460
rect 175307 345732 175627 345756
rect 175307 345460 175331 345732
rect 175603 345460 175627 345732
rect 175307 345436 175627 345460
rect 178307 345732 178627 345756
rect 178307 345460 178331 345732
rect 178603 345460 178627 345732
rect 178307 345436 178627 345460
rect 181307 345732 181627 345756
rect 181307 345460 181331 345732
rect 181603 345460 181627 345732
rect 181307 345436 181627 345460
rect 184307 345732 184627 345756
rect 184307 345460 184331 345732
rect 184603 345460 184627 345732
rect 184307 345436 184627 345460
rect 187307 345732 187627 345756
rect 187307 345460 187331 345732
rect 187603 345460 187627 345732
rect 187307 345436 187627 345460
rect 190307 345732 190627 345756
rect 190307 345460 190331 345732
rect 190603 345460 190627 345732
rect 190307 345436 190627 345460
rect 193307 345732 193627 345756
rect 193307 345460 193331 345732
rect 193603 345460 193627 345732
rect 193307 345436 193627 345460
rect 196307 345732 196627 345756
rect 196307 345460 196331 345732
rect 196603 345460 196627 345732
rect 196307 345436 196627 345460
rect 199307 345732 199627 345756
rect 199307 345460 199331 345732
rect 199603 345460 199627 345732
rect 199307 345436 199627 345460
rect 202307 345732 202627 345756
rect 202307 345460 202331 345732
rect 202603 345460 202627 345732
rect 202307 345436 202627 345460
rect 205307 345732 205627 345756
rect 205307 345460 205331 345732
rect 205603 345460 205627 345732
rect 205307 345436 205627 345460
rect 208307 345732 208627 345756
rect 208307 345460 208331 345732
rect 208603 345460 208627 345732
rect 208307 345436 208627 345460
rect 211307 345732 211627 345756
rect 211307 345460 211331 345732
rect 211603 345460 211627 345732
rect 211307 345436 211627 345460
rect 214307 345732 214627 345756
rect 214307 345460 214331 345732
rect 214603 345460 214627 345732
rect 214307 345436 214627 345460
rect 217307 345732 217627 345756
rect 217307 345460 217331 345732
rect 217603 345460 217627 345732
rect 217307 345436 217627 345460
rect 220307 345732 220627 345756
rect 220307 345460 220331 345732
rect 220603 345460 220627 345732
rect 220307 345436 220627 345460
rect 223307 345732 223627 345756
rect 223307 345460 223331 345732
rect 223603 345460 223627 345732
rect 223307 345436 223627 345460
rect 226307 345732 226627 345756
rect 226307 345460 226331 345732
rect 226603 345460 226627 345732
rect 226307 345436 226627 345460
rect 229307 345732 229627 345756
rect 229307 345460 229331 345732
rect 229603 345460 229627 345732
rect 229307 345436 229627 345460
rect 232307 345732 232627 345756
rect 232307 345460 232331 345732
rect 232603 345460 232627 345732
rect 232307 345436 232627 345460
rect 235307 345732 235627 345756
rect 235307 345460 235331 345732
rect 235603 345460 235627 345732
rect 235307 345436 235627 345460
rect 238307 345732 238627 345756
rect 238307 345460 238331 345732
rect 238603 345460 238627 345732
rect 238307 345436 238627 345460
rect 241307 345732 241627 345756
rect 241307 345460 241331 345732
rect 241603 345460 241627 345732
rect 241307 345436 241627 345460
rect 244307 345732 244627 345756
rect 244307 345460 244331 345732
rect 244603 345460 244627 345732
rect 244307 345436 244627 345460
rect 247307 345732 247627 345756
rect 247307 345460 247331 345732
rect 247603 345460 247627 345732
rect 247307 345436 247627 345460
rect 250307 345732 250627 345756
rect 250307 345460 250331 345732
rect 250603 345460 250627 345732
rect 250307 345436 250627 345460
rect 253307 345732 253627 345756
rect 253307 345460 253331 345732
rect 253603 345460 253627 345732
rect 253307 345436 253627 345460
rect 256307 345732 256627 345756
rect 256307 345460 256331 345732
rect 256603 345460 256627 345732
rect 256307 345436 256627 345460
rect 259307 345732 259627 345756
rect 259307 345460 259331 345732
rect 259603 345460 259627 345732
rect 259307 345436 259627 345460
rect 262307 345732 262627 345756
rect 262307 345460 262331 345732
rect 262603 345460 262627 345732
rect 262307 345436 262627 345460
rect 265307 345732 265627 345756
rect 265307 345460 265331 345732
rect 265603 345460 265627 345732
rect 265307 345436 265627 345460
rect 268307 345732 268627 345756
rect 268307 345460 268331 345732
rect 268603 345460 268627 345732
rect 268307 345436 268627 345460
rect 271307 345732 271627 345756
rect 271307 345460 271331 345732
rect 271603 345460 271627 345732
rect 271307 345436 271627 345460
rect 274307 345732 274627 345756
rect 274307 345460 274331 345732
rect 274603 345460 274627 345732
rect 274307 345436 274627 345460
rect 277307 345732 277627 345756
rect 277307 345460 277331 345732
rect 277603 345460 277627 345732
rect 277307 345436 277627 345460
rect 280307 345732 280627 345756
rect 280307 345460 280331 345732
rect 280603 345460 280627 345732
rect 280307 345436 280627 345460
rect 283307 345732 283627 345756
rect 283307 345460 283331 345732
rect 283603 345460 283627 345732
rect 283307 345436 283627 345460
rect 286307 345732 286627 345756
rect 286307 345460 286331 345732
rect 286603 345460 286627 345732
rect 286307 345436 286627 345460
rect 289307 345732 289627 345756
rect 289307 345460 289331 345732
rect 289603 345460 289627 345732
rect 289307 345436 289627 345460
rect 292307 345732 292627 345756
rect 292307 345460 292331 345732
rect 292603 345460 292627 345732
rect 292307 345436 292627 345460
rect 295307 345732 295627 345756
rect 295307 345460 295331 345732
rect 295603 345460 295627 345732
rect 295307 345436 295627 345460
rect 298307 345732 298627 345756
rect 298307 345460 298331 345732
rect 298603 345460 298627 345732
rect 298307 345436 298627 345460
rect 301307 345732 301627 345756
rect 301307 345460 301331 345732
rect 301603 345460 301627 345732
rect 301307 345436 301627 345460
rect 304307 345732 304627 345756
rect 304307 345460 304331 345732
rect 304603 345460 304627 345732
rect 304307 345436 304627 345460
rect 307307 345732 307627 345756
rect 307307 345460 307331 345732
rect 307603 345460 307627 345732
rect 307307 345436 307627 345460
rect 310307 345732 310627 345756
rect 310307 345460 310331 345732
rect 310603 345460 310627 345732
rect 310307 345436 310627 345460
rect 313307 345732 313627 345756
rect 313307 345460 313331 345732
rect 313603 345460 313627 345732
rect 313307 345436 313627 345460
rect 316307 345732 316627 345756
rect 316307 345460 316331 345732
rect 316603 345460 316627 345732
rect 316307 345436 316627 345460
rect 319307 345732 319627 345756
rect 319307 345460 319331 345732
rect 319603 345460 319627 345732
rect 319307 345436 319627 345460
rect 325307 345732 325627 345756
rect 325307 345460 325331 345732
rect 325603 345460 325627 345732
rect 325307 345436 325627 345460
rect 328307 345732 328627 345756
rect 328307 345460 328331 345732
rect 328603 345460 328627 345732
rect 328307 345436 328627 345460
rect 331307 345732 331627 345756
rect 331307 345460 331331 345732
rect 331603 345460 331627 345732
rect 331307 345436 331627 345460
rect 334307 345732 334627 345756
rect 334307 345460 334331 345732
rect 334603 345460 334627 345732
rect 334307 345436 334627 345460
rect 337307 345732 337627 345756
rect 337307 345460 337331 345732
rect 337603 345460 337627 345732
rect 337307 345436 337627 345460
rect 340307 345732 340627 345756
rect 340307 345460 340331 345732
rect 340603 345460 340627 345732
rect 340307 345436 340627 345460
rect 343307 345732 343627 345756
rect 343307 345460 343331 345732
rect 343603 345460 343627 345732
rect 343307 345436 343627 345460
rect 346307 345732 346627 345756
rect 346307 345460 346331 345732
rect 346603 345460 346627 345732
rect 346307 345436 346627 345460
rect 349307 345732 349627 345756
rect 349307 345460 349331 345732
rect 349603 345460 349627 345732
rect 349307 345436 349627 345460
rect 352307 345732 352627 345756
rect 352307 345460 352331 345732
rect 352603 345460 352627 345732
rect 352307 345436 352627 345460
rect 355307 345732 355627 345756
rect 355307 345460 355331 345732
rect 355603 345460 355627 345732
rect 355307 345436 355627 345460
rect 358307 345732 358627 345756
rect 358307 345460 358331 345732
rect 358603 345460 358627 345732
rect 358307 345436 358627 345460
rect 26558 344246 29084 344270
rect 26558 341774 26582 344246
rect 29042 341774 29084 344246
rect 26558 341750 29084 341774
rect 14675 337915 14740 340672
rect 17497 337915 20482 340672
rect 14675 324591 20482 337915
rect 26624 338142 29084 341750
rect 56876 338142 57196 345096
rect 59876 338142 60196 345096
rect 62876 338142 63196 345096
rect 65876 338142 66196 345096
rect 68876 338142 69196 345096
rect 71876 338142 72196 345096
rect 74876 338142 75196 345096
rect 77876 338142 78196 345096
rect 80876 338142 81196 345096
rect 83876 338142 84196 345096
rect 86876 338142 87196 345096
rect 89876 338142 90196 345096
rect 92876 338142 93196 345096
rect 95876 338142 96196 345096
rect 98876 338142 99196 345096
rect 101876 338142 102196 345096
rect 104876 338142 105196 345096
rect 107876 338142 108196 345096
rect 110876 338142 111196 345096
rect 113876 338142 114196 345096
rect 116876 338142 117196 345096
rect 119876 338142 120196 345096
rect 122876 338142 123196 345096
rect 125876 338142 126196 345096
rect 128876 338142 129196 345096
rect 131876 338142 132196 345096
rect 134876 338142 135196 345096
rect 137876 338142 138196 345096
rect 140876 338142 141196 345096
rect 143876 338142 144196 345096
rect 146876 338142 147196 345096
rect 149876 338142 150196 345096
rect 152876 338142 153196 345096
rect 155876 338142 156196 345096
rect 158876 338142 159196 345096
rect 161876 338142 162196 345096
rect 164876 338142 165196 345096
rect 167876 338142 168196 345096
rect 170876 338142 171196 345096
rect 173876 338142 174196 345096
rect 176876 338142 177196 345096
rect 179876 338142 180196 345096
rect 182876 338142 183196 345096
rect 185876 338142 186196 345096
rect 188876 338142 189196 345096
rect 191876 338142 192196 345096
rect 194876 338142 195196 345096
rect 197876 338142 198196 345096
rect 200876 338142 201196 345096
rect 203876 338142 204196 345096
rect 206876 338142 207196 345096
rect 209876 338142 210196 345096
rect 212876 338142 213196 345096
rect 215876 338142 216196 345096
rect 218876 338142 219196 345096
rect 221876 338142 222196 345096
rect 224876 338142 225196 345096
rect 227876 338142 228196 345096
rect 230876 338142 231196 345096
rect 233876 338142 234196 345096
rect 236876 338142 237196 345096
rect 239876 338142 240196 345096
rect 242876 338142 243196 345096
rect 245876 338142 246196 345096
rect 248876 338142 249196 345096
rect 251876 338142 252196 345096
rect 254876 338142 255196 345096
rect 257876 338142 258196 345096
rect 260876 338142 261196 345096
rect 263876 338142 264196 345096
rect 266876 338142 267196 345096
rect 269876 338142 270196 345096
rect 272876 338142 273196 345096
rect 275876 338142 276196 345096
rect 278876 338142 279196 345096
rect 281876 338142 282196 345096
rect 284876 338142 285196 345096
rect 287876 338142 288196 345096
rect 290876 338142 291196 345096
rect 293876 338142 294196 345096
rect 296876 338142 297196 345096
rect 299876 338142 300196 345096
rect 302876 338142 303196 345096
rect 305876 338142 306196 345096
rect 308876 338142 309196 345096
rect 311876 338142 312196 345096
rect 314876 338142 315196 345096
rect 317876 338142 318196 345096
rect 320876 338142 321196 345096
rect 323876 338142 324196 345096
rect 326876 338142 327196 345096
rect 329876 338142 330196 345096
rect 332876 338142 333196 345096
rect 335876 338142 336196 345096
rect 338876 338142 339196 345096
rect 341876 338142 342196 345096
rect 344876 338142 345196 345096
rect 347876 338142 348196 345096
rect 350876 338142 351196 345096
rect 353876 338142 354196 345096
rect 356876 338142 357196 345096
rect 359876 338142 360196 345096
rect 402810 338142 407019 359709
rect 26624 336914 407019 338142
rect 26624 336594 372476 336914
rect 372796 336594 375476 336914
rect 375796 336594 378476 336914
rect 378796 336594 381476 336914
rect 381796 336594 384476 336914
rect 384796 336594 387476 336914
rect 387796 336594 390476 336914
rect 390796 336594 393476 336914
rect 393796 336594 396476 336914
rect 396796 336594 407019 336914
rect 26624 335682 407019 336594
rect 413052 399771 415512 433462
rect 413052 397359 413076 399771
rect 415488 397359 415512 399771
rect 413052 385744 415512 397359
rect 413052 383332 413076 385744
rect 415488 383332 415512 385744
rect 413052 377777 415512 383332
rect 413052 377457 414088 377777
rect 414408 377457 415512 377777
rect 413052 377090 415512 377457
rect 413052 376770 413980 377090
rect 414300 376770 415512 377090
rect 413052 376223 415512 376770
rect 413052 375903 414233 376223
rect 414553 375903 415512 376223
rect 413052 374668 415512 375903
rect 413052 374348 414016 374668
rect 414336 374348 415512 374668
rect 413052 374069 415512 374348
rect 413052 373749 413984 374069
rect 414304 373749 415512 374069
rect 413052 373209 415512 373749
rect 413052 372889 414342 373209
rect 414662 372889 415512 373209
rect 413052 372492 415512 372889
rect 413052 372172 414235 372492
rect 414555 372172 415512 372492
rect 413052 371847 415512 372172
rect 413052 371527 414342 371847
rect 414662 371527 415512 371847
rect 413052 371310 415512 371527
rect 413052 370990 414766 371310
rect 415086 370990 415512 371310
rect 413052 370719 415512 370990
rect 413052 370399 413762 370719
rect 414082 370399 415512 370719
rect 413052 324591 415512 370399
rect 14675 323421 415512 324591
rect 14675 323101 55301 323421
rect 55633 323101 58301 323421
rect 58633 323101 61301 323421
rect 61633 323101 64301 323421
rect 64633 323101 67301 323421
rect 67633 323101 70301 323421
rect 70633 323101 73301 323421
rect 73633 323101 76301 323421
rect 76633 323101 79301 323421
rect 79633 323101 82301 323421
rect 82633 323101 85301 323421
rect 85633 323101 88301 323421
rect 88633 323101 91301 323421
rect 91633 323101 94301 323421
rect 94633 323101 97301 323421
rect 97633 323101 100301 323421
rect 100633 323101 103301 323421
rect 103633 323101 106301 323421
rect 106633 323101 109301 323421
rect 109633 323101 112301 323421
rect 112633 323101 115301 323421
rect 115633 323101 118301 323421
rect 118633 323101 121301 323421
rect 121633 323101 124301 323421
rect 124633 323101 127301 323421
rect 127633 323101 130301 323421
rect 130633 323101 133301 323421
rect 133633 323101 136301 323421
rect 136633 323101 139301 323421
rect 139633 323101 142301 323421
rect 142633 323101 145301 323421
rect 145633 323101 148301 323421
rect 148633 323101 151301 323421
rect 151633 323101 154301 323421
rect 154633 323101 157301 323421
rect 157633 323101 160301 323421
rect 160633 323101 163301 323421
rect 163633 323101 166301 323421
rect 166633 323101 169301 323421
rect 169633 323101 172301 323421
rect 172633 323101 175301 323421
rect 175633 323101 178301 323421
rect 178633 323101 181301 323421
rect 181633 323101 184301 323421
rect 184633 323101 187301 323421
rect 187633 323101 190301 323421
rect 190633 323101 193301 323421
rect 193633 323101 196301 323421
rect 196633 323101 199301 323421
rect 199633 323101 202301 323421
rect 202633 323101 205301 323421
rect 205633 323101 208301 323421
rect 208633 323101 211301 323421
rect 211633 323101 214301 323421
rect 214633 323101 217301 323421
rect 217633 323101 220301 323421
rect 220633 323101 223301 323421
rect 223633 323101 226301 323421
rect 226633 323101 228301 323421
rect 228633 323101 229301 323421
rect 229633 323101 232301 323421
rect 232633 323101 235301 323421
rect 235633 323101 238301 323421
rect 238633 323101 241301 323421
rect 241633 323101 244301 323421
rect 244633 323101 247301 323421
rect 247633 323101 250301 323421
rect 250633 323101 253301 323421
rect 253633 323101 256301 323421
rect 256633 323101 258301 323421
rect 258633 323101 259301 323421
rect 259633 323101 262301 323421
rect 262633 323101 265301 323421
rect 265633 323101 268301 323421
rect 268633 323101 269301 323421
rect 269633 323101 271301 323421
rect 271633 323101 274301 323421
rect 274633 323101 277301 323421
rect 277633 323101 278301 323421
rect 278633 323101 279301 323421
rect 279633 323101 280301 323421
rect 280633 323101 283301 323421
rect 283633 323101 286301 323421
rect 286633 323101 288301 323421
rect 288633 323101 289301 323421
rect 289633 323101 292301 323421
rect 292633 323101 295301 323421
rect 295633 323101 298301 323421
rect 298633 323101 299301 323421
rect 299633 323101 301301 323421
rect 301633 323101 304301 323421
rect 304633 323101 307301 323421
rect 307633 323101 310301 323421
rect 310633 323101 313301 323421
rect 313633 323101 316301 323421
rect 316633 323101 318301 323421
rect 318633 323101 319301 323421
rect 319633 323101 325301 323421
rect 325633 323101 328301 323421
rect 328633 323101 329301 323421
rect 329633 323101 331301 323421
rect 331633 323101 334301 323421
rect 334633 323101 337301 323421
rect 337633 323101 338301 323421
rect 338633 323101 339301 323421
rect 339633 323101 340301 323421
rect 340633 323101 343301 323421
rect 343633 323101 346301 323421
rect 346633 323101 348301 323421
rect 348633 323101 349301 323421
rect 349633 323101 352301 323421
rect 352633 323101 355301 323421
rect 355633 323101 358301 323421
rect 358633 323101 415512 323421
rect 14675 322264 415512 323101
rect 18022 322131 415512 322264
rect 39918 315921 42426 315945
rect 39918 313449 39942 315921
rect 42402 315915 42426 315921
rect 42402 315891 146461 315915
rect 42402 313479 97448 315891
rect 99860 313479 120141 315891
rect 122553 313479 143560 315891
rect 145972 313479 146461 315891
rect 42402 313455 146461 313479
rect 42402 313449 42426 313455
rect 39918 313425 42426 313449
rect 6988 243835 7356 243859
rect 6988 243515 7012 243835
rect 7332 243515 7356 243835
rect 6988 243491 7356 243515
rect 86852 230726 89312 230750
rect 86852 228314 86876 230726
rect 89288 228314 89312 230726
rect 86852 196031 89312 228314
rect 151706 208108 153468 322131
rect 158597 208108 160359 322131
rect 161597 208108 163359 322131
rect 164597 208108 166359 322131
rect 167597 208108 169359 322131
rect 170597 208108 172359 322131
rect 176597 208108 178359 322131
rect 182597 208108 184359 322131
rect 217963 208108 220423 322131
rect 227963 208108 230423 322131
rect 237963 208108 240423 322131
rect 247963 208108 250423 322131
rect 257963 208108 260423 322131
rect 267963 208108 270423 322131
rect 277963 208108 280423 322131
rect 287963 208108 290423 322131
rect 297963 208108 300423 322131
rect 307963 208108 310423 322131
rect 317963 208108 320423 322131
rect 327963 208108 330423 322131
rect 337963 208108 340423 322131
rect 347963 208108 350423 322131
rect 357963 208108 360423 322131
rect 367963 208108 370423 322131
rect 377963 208108 380423 322131
rect 387963 208108 390423 322131
rect 397963 208108 400423 322131
rect 407963 208108 410423 322131
rect 451369 208108 456169 629759
rect 151706 207499 456169 208108
rect 151706 207381 173401 207499
rect 151706 207157 170811 207381
rect 151706 206837 167887 207157
rect 168209 207061 170811 207157
rect 171133 207179 173401 207381
rect 173723 207381 456169 207499
rect 173723 207179 176811 207381
rect 171133 207061 176811 207179
rect 177133 207310 182811 207381
rect 177133 207061 180906 207310
rect 168209 206990 180906 207061
rect 181226 207061 182811 207310
rect 183133 207310 456169 207381
rect 183133 207061 183906 207310
rect 181226 206990 183906 207061
rect 184226 206990 186906 207310
rect 187226 206990 189906 207310
rect 190226 206990 192906 207310
rect 193226 206990 195906 207310
rect 196226 206990 198906 207310
rect 199226 206990 201906 207310
rect 202226 206990 204906 207310
rect 205226 206990 456169 207310
rect 168209 206837 456169 206990
rect 151706 206346 456169 206837
rect 86852 194269 87328 196031
rect 89090 194269 89312 196031
rect 86852 177688 89312 194269
rect 142234 198033 142554 198057
rect 142234 197761 142258 198033
rect 142530 197761 142554 198033
rect 142234 191061 142554 197761
rect 142210 191037 142578 191061
rect 142210 190717 142234 191037
rect 142554 190717 142578 191037
rect 142210 190693 142578 190717
rect 151706 188999 153468 206346
rect 163189 205852 163509 206346
rect 216497 205955 220423 206346
rect 227963 205955 230423 206346
rect 237963 205955 240423 206346
rect 247963 205955 250423 206346
rect 257963 205955 260423 206346
rect 267963 205955 270423 206346
rect 277963 205955 280423 206346
rect 287963 205955 290423 206346
rect 297963 205955 300423 206346
rect 307963 205955 310423 206346
rect 317963 205955 320423 206346
rect 327963 205955 330423 206346
rect 337963 205955 340423 206346
rect 347963 205955 350423 206346
rect 357963 205955 360423 206346
rect 367963 205955 370423 206346
rect 377963 205955 380423 206346
rect 387963 205955 390423 206346
rect 397963 205955 400423 206346
rect 407963 205955 410423 206346
rect 163165 205828 163533 205852
rect 163165 205508 163189 205828
rect 163509 205508 163533 205828
rect 163165 205484 163533 205508
rect 151706 188679 152727 188999
rect 153047 188679 153468 188999
rect 151706 185846 153468 188679
rect 151706 185526 152760 185846
rect 153080 185526 153468 185846
rect 151706 183154 153468 185526
rect 151706 182834 152494 183154
rect 152814 182834 153468 183154
rect 151706 180627 153468 182834
rect 151706 180307 152719 180627
rect 153039 180307 153468 180627
rect 85191 172888 89994 177688
rect 85191 169097 89991 172888
rect 85191 168038 86590 169097
rect 86566 166635 86590 168038
rect 89050 168038 89991 169097
rect 151706 169070 153468 180307
rect 156179 203679 212769 203703
rect 156179 201965 156565 203679
rect 158279 201965 174334 203679
rect 176048 201965 178443 203679
rect 180157 201965 190981 203679
rect 192695 201965 207523 203679
rect 209237 201965 212769 203679
rect 156179 201941 212769 201965
rect 156179 196007 157941 201941
rect 156179 194293 156203 196007
rect 157917 194293 157941 196007
rect 156179 193227 157941 194293
rect 162363 193377 162683 201941
rect 165363 193377 165683 201941
rect 168363 193377 168683 201941
rect 171363 193377 171683 201941
rect 174363 193377 174683 201941
rect 156179 192907 162261 193227
rect 156179 190227 157941 192907
rect 163189 192163 163509 192187
rect 163189 191891 163213 192163
rect 163485 191891 163509 192163
rect 163189 191867 163509 191891
rect 167888 192163 168208 192187
rect 167888 191891 167912 192163
rect 168184 191891 168208 192163
rect 167888 191867 168208 191891
rect 170812 192163 171132 192187
rect 170812 191891 170836 192163
rect 171108 191891 171132 192163
rect 170812 191867 171132 191891
rect 173402 192163 173722 192187
rect 173402 191891 173426 192163
rect 173698 191891 173722 192163
rect 173402 191867 173722 191891
rect 163693 191013 164013 191037
rect 163693 190741 163717 191013
rect 163989 190741 164013 191013
rect 163693 190717 164013 190741
rect 156179 189907 162261 190227
rect 156179 187227 157941 189907
rect 162811 188975 163131 188999
rect 162811 188703 162835 188975
rect 163107 188703 163131 188975
rect 162811 188679 163131 188703
rect 156179 186907 162261 187227
rect 156179 184227 157941 186907
rect 162811 185822 163131 185846
rect 162811 185550 162835 185822
rect 163107 185550 163131 185822
rect 162811 185526 163131 185550
rect 156179 183907 162261 184227
rect 156179 181227 157941 183907
rect 162811 183130 163131 183154
rect 162811 182858 162835 183130
rect 163107 182858 163131 183130
rect 162811 182834 163131 182858
rect 156179 180907 162261 181227
rect 156179 173279 157941 180907
rect 162841 180603 163161 180627
rect 162841 180331 162865 180603
rect 163137 180331 163161 180603
rect 162841 180307 163161 180331
rect 164431 180603 164751 180627
rect 164431 180331 164455 180603
rect 164727 180331 164751 180603
rect 164431 180307 164751 180331
rect 167772 180603 168092 180627
rect 167772 180331 167796 180603
rect 168068 180331 168092 180603
rect 167772 180307 168092 180331
rect 170722 180603 171042 180627
rect 170722 180331 170746 180603
rect 171018 180331 171042 180603
rect 170722 180307 171042 180331
rect 173032 180603 173352 180627
rect 173032 180331 173056 180603
rect 173328 180331 173352 180603
rect 173032 180307 173352 180331
rect 175008 180603 175328 180627
rect 175008 180331 175032 180603
rect 175304 180331 175328 180603
rect 175008 180307 175328 180331
rect 156179 171565 156203 173279
rect 157917 173070 157941 173279
rect 162435 173070 162755 179597
rect 165435 173070 165755 179597
rect 168435 173070 168755 179597
rect 171435 173070 171755 179597
rect 174435 173070 174755 179597
rect 211007 173070 212769 201941
rect 157917 173046 212769 173070
rect 157917 171565 162536 173046
rect 156179 171332 162536 171565
rect 164250 171332 177721 173046
rect 179435 172824 196503 173046
rect 179435 172504 180867 172824
rect 181187 172504 183867 172824
rect 184187 172504 186867 172824
rect 187187 172504 189867 172824
rect 190187 172504 192867 172824
rect 193187 172504 195867 172824
rect 196187 172504 196503 172824
rect 179435 171332 196503 172504
rect 198217 172824 207692 173046
rect 198217 172504 198867 172824
rect 199187 172504 201867 172824
rect 202187 172504 204867 172824
rect 205187 172504 207692 172824
rect 198217 171332 207692 172504
rect 209406 171332 212769 173046
rect 156179 171308 212769 171332
rect 216497 200014 218259 205955
rect 451369 200014 456169 206346
rect 216497 195214 456169 200014
rect 216497 180548 218259 195214
rect 451369 180548 456169 195214
rect 216497 175748 456169 180548
rect 156179 170901 157941 171308
rect 216497 169070 218259 175748
rect 451369 169070 456169 175748
rect 460694 169070 465494 629759
rect 151638 168528 465494 169070
rect 151638 168315 170721 168528
rect 89050 166635 89312 168038
rect 151638 167995 164430 168315
rect 164752 168208 170721 168315
rect 171043 168246 465494 168528
rect 171043 168244 175009 168246
rect 171043 168208 173031 168244
rect 164752 168173 173031 168208
rect 164752 167995 167771 168173
rect 151638 167853 167771 167995
rect 168093 167924 173031 168173
rect 173353 167924 175009 168244
rect 175329 167924 465494 168246
rect 168093 167853 465494 167924
rect 151638 167308 465494 167853
rect 501550 222136 504010 668401
rect 573820 222137 578668 222161
rect 573820 222136 573844 222137
rect 501550 217336 573844 222136
rect 501550 204057 504010 217336
rect 573820 217335 573844 217336
rect 578644 217335 578668 222137
rect 573820 217311 578668 217335
rect 573845 204082 578645 217311
rect 573845 204058 579092 204082
rect 573845 204057 574268 204058
rect 501550 199257 574268 204057
rect 501550 196255 504010 199257
rect 573845 199256 574268 199257
rect 579068 199256 579092 204058
rect 573845 199232 579092 199256
rect 501550 196231 504563 196255
rect 501550 193769 502079 196231
rect 504539 193915 504563 196231
rect 504539 193891 504585 193915
rect 501550 191429 502101 193769
rect 504561 191429 504585 193891
rect 573845 191430 579069 199232
rect 501550 191405 504585 191429
rect 501550 186255 504010 191405
rect 501550 186231 504874 186255
rect 501550 183769 502390 186231
rect 504850 183915 504874 186231
rect 504850 183891 505038 183915
rect 501550 181429 502554 183769
rect 505014 181429 505038 183891
rect 501550 181405 505038 181429
rect 501550 167476 504010 181405
rect 573820 167477 578668 167501
rect 573820 167476 573844 167477
rect 86566 166611 89312 166635
rect 86852 165373 89312 166611
rect 86421 165349 89312 165373
rect 86421 162887 86445 165349
rect 88905 162887 89312 165349
rect 151706 164937 153468 167308
rect 86421 162863 89312 162887
rect 86852 154479 89312 162863
rect 86699 154455 89312 154479
rect 86699 151993 86723 154455
rect 89183 151993 89312 154455
rect 86699 151969 89312 151993
rect 86852 136534 89312 151969
rect 159987 145835 161749 167308
rect 177972 145835 179734 167308
rect 189716 145835 191478 167308
rect 203103 145835 204865 167308
rect 214682 145835 216444 167308
rect 451369 165690 456169 167308
rect 460694 145835 465494 167308
rect 501529 162676 573844 167476
rect 154774 141035 465494 145835
rect 501550 149372 504010 162676
rect 573820 162675 573844 162676
rect 578644 162675 578668 167477
rect 573820 162651 578668 162675
rect 501550 149348 504304 149372
rect 501550 146886 501820 149348
rect 504280 146886 504304 149348
rect 501550 146862 504304 146886
rect 86699 136510 89312 136534
rect 86699 134048 86723 136510
rect 89183 134048 89312 136510
rect 86699 134024 89312 134048
rect 13357 124806 15865 124830
rect 86852 124806 89312 134024
rect 501550 139315 504010 146862
rect 501550 139291 504527 139315
rect 501550 136829 502043 139291
rect 504503 136829 504527 139291
rect 501550 136805 504527 136829
rect 13357 122346 13381 124806
rect 15841 122346 89377 124806
rect 13357 122322 15865 122346
rect 86852 118008 89312 122346
rect 287934 118952 290454 118976
rect 287934 118008 287958 118952
rect 86852 117757 287958 118008
rect 86852 115995 156179 117757
rect 157941 117557 287958 117757
rect 157941 117457 207668 117557
rect 157941 115995 162512 117457
rect 86852 115695 162512 115995
rect 164274 117058 196479 117457
rect 164274 115695 177697 117058
rect 86852 115548 177697 115695
rect 177673 115296 177697 115548
rect 179459 115695 196479 117058
rect 198241 115795 207668 117457
rect 209430 116492 287958 117557
rect 290430 118008 290454 118952
rect 501550 118008 504010 136805
rect 290430 116492 504010 118008
rect 209430 115795 504010 116492
rect 198241 115695 504010 115795
rect 179459 115548 504010 115695
rect 179459 115296 179483 115548
rect 177673 115272 179483 115296
use array_SR  array_SR_0
timestamp 1663269944
transform 1 0 54469 0 1 344190
box -21076 586 308046 327367
use bias  bias_0
timestamp 1655248036
transform 1 0 145381 0 1 675880
box 790 -2236 7180 -220
use opamp_wrapper  opamp_wrapper_0
timestamp 1655248036
transform 1 0 369481 0 1 359134
box -2280 -1640 26995 13665
use opamp_wrapper  opamp_wrapper_1
timestamp 1655248036
transform 1 0 179353 0 1 180877
box -2280 -1640 26995 13665
use pixel_array  pixel_array_0
timestamp 1655251226
transform 1 0 165661 0 1 187877
box -3720 -8600 11230 5820
<< labels >>
flabel metal3 s -800 381864 480 381976 0 FreeSans 1400 0 0 0 gpio_analog[10]
port 2 nsew
flabel metal3 s -800 338642 480 338754 0 FreeSans 1400 0 0 0 gpio_analog[11]
port 3 nsew
flabel metal3 s -800 295420 480 295532 0 FreeSans 1400 0 0 0 gpio_analog[12]
port 4 nsew
flabel metal3 s -800 252398 480 252510 0 FreeSans 1400 0 0 0 gpio_analog[13]
port 5 nsew
flabel metal3 s -800 124776 480 124888 0 FreeSans 1400 0 0 0 gpio_analog[14]
port 6 nsew
flabel metal3 s -800 81554 480 81666 0 FreeSans 1400 0 0 0 gpio_analog[15]
port 7 nsew
flabel metal3 s -800 38332 480 38444 0 FreeSans 1400 0 0 0 gpio_analog[16]
port 8 nsew
flabel metal3 s -800 16910 480 17022 0 FreeSans 1400 0 0 0 gpio_analog[17]
port 9 nsew
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1400 0 0 0 gpio_analog[3]
port 12 nsew
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1400 0 0 0 gpio_analog[4]
port 13 nsew
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1400 0 0 0 gpio_analog[5]
port 14 nsew
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1400 0 0 0 gpio_analog[6]
port 15 nsew
flabel metal3 s -800 511530 480 511642 0 FreeSans 1400 0 0 0 gpio_analog[7]
port 16 nsew
flabel metal3 s -800 468308 480 468420 0 FreeSans 1400 0 0 0 gpio_analog[8]
port 17 nsew
flabel metal3 s -800 425086 480 425198 0 FreeSans 1400 0 0 0 gpio_analog[9]
port 18 nsew
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1400 0 0 0 gpio_noesd[0]
port 19 nsew
flabel metal3 s -800 380682 480 380794 0 FreeSans 1400 0 0 0 gpio_noesd[10]
port 20 nsew
flabel metal3 s -800 337460 480 337572 0 FreeSans 1400 0 0 0 gpio_noesd[11]
port 21 nsew
flabel metal3 s -800 294238 480 294350 0 FreeSans 1400 0 0 0 gpio_noesd[12]
port 22 nsew
flabel metal3 s -800 251216 480 251328 0 FreeSans 1400 0 0 0 gpio_noesd[13]
port 23 nsew
flabel metal3 s -800 123594 480 123706 0 FreeSans 1400 0 0 0 gpio_noesd[14]
port 24 nsew
flabel metal3 s -800 80372 480 80484 0 FreeSans 1400 0 0 0 gpio_noesd[15]
port 25 nsew
flabel metal3 s -800 37150 480 37262 0 FreeSans 1400 0 0 0 gpio_noesd[16]
port 26 nsew
flabel metal3 s -800 15728 480 15840 0 FreeSans 1400 0 0 0 gpio_noesd[17]
port 27 nsew
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1400 0 0 0 gpio_noesd[1]
port 28 nsew
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1400 0 0 0 gpio_noesd[2]
port 29 nsew
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1400 0 0 0 gpio_noesd[3]
port 30 nsew
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1400 0 0 0 gpio_noesd[4]
port 31 nsew
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1400 0 0 0 gpio_noesd[5]
port 32 nsew
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1400 0 0 0 gpio_noesd[6]
port 33 nsew
flabel metal3 s -800 510348 480 510460 0 FreeSans 1400 0 0 0 gpio_noesd[7]
port 34 nsew
flabel metal3 s -800 467126 480 467238 0 FreeSans 1400 0 0 0 gpio_noesd[8]
port 35 nsew
flabel metal3 s -800 423904 480 424016 0 FreeSans 1400 0 0 0 gpio_noesd[9]
port 36 nsew
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1400 0 0 0 io_analog[0]
port 37 nsew
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1400 0 0 0 io_analog[10]
port 38 nsew
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 2400 180 0 0 io_analog[1]
port 39 nsew
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 2400 180 0 0 io_analog[2]
port 40 nsew
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 2400 180 0 0 io_analog[3]
port 41 nsew
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 2400 180 0 0 io_analog[7]
port 45 nsew
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 2400 180 0 0 io_analog[8]
port 46 nsew
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 2400 180 0 0 io_analog[9]
port 47 nsew
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 2400 180 0 0 io_clamp_high[0]
port 48 nsew
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 2400 180 0 0 io_clamp_high[1]
port 49 nsew
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 2400 180 0 0 io_clamp_high[2]
port 50 nsew
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 2400 180 0 0 io_clamp_low[0]
port 51 nsew
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 2400 180 0 0 io_clamp_low[1]
port 52 nsew
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 2400 180 0 0 io_clamp_low[2]
port 53 nsew
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1400 0 0 0 io_in[0]
port 54 nsew
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1400 0 0 0 io_in[10]
port 55 nsew
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1400 0 0 0 io_in[11]
port 56 nsew
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1400 0 0 0 io_in[12]
port 57 nsew
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1400 0 0 0 io_in[13]
port 58 nsew
flabel metal3 s -800 507984 480 508096 0 FreeSans 1400 0 0 0 io_in[14]
port 59 nsew
flabel metal3 s -800 464762 480 464874 0 FreeSans 1400 0 0 0 io_in[15]
port 60 nsew
flabel metal3 s -800 421540 480 421652 0 FreeSans 1400 0 0 0 io_in[16]
port 61 nsew
flabel metal3 s -800 378318 480 378430 0 FreeSans 1400 0 0 0 io_in[17]
port 62 nsew
flabel metal3 s -800 335096 480 335208 0 FreeSans 1400 0 0 0 io_in[18]
port 63 nsew
flabel metal3 s -800 291874 480 291986 0 FreeSans 1400 0 0 0 io_in[19]
port 64 nsew
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1400 0 0 0 io_in[1]
port 65 nsew
flabel metal3 s -800 248852 480 248964 0 FreeSans 1400 0 0 0 io_in[20]
port 66 nsew
flabel metal3 s -800 121230 480 121342 0 FreeSans 1400 0 0 0 io_in[21]
port 67 nsew
flabel metal3 s -800 78008 480 78120 0 FreeSans 1400 0 0 0 io_in[22]
port 68 nsew
flabel metal3 s -800 34786 480 34898 0 FreeSans 1400 0 0 0 io_in[23]
port 69 nsew
flabel metal3 s -800 13364 480 13476 0 FreeSans 1400 0 0 0 io_in[24]
port 70 nsew
flabel metal3 s -800 8636 480 8748 0 FreeSans 1400 0 0 0 io_in[25]
port 71 nsew
flabel metal3 s -800 3908 480 4020 0 FreeSans 1400 0 0 0 io_in[26]
port 72 nsew
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1400 0 0 0 io_in[2]
port 73 nsew
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1400 0 0 0 io_in[3]
port 74 nsew
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1400 0 0 0 io_in[4]
port 75 nsew
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1400 0 0 0 io_in[5]
port 76 nsew
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1400 0 0 0 io_in[6]
port 77 nsew
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1400 0 0 0 io_in[7]
port 78 nsew
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1400 0 0 0 io_in[8]
port 79 nsew
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1400 0 0 0 io_in[9]
port 80 nsew
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1400 0 0 0 io_in_3v3[0]
port 81 nsew
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1400 0 0 0 io_in_3v3[10]
port 82 nsew
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1400 0 0 0 io_in_3v3[11]
port 83 nsew
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1400 0 0 0 io_in_3v3[12]
port 84 nsew
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1400 0 0 0 io_in_3v3[13]
port 85 nsew
flabel metal3 s -800 509166 480 509278 0 FreeSans 1400 0 0 0 io_in_3v3[14]
port 86 nsew
flabel metal3 s -800 465944 480 466056 0 FreeSans 1400 0 0 0 io_in_3v3[15]
port 87 nsew
flabel metal3 s -800 422722 480 422834 0 FreeSans 1400 0 0 0 io_in_3v3[16]
port 88 nsew
flabel metal3 s -800 379500 480 379612 0 FreeSans 1400 0 0 0 io_in_3v3[17]
port 89 nsew
flabel metal3 s -800 336278 480 336390 0 FreeSans 1400 0 0 0 io_in_3v3[18]
port 90 nsew
flabel metal3 s -800 293056 480 293168 0 FreeSans 1400 0 0 0 io_in_3v3[19]
port 91 nsew
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1400 0 0 0 io_in_3v3[1]
port 92 nsew
flabel metal3 s -800 250034 480 250146 0 FreeSans 1400 0 0 0 io_in_3v3[20]
port 93 nsew
flabel metal3 s -800 122412 480 122524 0 FreeSans 1400 0 0 0 io_in_3v3[21]
port 94 nsew
flabel metal3 s -800 79190 480 79302 0 FreeSans 1400 0 0 0 io_in_3v3[22]
port 95 nsew
flabel metal3 s -800 35968 480 36080 0 FreeSans 1400 0 0 0 io_in_3v3[23]
port 96 nsew
flabel metal3 s -800 14546 480 14658 0 FreeSans 1400 0 0 0 io_in_3v3[24]
port 97 nsew
flabel metal3 s -800 9818 480 9930 0 FreeSans 1400 0 0 0 io_in_3v3[25]
port 98 nsew
flabel metal3 s -800 5090 480 5202 0 FreeSans 1400 0 0 0 io_in_3v3[26]
port 99 nsew
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1400 0 0 0 io_in_3v3[2]
port 100 nsew
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1400 0 0 0 io_in_3v3[3]
port 101 nsew
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1400 0 0 0 io_in_3v3[4]
port 102 nsew
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1400 0 0 0 io_in_3v3[5]
port 103 nsew
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1400 0 0 0 io_in_3v3[6]
port 104 nsew
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1400 0 0 0 io_in_3v3[7]
port 105 nsew
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1400 0 0 0 io_in_3v3[8]
port 106 nsew
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1400 0 0 0 io_in_3v3[9]
port 107 nsew
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1400 0 0 0 io_oeb[0]
port 108 nsew
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1400 0 0 0 io_oeb[10]
port 109 nsew
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1400 0 0 0 io_oeb[11]
port 110 nsew
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1400 0 0 0 io_oeb[12]
port 111 nsew
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1400 0 0 0 io_oeb[13]
port 112 nsew
flabel metal3 s -800 505620 480 505732 0 FreeSans 1400 0 0 0 io_oeb[14]
port 113 nsew
flabel metal3 s -800 462398 480 462510 0 FreeSans 1400 0 0 0 io_oeb[15]
port 114 nsew
flabel metal3 s -800 419176 480 419288 0 FreeSans 1400 0 0 0 io_oeb[16]
port 115 nsew
flabel metal3 s -800 375954 480 376066 0 FreeSans 1400 0 0 0 io_oeb[17]
port 116 nsew
flabel metal3 s -800 332732 480 332844 0 FreeSans 1400 0 0 0 io_oeb[18]
port 117 nsew
flabel metal3 s -800 289510 480 289622 0 FreeSans 1400 0 0 0 io_oeb[19]
port 118 nsew
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1400 0 0 0 io_oeb[1]
port 119 nsew
flabel metal3 s -800 246488 480 246600 0 FreeSans 1400 0 0 0 io_oeb[20]
port 120 nsew
flabel metal3 s -800 118866 480 118978 0 FreeSans 1400 0 0 0 io_oeb[21]
port 121 nsew
flabel metal3 s -800 75644 480 75756 0 FreeSans 1400 0 0 0 io_oeb[22]
port 122 nsew
flabel metal3 s -800 32422 480 32534 0 FreeSans 1400 0 0 0 io_oeb[23]
port 123 nsew
flabel metal3 s -800 11000 480 11112 0 FreeSans 1400 0 0 0 io_oeb[24]
port 124 nsew
flabel metal3 s -800 6272 480 6384 0 FreeSans 1400 0 0 0 io_oeb[25]
port 125 nsew
flabel metal3 s -800 1544 480 1656 0 FreeSans 1400 0 0 0 io_oeb[26]
port 126 nsew
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1400 0 0 0 io_oeb[2]
port 127 nsew
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1400 0 0 0 io_oeb[3]
port 128 nsew
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1400 0 0 0 io_oeb[4]
port 129 nsew
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1400 0 0 0 io_oeb[5]
port 130 nsew
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1400 0 0 0 io_oeb[6]
port 131 nsew
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1400 0 0 0 io_oeb[7]
port 132 nsew
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1400 0 0 0 io_oeb[8]
port 133 nsew
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1400 0 0 0 io_oeb[9]
port 134 nsew
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1400 0 0 0 io_out[0]
port 135 nsew
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1400 0 0 0 io_out[10]
port 136 nsew
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1400 0 0 0 io_out[11]
port 137 nsew
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1400 0 0 0 io_out[12]
port 138 nsew
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1400 0 0 0 io_out[13]
port 139 nsew
flabel metal3 s -800 506802 480 506914 0 FreeSans 1400 0 0 0 io_out[14]
port 140 nsew
flabel metal3 s -800 463580 480 463692 0 FreeSans 1400 0 0 0 io_out[15]
port 141 nsew
flabel metal3 s -800 420358 480 420470 0 FreeSans 1400 0 0 0 io_out[16]
port 142 nsew
flabel metal3 s -800 377136 480 377248 0 FreeSans 1400 0 0 0 io_out[17]
port 143 nsew
flabel metal3 s -800 333914 480 334026 0 FreeSans 1400 0 0 0 io_out[18]
port 144 nsew
flabel metal3 s -800 290692 480 290804 0 FreeSans 1400 0 0 0 io_out[19]
port 145 nsew
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1400 0 0 0 io_out[1]
port 146 nsew
flabel metal3 s -800 247670 480 247782 0 FreeSans 1400 0 0 0 io_out[20]
port 147 nsew
flabel metal3 s -800 120048 480 120160 0 FreeSans 1400 0 0 0 io_out[21]
port 148 nsew
flabel metal3 s -800 76826 480 76938 0 FreeSans 1400 0 0 0 io_out[22]
port 149 nsew
flabel metal3 s -800 33604 480 33716 0 FreeSans 1400 0 0 0 io_out[23]
port 150 nsew
flabel metal3 s -800 12182 480 12294 0 FreeSans 1400 0 0 0 io_out[24]
port 151 nsew
flabel metal3 s -800 7454 480 7566 0 FreeSans 1400 0 0 0 io_out[25]
port 152 nsew
flabel metal3 s -800 2726 480 2838 0 FreeSans 1400 0 0 0 io_out[26]
port 153 nsew
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1400 0 0 0 io_out[2]
port 154 nsew
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1400 0 0 0 io_out[3]
port 155 nsew
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1400 0 0 0 io_out[4]
port 156 nsew
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1400 0 0 0 io_out[5]
port 157 nsew
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1400 0 0 0 io_out[6]
port 158 nsew
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1400 0 0 0 io_out[7]
port 159 nsew
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1400 0 0 0 io_out[8]
port 160 nsew
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1400 0 0 0 io_out[9]
port 161 nsew
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1400 90 0 0 la_data_in[0]
port 162 nsew
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1400 90 0 0 la_data_in[100]
port 163 nsew
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1400 90 0 0 la_data_in[101]
port 164 nsew
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1400 90 0 0 la_data_in[102]
port 165 nsew
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1400 90 0 0 la_data_in[103]
port 166 nsew
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1400 90 0 0 la_data_in[104]
port 167 nsew
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1400 90 0 0 la_data_in[105]
port 168 nsew
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1400 90 0 0 la_data_in[106]
port 169 nsew
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1400 90 0 0 la_data_in[107]
port 170 nsew
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1400 90 0 0 la_data_in[108]
port 171 nsew
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1400 90 0 0 la_data_in[109]
port 172 nsew
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1400 90 0 0 la_data_in[10]
port 173 nsew
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1400 90 0 0 la_data_in[110]
port 174 nsew
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1400 90 0 0 la_data_in[111]
port 175 nsew
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1400 90 0 0 la_data_in[112]
port 176 nsew
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1400 90 0 0 la_data_in[113]
port 177 nsew
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1400 90 0 0 la_data_in[114]
port 178 nsew
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1400 90 0 0 la_data_in[115]
port 179 nsew
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1400 90 0 0 la_data_in[116]
port 180 nsew
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1400 90 0 0 la_data_in[117]
port 181 nsew
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1400 90 0 0 la_data_in[118]
port 182 nsew
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1400 90 0 0 la_data_in[119]
port 183 nsew
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1400 90 0 0 la_data_in[11]
port 184 nsew
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1400 90 0 0 la_data_in[120]
port 185 nsew
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1400 90 0 0 la_data_in[121]
port 186 nsew
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1400 90 0 0 la_data_in[122]
port 187 nsew
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1400 90 0 0 la_data_in[123]
port 188 nsew
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1400 90 0 0 la_data_in[124]
port 189 nsew
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1400 90 0 0 la_data_in[125]
port 190 nsew
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1400 90 0 0 la_data_in[126]
port 191 nsew
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1400 90 0 0 la_data_in[127]
port 192 nsew
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1400 90 0 0 la_data_in[12]
port 193 nsew
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1400 90 0 0 la_data_in[13]
port 194 nsew
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1400 90 0 0 la_data_in[14]
port 195 nsew
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1400 90 0 0 la_data_in[15]
port 196 nsew
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1400 90 0 0 la_data_in[16]
port 197 nsew
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1400 90 0 0 la_data_in[17]
port 198 nsew
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1400 90 0 0 la_data_in[18]
port 199 nsew
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1400 90 0 0 la_data_in[19]
port 200 nsew
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1400 90 0 0 la_data_in[1]
port 201 nsew
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1400 90 0 0 la_data_in[20]
port 202 nsew
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1400 90 0 0 la_data_in[21]
port 203 nsew
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1400 90 0 0 la_data_in[22]
port 204 nsew
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1400 90 0 0 la_data_in[23]
port 205 nsew
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1400 90 0 0 la_data_in[24]
port 206 nsew
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1400 90 0 0 la_data_in[25]
port 207 nsew
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1400 90 0 0 la_data_in[26]
port 208 nsew
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1400 90 0 0 la_data_in[27]
port 209 nsew
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1400 90 0 0 la_data_in[28]
port 210 nsew
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1400 90 0 0 la_data_in[29]
port 211 nsew
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1400 90 0 0 la_data_in[2]
port 212 nsew
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1400 90 0 0 la_data_in[30]
port 213 nsew
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1400 90 0 0 la_data_in[31]
port 214 nsew
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1400 90 0 0 la_data_in[32]
port 215 nsew
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1400 90 0 0 la_data_in[33]
port 216 nsew
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1400 90 0 0 la_data_in[34]
port 217 nsew
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1400 90 0 0 la_data_in[35]
port 218 nsew
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1400 90 0 0 la_data_in[36]
port 219 nsew
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1400 90 0 0 la_data_in[37]
port 220 nsew
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1400 90 0 0 la_data_in[38]
port 221 nsew
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1400 90 0 0 la_data_in[39]
port 222 nsew
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1400 90 0 0 la_data_in[3]
port 223 nsew
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1400 90 0 0 la_data_in[40]
port 224 nsew
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1400 90 0 0 la_data_in[41]
port 225 nsew
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1400 90 0 0 la_data_in[42]
port 226 nsew
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1400 90 0 0 la_data_in[43]
port 227 nsew
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1400 90 0 0 la_data_in[44]
port 228 nsew
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1400 90 0 0 la_data_in[45]
port 229 nsew
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1400 90 0 0 la_data_in[46]
port 230 nsew
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1400 90 0 0 la_data_in[47]
port 231 nsew
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1400 90 0 0 la_data_in[48]
port 232 nsew
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1400 90 0 0 la_data_in[49]
port 233 nsew
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1400 90 0 0 la_data_in[4]
port 234 nsew
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1400 90 0 0 la_data_in[50]
port 235 nsew
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1400 90 0 0 la_data_in[51]
port 236 nsew
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1400 90 0 0 la_data_in[52]
port 237 nsew
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1400 90 0 0 la_data_in[53]
port 238 nsew
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1400 90 0 0 la_data_in[54]
port 239 nsew
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1400 90 0 0 la_data_in[55]
port 240 nsew
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1400 90 0 0 la_data_in[56]
port 241 nsew
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1400 90 0 0 la_data_in[57]
port 242 nsew
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1400 90 0 0 la_data_in[58]
port 243 nsew
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1400 90 0 0 la_data_in[59]
port 244 nsew
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1400 90 0 0 la_data_in[5]
port 245 nsew
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1400 90 0 0 la_data_in[60]
port 246 nsew
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1400 90 0 0 la_data_in[61]
port 247 nsew
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1400 90 0 0 la_data_in[62]
port 248 nsew
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1400 90 0 0 la_data_in[63]
port 249 nsew
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1400 90 0 0 la_data_in[64]
port 250 nsew
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1400 90 0 0 la_data_in[65]
port 251 nsew
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1400 90 0 0 la_data_in[66]
port 252 nsew
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1400 90 0 0 la_data_in[67]
port 253 nsew
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1400 90 0 0 la_data_in[68]
port 254 nsew
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1400 90 0 0 la_data_in[69]
port 255 nsew
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1400 90 0 0 la_data_in[6]
port 256 nsew
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1400 90 0 0 la_data_in[70]
port 257 nsew
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1400 90 0 0 la_data_in[71]
port 258 nsew
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1400 90 0 0 la_data_in[72]
port 259 nsew
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1400 90 0 0 la_data_in[73]
port 260 nsew
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1400 90 0 0 la_data_in[74]
port 261 nsew
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1400 90 0 0 la_data_in[75]
port 262 nsew
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1400 90 0 0 la_data_in[76]
port 263 nsew
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1400 90 0 0 la_data_in[77]
port 264 nsew
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1400 90 0 0 la_data_in[78]
port 265 nsew
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1400 90 0 0 la_data_in[79]
port 266 nsew
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1400 90 0 0 la_data_in[7]
port 267 nsew
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1400 90 0 0 la_data_in[80]
port 268 nsew
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1400 90 0 0 la_data_in[81]
port 269 nsew
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1400 90 0 0 la_data_in[82]
port 270 nsew
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1400 90 0 0 la_data_in[83]
port 271 nsew
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1400 90 0 0 la_data_in[84]
port 272 nsew
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1400 90 0 0 la_data_in[85]
port 273 nsew
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1400 90 0 0 la_data_in[86]
port 274 nsew
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1400 90 0 0 la_data_in[87]
port 275 nsew
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1400 90 0 0 la_data_in[88]
port 276 nsew
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1400 90 0 0 la_data_in[89]
port 277 nsew
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1400 90 0 0 la_data_in[8]
port 278 nsew
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1400 90 0 0 la_data_in[90]
port 279 nsew
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1400 90 0 0 la_data_in[91]
port 280 nsew
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1400 90 0 0 la_data_in[92]
port 281 nsew
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1400 90 0 0 la_data_in[93]
port 282 nsew
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1400 90 0 0 la_data_in[94]
port 283 nsew
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1400 90 0 0 la_data_in[95]
port 284 nsew
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1400 90 0 0 la_data_in[96]
port 285 nsew
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1400 90 0 0 la_data_in[97]
port 286 nsew
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1400 90 0 0 la_data_in[98]
port 287 nsew
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1400 90 0 0 la_data_in[99]
port 288 nsew
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1400 90 0 0 la_data_in[9]
port 289 nsew
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1400 90 0 0 la_data_out[0]
port 290 nsew
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1400 90 0 0 la_data_out[100]
port 291 nsew
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1400 90 0 0 la_data_out[101]
port 292 nsew
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1400 90 0 0 la_data_out[102]
port 293 nsew
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1400 90 0 0 la_data_out[103]
port 294 nsew
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1400 90 0 0 la_data_out[104]
port 295 nsew
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1400 90 0 0 la_data_out[105]
port 296 nsew
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1400 90 0 0 la_data_out[106]
port 297 nsew
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1400 90 0 0 la_data_out[107]
port 298 nsew
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1400 90 0 0 la_data_out[108]
port 299 nsew
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1400 90 0 0 la_data_out[109]
port 300 nsew
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1400 90 0 0 la_data_out[10]
port 301 nsew
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1400 90 0 0 la_data_out[110]
port 302 nsew
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1400 90 0 0 la_data_out[111]
port 303 nsew
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1400 90 0 0 la_data_out[112]
port 304 nsew
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1400 90 0 0 la_data_out[113]
port 305 nsew
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1400 90 0 0 la_data_out[114]
port 306 nsew
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1400 90 0 0 la_data_out[115]
port 307 nsew
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1400 90 0 0 la_data_out[116]
port 308 nsew
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1400 90 0 0 la_data_out[117]
port 309 nsew
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1400 90 0 0 la_data_out[118]
port 310 nsew
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1400 90 0 0 la_data_out[119]
port 311 nsew
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1400 90 0 0 la_data_out[11]
port 312 nsew
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1400 90 0 0 la_data_out[120]
port 313 nsew
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1400 90 0 0 la_data_out[121]
port 314 nsew
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1400 90 0 0 la_data_out[122]
port 315 nsew
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1400 90 0 0 la_data_out[123]
port 316 nsew
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1400 90 0 0 la_data_out[124]
port 317 nsew
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1400 90 0 0 la_data_out[125]
port 318 nsew
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1400 90 0 0 la_data_out[126]
port 319 nsew
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1400 90 0 0 la_data_out[127]
port 320 nsew
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1400 90 0 0 la_data_out[12]
port 321 nsew
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1400 90 0 0 la_data_out[13]
port 322 nsew
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1400 90 0 0 la_data_out[14]
port 323 nsew
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1400 90 0 0 la_data_out[15]
port 324 nsew
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1400 90 0 0 la_data_out[16]
port 325 nsew
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1400 90 0 0 la_data_out[17]
port 326 nsew
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1400 90 0 0 la_data_out[18]
port 327 nsew
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1400 90 0 0 la_data_out[19]
port 328 nsew
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1400 90 0 0 la_data_out[1]
port 329 nsew
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1400 90 0 0 la_data_out[20]
port 330 nsew
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1400 90 0 0 la_data_out[21]
port 331 nsew
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1400 90 0 0 la_data_out[22]
port 332 nsew
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1400 90 0 0 la_data_out[23]
port 333 nsew
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1400 90 0 0 la_data_out[24]
port 334 nsew
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1400 90 0 0 la_data_out[25]
port 335 nsew
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1400 90 0 0 la_data_out[26]
port 336 nsew
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1400 90 0 0 la_data_out[27]
port 337 nsew
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1400 90 0 0 la_data_out[28]
port 338 nsew
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1400 90 0 0 la_data_out[29]
port 339 nsew
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1400 90 0 0 la_data_out[2]
port 340 nsew
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1400 90 0 0 la_data_out[30]
port 341 nsew
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1400 90 0 0 la_data_out[31]
port 342 nsew
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1400 90 0 0 la_data_out[32]
port 343 nsew
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1400 90 0 0 la_data_out[33]
port 344 nsew
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1400 90 0 0 la_data_out[34]
port 345 nsew
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1400 90 0 0 la_data_out[35]
port 346 nsew
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1400 90 0 0 la_data_out[36]
port 347 nsew
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1400 90 0 0 la_data_out[37]
port 348 nsew
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1400 90 0 0 la_data_out[38]
port 349 nsew
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1400 90 0 0 la_data_out[39]
port 350 nsew
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1400 90 0 0 la_data_out[3]
port 351 nsew
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1400 90 0 0 la_data_out[40]
port 352 nsew
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1400 90 0 0 la_data_out[41]
port 353 nsew
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1400 90 0 0 la_data_out[42]
port 354 nsew
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1400 90 0 0 la_data_out[43]
port 355 nsew
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1400 90 0 0 la_data_out[44]
port 356 nsew
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1400 90 0 0 la_data_out[45]
port 357 nsew
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1400 90 0 0 la_data_out[46]
port 358 nsew
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1400 90 0 0 la_data_out[47]
port 359 nsew
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1400 90 0 0 la_data_out[48]
port 360 nsew
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1400 90 0 0 la_data_out[49]
port 361 nsew
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1400 90 0 0 la_data_out[4]
port 362 nsew
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1400 90 0 0 la_data_out[50]
port 363 nsew
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1400 90 0 0 la_data_out[51]
port 364 nsew
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1400 90 0 0 la_data_out[52]
port 365 nsew
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1400 90 0 0 la_data_out[53]
port 366 nsew
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1400 90 0 0 la_data_out[54]
port 367 nsew
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1400 90 0 0 la_data_out[55]
port 368 nsew
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1400 90 0 0 la_data_out[56]
port 369 nsew
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1400 90 0 0 la_data_out[57]
port 370 nsew
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1400 90 0 0 la_data_out[58]
port 371 nsew
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1400 90 0 0 la_data_out[59]
port 372 nsew
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1400 90 0 0 la_data_out[5]
port 373 nsew
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1400 90 0 0 la_data_out[60]
port 374 nsew
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1400 90 0 0 la_data_out[61]
port 375 nsew
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1400 90 0 0 la_data_out[62]
port 376 nsew
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1400 90 0 0 la_data_out[63]
port 377 nsew
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1400 90 0 0 la_data_out[64]
port 378 nsew
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1400 90 0 0 la_data_out[65]
port 379 nsew
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1400 90 0 0 la_data_out[66]
port 380 nsew
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1400 90 0 0 la_data_out[67]
port 381 nsew
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1400 90 0 0 la_data_out[68]
port 382 nsew
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1400 90 0 0 la_data_out[69]
port 383 nsew
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1400 90 0 0 la_data_out[6]
port 384 nsew
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1400 90 0 0 la_data_out[70]
port 385 nsew
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1400 90 0 0 la_data_out[71]
port 386 nsew
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1400 90 0 0 la_data_out[72]
port 387 nsew
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1400 90 0 0 la_data_out[73]
port 388 nsew
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1400 90 0 0 la_data_out[74]
port 389 nsew
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1400 90 0 0 la_data_out[75]
port 390 nsew
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1400 90 0 0 la_data_out[76]
port 391 nsew
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1400 90 0 0 la_data_out[77]
port 392 nsew
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1400 90 0 0 la_data_out[78]
port 393 nsew
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1400 90 0 0 la_data_out[79]
port 394 nsew
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1400 90 0 0 la_data_out[7]
port 395 nsew
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1400 90 0 0 la_data_out[80]
port 396 nsew
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1400 90 0 0 la_data_out[81]
port 397 nsew
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1400 90 0 0 la_data_out[82]
port 398 nsew
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1400 90 0 0 la_data_out[83]
port 399 nsew
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1400 90 0 0 la_data_out[84]
port 400 nsew
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1400 90 0 0 la_data_out[85]
port 401 nsew
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1400 90 0 0 la_data_out[86]
port 402 nsew
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1400 90 0 0 la_data_out[87]
port 403 nsew
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1400 90 0 0 la_data_out[88]
port 404 nsew
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1400 90 0 0 la_data_out[89]
port 405 nsew
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1400 90 0 0 la_data_out[8]
port 406 nsew
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1400 90 0 0 la_data_out[90]
port 407 nsew
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1400 90 0 0 la_data_out[91]
port 408 nsew
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1400 90 0 0 la_data_out[92]
port 409 nsew
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1400 90 0 0 la_data_out[93]
port 410 nsew
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1400 90 0 0 la_data_out[94]
port 411 nsew
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1400 90 0 0 la_data_out[95]
port 412 nsew
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1400 90 0 0 la_data_out[96]
port 413 nsew
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1400 90 0 0 la_data_out[97]
port 414 nsew
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1400 90 0 0 la_data_out[98]
port 415 nsew
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1400 90 0 0 la_data_out[99]
port 416 nsew
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1400 90 0 0 la_data_out[9]
port 417 nsew
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1400 90 0 0 la_oenb[0]
port 418 nsew
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1400 90 0 0 la_oenb[100]
port 419 nsew
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1400 90 0 0 la_oenb[101]
port 420 nsew
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1400 90 0 0 la_oenb[102]
port 421 nsew
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1400 90 0 0 la_oenb[103]
port 422 nsew
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1400 90 0 0 la_oenb[104]
port 423 nsew
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1400 90 0 0 la_oenb[105]
port 424 nsew
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1400 90 0 0 la_oenb[106]
port 425 nsew
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1400 90 0 0 la_oenb[107]
port 426 nsew
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1400 90 0 0 la_oenb[108]
port 427 nsew
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1400 90 0 0 la_oenb[109]
port 428 nsew
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1400 90 0 0 la_oenb[10]
port 429 nsew
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1400 90 0 0 la_oenb[110]
port 430 nsew
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1400 90 0 0 la_oenb[111]
port 431 nsew
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1400 90 0 0 la_oenb[112]
port 432 nsew
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1400 90 0 0 la_oenb[113]
port 433 nsew
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1400 90 0 0 la_oenb[114]
port 434 nsew
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1400 90 0 0 la_oenb[115]
port 435 nsew
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1400 90 0 0 la_oenb[116]
port 436 nsew
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1400 90 0 0 la_oenb[117]
port 437 nsew
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1400 90 0 0 la_oenb[118]
port 438 nsew
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1400 90 0 0 la_oenb[119]
port 439 nsew
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1400 90 0 0 la_oenb[11]
port 440 nsew
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1400 90 0 0 la_oenb[120]
port 441 nsew
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1400 90 0 0 la_oenb[121]
port 442 nsew
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1400 90 0 0 la_oenb[122]
port 443 nsew
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1400 90 0 0 la_oenb[123]
port 444 nsew
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1400 90 0 0 la_oenb[124]
port 445 nsew
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1400 90 0 0 la_oenb[125]
port 446 nsew
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1400 90 0 0 la_oenb[126]
port 447 nsew
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1400 90 0 0 la_oenb[127]
port 448 nsew
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1400 90 0 0 la_oenb[12]
port 449 nsew
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1400 90 0 0 la_oenb[13]
port 450 nsew
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1400 90 0 0 la_oenb[14]
port 451 nsew
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1400 90 0 0 la_oenb[15]
port 452 nsew
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1400 90 0 0 la_oenb[16]
port 453 nsew
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1400 90 0 0 la_oenb[17]
port 454 nsew
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1400 90 0 0 la_oenb[18]
port 455 nsew
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1400 90 0 0 la_oenb[19]
port 456 nsew
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1400 90 0 0 la_oenb[1]
port 457 nsew
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1400 90 0 0 la_oenb[20]
port 458 nsew
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1400 90 0 0 la_oenb[21]
port 459 nsew
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1400 90 0 0 la_oenb[22]
port 460 nsew
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1400 90 0 0 la_oenb[23]
port 461 nsew
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1400 90 0 0 la_oenb[24]
port 462 nsew
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1400 90 0 0 la_oenb[25]
port 463 nsew
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1400 90 0 0 la_oenb[26]
port 464 nsew
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1400 90 0 0 la_oenb[27]
port 465 nsew
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1400 90 0 0 la_oenb[28]
port 466 nsew
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1400 90 0 0 la_oenb[29]
port 467 nsew
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1400 90 0 0 la_oenb[2]
port 468 nsew
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1400 90 0 0 la_oenb[30]
port 469 nsew
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1400 90 0 0 la_oenb[31]
port 470 nsew
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1400 90 0 0 la_oenb[32]
port 471 nsew
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1400 90 0 0 la_oenb[33]
port 472 nsew
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1400 90 0 0 la_oenb[34]
port 473 nsew
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1400 90 0 0 la_oenb[35]
port 474 nsew
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1400 90 0 0 la_oenb[36]
port 475 nsew
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1400 90 0 0 la_oenb[37]
port 476 nsew
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1400 90 0 0 la_oenb[38]
port 477 nsew
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1400 90 0 0 la_oenb[39]
port 478 nsew
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1400 90 0 0 la_oenb[3]
port 479 nsew
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1400 90 0 0 la_oenb[40]
port 480 nsew
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1400 90 0 0 la_oenb[41]
port 481 nsew
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1400 90 0 0 la_oenb[42]
port 482 nsew
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1400 90 0 0 la_oenb[43]
port 483 nsew
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1400 90 0 0 la_oenb[44]
port 484 nsew
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1400 90 0 0 la_oenb[45]
port 485 nsew
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1400 90 0 0 la_oenb[46]
port 486 nsew
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1400 90 0 0 la_oenb[47]
port 487 nsew
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1400 90 0 0 la_oenb[48]
port 488 nsew
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1400 90 0 0 la_oenb[49]
port 489 nsew
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1400 90 0 0 la_oenb[4]
port 490 nsew
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1400 90 0 0 la_oenb[50]
port 491 nsew
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1400 90 0 0 la_oenb[51]
port 492 nsew
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1400 90 0 0 la_oenb[52]
port 493 nsew
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1400 90 0 0 la_oenb[53]
port 494 nsew
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1400 90 0 0 la_oenb[54]
port 495 nsew
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1400 90 0 0 la_oenb[55]
port 496 nsew
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1400 90 0 0 la_oenb[56]
port 497 nsew
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1400 90 0 0 la_oenb[57]
port 498 nsew
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1400 90 0 0 la_oenb[58]
port 499 nsew
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1400 90 0 0 la_oenb[59]
port 500 nsew
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1400 90 0 0 la_oenb[5]
port 501 nsew
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1400 90 0 0 la_oenb[60]
port 502 nsew
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1400 90 0 0 la_oenb[61]
port 503 nsew
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1400 90 0 0 la_oenb[62]
port 504 nsew
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1400 90 0 0 la_oenb[63]
port 505 nsew
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1400 90 0 0 la_oenb[64]
port 506 nsew
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1400 90 0 0 la_oenb[65]
port 507 nsew
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1400 90 0 0 la_oenb[66]
port 508 nsew
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1400 90 0 0 la_oenb[67]
port 509 nsew
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1400 90 0 0 la_oenb[68]
port 510 nsew
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1400 90 0 0 la_oenb[69]
port 511 nsew
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1400 90 0 0 la_oenb[6]
port 512 nsew
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1400 90 0 0 la_oenb[70]
port 513 nsew
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1400 90 0 0 la_oenb[71]
port 514 nsew
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1400 90 0 0 la_oenb[72]
port 515 nsew
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1400 90 0 0 la_oenb[73]
port 516 nsew
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1400 90 0 0 la_oenb[74]
port 517 nsew
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1400 90 0 0 la_oenb[75]
port 518 nsew
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1400 90 0 0 la_oenb[76]
port 519 nsew
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1400 90 0 0 la_oenb[77]
port 520 nsew
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1400 90 0 0 la_oenb[78]
port 521 nsew
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1400 90 0 0 la_oenb[79]
port 522 nsew
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1400 90 0 0 la_oenb[7]
port 523 nsew
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1400 90 0 0 la_oenb[80]
port 524 nsew
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1400 90 0 0 la_oenb[81]
port 525 nsew
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1400 90 0 0 la_oenb[82]
port 526 nsew
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1400 90 0 0 la_oenb[83]
port 527 nsew
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1400 90 0 0 la_oenb[84]
port 528 nsew
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1400 90 0 0 la_oenb[85]
port 529 nsew
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1400 90 0 0 la_oenb[86]
port 530 nsew
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1400 90 0 0 la_oenb[87]
port 531 nsew
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1400 90 0 0 la_oenb[88]
port 532 nsew
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1400 90 0 0 la_oenb[89]
port 533 nsew
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1400 90 0 0 la_oenb[8]
port 534 nsew
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1400 90 0 0 la_oenb[90]
port 535 nsew
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1400 90 0 0 la_oenb[91]
port 536 nsew
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1400 90 0 0 la_oenb[92]
port 537 nsew
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1400 90 0 0 la_oenb[93]
port 538 nsew
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1400 90 0 0 la_oenb[94]
port 539 nsew
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1400 90 0 0 la_oenb[95]
port 540 nsew
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1400 90 0 0 la_oenb[96]
port 541 nsew
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1400 90 0 0 la_oenb[97]
port 542 nsew
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1400 90 0 0 la_oenb[98]
port 543 nsew
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1400 90 0 0 la_oenb[99]
port 544 nsew
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1400 90 0 0 la_oenb[9]
port 545 nsew
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1400 90 0 0 user_clock2
port 546 nsew
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1400 90 0 0 user_irq[0]
port 547 nsew
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1400 90 0 0 user_irq[1]
port 548 nsew
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1400 90 0 0 user_irq[2]
port 549 nsew
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1400 0 0 0 vccd1
port 550 nsew
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1400 0 0 0 vccd1
port 550 nsew
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1400 0 0 0 vccd2
port 551 nsew
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1400 0 0 0 vccd2
port 551 nsew
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1400 0 0 0 vdda2
port 553 nsew
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1400 0 0 0 vdda2
port 553 nsew
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1400 0 0 0 vssd1
port 556 nsew
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1400 0 0 0 vssd1
port 556 nsew
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1400 0 0 0 vssd2
port 557 nsew
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1400 0 0 0 vssd2
port 557 nsew
flabel metal2 s 524 -800 636 480 0 FreeSans 1400 90 0 0 wb_clk_i
port 558 nsew
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1400 90 0 0 wb_rst_i
port 559 nsew
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1400 90 0 0 wbs_ack_o
port 560 nsew
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1400 90 0 0 wbs_adr_i[0]
port 561 nsew
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1400 90 0 0 wbs_adr_i[10]
port 562 nsew
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1400 90 0 0 wbs_adr_i[11]
port 563 nsew
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1400 90 0 0 wbs_adr_i[12]
port 564 nsew
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1400 90 0 0 wbs_adr_i[13]
port 565 nsew
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1400 90 0 0 wbs_adr_i[14]
port 566 nsew
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1400 90 0 0 wbs_adr_i[15]
port 567 nsew
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1400 90 0 0 wbs_adr_i[16]
port 568 nsew
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1400 90 0 0 wbs_adr_i[17]
port 569 nsew
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1400 90 0 0 wbs_adr_i[18]
port 570 nsew
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1400 90 0 0 wbs_adr_i[19]
port 571 nsew
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1400 90 0 0 wbs_adr_i[1]
port 572 nsew
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1400 90 0 0 wbs_adr_i[20]
port 573 nsew
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1400 90 0 0 wbs_adr_i[21]
port 574 nsew
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1400 90 0 0 wbs_adr_i[22]
port 575 nsew
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1400 90 0 0 wbs_adr_i[23]
port 576 nsew
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1400 90 0 0 wbs_adr_i[24]
port 577 nsew
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1400 90 0 0 wbs_adr_i[25]
port 578 nsew
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1400 90 0 0 wbs_adr_i[26]
port 579 nsew
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1400 90 0 0 wbs_adr_i[27]
port 580 nsew
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1400 90 0 0 wbs_adr_i[28]
port 581 nsew
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1400 90 0 0 wbs_adr_i[29]
port 582 nsew
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1400 90 0 0 wbs_adr_i[2]
port 583 nsew
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1400 90 0 0 wbs_adr_i[30]
port 584 nsew
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1400 90 0 0 wbs_adr_i[31]
port 585 nsew
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1400 90 0 0 wbs_adr_i[3]
port 586 nsew
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1400 90 0 0 wbs_adr_i[4]
port 587 nsew
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1400 90 0 0 wbs_adr_i[5]
port 588 nsew
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1400 90 0 0 wbs_adr_i[6]
port 589 nsew
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1400 90 0 0 wbs_adr_i[7]
port 590 nsew
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1400 90 0 0 wbs_adr_i[8]
port 591 nsew
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1400 90 0 0 wbs_adr_i[9]
port 592 nsew
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1400 90 0 0 wbs_cyc_i
port 593 nsew
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1400 90 0 0 wbs_dat_i[0]
port 594 nsew
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1400 90 0 0 wbs_dat_i[10]
port 595 nsew
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1400 90 0 0 wbs_dat_i[11]
port 596 nsew
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1400 90 0 0 wbs_dat_i[12]
port 597 nsew
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1400 90 0 0 wbs_dat_i[13]
port 598 nsew
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1400 90 0 0 wbs_dat_i[14]
port 599 nsew
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1400 90 0 0 wbs_dat_i[15]
port 600 nsew
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1400 90 0 0 wbs_dat_i[16]
port 601 nsew
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1400 90 0 0 wbs_dat_i[17]
port 602 nsew
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1400 90 0 0 wbs_dat_i[18]
port 603 nsew
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1400 90 0 0 wbs_dat_i[19]
port 604 nsew
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1400 90 0 0 wbs_dat_i[1]
port 605 nsew
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1400 90 0 0 wbs_dat_i[20]
port 606 nsew
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1400 90 0 0 wbs_dat_i[21]
port 607 nsew
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1400 90 0 0 wbs_dat_i[22]
port 608 nsew
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1400 90 0 0 wbs_dat_i[23]
port 609 nsew
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1400 90 0 0 wbs_dat_i[24]
port 610 nsew
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1400 90 0 0 wbs_dat_i[25]
port 611 nsew
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1400 90 0 0 wbs_dat_i[26]
port 612 nsew
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1400 90 0 0 wbs_dat_i[27]
port 613 nsew
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1400 90 0 0 wbs_dat_i[28]
port 614 nsew
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1400 90 0 0 wbs_dat_i[29]
port 615 nsew
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1400 90 0 0 wbs_dat_i[2]
port 616 nsew
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1400 90 0 0 wbs_dat_i[30]
port 617 nsew
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1400 90 0 0 wbs_dat_i[31]
port 618 nsew
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1400 90 0 0 wbs_dat_i[3]
port 619 nsew
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1400 90 0 0 wbs_dat_i[4]
port 620 nsew
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1400 90 0 0 wbs_dat_i[5]
port 621 nsew
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1400 90 0 0 wbs_dat_i[6]
port 622 nsew
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1400 90 0 0 wbs_dat_i[7]
port 623 nsew
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1400 90 0 0 wbs_dat_i[8]
port 624 nsew
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1400 90 0 0 wbs_dat_i[9]
port 625 nsew
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1400 90 0 0 wbs_dat_o[0]
port 626 nsew
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1400 90 0 0 wbs_dat_o[10]
port 627 nsew
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1400 90 0 0 wbs_dat_o[11]
port 628 nsew
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1400 90 0 0 wbs_dat_o[12]
port 629 nsew
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1400 90 0 0 wbs_dat_o[13]
port 630 nsew
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1400 90 0 0 wbs_dat_o[14]
port 631 nsew
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1400 90 0 0 wbs_dat_o[15]
port 632 nsew
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1400 90 0 0 wbs_dat_o[16]
port 633 nsew
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1400 90 0 0 wbs_dat_o[17]
port 634 nsew
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1400 90 0 0 wbs_dat_o[18]
port 635 nsew
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1400 90 0 0 wbs_dat_o[19]
port 636 nsew
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1400 90 0 0 wbs_dat_o[1]
port 637 nsew
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1400 90 0 0 wbs_dat_o[20]
port 638 nsew
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1400 90 0 0 wbs_dat_o[21]
port 639 nsew
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1400 90 0 0 wbs_dat_o[22]
port 640 nsew
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1400 90 0 0 wbs_dat_o[23]
port 641 nsew
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1400 90 0 0 wbs_dat_o[24]
port 642 nsew
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1400 90 0 0 wbs_dat_o[25]
port 643 nsew
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1400 90 0 0 wbs_dat_o[26]
port 644 nsew
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1400 90 0 0 wbs_dat_o[27]
port 645 nsew
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1400 90 0 0 wbs_dat_o[28]
port 646 nsew
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1400 90 0 0 wbs_dat_o[29]
port 647 nsew
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1400 90 0 0 wbs_dat_o[2]
port 648 nsew
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1400 90 0 0 wbs_dat_o[30]
port 649 nsew
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1400 90 0 0 wbs_dat_o[31]
port 650 nsew
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1400 90 0 0 wbs_dat_o[3]
port 651 nsew
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1400 90 0 0 wbs_dat_o[4]
port 652 nsew
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1400 90 0 0 wbs_dat_o[5]
port 653 nsew
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1400 90 0 0 wbs_dat_o[6]
port 654 nsew
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1400 90 0 0 wbs_dat_o[7]
port 655 nsew
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1400 90 0 0 wbs_dat_o[8]
port 656 nsew
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1400 90 0 0 wbs_dat_o[9]
port 657 nsew
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1400 90 0 0 wbs_sel_i[0]
port 658 nsew
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1400 90 0 0 wbs_sel_i[1]
port 659 nsew
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1400 90 0 0 wbs_sel_i[2]
port 660 nsew
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1400 90 0 0 wbs_sel_i[3]
port 661 nsew
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1400 90 0 0 wbs_stb_i
port 662 nsew
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1400 90 0 0 wbs_we_i
port 663 nsew
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1400 0 0 0 gpio_analog[0]
port 1 nsew
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1400 0 0 0 gpio_analog[1]
port 10 nsew
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1400 0 0 0 gpio_analog[2]
port 11 nsew
rlabel space 168881 180777 169101 181177 1 COL_SEL0
port 253 n
rlabel space 171881 180777 172101 181177 1 COL_SEL0
port 253 n
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 2400 180 0 0 vssa1
port 554 nsew
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1400 0 0 0 vssa1
port 554 nsew
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1400 0 0 0 vssa1
port 554 nsew
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 2400 180 0 0 vssa1
port 554 nsew
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1400 0 0 0 vssa2
port 555 nsew
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1400 0 0 0 vssa2
port 555 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
